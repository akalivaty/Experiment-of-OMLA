//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 1 0 0 0 1 1 0 1 0 0 0 1 1 1 1 1 1 0 1 1 0 0 1 1 1 0 0 0 0 1 0 1 1 1 0 1 0 0 1 1 1 1 0 1 0 0 1 1 0 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:12 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n703, new_n704, new_n705, new_n706,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n755, new_n756, new_n757, new_n758, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039;
  INV_X1    g000(.A(G221), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT9), .B(G234), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G902), .ZN(new_n190));
  AOI21_X1  g004(.A(new_n187), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G469), .ZN(new_n192));
  XNOR2_X1  g006(.A(G110), .B(G140), .ZN(new_n193));
  INV_X1    g007(.A(G953), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G227), .ZN(new_n195));
  XOR2_X1   g009(.A(new_n193), .B(new_n195), .Z(new_n196));
  INV_X1    g010(.A(G128), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n197), .A2(KEYINPUT1), .ZN(new_n198));
  INV_X1    g012(.A(G146), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G143), .ZN(new_n200));
  INV_X1    g014(.A(G143), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G146), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n198), .A2(new_n200), .A3(new_n202), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n197), .B1(new_n200), .B2(KEYINPUT1), .ZN(new_n204));
  XNOR2_X1  g018(.A(G143), .B(G146), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n203), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G101), .ZN(new_n207));
  INV_X1    g021(.A(G107), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(KEYINPUT71), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT71), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G107), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G104), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n208), .A2(G104), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n207), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  XNOR2_X1  g030(.A(KEYINPUT71), .B(G107), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n213), .A2(KEYINPUT3), .ZN(new_n218));
  AOI22_X1  g032(.A1(new_n217), .A2(new_n218), .B1(KEYINPUT3), .B2(new_n215), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT72), .ZN(new_n220));
  AOI21_X1  g034(.A(G101), .B1(new_n213), .B2(G107), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n218), .A2(new_n209), .A3(new_n211), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n215), .A2(KEYINPUT3), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n223), .A2(new_n224), .A3(new_n221), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(KEYINPUT72), .ZN(new_n226));
  AOI211_X1 g040(.A(KEYINPUT75), .B(new_n216), .C1(new_n222), .C2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT75), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n222), .A2(new_n226), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n214), .A2(new_n215), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G101), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n228), .B1(new_n229), .B2(new_n231), .ZN(new_n232));
  OAI211_X1 g046(.A(KEYINPUT10), .B(new_n206), .C1(new_n227), .C2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(KEYINPUT0), .A2(G128), .ZN(new_n234));
  OR2_X1    g048(.A1(KEYINPUT0), .A2(G128), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n201), .A2(G146), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n199), .A2(G143), .ZN(new_n237));
  OAI211_X1 g051(.A(new_n234), .B(new_n235), .C1(new_n236), .C2(new_n237), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n200), .A2(new_n202), .A3(KEYINPUT0), .A4(G128), .ZN(new_n239));
  AND2_X1   g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT4), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n219), .B1(G104), .B2(new_n208), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G101), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n241), .B1(new_n243), .B2(new_n229), .ZN(new_n244));
  AOI21_X1  g058(.A(KEYINPUT4), .B1(new_n242), .B2(G101), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n240), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT11), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n247), .A2(G137), .ZN(new_n248));
  AND2_X1   g062(.A1(KEYINPUT64), .A2(G134), .ZN(new_n249));
  NOR2_X1   g063(.A1(KEYINPUT64), .A2(G134), .ZN(new_n250));
  NOR3_X1   g064(.A1(new_n248), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(G137), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n252), .A2(KEYINPUT11), .A3(G134), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n247), .A2(G137), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NOR3_X1   g069(.A1(new_n251), .A2(G131), .A3(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(G131), .ZN(new_n257));
  AND2_X1   g071(.A1(new_n253), .A2(new_n254), .ZN(new_n258));
  OR2_X1    g072(.A1(KEYINPUT64), .A2(G134), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n252), .A2(KEYINPUT11), .ZN(new_n260));
  NAND2_X1  g074(.A1(KEYINPUT64), .A2(G134), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n259), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n257), .B1(new_n258), .B2(new_n262), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n256), .A2(new_n263), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n216), .B1(new_n222), .B2(new_n226), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n200), .A2(KEYINPUT1), .ZN(new_n266));
  AND2_X1   g080(.A1(new_n266), .A2(KEYINPUT74), .ZN(new_n267));
  OAI21_X1  g081(.A(G128), .B1(new_n266), .B2(KEYINPUT74), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n269), .A2(new_n205), .ZN(new_n270));
  XNOR2_X1  g084(.A(new_n203), .B(KEYINPUT73), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n265), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT10), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n233), .A2(new_n246), .A3(new_n264), .A4(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n243), .A2(new_n241), .ZN(new_n277));
  AOI22_X1  g091(.A1(G101), .A2(new_n242), .B1(new_n222), .B2(new_n226), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n277), .B1(new_n278), .B2(new_n241), .ZN(new_n279));
  AOI22_X1  g093(.A1(new_n279), .A2(new_n240), .B1(new_n272), .B2(new_n273), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n264), .B1(new_n280), .B2(new_n233), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n196), .B1(new_n276), .B2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n196), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n220), .B1(new_n219), .B2(new_n221), .ZN(new_n284));
  AND4_X1   g098(.A1(new_n220), .A2(new_n223), .A3(new_n224), .A4(new_n221), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n231), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(KEYINPUT75), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n265), .A2(new_n228), .ZN(new_n288));
  INV_X1    g102(.A(new_n206), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n287), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(new_n272), .ZN(new_n291));
  INV_X1    g105(.A(new_n264), .ZN(new_n292));
  AOI21_X1  g106(.A(KEYINPUT12), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT12), .ZN(new_n294));
  AOI211_X1 g108(.A(new_n294), .B(new_n264), .C1(new_n290), .C2(new_n272), .ZN(new_n295));
  OAI211_X1 g109(.A(new_n275), .B(new_n283), .C1(new_n293), .C2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT76), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n282), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n291), .A2(new_n292), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(new_n294), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n291), .A2(KEYINPUT12), .A3(new_n292), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n275), .A2(new_n283), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(KEYINPUT76), .B1(new_n302), .B2(new_n304), .ZN(new_n305));
  OAI211_X1 g119(.A(new_n192), .B(new_n190), .C1(new_n298), .C2(new_n305), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n192), .A2(new_n190), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n303), .A2(new_n281), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n275), .B1(new_n293), .B2(new_n295), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n308), .B1(new_n196), .B2(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n307), .B1(new_n310), .B2(G469), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n191), .B1(new_n306), .B2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(G119), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(G116), .ZN(new_n314));
  OAI21_X1  g128(.A(G113), .B1(new_n314), .B2(KEYINPUT5), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(G116), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(G119), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n314), .A2(new_n318), .A3(KEYINPUT5), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n316), .A2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT2), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n321), .A2(G113), .ZN(new_n322));
  INV_X1    g136(.A(G113), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n323), .A2(KEYINPUT2), .ZN(new_n324));
  OAI211_X1 g138(.A(new_n314), .B(new_n318), .C1(new_n322), .C2(new_n324), .ZN(new_n325));
  AND2_X1   g139(.A1(new_n320), .A2(new_n325), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n326), .B1(new_n227), .B2(new_n232), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n314), .A2(new_n318), .ZN(new_n328));
  XNOR2_X1  g142(.A(KEYINPUT2), .B(G113), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n325), .A2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT65), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n325), .A2(new_n330), .A3(KEYINPUT65), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n335), .B1(new_n244), .B2(new_n245), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n327), .A2(new_n336), .ZN(new_n337));
  XNOR2_X1  g151(.A(G110), .B(G122), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n327), .A2(new_n336), .A3(new_n338), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n340), .A2(KEYINPUT6), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n238), .A2(new_n239), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(G125), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n344), .B1(G125), .B2(new_n206), .ZN(new_n345));
  INV_X1    g159(.A(G224), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n346), .A2(G953), .ZN(new_n347));
  XNOR2_X1  g161(.A(new_n347), .B(KEYINPUT77), .ZN(new_n348));
  XNOR2_X1  g162(.A(new_n345), .B(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT6), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n337), .A2(new_n350), .A3(new_n339), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n342), .A2(new_n349), .A3(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT78), .ZN(new_n353));
  XOR2_X1   g167(.A(new_n338), .B(KEYINPUT8), .Z(new_n354));
  NOR2_X1   g168(.A1(new_n265), .A2(new_n326), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n354), .B1(new_n327), .B2(new_n356), .ZN(new_n357));
  OAI21_X1  g171(.A(KEYINPUT7), .B1(new_n346), .B2(G953), .ZN(new_n358));
  XOR2_X1   g172(.A(new_n345), .B(new_n358), .Z(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n353), .B1(new_n357), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n287), .A2(new_n288), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n355), .B1(new_n362), .B2(new_n326), .ZN(new_n363));
  OAI211_X1 g177(.A(KEYINPUT78), .B(new_n359), .C1(new_n363), .C2(new_n354), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n361), .A2(new_n364), .A3(new_n341), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n352), .A2(new_n190), .A3(new_n365), .ZN(new_n366));
  OAI21_X1  g180(.A(G210), .B1(G237), .B2(G902), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  NAND4_X1  g183(.A1(new_n352), .A2(new_n365), .A3(new_n190), .A4(new_n367), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  OAI21_X1  g185(.A(G214), .B1(G237), .B2(G902), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n197), .A2(G143), .ZN(new_n373));
  XOR2_X1   g187(.A(KEYINPUT83), .B(KEYINPUT13), .Z(new_n374));
  INV_X1    g188(.A(KEYINPUT82), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n375), .B1(new_n197), .B2(G143), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n201), .A2(KEYINPUT82), .A3(G128), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n373), .B1(new_n374), .B2(new_n378), .ZN(new_n379));
  XNOR2_X1  g193(.A(KEYINPUT83), .B(KEYINPUT13), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n380), .B1(new_n376), .B2(new_n377), .ZN(new_n381));
  OAI21_X1  g195(.A(G134), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  XNOR2_X1  g196(.A(G116), .B(G122), .ZN(new_n383));
  OR2_X1    g197(.A1(new_n217), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n217), .A2(new_n383), .ZN(new_n385));
  AOI22_X1  g199(.A1(new_n376), .A2(new_n377), .B1(new_n197), .B2(G143), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n259), .A2(new_n261), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  AOI22_X1  g202(.A1(new_n384), .A2(new_n385), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n382), .A2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT14), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n383), .A2(new_n391), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n317), .A2(KEYINPUT14), .A3(G122), .ZN(new_n393));
  AND2_X1   g207(.A1(new_n393), .A2(G107), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n378), .A2(new_n373), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n396), .A2(new_n387), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n386), .A2(new_n388), .ZN(new_n398));
  OAI211_X1 g212(.A(new_n385), .B(new_n395), .C1(new_n397), .C2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(G217), .ZN(new_n400));
  NOR3_X1   g214(.A1(new_n188), .A2(new_n400), .A3(G953), .ZN(new_n401));
  AND3_X1   g215(.A1(new_n390), .A2(new_n399), .A3(new_n401), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n401), .B1(new_n390), .B2(new_n399), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n190), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(G478), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n405), .A2(KEYINPUT15), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  XNOR2_X1  g221(.A(new_n404), .B(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(G234), .ZN(new_n409));
  INV_X1    g223(.A(G237), .ZN(new_n410));
  OAI211_X1 g224(.A(G952), .B(new_n194), .C1(new_n409), .C2(new_n410), .ZN(new_n411));
  XNOR2_X1  g225(.A(KEYINPUT21), .B(G898), .ZN(new_n412));
  XOR2_X1   g226(.A(new_n412), .B(KEYINPUT84), .Z(new_n413));
  OAI211_X1 g227(.A(G902), .B(G953), .C1(new_n409), .C2(new_n410), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n411), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  AND2_X1   g229(.A1(new_n408), .A2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(G140), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(G125), .ZN(new_n418));
  INV_X1    g232(.A(G125), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(G140), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT69), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n418), .A2(new_n420), .A3(KEYINPUT69), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n423), .A2(new_n199), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n421), .A2(G146), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NOR2_X1   g241(.A1(G237), .A2(G953), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(G214), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(new_n201), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n428), .A2(G143), .A3(G214), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT18), .ZN(new_n432));
  OAI211_X1 g246(.A(new_n430), .B(new_n431), .C1(new_n432), .C2(new_n257), .ZN(new_n433));
  INV_X1    g247(.A(new_n431), .ZN(new_n434));
  AOI21_X1  g248(.A(G143), .B1(new_n428), .B2(G214), .ZN(new_n435));
  OAI211_X1 g249(.A(KEYINPUT18), .B(G131), .C1(new_n434), .C2(new_n435), .ZN(new_n436));
  AND3_X1   g250(.A1(new_n427), .A2(new_n433), .A3(new_n436), .ZN(new_n437));
  NOR3_X1   g251(.A1(new_n419), .A2(KEYINPUT16), .A3(G140), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n418), .A2(new_n420), .A3(KEYINPUT16), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(new_n199), .ZN(new_n442));
  OAI211_X1 g256(.A(KEYINPUT17), .B(G131), .C1(new_n434), .C2(new_n435), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n439), .A2(new_n440), .A3(G146), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n442), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  OAI21_X1  g259(.A(G131), .B1(new_n434), .B2(new_n435), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n430), .A2(new_n257), .A3(new_n431), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT17), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n446), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n445), .B1(KEYINPUT81), .B2(new_n449), .ZN(new_n450));
  OR2_X1    g264(.A1(new_n449), .A2(KEYINPUT81), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n437), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  XNOR2_X1  g266(.A(G113), .B(G122), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n453), .B(new_n213), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n452), .A2(new_n454), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n190), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(G475), .ZN(new_n459));
  NOR2_X1   g273(.A1(G475), .A2(G902), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT19), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n423), .A2(new_n462), .A3(new_n424), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n421), .A2(KEYINPUT19), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n463), .A2(new_n199), .A3(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT79), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND4_X1  g281(.A1(new_n463), .A2(KEYINPUT79), .A3(new_n199), .A4(new_n464), .ZN(new_n468));
  XNOR2_X1  g282(.A(G125), .B(G140), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n438), .B1(new_n469), .B2(KEYINPUT16), .ZN(new_n470));
  AOI22_X1  g284(.A1(new_n446), .A2(new_n447), .B1(new_n470), .B2(G146), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n467), .A2(new_n468), .A3(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n427), .A2(new_n433), .A3(new_n436), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n454), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT80), .ZN(new_n475));
  AOI22_X1  g289(.A1(new_n474), .A2(new_n475), .B1(new_n452), .B2(new_n454), .ZN(new_n476));
  AND2_X1   g290(.A1(new_n468), .A2(new_n471), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n437), .B1(new_n477), .B2(new_n467), .ZN(new_n478));
  OAI21_X1  g292(.A(KEYINPUT80), .B1(new_n478), .B2(new_n454), .ZN(new_n479));
  AOI211_X1 g293(.A(KEYINPUT20), .B(new_n461), .C1(new_n476), .C2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT20), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n472), .A2(new_n473), .ZN(new_n482));
  INV_X1    g296(.A(new_n454), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n482), .A2(new_n475), .A3(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n479), .A2(new_n455), .A3(new_n484), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n481), .B1(new_n485), .B2(new_n460), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n416), .B(new_n459), .C1(new_n480), .C2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  AND3_X1   g302(.A1(new_n371), .A2(new_n372), .A3(new_n488), .ZN(new_n489));
  NOR2_X1   g303(.A1(G472), .A2(G902), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  OAI21_X1  g305(.A(G131), .B1(new_n251), .B2(new_n255), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n262), .A2(new_n257), .A3(new_n253), .A4(new_n254), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n343), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n257), .B1(G134), .B2(G137), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n495), .B1(new_n387), .B2(G137), .ZN(new_n496));
  AND3_X1   g310(.A1(new_n206), .A2(new_n493), .A3(new_n496), .ZN(new_n497));
  NOR3_X1   g311(.A1(new_n494), .A2(new_n497), .A3(KEYINPUT30), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT30), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n240), .B1(new_n256), .B2(new_n263), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n206), .A2(new_n493), .A3(new_n496), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n335), .B1(new_n498), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n428), .A2(G210), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n504), .B(KEYINPUT27), .ZN(new_n505));
  XNOR2_X1  g319(.A(KEYINPUT26), .B(G101), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n505), .B(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n334), .ZN(new_n508));
  AOI21_X1  g322(.A(KEYINPUT65), .B1(new_n325), .B2(new_n330), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n510), .A2(new_n500), .A3(new_n501), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n503), .A2(new_n507), .A3(new_n511), .ZN(new_n512));
  NOR3_X1   g326(.A1(new_n335), .A2(new_n494), .A3(new_n497), .ZN(new_n513));
  AOI22_X1  g327(.A1(new_n500), .A2(new_n501), .B1(new_n333), .B2(new_n334), .ZN(new_n514));
  OAI21_X1  g328(.A(KEYINPUT28), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT28), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n511), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n507), .ZN(new_n519));
  AOI22_X1  g333(.A1(KEYINPUT31), .A2(new_n512), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  OAI21_X1  g334(.A(KEYINPUT30), .B1(new_n494), .B2(new_n497), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n500), .A2(new_n499), .A3(new_n501), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n513), .B1(new_n523), .B2(new_n335), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT31), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n524), .A2(new_n525), .A3(new_n507), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n491), .B1(new_n520), .B2(new_n526), .ZN(new_n527));
  OAI21_X1  g341(.A(KEYINPUT66), .B1(new_n527), .B2(KEYINPUT32), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n512), .A2(KEYINPUT31), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n335), .B1(new_n494), .B2(new_n497), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n516), .B1(new_n511), .B2(new_n530), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n494), .A2(new_n497), .ZN(new_n532));
  AOI21_X1  g346(.A(KEYINPUT28), .B1(new_n532), .B2(new_n510), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n519), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n529), .A2(new_n526), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(new_n490), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT66), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT32), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  NOR3_X1   g353(.A1(new_n531), .A2(new_n533), .A3(new_n519), .ZN(new_n540));
  AOI21_X1  g354(.A(G902), .B1(new_n540), .B2(KEYINPUT29), .ZN(new_n541));
  NAND4_X1  g355(.A1(new_n515), .A2(KEYINPUT67), .A3(new_n507), .A4(new_n517), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT29), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n510), .B1(new_n521), .B2(new_n522), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n519), .B1(new_n544), .B2(new_n513), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n542), .A2(new_n543), .A3(new_n545), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n540), .A2(KEYINPUT67), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n541), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(G472), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n535), .A2(KEYINPUT32), .A3(new_n490), .ZN(new_n550));
  NAND4_X1  g364(.A1(new_n528), .A2(new_n539), .A3(new_n549), .A4(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n400), .B1(G234), .B2(new_n190), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n442), .A2(new_n444), .ZN(new_n554));
  OAI21_X1  g368(.A(KEYINPUT68), .B1(new_n313), .B2(G128), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT68), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n556), .A2(new_n197), .A3(G119), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n313), .A2(G128), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n555), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  XNOR2_X1  g373(.A(KEYINPUT24), .B(G110), .ZN(new_n560));
  OR2_X1    g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n197), .A2(KEYINPUT23), .A3(G119), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n313), .A2(G128), .ZN(new_n563));
  OAI211_X1 g377(.A(new_n558), .B(new_n562), .C1(new_n563), .C2(KEYINPUT23), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(G110), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n554), .A2(new_n561), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n559), .A2(new_n560), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n567), .B1(G110), .B2(new_n564), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n568), .A2(new_n425), .A3(new_n444), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n566), .A2(new_n569), .ZN(new_n570));
  XNOR2_X1  g384(.A(KEYINPUT22), .B(G137), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n194), .A2(G221), .A3(G234), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n571), .B(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n570), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n566), .A2(new_n569), .A3(new_n573), .ZN(new_n576));
  AND2_X1   g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n577), .A2(KEYINPUT25), .A3(new_n190), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n575), .A2(new_n190), .A3(new_n576), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT25), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n553), .B1(new_n578), .B2(new_n581), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n552), .A2(G902), .ZN(new_n583));
  AND2_X1   g397(.A1(new_n577), .A2(new_n583), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  AND3_X1   g399(.A1(new_n551), .A2(KEYINPUT70), .A3(new_n585), .ZN(new_n586));
  AOI21_X1  g400(.A(KEYINPUT70), .B1(new_n551), .B2(new_n585), .ZN(new_n587));
  OAI211_X1 g401(.A(new_n312), .B(new_n489), .C1(new_n586), .C2(new_n587), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n588), .B(G101), .ZN(G3));
  NAND2_X1  g403(.A1(new_n535), .A2(new_n190), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(G472), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(new_n536), .ZN(new_n592));
  INV_X1    g406(.A(new_n585), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n312), .A2(new_n594), .ZN(new_n595));
  XOR2_X1   g409(.A(new_n595), .B(KEYINPUT85), .Z(new_n596));
  INV_X1    g410(.A(new_n372), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n597), .B1(new_n369), .B2(new_n370), .ZN(new_n598));
  NAND2_X1  g412(.A1(KEYINPUT86), .A2(KEYINPUT33), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n599), .B1(new_n402), .B2(new_n403), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n390), .A2(new_n399), .ZN(new_n601));
  INV_X1    g415(.A(new_n401), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n390), .A2(new_n399), .A3(new_n401), .ZN(new_n604));
  XNOR2_X1  g418(.A(KEYINPUT86), .B(KEYINPUT33), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n405), .A2(G902), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n600), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT87), .ZN(new_n609));
  AND2_X1   g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n600), .A2(new_n606), .A3(KEYINPUT87), .A4(new_n607), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n404), .A2(new_n405), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g427(.A(KEYINPUT88), .B1(new_n610), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n608), .A2(new_n609), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT88), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n615), .A2(new_n616), .A3(new_n612), .A4(new_n611), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n614), .A2(new_n617), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n459), .B1(new_n480), .B2(new_n486), .ZN(new_n619));
  AND3_X1   g433(.A1(new_n618), .A2(new_n619), .A3(new_n415), .ZN(new_n620));
  AND2_X1   g434(.A1(new_n598), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n596), .A2(new_n621), .ZN(new_n622));
  XOR2_X1   g436(.A(KEYINPUT34), .B(G104), .Z(new_n623));
  XNOR2_X1  g437(.A(new_n622), .B(new_n623), .ZN(G6));
  NAND3_X1  g438(.A1(new_n485), .A2(new_n481), .A3(new_n460), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT89), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n480), .A2(new_n486), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n627), .B1(new_n628), .B2(new_n626), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT91), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n408), .B1(G475), .B2(new_n458), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n415), .B(KEYINPUT90), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n629), .A2(new_n630), .A3(new_n631), .A4(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n485), .A2(new_n460), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(KEYINPUT20), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n635), .A2(new_n626), .A3(new_n625), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n480), .A2(KEYINPUT89), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n636), .A2(new_n637), .A3(new_n631), .A4(new_n632), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(KEYINPUT91), .ZN(new_n639));
  AND3_X1   g453(.A1(new_n633), .A2(new_n598), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n596), .A2(new_n640), .ZN(new_n641));
  XOR2_X1   g455(.A(KEYINPUT35), .B(G107), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G9));
  NAND2_X1  g457(.A1(new_n578), .A2(new_n581), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(new_n552), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n574), .A2(KEYINPUT36), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n570), .B(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n583), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n645), .A2(KEYINPUT92), .A3(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT92), .ZN(new_n650));
  INV_X1    g464(.A(new_n648), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n650), .B1(new_n582), .B2(new_n651), .ZN(new_n652));
  AND2_X1   g466(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n653), .A2(new_n592), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n489), .A2(new_n312), .A3(new_n654), .ZN(new_n655));
  XOR2_X1   g469(.A(KEYINPUT37), .B(G110), .Z(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G12));
  NAND2_X1  g471(.A1(new_n649), .A2(new_n652), .ZN(new_n658));
  AND2_X1   g472(.A1(new_n551), .A2(new_n658), .ZN(new_n659));
  XOR2_X1   g473(.A(KEYINPUT93), .B(G900), .Z(new_n660));
  OAI21_X1  g474(.A(new_n411), .B1(new_n660), .B2(new_n414), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n629), .A2(new_n631), .A3(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n659), .A2(new_n663), .A3(new_n312), .A4(new_n598), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(G128), .ZN(G30));
  XNOR2_X1  g479(.A(new_n661), .B(KEYINPUT39), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n312), .A2(new_n666), .ZN(new_n667));
  XOR2_X1   g481(.A(new_n667), .B(KEYINPUT40), .Z(new_n668));
  INV_X1    g482(.A(new_n371), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(KEYINPUT38), .ZN(new_n670));
  INV_X1    g484(.A(new_n619), .ZN(new_n671));
  NOR4_X1   g485(.A1(new_n671), .A2(new_n658), .A3(new_n597), .A4(new_n408), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT38), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n371), .A2(new_n673), .ZN(new_n674));
  AND2_X1   g488(.A1(new_n528), .A2(new_n539), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n507), .B1(new_n544), .B2(new_n513), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n511), .A2(new_n530), .ZN(new_n677));
  OAI211_X1 g491(.A(new_n676), .B(new_n190), .C1(new_n507), .C2(new_n677), .ZN(new_n678));
  AOI22_X1  g492(.A1(new_n527), .A2(KEYINPUT32), .B1(G472), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n675), .A2(new_n679), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n670), .A2(new_n672), .A3(new_n674), .A4(new_n680), .ZN(new_n681));
  OR2_X1    g495(.A1(new_n681), .A2(KEYINPUT94), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n681), .A2(KEYINPUT94), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n668), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G143), .ZN(G45));
  AND3_X1   g499(.A1(new_n618), .A2(new_n619), .A3(new_n661), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n659), .A2(new_n312), .A3(new_n598), .A4(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G146), .ZN(G48));
  OAI21_X1  g502(.A(new_n190), .B1(new_n298), .B2(new_n305), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(G469), .ZN(new_n690));
  INV_X1    g504(.A(new_n191), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n690), .A2(new_n691), .A3(new_n306), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(KEYINPUT95), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n551), .A2(new_n585), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT95), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n690), .A2(new_n696), .A3(new_n691), .A4(new_n306), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n693), .A2(new_n695), .A3(new_n621), .A4(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(KEYINPUT41), .B(G113), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n698), .B(new_n699), .ZN(G15));
  NAND4_X1  g514(.A1(new_n693), .A2(new_n640), .A3(new_n695), .A4(new_n697), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G116), .ZN(G18));
  INV_X1    g516(.A(new_n692), .ZN(new_n703));
  AND3_X1   g517(.A1(new_n598), .A2(new_n551), .A3(new_n658), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n703), .A2(new_n704), .A3(new_n488), .ZN(new_n705));
  XNOR2_X1  g519(.A(KEYINPUT96), .B(G119), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n705), .B(new_n706), .ZN(G21));
  NOR2_X1   g521(.A1(new_n671), .A2(new_n408), .ZN(new_n708));
  AND4_X1   g522(.A1(new_n598), .A2(new_n594), .A3(new_n632), .A4(new_n708), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n693), .A2(new_n709), .A3(new_n697), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT97), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n693), .A2(new_n709), .A3(KEYINPUT97), .A4(new_n697), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G122), .ZN(G24));
  INV_X1    g529(.A(new_n306), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n296), .A2(new_n297), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n302), .A2(KEYINPUT76), .A3(new_n304), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n717), .A2(new_n718), .A3(new_n282), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n192), .B1(new_n719), .B2(new_n190), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n716), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n618), .A2(new_n619), .A3(new_n661), .ZN(new_n722));
  NOR3_X1   g536(.A1(new_n722), .A2(new_n653), .A3(new_n592), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n721), .A2(new_n723), .A3(new_n691), .A4(new_n598), .ZN(new_n724));
  XOR2_X1   g538(.A(KEYINPUT98), .B(G125), .Z(new_n725));
  XNOR2_X1  g539(.A(new_n724), .B(new_n725), .ZN(G27));
  INV_X1    g540(.A(KEYINPUT42), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n276), .B1(new_n300), .B2(new_n301), .ZN(new_n728));
  OAI21_X1  g542(.A(KEYINPUT99), .B1(new_n728), .B2(new_n283), .ZN(new_n729));
  OR2_X1    g543(.A1(new_n303), .A2(new_n281), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT99), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n309), .A2(new_n731), .A3(new_n196), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n729), .A2(G469), .A3(new_n730), .A4(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(new_n307), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n306), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n191), .A2(new_n597), .ZN(new_n736));
  AND3_X1   g550(.A1(new_n369), .A2(new_n370), .A3(new_n736), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n735), .A2(new_n737), .A3(new_n551), .A4(new_n585), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n727), .B1(new_n738), .B2(new_n722), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT101), .ZN(new_n740));
  AND2_X1   g554(.A1(new_n735), .A2(new_n737), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n550), .A2(KEYINPUT100), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n536), .A2(new_n538), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT100), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n535), .A2(new_n744), .A3(KEYINPUT32), .A4(new_n490), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n742), .A2(new_n549), .A3(new_n743), .A4(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(new_n585), .ZN(new_n747));
  NOR3_X1   g561(.A1(new_n747), .A2(new_n727), .A3(new_n722), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n740), .B1(new_n741), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n735), .A2(new_n737), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n686), .A2(KEYINPUT42), .A3(new_n585), .A4(new_n746), .ZN(new_n751));
  NOR3_X1   g565(.A1(new_n750), .A2(new_n751), .A3(KEYINPUT101), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n739), .B1(new_n749), .B2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G131), .ZN(G33));
  INV_X1    g568(.A(KEYINPUT102), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n755), .B1(new_n738), .B2(new_n662), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n741), .A2(KEYINPUT102), .A3(new_n695), .A4(new_n663), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G134), .ZN(G36));
  OR2_X1    g573(.A1(new_n619), .A2(KEYINPUT103), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n619), .A2(KEYINPUT103), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n760), .A2(new_n618), .A3(new_n761), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n619), .A2(KEYINPUT43), .ZN(new_n763));
  AOI22_X1  g577(.A1(new_n762), .A2(KEYINPUT43), .B1(new_n618), .B2(new_n763), .ZN(new_n764));
  AND2_X1   g578(.A1(new_n592), .A2(new_n658), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT44), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n371), .A2(new_n597), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n764), .A2(KEYINPUT44), .A3(new_n765), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n768), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT46), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n730), .B1(new_n728), .B2(new_n283), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT45), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n192), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n729), .A2(KEYINPUT45), .A3(new_n730), .A4(new_n732), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(new_n777), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n772), .B1(new_n778), .B2(new_n307), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n307), .A2(new_n772), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n716), .B1(new_n777), .B2(new_n780), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n191), .B1(new_n779), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(new_n666), .ZN(new_n783));
  OR2_X1    g597(.A1(new_n771), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(KEYINPUT104), .B(G137), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n784), .B(new_n785), .ZN(G39));
  INV_X1    g600(.A(new_n769), .ZN(new_n787));
  NOR4_X1   g601(.A1(new_n787), .A2(new_n551), .A3(new_n585), .A4(new_n722), .ZN(new_n788));
  XNOR2_X1  g602(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n789));
  AND2_X1   g603(.A1(new_n782), .A2(new_n789), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n782), .A2(new_n789), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n788), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G140), .ZN(G42));
  INV_X1    g607(.A(KEYINPUT117), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT115), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n372), .B1(new_n670), .B2(new_n674), .ZN(new_n796));
  NOR3_X1   g610(.A1(new_n592), .A2(new_n411), .A3(new_n593), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n796), .A2(new_n764), .A3(new_n703), .A4(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT113), .ZN(new_n799));
  AOI21_X1  g613(.A(KEYINPUT50), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n764), .A2(new_n797), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n801), .A2(KEYINPUT113), .A3(new_n703), .A4(new_n796), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT114), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT50), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n804), .B1(new_n798), .B2(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n803), .A2(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n800), .A2(KEYINPUT114), .A3(new_n802), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n795), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(new_n737), .ZN(new_n811));
  NOR4_X1   g625(.A1(new_n811), .A2(new_n716), .A3(new_n411), .A4(new_n720), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n680), .A2(new_n593), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n618), .A2(new_n619), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n812), .A2(new_n654), .A3(new_n764), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n801), .A2(new_n769), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(KEYINPUT111), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n721), .A2(new_n191), .ZN(new_n822));
  XOR2_X1   g636(.A(new_n822), .B(KEYINPUT112), .Z(new_n823));
  NOR3_X1   g637(.A1(new_n790), .A2(new_n823), .A3(new_n791), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n819), .B1(new_n821), .B2(new_n824), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n810), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n808), .A2(new_n795), .A3(new_n809), .ZN(new_n827));
  AOI21_X1  g641(.A(KEYINPUT51), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n812), .A2(new_n585), .A3(new_n746), .A4(new_n764), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n829), .B(KEYINPUT48), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n814), .A2(new_n619), .A3(new_n618), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n801), .A2(new_n598), .A3(new_n703), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n194), .A2(G952), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n833), .B(KEYINPUT116), .ZN(new_n834));
  AND3_X1   g648(.A1(new_n831), .A2(new_n832), .A3(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(new_n822), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n790), .A2(new_n791), .A3(new_n836), .ZN(new_n837));
  OAI211_X1 g651(.A(new_n819), .B(KEYINPUT51), .C1(new_n821), .C2(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n808), .A2(new_n809), .ZN(new_n839));
  OAI211_X1 g653(.A(new_n830), .B(new_n835), .C1(new_n838), .C2(new_n839), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n794), .B1(new_n828), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n839), .A2(KEYINPUT115), .ZN(new_n842));
  INV_X1    g656(.A(new_n824), .ZN(new_n843));
  XOR2_X1   g657(.A(new_n820), .B(KEYINPUT111), .Z(new_n844));
  AOI21_X1  g658(.A(new_n818), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n842), .A2(new_n845), .A3(new_n827), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT51), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(new_n840), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n848), .A2(new_n849), .A3(KEYINPUT117), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n841), .A2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT53), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n645), .A2(new_n691), .A3(new_n648), .A4(new_n661), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n853), .B1(new_n675), .B2(new_n679), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n854), .A2(new_n598), .A3(new_n708), .A4(new_n735), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n664), .A2(new_n724), .A3(new_n855), .A4(new_n687), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(KEYINPUT109), .ZN(new_n857));
  OAI211_X1 g671(.A(new_n704), .B(new_n312), .C1(new_n663), .C2(new_n686), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT109), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n858), .A2(new_n859), .A3(new_n724), .A4(new_n855), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT52), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n618), .A2(new_n619), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n864), .A2(KEYINPUT106), .ZN(new_n865));
  OR2_X1    g679(.A1(new_n619), .A2(new_n408), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT106), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n618), .A2(new_n867), .A3(new_n619), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n865), .A2(new_n866), .A3(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(new_n632), .ZN(new_n870));
  AOI211_X1 g684(.A(new_n597), .B(new_n870), .C1(new_n369), .C2(new_n370), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n869), .A2(new_n871), .A3(new_n312), .A4(new_n594), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n588), .A2(new_n655), .A3(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT107), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  AND3_X1   g689(.A1(new_n312), .A2(new_n598), .A3(new_n488), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT70), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n694), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n551), .A2(KEYINPUT70), .A3(new_n585), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n876), .B1(new_n880), .B2(new_n654), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n881), .A2(KEYINPUT107), .A3(new_n872), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n875), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n701), .A2(new_n698), .A3(new_n705), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n884), .B1(new_n712), .B2(new_n713), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT108), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n654), .A2(new_n686), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n886), .B1(new_n750), .B2(new_n887), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n723), .A2(new_n735), .A3(new_n737), .A4(KEYINPUT108), .ZN(new_n889));
  AND3_X1   g703(.A1(new_n459), .A2(new_n408), .A3(new_n661), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n551), .A2(new_n629), .A3(new_n658), .A4(new_n890), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n787), .A2(new_n891), .ZN(new_n892));
  AOI22_X1  g706(.A1(new_n888), .A2(new_n889), .B1(new_n892), .B2(new_n312), .ZN(new_n893));
  AND3_X1   g707(.A1(new_n753), .A2(new_n893), .A3(new_n758), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n863), .A2(new_n883), .A3(new_n885), .A4(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n856), .A2(KEYINPUT52), .ZN(new_n896));
  INV_X1    g710(.A(new_n896), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n852), .B1(new_n895), .B2(new_n897), .ZN(new_n898));
  AND3_X1   g712(.A1(new_n701), .A2(new_n698), .A3(new_n705), .ZN(new_n899));
  AOI21_X1  g713(.A(KEYINPUT107), .B1(new_n881), .B2(new_n872), .ZN(new_n900));
  AND4_X1   g714(.A1(KEYINPUT107), .A2(new_n588), .A3(new_n655), .A4(new_n872), .ZN(new_n901));
  OAI211_X1 g715(.A(new_n714), .B(new_n899), .C1(new_n900), .C2(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(KEYINPUT52), .B1(new_n857), .B2(new_n860), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n753), .A2(new_n893), .A3(new_n758), .ZN(new_n904));
  NOR3_X1   g718(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n861), .A2(new_n862), .ZN(new_n906));
  INV_X1    g720(.A(new_n906), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n905), .A2(KEYINPUT53), .A3(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n898), .A2(new_n908), .A3(KEYINPUT110), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT110), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n905), .A2(new_n910), .A3(KEYINPUT53), .A4(new_n907), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n909), .A2(new_n911), .A3(KEYINPUT54), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n852), .B1(new_n895), .B2(new_n906), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n905), .A2(KEYINPUT53), .A3(new_n896), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT54), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n913), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n912), .A2(new_n916), .ZN(new_n917));
  OAI22_X1  g731(.A1(new_n851), .A2(new_n917), .B1(G952), .B2(G953), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n721), .B(KEYINPUT49), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n670), .A2(new_n674), .ZN(new_n920));
  NOR3_X1   g734(.A1(new_n762), .A2(new_n191), .A3(new_n597), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n919), .A2(new_n920), .A3(new_n813), .A4(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n918), .A2(new_n922), .ZN(G75));
  NOR2_X1   g737(.A1(new_n194), .A2(G952), .ZN(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n190), .B1(new_n913), .B2(new_n914), .ZN(new_n926));
  AOI21_X1  g740(.A(KEYINPUT56), .B1(new_n926), .B2(G210), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n342), .A2(new_n351), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(new_n349), .ZN(new_n929));
  XNOR2_X1  g743(.A(KEYINPUT118), .B(KEYINPUT55), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n929), .B(new_n930), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n925), .B1(new_n927), .B2(new_n931), .ZN(new_n932));
  AOI21_X1  g746(.A(KEYINPUT53), .B1(new_n905), .B2(new_n907), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n894), .A2(new_n885), .A3(new_n883), .ZN(new_n934));
  NOR4_X1   g748(.A1(new_n934), .A2(new_n852), .A3(new_n903), .A4(new_n897), .ZN(new_n935));
  OAI21_X1  g749(.A(G902), .B1(new_n933), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(KEYINPUT119), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n913), .A2(new_n914), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT119), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n938), .A2(new_n939), .A3(G902), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n937), .A2(new_n368), .A3(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT56), .ZN(new_n942));
  AND2_X1   g756(.A1(new_n931), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n932), .B1(new_n941), .B2(new_n943), .ZN(G51));
  INV_X1    g758(.A(new_n916), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n915), .B1(new_n913), .B2(new_n914), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n307), .B(KEYINPUT57), .Z(new_n948));
  OAI21_X1  g762(.A(new_n719), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n937), .A2(new_n778), .A3(new_n940), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n924), .B1(new_n949), .B2(new_n950), .ZN(G54));
  AND2_X1   g765(.A1(KEYINPUT58), .A2(G475), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n937), .A2(new_n940), .A3(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(new_n485), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n937), .A2(new_n485), .A3(new_n940), .A4(new_n952), .ZN(new_n956));
  AND3_X1   g770(.A1(new_n955), .A2(new_n925), .A3(new_n956), .ZN(G60));
  NAND2_X1  g771(.A1(G478), .A2(G902), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n958), .B(KEYINPUT59), .Z(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n600), .A2(new_n606), .A3(new_n960), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n925), .B1(new_n947), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n917), .A2(new_n960), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n600), .A2(new_n606), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n962), .B1(new_n963), .B2(new_n964), .ZN(G63));
  NAND2_X1  g779(.A1(G217), .A2(G902), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n966), .B(KEYINPUT120), .Z(new_n967));
  XOR2_X1   g781(.A(new_n967), .B(KEYINPUT60), .Z(new_n968));
  NAND2_X1  g782(.A1(new_n938), .A2(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(new_n577), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n924), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT121), .ZN(new_n972));
  INV_X1    g786(.A(KEYINPUT61), .ZN(new_n973));
  INV_X1    g787(.A(new_n968), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n974), .B1(new_n913), .B2(new_n914), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n975), .A2(new_n647), .ZN(new_n976));
  NAND4_X1  g790(.A1(new_n971), .A2(new_n972), .A3(new_n973), .A4(new_n976), .ZN(new_n977));
  NAND2_X1  g791(.A1(KEYINPUT121), .A2(KEYINPUT61), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n972), .A2(new_n973), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n925), .B1(new_n975), .B2(new_n577), .ZN(new_n980));
  AND3_X1   g794(.A1(new_n938), .A2(new_n647), .A3(new_n968), .ZN(new_n981));
  OAI211_X1 g795(.A(new_n978), .B(new_n979), .C1(new_n980), .C2(new_n981), .ZN(new_n982));
  AND2_X1   g796(.A1(new_n977), .A2(new_n982), .ZN(G66));
  INV_X1    g797(.A(new_n413), .ZN(new_n984));
  OAI21_X1  g798(.A(G953), .B1(new_n984), .B2(new_n346), .ZN(new_n985));
  INV_X1    g799(.A(new_n902), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n985), .B1(new_n986), .B2(G953), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n928), .B1(G898), .B2(new_n194), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n987), .B(new_n988), .ZN(G69));
  AOI21_X1  g803(.A(new_n194), .B1(G227), .B2(G900), .ZN(new_n990));
  INV_X1    g804(.A(KEYINPUT127), .ZN(new_n991));
  AND2_X1   g805(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NOR2_X1   g806(.A1(new_n990), .A2(new_n991), .ZN(new_n993));
  AND4_X1   g807(.A1(new_n598), .A2(new_n585), .A3(new_n708), .A4(new_n746), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n782), .A2(new_n666), .A3(new_n994), .ZN(new_n995));
  OR2_X1    g809(.A1(new_n995), .A2(KEYINPUT125), .ZN(new_n996));
  AND2_X1   g810(.A1(new_n753), .A2(new_n758), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n995), .A2(KEYINPUT125), .ZN(new_n998));
  AND4_X1   g812(.A1(new_n792), .A2(new_n996), .A3(new_n997), .A4(new_n998), .ZN(new_n999));
  AND2_X1   g813(.A1(new_n858), .A2(new_n724), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n1000), .B1(new_n771), .B2(new_n783), .ZN(new_n1001));
  INV_X1    g815(.A(KEYINPUT124), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  OAI211_X1 g817(.A(KEYINPUT124), .B(new_n1000), .C1(new_n771), .C2(new_n783), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g819(.A(G953), .B1(new_n999), .B2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g820(.A1(new_n194), .A2(G900), .ZN(new_n1007));
  OAI21_X1  g821(.A(KEYINPUT126), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g822(.A(KEYINPUT126), .ZN(new_n1009));
  INV_X1    g823(.A(new_n1007), .ZN(new_n1010));
  NAND4_X1  g824(.A1(new_n792), .A2(new_n996), .A3(new_n997), .A4(new_n998), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n1011), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1012));
  OAI211_X1 g826(.A(new_n1009), .B(new_n1010), .C1(new_n1012), .C2(G953), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n463), .A2(new_n464), .ZN(new_n1014));
  XNOR2_X1  g828(.A(new_n1014), .B(KEYINPUT122), .ZN(new_n1015));
  XNOR2_X1  g829(.A(new_n523), .B(new_n1015), .ZN(new_n1016));
  NAND3_X1  g830(.A1(new_n1008), .A2(new_n1013), .A3(new_n1016), .ZN(new_n1017));
  NAND3_X1  g831(.A1(new_n880), .A2(new_n769), .A3(new_n869), .ZN(new_n1018));
  OR2_X1    g832(.A1(new_n1018), .A2(new_n667), .ZN(new_n1019));
  AND2_X1   g833(.A1(new_n784), .A2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g834(.A(KEYINPUT62), .B1(new_n684), .B2(new_n1000), .ZN(new_n1021));
  AND3_X1   g835(.A1(new_n684), .A2(KEYINPUT62), .A3(new_n1000), .ZN(new_n1022));
  OAI211_X1 g836(.A(new_n1020), .B(new_n792), .C1(new_n1021), .C2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n1023), .A2(new_n194), .ZN(new_n1024));
  XOR2_X1   g838(.A(new_n1016), .B(KEYINPUT123), .Z(new_n1025));
  NAND2_X1  g839(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  AOI211_X1 g840(.A(new_n992), .B(new_n993), .C1(new_n1017), .C2(new_n1026), .ZN(new_n1027));
  AND4_X1   g841(.A1(new_n991), .A2(new_n1017), .A3(new_n990), .A4(new_n1026), .ZN(new_n1028));
  NOR2_X1   g842(.A1(new_n1027), .A2(new_n1028), .ZN(G72));
  NAND2_X1  g843(.A1(new_n524), .A2(new_n519), .ZN(new_n1030));
  NAND2_X1  g844(.A1(G472), .A2(G902), .ZN(new_n1031));
  XOR2_X1   g845(.A(new_n1031), .B(KEYINPUT63), .Z(new_n1032));
  INV_X1    g846(.A(new_n1032), .ZN(new_n1033));
  AOI21_X1  g847(.A(new_n1033), .B1(new_n1012), .B2(new_n986), .ZN(new_n1034));
  NOR2_X1   g848(.A1(new_n1023), .A2(new_n902), .ZN(new_n1035));
  NOR2_X1   g849(.A1(new_n1035), .A2(new_n1033), .ZN(new_n1036));
  OAI221_X1 g850(.A(new_n925), .B1(new_n1030), .B2(new_n1034), .C1(new_n1036), .C2(new_n676), .ZN(new_n1037));
  AND2_X1   g851(.A1(new_n909), .A2(new_n911), .ZN(new_n1038));
  AND3_X1   g852(.A1(new_n1030), .A2(new_n676), .A3(new_n1032), .ZN(new_n1039));
  AOI21_X1  g853(.A(new_n1037), .B1(new_n1038), .B2(new_n1039), .ZN(G57));
endmodule


