//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 0 0 0 0 0 0 1 1 1 1 0 0 1 1 0 0 1 1 0 0 0 1 1 0 1 0 0 0 1 1 0 1 0 1 0 1 0 1 1 1 1 0 0 1 0 0 0 1 1 1 0 0 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:35 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1235, new_n1236, new_n1237,
    new_n1238, new_n1239, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n203), .A2(G50), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n207), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(KEYINPUT1), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n222));
  NAND4_X1  g0022(.A1(new_n219), .A2(new_n220), .A3(new_n221), .A4(new_n222), .ZN(new_n223));
  AND2_X1   g0023(.A1(new_n223), .A2(new_n209), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n212), .B(new_n217), .C1(new_n218), .C2(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(new_n218), .ZN(new_n226));
  XOR2_X1   g0026(.A(new_n226), .B(KEYINPUT64), .Z(new_n227));
  NOR2_X1   g0027(.A1(new_n225), .A2(new_n227), .ZN(G361));
  XOR2_X1   g0028(.A(G238), .B(G244), .Z(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G226), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XNOR2_X1  g0037(.A(G50), .B(G68), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G58), .B(G77), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n238), .B(new_n239), .Z(new_n240));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XOR2_X1   g0041(.A(G107), .B(G116), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n240), .B(new_n243), .Z(G351));
  NAND3_X1  g0044(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n245), .A2(new_n215), .ZN(new_n246));
  OAI21_X1  g0046(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n247));
  INV_X1    g0047(.A(G150), .ZN(new_n248));
  NOR2_X1   g0048(.A1(G20), .A2(G33), .ZN(new_n249));
  INV_X1    g0049(.A(new_n249), .ZN(new_n250));
  OAI21_X1  g0050(.A(new_n247), .B1(new_n248), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(KEYINPUT8), .A2(G58), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  NOR2_X1   g0053(.A1(KEYINPUT8), .A2(G58), .ZN(new_n254));
  INV_X1    g0054(.A(G33), .ZN(new_n255));
  NOR4_X1   g0055(.A1(new_n253), .A2(new_n254), .A3(G20), .A4(new_n255), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n246), .B1(new_n251), .B2(new_n256), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n259), .A2(new_n246), .ZN(new_n260));
  INV_X1    g0060(.A(G50), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n261), .B1(new_n206), .B2(G20), .ZN(new_n262));
  AOI22_X1  g0062(.A1(new_n260), .A2(new_n262), .B1(new_n261), .B2(new_n259), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n257), .A2(new_n263), .ZN(new_n264));
  XNOR2_X1  g0064(.A(new_n264), .B(KEYINPUT9), .ZN(new_n265));
  XNOR2_X1  g0065(.A(KEYINPUT3), .B(G33), .ZN(new_n266));
  INV_X1    g0066(.A(G1698), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n266), .A2(G222), .A3(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G77), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n266), .A2(G1698), .ZN(new_n270));
  INV_X1    g0070(.A(G223), .ZN(new_n271));
  OAI221_X1 g0071(.A(new_n268), .B1(new_n269), .B2(new_n266), .C1(new_n270), .C2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(G33), .A2(G41), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n273), .A2(G1), .A3(G13), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n272), .A2(new_n275), .ZN(new_n276));
  OAI211_X1 g0076(.A(new_n206), .B(G274), .C1(G41), .C2(G45), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n279));
  AND2_X1   g0079(.A1(new_n274), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n278), .B1(new_n280), .B2(G226), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n276), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G200), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n265), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G190), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n282), .A2(new_n285), .ZN(new_n286));
  OAI21_X1  g0086(.A(KEYINPUT10), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  XNOR2_X1  g0087(.A(KEYINPUT68), .B(KEYINPUT10), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT67), .ZN(new_n289));
  OAI221_X1 g0089(.A(new_n288), .B1(new_n285), .B2(new_n282), .C1(new_n265), .C2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n265), .A2(new_n289), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n283), .A2(KEYINPUT69), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT69), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n282), .A2(new_n293), .A3(G200), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n291), .A2(new_n292), .A3(new_n294), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n287), .B1(new_n290), .B2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n282), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n264), .B1(new_n297), .B2(G169), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n282), .A2(G179), .ZN(new_n299));
  OR2_X1    g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n296), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT72), .ZN(new_n303));
  INV_X1    g0103(.A(G169), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n255), .A2(KEYINPUT3), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT3), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(G33), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n305), .A2(new_n307), .A3(G226), .A4(new_n267), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT70), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND4_X1  g0110(.A1(new_n266), .A2(KEYINPUT70), .A3(G226), .A4(new_n267), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n305), .A2(new_n307), .A3(G232), .A4(G1698), .ZN(new_n313));
  NAND2_X1  g0113(.A1(G33), .A2(G97), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n274), .B1(new_n312), .B2(new_n316), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n274), .A2(G238), .A3(new_n279), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT71), .ZN(new_n319));
  AND3_X1   g0119(.A1(new_n318), .A2(new_n319), .A3(new_n277), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n319), .B1(new_n318), .B2(new_n277), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  OAI21_X1  g0122(.A(KEYINPUT13), .B1(new_n317), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n318), .A2(new_n277), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(KEYINPUT71), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n318), .A2(new_n319), .A3(new_n277), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT13), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n315), .B1(new_n310), .B2(new_n311), .ZN(new_n329));
  OAI211_X1 g0129(.A(new_n327), .B(new_n328), .C1(new_n274), .C2(new_n329), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n304), .B1(new_n323), .B2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT14), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n323), .A2(new_n330), .ZN(new_n333));
  INV_X1    g0133(.A(G179), .ZN(new_n334));
  OAI22_X1  g0134(.A1(new_n331), .A2(new_n332), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  AOI211_X1 g0135(.A(KEYINPUT14), .B(new_n304), .C1(new_n323), .C2(new_n330), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n303), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  AND2_X1   g0137(.A1(new_n323), .A2(new_n330), .ZN(new_n338));
  OAI21_X1  g0138(.A(KEYINPUT14), .B1(new_n338), .B2(new_n304), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n331), .A2(new_n332), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n338), .A2(G179), .ZN(new_n341));
  NAND4_X1  g0141(.A1(new_n339), .A2(KEYINPUT72), .A3(new_n340), .A4(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n337), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n259), .A2(KEYINPUT66), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT66), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n258), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n348), .A2(KEYINPUT12), .A3(new_n202), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n349), .B1(KEYINPUT12), .B2(new_n259), .ZN(new_n350));
  INV_X1    g0150(.A(new_n246), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n255), .A2(G20), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n352), .A2(G77), .B1(G20), .B2(new_n202), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n249), .A2(G50), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n351), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  XNOR2_X1  g0155(.A(new_n355), .B(KEYINPUT11), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n206), .A2(G20), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n347), .A2(new_n351), .A3(new_n357), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n202), .B1(new_n358), .B2(KEYINPUT12), .ZN(new_n359));
  NOR3_X1   g0159(.A1(new_n350), .A2(new_n356), .A3(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n343), .A2(new_n361), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n361), .B1(G190), .B2(new_n338), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n333), .A2(G200), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  XNOR2_X1  g0165(.A(KEYINPUT15), .B(G87), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  AOI22_X1  g0167(.A1(new_n367), .A2(new_n352), .B1(G20), .B2(G77), .ZN(new_n368));
  OR2_X1    g0168(.A1(new_n253), .A2(new_n254), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n368), .B1(new_n250), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(new_n246), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n348), .A2(new_n269), .ZN(new_n372));
  OAI211_X1 g0172(.A(new_n371), .B(new_n372), .C1(new_n269), .C2(new_n358), .ZN(new_n373));
  AND2_X1   g0173(.A1(new_n280), .A2(G244), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n266), .A2(G232), .A3(new_n267), .ZN(new_n375));
  INV_X1    g0175(.A(G107), .ZN(new_n376));
  INV_X1    g0176(.A(G238), .ZN(new_n377));
  OAI221_X1 g0177(.A(new_n375), .B1(new_n376), .B2(new_n266), .C1(new_n270), .C2(new_n377), .ZN(new_n378));
  AOI211_X1 g0178(.A(new_n278), .B(new_n374), .C1(new_n378), .C2(new_n275), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n373), .B1(new_n379), .B2(G169), .ZN(new_n380));
  AND2_X1   g0180(.A1(new_n379), .A2(new_n334), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n373), .B1(new_n379), .B2(G190), .ZN(new_n384));
  INV_X1    g0184(.A(G200), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n384), .B1(new_n385), .B2(new_n379), .ZN(new_n386));
  AND2_X1   g0186(.A1(new_n383), .A2(new_n386), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n302), .A2(new_n362), .A3(new_n365), .A4(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n203), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n201), .A2(new_n202), .ZN(new_n390));
  OAI21_X1  g0190(.A(G20), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n249), .A2(G159), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n306), .A2(KEYINPUT73), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT73), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(KEYINPUT3), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n395), .A2(new_n397), .A3(G33), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(new_n305), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT7), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n399), .A2(new_n400), .A3(new_n207), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(G68), .ZN(new_n402));
  AOI21_X1  g0202(.A(G20), .B1(new_n398), .B2(new_n305), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n403), .A2(new_n400), .ZN(new_n404));
  OAI211_X1 g0204(.A(KEYINPUT16), .B(new_n394), .C1(new_n402), .C2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT16), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n400), .A2(G20), .ZN(new_n407));
  AOI21_X1  g0207(.A(G33), .B1(new_n395), .B2(new_n397), .ZN(new_n408));
  INV_X1    g0208(.A(new_n307), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n407), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n400), .B1(new_n266), .B2(G20), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n202), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n406), .B1(new_n412), .B2(new_n393), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n405), .A2(new_n413), .A3(new_n246), .ZN(new_n414));
  INV_X1    g0214(.A(new_n369), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(new_n357), .ZN(new_n416));
  INV_X1    g0216(.A(new_n260), .ZN(new_n417));
  OAI22_X1  g0217(.A1(new_n416), .A2(new_n417), .B1(new_n258), .B2(new_n415), .ZN(new_n418));
  INV_X1    g0218(.A(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n414), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(KEYINPUT74), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT74), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n414), .A2(new_n422), .A3(new_n419), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n274), .A2(G232), .A3(new_n279), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(KEYINPUT75), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT75), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n274), .A2(new_n279), .A3(new_n426), .A4(G232), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(new_n277), .ZN(new_n429));
  MUX2_X1   g0229(.A(G223), .B(G226), .S(G1698), .Z(new_n430));
  NAND3_X1  g0230(.A1(new_n430), .A2(new_n398), .A3(new_n305), .ZN(new_n431));
  NAND2_X1  g0231(.A1(G33), .A2(G87), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n274), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(G169), .B1(new_n429), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n431), .A2(new_n432), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(new_n275), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n278), .B1(new_n425), .B2(new_n427), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n436), .A2(G179), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n434), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n421), .A2(new_n423), .A3(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT18), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n421), .A2(KEYINPUT18), .A3(new_n439), .A4(new_n423), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n442), .A2(KEYINPUT76), .A3(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT76), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n440), .A2(new_n445), .A3(new_n441), .ZN(new_n446));
  NOR3_X1   g0246(.A1(new_n429), .A2(new_n285), .A3(new_n433), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n385), .B1(new_n436), .B2(new_n437), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n449), .A2(new_n414), .A3(new_n419), .ZN(new_n450));
  XNOR2_X1  g0250(.A(new_n450), .B(KEYINPUT17), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n444), .A2(new_n446), .A3(new_n451), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n388), .A2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT25), .ZN(new_n454));
  AOI211_X1 g0254(.A(G107), .B(new_n258), .C1(KEYINPUT83), .C2(new_n454), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n454), .A2(KEYINPUT83), .ZN(new_n456));
  XNOR2_X1  g0256(.A(new_n455), .B(new_n456), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n417), .B1(new_n206), .B2(G33), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(G107), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(new_n305), .ZN(new_n461));
  XNOR2_X1  g0261(.A(KEYINPUT73), .B(KEYINPUT3), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n461), .B1(new_n462), .B2(G33), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n463), .A2(KEYINPUT22), .A3(new_n207), .A4(G87), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT22), .ZN(new_n465));
  INV_X1    g0265(.A(new_n266), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n207), .A2(G87), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(G33), .A2(G116), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n469), .A2(G20), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT23), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n471), .B1(new_n207), .B2(G107), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n376), .A2(KEYINPUT23), .A3(G20), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n470), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n464), .A2(new_n468), .A3(new_n474), .ZN(new_n475));
  XNOR2_X1  g0275(.A(new_n475), .B(KEYINPUT24), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n460), .B1(new_n476), .B2(new_n246), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT84), .ZN(new_n478));
  MUX2_X1   g0278(.A(G250), .B(G257), .S(G1698), .Z(new_n479));
  NAND3_X1  g0279(.A1(new_n479), .A2(new_n398), .A3(new_n305), .ZN(new_n480));
  INV_X1    g0280(.A(G294), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n255), .A2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n274), .B1(new_n480), .B2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT5), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT77), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n485), .B1(new_n486), .B2(G41), .ZN(new_n487));
  INV_X1    g0287(.A(G45), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n488), .A2(G1), .ZN(new_n489));
  INV_X1    g0289(.A(G41), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n490), .A2(KEYINPUT77), .A3(KEYINPUT5), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n487), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n492), .A2(G264), .A3(new_n274), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n478), .B1(new_n484), .B2(new_n494), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n482), .B1(new_n463), .B2(new_n479), .ZN(new_n496));
  OAI211_X1 g0296(.A(KEYINPUT84), .B(new_n493), .C1(new_n496), .C2(new_n274), .ZN(new_n497));
  AND2_X1   g0297(.A1(new_n489), .A2(G274), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n498), .A2(new_n274), .A3(new_n487), .A4(new_n491), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n495), .A2(new_n497), .A3(new_n499), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n500), .A2(KEYINPUT85), .A3(new_n385), .ZN(new_n501));
  INV_X1    g0301(.A(new_n499), .ZN(new_n502));
  NOR3_X1   g0302(.A1(new_n484), .A2(new_n494), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(new_n285), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n501), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(KEYINPUT85), .B1(new_n500), .B2(new_n385), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n477), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(KEYINPUT86), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT86), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n509), .B(new_n477), .C1(new_n505), .C2(new_n506), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT24), .ZN(new_n512));
  XNOR2_X1  g0312(.A(new_n475), .B(new_n512), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n459), .B(new_n457), .C1(new_n513), .C2(new_n351), .ZN(new_n514));
  OAI22_X1  g0314(.A1(new_n500), .A2(new_n334), .B1(new_n503), .B2(new_n304), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n511), .A2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT80), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT19), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n352), .A2(new_n520), .A3(G97), .ZN(new_n521));
  NOR2_X1   g0321(.A1(G97), .A2(G107), .ZN(new_n522));
  INV_X1    g0322(.A(G87), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n522), .A2(new_n523), .B1(new_n314), .B2(new_n207), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n521), .B1(new_n524), .B2(new_n520), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n398), .A2(new_n207), .A3(G68), .A4(new_n305), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(KEYINPUT79), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT79), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n525), .A2(new_n526), .A3(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n528), .A2(new_n246), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n348), .A2(new_n366), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n458), .A2(G87), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n398), .A2(G238), .A3(new_n267), .A4(new_n305), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n398), .A2(G244), .A3(G1698), .A4(new_n305), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n535), .A2(new_n536), .A3(new_n469), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(new_n275), .ZN(new_n538));
  INV_X1    g0338(.A(G250), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n489), .A2(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n498), .B1(new_n540), .B2(new_n274), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n385), .B1(new_n538), .B2(new_n541), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n519), .B1(new_n534), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n538), .A2(new_n541), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(G200), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n351), .B1(new_n527), .B2(KEYINPUT79), .ZN(new_n546));
  AOI22_X1  g0346(.A1(new_n546), .A2(new_n530), .B1(new_n348), .B2(new_n366), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n545), .A2(new_n547), .A3(KEYINPUT80), .A4(new_n533), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n538), .A2(G190), .A3(new_n541), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n543), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n458), .A2(new_n367), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n531), .A2(new_n551), .A3(new_n532), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n544), .A2(new_n304), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n538), .A2(new_n334), .A3(new_n541), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n550), .A2(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(G116), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n557), .B1(new_n206), .B2(G33), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n347), .A2(new_n351), .A3(new_n558), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n344), .A2(new_n557), .A3(new_n346), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  AOI22_X1  g0361(.A1(new_n245), .A2(new_n215), .B1(G20), .B2(new_n557), .ZN(new_n562));
  NAND2_X1  g0362(.A1(G33), .A2(G283), .ZN(new_n563));
  INV_X1    g0363(.A(G97), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n563), .B(new_n207), .C1(G33), .C2(new_n564), .ZN(new_n565));
  AND3_X1   g0365(.A1(new_n562), .A2(KEYINPUT20), .A3(new_n565), .ZN(new_n566));
  AOI21_X1  g0366(.A(KEYINPUT20), .B1(new_n562), .B2(new_n565), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  OAI21_X1  g0368(.A(G169), .B1(new_n561), .B2(new_n568), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n492), .A2(G270), .A3(new_n274), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n499), .ZN(new_n571));
  AND2_X1   g0371(.A1(G264), .A2(G1698), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n398), .A2(new_n305), .A3(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT81), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n466), .A2(G303), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n398), .A2(G257), .A3(new_n267), .A4(new_n305), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n398), .A2(KEYINPUT81), .A3(new_n305), .A4(new_n572), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n575), .A2(new_n576), .A3(new_n577), .A4(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n571), .B1(new_n579), .B2(new_n275), .ZN(new_n580));
  OAI21_X1  g0380(.A(KEYINPUT82), .B1(new_n569), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(KEYINPUT21), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n580), .A2(G190), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n561), .A2(new_n568), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n583), .B(new_n584), .C1(new_n385), .C2(new_n580), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT21), .ZN(new_n586));
  OAI211_X1 g0386(.A(KEYINPUT82), .B(new_n586), .C1(new_n569), .C2(new_n580), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n580), .B(G179), .C1(new_n568), .C2(new_n561), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n582), .A2(new_n585), .A3(new_n587), .A4(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n492), .A2(G257), .A3(new_n274), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n499), .A2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(new_n591), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n305), .A2(new_n307), .A3(G250), .A4(G1698), .ZN(new_n593));
  AND2_X1   g0393(.A1(KEYINPUT4), .A2(G244), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n305), .A2(new_n307), .A3(new_n594), .A4(new_n267), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n593), .A2(new_n595), .A3(new_n563), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT4), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n398), .A2(G244), .A3(new_n267), .A4(new_n305), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n596), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n592), .B(new_n334), .C1(new_n599), .C2(new_n274), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(KEYINPUT78), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n598), .A2(new_n597), .ZN(new_n602));
  INV_X1    g0402(.A(new_n596), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(new_n275), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT78), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n605), .A2(new_n606), .A3(new_n334), .A4(new_n592), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n601), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n592), .B1(new_n599), .B2(new_n274), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n258), .A2(G97), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n610), .B1(new_n458), .B2(G97), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n376), .B1(new_n410), .B2(new_n411), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT6), .ZN(new_n613));
  NOR3_X1   g0413(.A1(new_n613), .A2(new_n564), .A3(G107), .ZN(new_n614));
  XNOR2_X1  g0414(.A(G97), .B(G107), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n614), .B1(new_n613), .B2(new_n615), .ZN(new_n616));
  OAI22_X1  g0416(.A1(new_n616), .A2(new_n207), .B1(new_n269), .B2(new_n250), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n246), .B1(new_n612), .B2(new_n617), .ZN(new_n618));
  AOI22_X1  g0418(.A1(new_n304), .A2(new_n609), .B1(new_n611), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n608), .A2(new_n619), .ZN(new_n620));
  AND2_X1   g0420(.A1(new_n611), .A2(new_n618), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n609), .A2(G200), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n621), .B(new_n622), .C1(new_n285), .C2(new_n609), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n620), .A2(new_n623), .ZN(new_n624));
  NOR3_X1   g0424(.A1(new_n556), .A2(new_n589), .A3(new_n624), .ZN(new_n625));
  AND3_X1   g0425(.A1(new_n453), .A2(new_n518), .A3(new_n625), .ZN(G372));
  INV_X1    g0426(.A(KEYINPUT88), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT87), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n365), .A2(new_n382), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n362), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n360), .B1(new_n337), .B2(new_n342), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n383), .B1(new_n363), .B2(new_n364), .ZN(new_n632));
  OAI21_X1  g0432(.A(KEYINPUT87), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n630), .A2(new_n451), .A3(new_n633), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n202), .B1(new_n403), .B2(new_n400), .ZN(new_n635));
  OAI21_X1  g0435(.A(KEYINPUT7), .B1(new_n463), .B2(G20), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n393), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n351), .B1(new_n637), .B2(KEYINPUT16), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n418), .B1(new_n638), .B2(new_n413), .ZN(new_n639));
  INV_X1    g0439(.A(new_n439), .ZN(new_n640));
  OAI21_X1  g0440(.A(KEYINPUT18), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  AOI22_X1  g0441(.A1(new_n414), .A2(new_n419), .B1(new_n438), .B2(new_n434), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(new_n441), .ZN(new_n643));
  AND2_X1   g0443(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n634), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(new_n296), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n627), .B1(new_n646), .B2(new_n300), .ZN(new_n647));
  INV_X1    g0447(.A(new_n296), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n648), .B1(new_n634), .B2(new_n644), .ZN(new_n649));
  INV_X1    g0449(.A(new_n300), .ZN(new_n650));
  NOR3_X1   g0450(.A1(new_n649), .A2(KEYINPUT88), .A3(new_n650), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n647), .A2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  AND2_X1   g0453(.A1(new_n587), .A2(new_n588), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n516), .A2(new_n654), .A3(new_n582), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n545), .A2(new_n547), .A3(new_n533), .A4(new_n549), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(new_n555), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n624), .A2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n510), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n500), .A2(new_n385), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT85), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n662), .A2(new_n501), .A3(new_n504), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n509), .B1(new_n663), .B2(new_n477), .ZN(new_n664));
  OAI211_X1 g0464(.A(new_n655), .B(new_n658), .C1(new_n659), .C2(new_n664), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n656), .A2(new_n555), .A3(new_n608), .A4(new_n619), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n555), .B1(new_n666), .B2(KEYINPUT26), .ZN(new_n667));
  INV_X1    g0467(.A(new_n620), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n668), .A2(new_n550), .A3(new_n555), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n667), .B1(KEYINPUT26), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n665), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n453), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n653), .A2(new_n672), .ZN(G369));
  NAND3_X1  g0473(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n674));
  OR2_X1    g0474(.A1(new_n674), .A2(KEYINPUT27), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(G213), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n676), .B1(KEYINPUT27), .B2(new_n674), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(G343), .ZN(new_n678));
  XNOR2_X1  g0478(.A(new_n678), .B(KEYINPUT89), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n477), .A2(new_n680), .ZN(new_n681));
  OAI22_X1  g0481(.A1(new_n517), .A2(new_n681), .B1(new_n516), .B2(new_n680), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n654), .A2(new_n582), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n680), .A2(new_n584), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n685), .B1(new_n589), .B2(new_n684), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(G330), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n682), .A2(new_n688), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n679), .B1(new_n654), .B2(new_n582), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n511), .A2(new_n690), .A3(new_n516), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n514), .A2(new_n515), .A3(new_n680), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n689), .A2(new_n694), .ZN(G399));
  INV_X1    g0495(.A(new_n210), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n696), .A2(G41), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n522), .A2(new_n523), .A3(new_n557), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n698), .A2(G1), .A3(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n701), .B1(new_n213), .B2(new_n698), .ZN(new_n702));
  XNOR2_X1  g0502(.A(new_n702), .B(KEYINPUT28), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n625), .A2(new_n511), .A3(new_n516), .A4(new_n680), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT31), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n680), .A2(new_n705), .ZN(new_n706));
  AND2_X1   g0506(.A1(new_n538), .A2(new_n541), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n591), .B1(new_n604), .B2(new_n275), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n707), .A2(new_n495), .A3(new_n497), .A4(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT30), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n580), .A2(G179), .ZN(new_n711));
  OR3_X1    g0511(.A1(new_n709), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n710), .B1(new_n709), .B2(new_n711), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n580), .A2(new_n708), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n714), .A2(new_n334), .A3(new_n500), .A4(new_n544), .ZN(new_n715));
  AND2_X1   g0515(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT90), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n712), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  AND3_X1   g0518(.A1(new_n713), .A2(new_n717), .A3(new_n715), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n706), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n716), .A2(new_n712), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(new_n679), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(new_n705), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n704), .A2(new_n720), .A3(new_n723), .ZN(new_n724));
  AND3_X1   g0524(.A1(new_n724), .A2(KEYINPUT91), .A3(G330), .ZN(new_n725));
  AOI21_X1  g0525(.A(KEYINPUT91), .B1(new_n724), .B2(G330), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  OR2_X1    g0527(.A1(new_n655), .A2(KEYINPUT92), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n655), .A2(KEYINPUT92), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n728), .A2(new_n511), .A3(new_n658), .A4(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n669), .A2(KEYINPUT26), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n666), .A2(KEYINPUT26), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(new_n555), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n679), .B1(new_n730), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(KEYINPUT29), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n679), .B1(new_n665), .B2(new_n670), .ZN(new_n737));
  OR2_X1    g0537(.A1(new_n737), .A2(KEYINPUT29), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n727), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n703), .B1(new_n741), .B2(G1), .ZN(G364));
  AND2_X1   g0542(.A1(new_n207), .A2(G13), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n206), .B1(new_n743), .B2(G45), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n697), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n688), .A2(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n747), .B1(G330), .B2(new_n686), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n696), .A2(new_n466), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(G355), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n750), .B1(G116), .B2(new_n210), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n696), .A2(new_n463), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n753), .B1(new_n488), .B2(new_n214), .ZN(new_n754));
  OR2_X1    g0554(.A1(new_n240), .A2(new_n488), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n751), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n215), .B1(G20), .B2(new_n304), .ZN(new_n757));
  OR2_X1    g0557(.A1(new_n757), .A2(KEYINPUT93), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(KEYINPUT93), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(G13), .A2(G33), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(G20), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n760), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n746), .B1(new_n756), .B2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n207), .A2(new_n285), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n334), .A2(G200), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  XOR2_X1   g0569(.A(new_n769), .B(KEYINPUT94), .Z(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(G58), .ZN(new_n772));
  NOR2_X1   g0572(.A1(G179), .A2(G200), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n207), .B1(new_n773), .B2(G190), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(new_n564), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n385), .A2(G179), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n767), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  AOI211_X1 g0578(.A(new_n466), .B(new_n775), .C1(G87), .C2(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n207), .A2(G190), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(new_n773), .ZN(new_n781));
  INV_X1    g0581(.A(G159), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n783), .B(KEYINPUT32), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n334), .A2(new_n385), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n767), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n780), .A2(new_n776), .ZN(new_n787));
  OAI22_X1  g0587(.A1(new_n786), .A2(new_n261), .B1(new_n787), .B2(new_n376), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n785), .A2(new_n780), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n768), .A2(new_n780), .ZN(new_n790));
  OAI22_X1  g0590(.A1(new_n789), .A2(new_n202), .B1(new_n790), .B2(new_n269), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n788), .A2(new_n791), .ZN(new_n792));
  NAND4_X1  g0592(.A1(new_n772), .A2(new_n779), .A3(new_n784), .A4(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n789), .ZN(new_n794));
  XNOR2_X1  g0594(.A(KEYINPUT33), .B(G317), .ZN(new_n795));
  INV_X1    g0595(.A(new_n769), .ZN(new_n796));
  AOI22_X1  g0596(.A1(new_n794), .A2(new_n795), .B1(new_n796), .B2(G322), .ZN(new_n797));
  XNOR2_X1  g0597(.A(new_n797), .B(KEYINPUT95), .ZN(new_n798));
  INV_X1    g0598(.A(new_n781), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n266), .B1(new_n799), .B2(G329), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n800), .B1(new_n481), .B2(new_n774), .ZN(new_n801));
  INV_X1    g0601(.A(G326), .ZN(new_n802));
  INV_X1    g0602(.A(G311), .ZN(new_n803));
  OAI22_X1  g0603(.A1(new_n786), .A2(new_n802), .B1(new_n790), .B2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(G303), .ZN(new_n805));
  INV_X1    g0605(.A(G283), .ZN(new_n806));
  OAI22_X1  g0606(.A1(new_n777), .A2(new_n805), .B1(new_n787), .B2(new_n806), .ZN(new_n807));
  OR3_X1    g0607(.A1(new_n801), .A2(new_n804), .A3(new_n807), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n793), .B1(new_n798), .B2(new_n808), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n766), .B1(new_n809), .B2(new_n760), .ZN(new_n810));
  INV_X1    g0610(.A(new_n763), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n810), .B1(new_n686), .B2(new_n811), .ZN(new_n812));
  AND2_X1   g0612(.A1(new_n748), .A2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(G396));
  INV_X1    g0614(.A(new_n760), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n815), .A2(new_n762), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n746), .B1(new_n816), .B2(G77), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n790), .A2(new_n782), .ZN(new_n818));
  INV_X1    g0618(.A(G137), .ZN(new_n819));
  OAI22_X1  g0619(.A1(new_n786), .A2(new_n819), .B1(new_n789), .B2(new_n248), .ZN(new_n820));
  AOI211_X1 g0620(.A(new_n818), .B(new_n820), .C1(new_n771), .C2(G143), .ZN(new_n821));
  OR2_X1    g0621(.A1(new_n821), .A2(KEYINPUT34), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n821), .A2(KEYINPUT34), .ZN(new_n823));
  INV_X1    g0623(.A(new_n787), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(G68), .ZN(new_n825));
  INV_X1    g0625(.A(G132), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n825), .B1(new_n261), .B2(new_n777), .C1(new_n826), .C2(new_n781), .ZN(new_n827));
  INV_X1    g0627(.A(new_n774), .ZN(new_n828));
  AOI211_X1 g0628(.A(new_n399), .B(new_n827), .C1(G58), .C2(new_n828), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n822), .A2(new_n823), .A3(new_n829), .ZN(new_n830));
  OAI22_X1  g0630(.A1(new_n786), .A2(new_n805), .B1(new_n789), .B2(new_n806), .ZN(new_n831));
  AOI211_X1 g0631(.A(new_n266), .B(new_n831), .C1(G294), .C2(new_n796), .ZN(new_n832));
  INV_X1    g0632(.A(new_n775), .ZN(new_n833));
  AOI22_X1  g0633(.A1(G87), .A2(new_n824), .B1(new_n799), .B2(G311), .ZN(new_n834));
  INV_X1    g0634(.A(new_n790), .ZN(new_n835));
  AOI22_X1  g0635(.A1(G107), .A2(new_n778), .B1(new_n835), .B2(G116), .ZN(new_n836));
  NAND4_X1  g0636(.A1(new_n832), .A2(new_n833), .A3(new_n834), .A4(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n830), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n817), .B1(new_n838), .B2(new_n760), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n679), .A2(new_n373), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n386), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(new_n383), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n382), .A2(new_n680), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n839), .B1(new_n845), .B2(new_n762), .ZN(new_n846));
  AND4_X1   g0646(.A1(KEYINPUT96), .A2(new_n671), .A3(new_n680), .A4(new_n845), .ZN(new_n847));
  AOI21_X1  g0647(.A(KEYINPUT96), .B1(new_n737), .B2(new_n845), .ZN(new_n848));
  OAI22_X1  g0648(.A1(new_n847), .A2(new_n848), .B1(new_n737), .B2(new_n845), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n746), .B1(new_n727), .B2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n727), .A2(new_n849), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n846), .B1(new_n851), .B2(new_n852), .ZN(G384));
  INV_X1    g0653(.A(new_n616), .ZN(new_n854));
  OR2_X1    g0654(.A1(new_n854), .A2(KEYINPUT35), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n854), .A2(KEYINPUT35), .ZN(new_n856));
  NAND4_X1  g0656(.A1(new_n855), .A2(G116), .A3(new_n216), .A4(new_n856), .ZN(new_n857));
  XOR2_X1   g0657(.A(new_n857), .B(KEYINPUT36), .Z(new_n858));
  OR3_X1    g0658(.A1(new_n213), .A2(new_n269), .A3(new_n390), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n261), .A2(G68), .ZN(new_n860));
  AOI211_X1 g0660(.A(new_n206), .B(G13), .C1(new_n859), .C2(new_n860), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n858), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n736), .A2(new_n453), .A3(new_n738), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n652), .A2(new_n864), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n843), .B1(new_n847), .B2(new_n848), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT38), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n405), .A2(new_n246), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n637), .A2(KEYINPUT16), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n419), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(new_n677), .ZN(new_n871));
  AND2_X1   g0671(.A1(new_n446), .A2(new_n451), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n871), .B1(new_n872), .B2(new_n444), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT37), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n450), .A2(new_n874), .ZN(new_n875));
  AND3_X1   g0675(.A1(new_n414), .A2(new_n422), .A3(new_n419), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n422), .B1(new_n414), .B2(new_n419), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n875), .B1(new_n878), .B2(new_n439), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n421), .A2(new_n423), .A3(new_n677), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n870), .A2(new_n439), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n881), .A2(new_n871), .A3(new_n450), .ZN(new_n882));
  AOI22_X1  g0682(.A1(new_n879), .A2(new_n880), .B1(KEYINPUT37), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n867), .B1(new_n873), .B2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(new_n871), .ZN(new_n885));
  AOI21_X1  g0685(.A(KEYINPUT18), .B1(new_n878), .B2(new_n439), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n443), .A2(KEYINPUT76), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n446), .A2(new_n451), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n885), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n883), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n890), .A2(KEYINPUT38), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n884), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n361), .A2(new_n679), .ZN(new_n894));
  AOI22_X1  g0694(.A1(new_n343), .A2(new_n361), .B1(new_n365), .B2(new_n894), .ZN(new_n895));
  AOI211_X1 g0695(.A(new_n360), .B(new_n679), .C1(new_n337), .C2(new_n342), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n866), .A2(new_n893), .A3(new_n897), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n884), .A2(KEYINPUT39), .A3(new_n892), .ZN(new_n899));
  AND3_X1   g0699(.A1(new_n449), .A2(new_n414), .A3(new_n419), .ZN(new_n900));
  OAI21_X1  g0700(.A(KEYINPUT97), .B1(new_n900), .B2(new_n642), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT97), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n450), .B(new_n902), .C1(new_n639), .C2(new_n640), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n901), .A2(new_n880), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(KEYINPUT37), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n879), .A2(new_n880), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n880), .B1(new_n644), .B2(new_n451), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  AOI21_X1  g0709(.A(KEYINPUT38), .B1(new_n907), .B2(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n883), .B1(new_n452), .B2(new_n885), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n910), .B1(KEYINPUT38), .B2(new_n911), .ZN(new_n912));
  OAI211_X1 g0712(.A(new_n899), .B(new_n896), .C1(KEYINPUT39), .C2(new_n912), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n644), .A2(new_n677), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  AND3_X1   g0715(.A1(new_n898), .A2(new_n913), .A3(new_n915), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n865), .B(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(G330), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n721), .A2(KEYINPUT31), .A3(new_n679), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n704), .A2(new_n723), .A3(new_n919), .ZN(new_n920));
  NOR3_X1   g0720(.A1(new_n895), .A2(new_n896), .A3(new_n844), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(KEYINPUT40), .B1(new_n912), .B2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT40), .ZN(new_n924));
  AND3_X1   g0724(.A1(new_n920), .A2(new_n921), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(new_n893), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n923), .A2(new_n926), .ZN(new_n927));
  AND2_X1   g0727(.A1(new_n453), .A2(new_n920), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n918), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n929), .B1(new_n928), .B2(new_n927), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n917), .A2(KEYINPUT98), .A3(new_n930), .ZN(new_n931));
  OAI221_X1 g0731(.A(new_n931), .B1(new_n206), .B2(new_n743), .C1(new_n917), .C2(new_n930), .ZN(new_n932));
  AOI21_X1  g0732(.A(KEYINPUT98), .B1(new_n917), .B2(new_n930), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n862), .B1(new_n932), .B2(new_n933), .ZN(G367));
  OAI21_X1  g0734(.A(new_n764), .B1(new_n210), .B2(new_n366), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n753), .A2(new_n236), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n746), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n770), .A2(new_n805), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n787), .A2(new_n564), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n939), .B1(G294), .B2(new_n794), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n803), .B2(new_n786), .ZN(new_n941));
  INV_X1    g0741(.A(G317), .ZN(new_n942));
  OAI221_X1 g0742(.A(new_n399), .B1(new_n806), .B2(new_n790), .C1(new_n942), .C2(new_n781), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n778), .A2(KEYINPUT46), .A3(G116), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT46), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n945), .B1(new_n777), .B2(new_n557), .ZN(new_n946));
  OAI211_X1 g0746(.A(new_n944), .B(new_n946), .C1(new_n376), .C2(new_n774), .ZN(new_n947));
  NOR4_X1   g0747(.A1(new_n938), .A2(new_n941), .A3(new_n943), .A4(new_n947), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n774), .A2(new_n202), .ZN(new_n949));
  AOI211_X1 g0749(.A(new_n466), .B(new_n949), .C1(G50), .C2(new_n835), .ZN(new_n950));
  INV_X1    g0750(.A(G143), .ZN(new_n951));
  OAI22_X1  g0751(.A1(new_n786), .A2(new_n951), .B1(new_n769), .B2(new_n248), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  AOI22_X1  g0753(.A1(G159), .A2(new_n794), .B1(new_n824), .B2(G77), .ZN(new_n954));
  AND3_X1   g0754(.A1(new_n950), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  OAI22_X1  g0755(.A1(new_n777), .A2(new_n201), .B1(new_n781), .B2(new_n819), .ZN(new_n956));
  XOR2_X1   g0756(.A(new_n956), .B(KEYINPUT104), .Z(new_n957));
  AOI21_X1  g0757(.A(new_n948), .B1(new_n955), .B2(new_n957), .ZN(new_n958));
  OR2_X1    g0758(.A1(new_n958), .A2(KEYINPUT47), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n815), .B1(new_n958), .B2(KEYINPUT47), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n937), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n679), .A2(new_n534), .ZN(new_n962));
  MUX2_X1   g0762(.A(new_n555), .B(new_n657), .S(new_n962), .Z(new_n963));
  XOR2_X1   g0763(.A(new_n963), .B(KEYINPUT99), .Z(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n961), .B1(new_n965), .B2(new_n811), .ZN(new_n966));
  XOR2_X1   g0766(.A(new_n966), .B(KEYINPUT105), .Z(new_n967));
  INV_X1    g0767(.A(KEYINPUT103), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n691), .B1(new_n682), .B2(new_n690), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(new_n688), .ZN(new_n970));
  OAI211_X1 g0770(.A(new_n687), .B(new_n691), .C1(new_n682), .C2(new_n690), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n972), .A2(new_n727), .A3(new_n739), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(KEYINPUT102), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT102), .ZN(new_n975));
  NAND4_X1  g0775(.A1(new_n972), .A2(new_n727), .A3(new_n975), .A4(new_n739), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT44), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n668), .A2(new_n679), .ZN(new_n979));
  OAI211_X1 g0779(.A(new_n620), .B(new_n623), .C1(new_n621), .C2(new_n680), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n978), .B1(new_n694), .B2(new_n981), .ZN(new_n982));
  NAND4_X1  g0782(.A1(new_n693), .A2(KEYINPUT44), .A3(new_n980), .A4(new_n979), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n691), .A2(new_n692), .A3(new_n981), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT45), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n985), .B(new_n986), .ZN(new_n987));
  AND3_X1   g0787(.A1(new_n984), .A2(new_n689), .A3(new_n987), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n689), .B1(new_n984), .B2(new_n987), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n968), .B1(new_n977), .B2(new_n991), .ZN(new_n992));
  NAND4_X1  g0792(.A1(new_n990), .A2(new_n974), .A3(KEYINPUT103), .A4(new_n976), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(new_n741), .ZN(new_n995));
  XOR2_X1   g0795(.A(new_n697), .B(KEYINPUT41), .Z(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n745), .B1(new_n995), .B2(new_n997), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n518), .A2(new_n690), .A3(new_n981), .ZN(new_n999));
  OR2_X1    g0799(.A1(new_n999), .A2(KEYINPUT42), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(KEYINPUT42), .ZN(new_n1001));
  AND3_X1   g0801(.A1(new_n514), .A2(new_n623), .A3(new_n515), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n680), .B1(new_n1002), .B2(new_n668), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n1000), .A2(new_n1001), .A3(new_n1003), .ZN(new_n1004));
  OR2_X1    g0804(.A1(new_n1004), .A2(KEYINPUT100), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n965), .A2(KEYINPUT43), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1004), .A2(KEYINPUT100), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1005), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT101), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT100), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1004), .B(new_n1011), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1012), .A2(KEYINPUT101), .A3(new_n1006), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1010), .A2(new_n1013), .ZN(new_n1014));
  XOR2_X1   g0814(.A(new_n964), .B(KEYINPUT43), .Z(new_n1015));
  AOI21_X1  g0815(.A(new_n1015), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n1016), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n689), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(new_n1014), .A2(new_n1017), .B1(new_n1018), .B2(new_n981), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1018), .A2(new_n981), .ZN(new_n1020));
  AOI211_X1 g0820(.A(new_n1020), .B(new_n1016), .C1(new_n1010), .C2(new_n1013), .ZN(new_n1021));
  OR2_X1    g0821(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n967), .B1(new_n998), .B2(new_n1022), .ZN(G387));
  INV_X1    g0823(.A(new_n972), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n740), .A2(new_n1024), .ZN(new_n1025));
  XOR2_X1   g0825(.A(new_n1025), .B(KEYINPUT110), .Z(new_n1026));
  XNOR2_X1  g0826(.A(new_n697), .B(KEYINPUT109), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1026), .A2(new_n977), .A3(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n415), .A2(new_n261), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT50), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n700), .B(new_n488), .C1(new_n202), .C2(new_n269), .ZN(new_n1031));
  OAI221_X1 g0831(.A(new_n752), .B1(new_n1030), .B2(new_n1031), .C1(new_n233), .C2(new_n488), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n749), .A2(new_n699), .B1(new_n376), .B2(new_n696), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1032), .A2(KEYINPUT106), .A3(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1034), .A2(new_n764), .ZN(new_n1035));
  AOI21_X1  g0835(.A(KEYINPUT106), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n746), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  XOR2_X1   g0837(.A(new_n1037), .B(KEYINPUT107), .Z(new_n1038));
  OAI22_X1  g0838(.A1(new_n369), .A2(new_n789), .B1(new_n786), .B2(new_n782), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1039), .B1(G50), .B2(new_n796), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n939), .B1(G68), .B2(new_n835), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(G77), .A2(new_n778), .B1(new_n799), .B2(G150), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n774), .A2(new_n366), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n1043), .A2(new_n399), .ZN(new_n1044));
  NAND4_X1  g0844(.A1(new_n1040), .A2(new_n1041), .A3(new_n1042), .A4(new_n1044), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(G311), .A2(new_n794), .B1(new_n835), .B2(G303), .ZN(new_n1046));
  INV_X1    g0846(.A(G322), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1046), .B1(new_n1047), .B2(new_n786), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1048), .B1(G317), .B2(new_n771), .ZN(new_n1049));
  OR2_X1    g0849(.A1(new_n1049), .A2(KEYINPUT48), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n777), .A2(new_n481), .B1(new_n774), .B2(new_n806), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT108), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1052), .B1(new_n1049), .B2(KEYINPUT48), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1050), .A2(KEYINPUT49), .A3(new_n1053), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(G116), .A2(new_n824), .B1(new_n799), .B2(G326), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1054), .A2(new_n399), .A3(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(KEYINPUT49), .B1(new_n1050), .B2(new_n1053), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1045), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1058), .A2(new_n760), .ZN(new_n1059));
  OAI211_X1 g0859(.A(new_n1038), .B(new_n1059), .C1(new_n682), .C2(new_n811), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n1028), .B(new_n1060), .C1(new_n744), .C2(new_n1024), .ZN(G393));
  INV_X1    g0861(.A(new_n1027), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1062), .B1(new_n977), .B2(new_n991), .ZN(new_n1063));
  AND2_X1   g0863(.A1(new_n994), .A2(new_n1063), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n981), .A2(new_n811), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1065), .B(KEYINPUT111), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n765), .B1(G97), .B2(new_n696), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n752), .A2(new_n243), .ZN(new_n1068));
  AOI211_X1 g0868(.A(new_n697), .B(new_n745), .C1(new_n1067), .C2(new_n1068), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n463), .B1(new_n523), .B2(new_n787), .C1(new_n951), .C2(new_n781), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n415), .A2(new_n835), .B1(new_n794), .B2(G50), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1071), .B1(new_n202), .B2(new_n777), .ZN(new_n1072));
  AOI211_X1 g0872(.A(new_n1070), .B(new_n1072), .C1(G77), .C2(new_n828), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n786), .A2(new_n248), .B1(new_n769), .B2(new_n782), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n1074), .B(KEYINPUT51), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n786), .A2(new_n942), .B1(new_n769), .B2(new_n803), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT52), .ZN(new_n1077));
  OAI221_X1 g0877(.A(new_n466), .B1(new_n774), .B2(new_n557), .C1(new_n376), .C2(new_n787), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n789), .A2(new_n805), .B1(new_n790), .B2(new_n481), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n777), .A2(new_n806), .B1(new_n781), .B2(new_n1047), .ZN(new_n1080));
  NOR3_X1   g0880(.A1(new_n1078), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n1073), .A2(new_n1075), .B1(new_n1077), .B2(new_n1081), .ZN(new_n1082));
  OAI211_X1 g0882(.A(new_n1066), .B(new_n1069), .C1(new_n815), .C2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1083), .B1(new_n991), .B2(new_n744), .ZN(new_n1084));
  OR2_X1    g0884(.A1(new_n1064), .A2(new_n1084), .ZN(G390));
  INV_X1    g0885(.A(new_n896), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(KEYINPUT37), .A2(new_n904), .B1(new_n879), .B2(new_n880), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n867), .B1(new_n1087), .B2(new_n908), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n892), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n843), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(new_n735), .B2(new_n842), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n897), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n1086), .B(new_n1089), .C1(new_n1091), .C2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n896), .B1(new_n866), .B2(new_n897), .ZN(new_n1094));
  AOI21_X1  g0894(.A(KEYINPUT39), .B1(new_n892), .B2(new_n1088), .ZN(new_n1095));
  AND2_X1   g0895(.A1(new_n884), .A2(new_n892), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1095), .B1(new_n1096), .B2(KEYINPUT39), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1093), .B1(new_n1094), .B2(new_n1097), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n922), .A2(new_n918), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n845), .B(new_n897), .C1(new_n725), .C2(new_n726), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n1101), .B(new_n1093), .C1(new_n1094), .C2(new_n1097), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1100), .A2(new_n745), .A3(new_n1102), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n746), .B1(new_n816), .B2(new_n415), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n266), .B1(new_n787), .B2(new_n261), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(new_n1105), .B(KEYINPUT113), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n777), .A2(new_n248), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1107), .ZN(new_n1108));
  XOR2_X1   g0908(.A(KEYINPUT114), .B(KEYINPUT53), .Z(new_n1109));
  NAND2_X1  g0909(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(G125), .ZN(new_n1111));
  OAI221_X1 g0911(.A(new_n1110), .B1(new_n1111), .B2(new_n781), .C1(new_n826), .C2(new_n769), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(KEYINPUT54), .B(G143), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n835), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(G128), .ZN(new_n1116));
  OAI221_X1 g0916(.A(new_n1115), .B1(new_n1116), .B2(new_n786), .C1(new_n819), .C2(new_n789), .ZN(new_n1117));
  OAI22_X1  g0917(.A1(new_n1108), .A2(new_n1109), .B1(new_n782), .B2(new_n774), .ZN(new_n1118));
  NOR3_X1   g0918(.A1(new_n1112), .A2(new_n1117), .A3(new_n1118), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(G107), .A2(new_n794), .B1(new_n835), .B2(G97), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1120), .B1(new_n806), .B2(new_n786), .ZN(new_n1121));
  XNOR2_X1  g0921(.A(new_n1121), .B(KEYINPUT115), .ZN(new_n1122));
  OAI221_X1 g0922(.A(new_n466), .B1(new_n774), .B2(new_n269), .C1(new_n523), .C2(new_n777), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n825), .B1(new_n557), .B2(new_n769), .ZN(new_n1124));
  AOI211_X1 g0924(.A(new_n1123), .B(new_n1124), .C1(G294), .C2(new_n799), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n1106), .A2(new_n1119), .B1(new_n1122), .B2(new_n1125), .ZN(new_n1126));
  OR2_X1    g0926(.A1(new_n1126), .A2(KEYINPUT116), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n815), .B1(new_n1126), .B2(KEYINPUT116), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1104), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1129), .B1(new_n1097), .B2(new_n762), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT112), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n920), .A2(new_n1132), .A3(G330), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1133), .A2(new_n845), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1132), .B1(new_n920), .B2(G330), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1092), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1136), .A2(new_n1101), .A3(new_n1091), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n845), .B1(new_n725), .B2(new_n726), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1099), .B1(new_n1138), .B2(new_n1092), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n848), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n737), .A2(KEYINPUT96), .A3(new_n845), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1090), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1137), .B1(new_n1139), .B2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n453), .A2(G330), .A3(new_n920), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n863), .B(new_n1144), .C1(new_n647), .C2(new_n651), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1143), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1131), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n1100), .A2(new_n1102), .A3(new_n1146), .A4(new_n1143), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1150), .A2(new_n1027), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n1103), .B(new_n1130), .C1(new_n1149), .C2(new_n1151), .ZN(G378));
  NAND2_X1  g0952(.A1(new_n264), .A2(new_n677), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n301), .B(new_n1153), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(new_n1154), .B(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1158), .B1(new_n927), .B2(G330), .ZN(new_n1159));
  AOI211_X1 g0959(.A(new_n918), .B(new_n1157), .C1(new_n923), .C2(new_n926), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n898), .A2(new_n913), .A3(new_n915), .ZN(new_n1161));
  NOR3_X1   g0961(.A1(new_n1159), .A2(new_n1160), .A3(new_n1161), .ZN(new_n1162));
  AND2_X1   g0962(.A1(new_n920), .A2(new_n921), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1163), .A2(new_n1089), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(new_n1164), .A2(KEYINPUT40), .B1(new_n893), .B2(new_n925), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1157), .B1(new_n1165), .B2(new_n918), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n927), .A2(G330), .A3(new_n1158), .ZN(new_n1167));
  AND2_X1   g0967(.A1(new_n913), .A2(new_n915), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n1166), .A2(new_n1167), .B1(new_n1168), .B2(new_n898), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n745), .B1(new_n1162), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT119), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n746), .B1(new_n816), .B2(G50), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(G97), .A2(new_n794), .B1(new_n799), .B2(G283), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1173), .B1(new_n557), .B2(new_n786), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(G77), .A2(new_n778), .B1(new_n835), .B2(new_n367), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(G107), .A2(new_n796), .B1(new_n824), .B2(G58), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n399), .A2(new_n490), .ZN(new_n1178));
  NOR4_X1   g0978(.A1(new_n1174), .A2(new_n1177), .A3(new_n949), .A4(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  XOR2_X1   g0980(.A(KEYINPUT117), .B(KEYINPUT58), .Z(new_n1181));
  NAND2_X1  g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n1178), .B(new_n261), .C1(G33), .C2(G41), .ZN(new_n1183));
  AND2_X1   g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n786), .A2(new_n1111), .B1(new_n789), .B2(new_n826), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n778), .A2(new_n1114), .B1(new_n835), .B2(G137), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1186), .B1(new_n1116), .B2(new_n769), .ZN(new_n1187));
  AOI211_X1 g0987(.A(new_n1185), .B(new_n1187), .C1(G150), .C2(new_n828), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1189), .A2(KEYINPUT59), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n824), .A2(G159), .ZN(new_n1191));
  AOI211_X1 g0991(.A(G33), .B(G41), .C1(new_n799), .C2(G124), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1190), .A2(new_n1191), .A3(new_n1192), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n1189), .A2(KEYINPUT59), .ZN(new_n1194));
  OAI221_X1 g0994(.A(new_n1184), .B1(new_n1181), .B2(new_n1180), .C1(new_n1193), .C2(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1172), .B1(new_n1195), .B2(new_n760), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1196), .B1(new_n1158), .B2(new_n762), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(new_n1197), .B(KEYINPUT118), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1170), .A2(new_n1171), .A3(new_n1198), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1161), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n916), .A2(new_n1166), .A3(new_n1167), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n744), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1198), .ZN(new_n1203));
  OAI21_X1  g1003(.A(KEYINPUT119), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1199), .A2(new_n1204), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(new_n1150), .A2(new_n1146), .B1(new_n1201), .B2(new_n1200), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1027), .B1(new_n1206), .B2(KEYINPUT57), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1150), .A2(new_n1146), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1209));
  AND3_X1   g1009(.A1(new_n1208), .A2(KEYINPUT57), .A3(new_n1209), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1205), .B1(new_n1207), .B2(new_n1210), .ZN(G375));
  OAI211_X1 g1011(.A(new_n1145), .B(new_n1137), .C1(new_n1139), .C2(new_n1142), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1147), .A2(new_n997), .A3(new_n1212), .ZN(new_n1213));
  OAI22_X1  g1013(.A1(new_n786), .A2(new_n826), .B1(new_n781), .B2(new_n1116), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n789), .A2(new_n1113), .B1(new_n790), .B2(new_n248), .ZN(new_n1215));
  AOI211_X1 g1015(.A(new_n1214), .B(new_n1215), .C1(new_n771), .C2(G137), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n777), .A2(new_n782), .B1(new_n787), .B2(new_n201), .ZN(new_n1217));
  AOI211_X1 g1017(.A(new_n399), .B(new_n1217), .C1(G50), .C2(new_n828), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n786), .A2(new_n481), .B1(new_n777), .B2(new_n564), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n790), .A2(new_n376), .B1(new_n781), .B2(new_n805), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  OAI22_X1  g1021(.A1(new_n557), .A2(new_n789), .B1(new_n769), .B2(new_n806), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n466), .B1(new_n787), .B2(new_n269), .ZN(new_n1223));
  NOR3_X1   g1023(.A1(new_n1222), .A2(new_n1223), .A3(new_n1043), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n1216), .A2(new_n1218), .B1(new_n1221), .B2(new_n1224), .ZN(new_n1225));
  OAI221_X1 g1025(.A(new_n746), .B1(G68), .B2(new_n816), .C1(new_n1225), .C2(new_n815), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1226), .B1(new_n1092), .B2(new_n761), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1227), .B1(new_n1143), .B2(new_n745), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1213), .A2(new_n1228), .ZN(G381));
  INV_X1    g1029(.A(KEYINPUT120), .ZN(new_n1230));
  AOI21_X1  g1030(.A(G378), .B1(G375), .B2(new_n1230), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1231), .B1(new_n1230), .B2(G375), .ZN(new_n1232));
  OR4_X1    g1032(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1233));
  OR4_X1    g1033(.A1(G387), .A2(new_n1232), .A3(new_n1233), .A4(G381), .ZN(G407));
  INV_X1    g1034(.A(G343), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1235), .A2(G213), .ZN(new_n1236));
  OR2_X1    g1036(.A1(new_n1232), .A2(new_n1236), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(G407), .A2(G213), .A3(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT121), .ZN(new_n1239));
  XNOR2_X1  g1039(.A(new_n1238), .B(new_n1239), .ZN(G409));
  INV_X1    g1040(.A(KEYINPUT125), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1064), .A2(new_n1084), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1241), .B1(G387), .B2(new_n1242), .ZN(new_n1243));
  XNOR2_X1  g1043(.A(G393), .B(G396), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1244), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n996), .B1(new_n994), .B2(new_n741), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1246), .B1(new_n1247), .B2(new_n745), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(G390), .A2(new_n1248), .A3(new_n967), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(G390), .B1(new_n1248), .B2(new_n967), .ZN(new_n1251));
  OAI22_X1  g1051(.A1(new_n1243), .A2(new_n1245), .B1(new_n1250), .B2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(G387), .A2(new_n1242), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1253), .A2(new_n1241), .A3(new_n1249), .A4(new_n1244), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1252), .A2(new_n1254), .ZN(new_n1255));
  OAI211_X1 g1055(.A(new_n1205), .B(G378), .C1(new_n1207), .C2(new_n1210), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1257));
  OAI211_X1 g1057(.A(new_n1170), .B(new_n1198), .C1(new_n1257), .C2(new_n996), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1103), .A2(new_n1130), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1151), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1259), .B1(new_n1260), .B2(new_n1148), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1258), .A2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1256), .A2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1212), .A2(KEYINPUT122), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1264), .A2(KEYINPUT60), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT60), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1212), .A2(KEYINPUT122), .A3(new_n1266), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1265), .A2(new_n1027), .A3(new_n1147), .A4(new_n1267), .ZN(new_n1268));
  AND3_X1   g1068(.A1(new_n1268), .A2(G384), .A3(new_n1228), .ZN(new_n1269));
  AOI21_X1  g1069(.A(G384), .B1(new_n1268), .B2(new_n1228), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1263), .A2(new_n1236), .A3(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(KEYINPUT62), .ZN(new_n1273));
  AOI22_X1  g1073(.A1(new_n1256), .A2(new_n1262), .B1(G213), .B2(new_n1235), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT62), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1274), .A2(new_n1275), .A3(new_n1271), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1273), .A2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT126), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT61), .ZN(new_n1279));
  OAI21_X1  g1079(.A(KEYINPUT124), .B1(new_n1269), .B2(new_n1270), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1235), .A2(G213), .A3(G2897), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1281), .ZN(new_n1283));
  OAI211_X1 g1083(.A(KEYINPUT124), .B(new_n1283), .C1(new_n1269), .C2(new_n1270), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1270), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT124), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1268), .A2(G384), .A3(new_n1228), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1285), .A2(new_n1286), .A3(new_n1287), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1282), .A2(new_n1284), .A3(new_n1288), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1279), .B1(new_n1289), .B2(new_n1274), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1277), .B1(new_n1278), .B2(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1274), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1292), .A2(new_n1282), .A3(new_n1284), .A4(new_n1288), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1293), .A2(KEYINPUT126), .A3(new_n1279), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1255), .B1(new_n1291), .B2(new_n1294), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1274), .A2(KEYINPUT63), .A3(new_n1271), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1255), .A2(new_n1279), .A3(new_n1293), .A4(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT63), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1272), .A2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT123), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1272), .A2(KEYINPUT123), .A3(new_n1298), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  NOR2_X1   g1103(.A1(new_n1297), .A2(new_n1303), .ZN(new_n1304));
  OAI21_X1  g1104(.A(KEYINPUT127), .B1(new_n1295), .B2(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1290), .A2(new_n1278), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1277), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1306), .A2(new_n1294), .A3(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1255), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  OR2_X1    g1110(.A1(new_n1297), .A2(new_n1303), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT127), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1310), .A2(new_n1311), .A3(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1305), .A2(new_n1313), .ZN(G405));
  NAND2_X1  g1114(.A1(G375), .A2(new_n1261), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1315), .A2(new_n1256), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1309), .A2(new_n1316), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1255), .A2(new_n1256), .A3(new_n1315), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1319));
  XNOR2_X1  g1119(.A(new_n1319), .B(new_n1271), .ZN(G402));
endmodule


