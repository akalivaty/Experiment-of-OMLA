//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 1 1 0 0 1 0 0 0 1 0 0 0 0 1 0 0 0 1 0 1 1 1 0 0 0 1 1 1 0 0 0 0 1 0 0 1 0 1 1 0 1 0 0 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:25 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n452, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n582, new_n583, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n592, new_n596, new_n597,
    new_n598, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n628, new_n631, new_n633,
    new_n634, new_n635, new_n636, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n887, new_n888, new_n889, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1249, new_n1250, new_n1251;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT65), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT66), .B(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g021(.A(KEYINPUT67), .B(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT68), .ZN(G217));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT2), .ZN(new_n455));
  NOR4_X1   g030(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n455), .A2(new_n456), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n456), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n455), .ZN(new_n461));
  AOI21_X1  g036(.A(new_n460), .B1(new_n461), .B2(G2106), .ZN(G319));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  AND3_X1   g038(.A1(new_n463), .A2(KEYINPUT69), .A3(KEYINPUT3), .ZN(new_n464));
  AOI21_X1  g039(.A(KEYINPUT69), .B1(new_n463), .B2(KEYINPUT3), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  OAI21_X1  g042(.A(KEYINPUT70), .B1(new_n463), .B2(KEYINPUT3), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT70), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT3), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n469), .A2(new_n470), .A3(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  NAND4_X1  g047(.A1(new_n466), .A2(G137), .A3(new_n467), .A4(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n463), .A2(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G101), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(G113), .A2(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n470), .A2(G2104), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(G125), .ZN(new_n481));
  OAI21_X1  g056(.A(new_n477), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n476), .A2(new_n484), .ZN(G160));
  INV_X1    g060(.A(new_n465), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n463), .A2(KEYINPUT69), .A3(KEYINPUT3), .ZN(new_n487));
  AND3_X1   g062(.A1(new_n472), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n488), .A2(KEYINPUT72), .A3(G2105), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT72), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n472), .A2(new_n486), .A3(new_n487), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n490), .B1(new_n491), .B2(new_n467), .ZN(new_n492));
  AND2_X1   g067(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(G124), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n488), .A2(KEYINPUT71), .A3(new_n467), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT71), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n496), .B1(new_n491), .B2(G2105), .ZN(new_n497));
  AND2_X1   g072(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(G136), .ZN(new_n499));
  OR2_X1    g074(.A1(G100), .A2(G2105), .ZN(new_n500));
  OAI211_X1 g075(.A(new_n500), .B(G2104), .C1(G112), .C2(new_n467), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n494), .A2(new_n499), .A3(new_n501), .ZN(new_n502));
  OR2_X1    g077(.A1(new_n502), .A2(KEYINPUT73), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(KEYINPUT73), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(G162));
  NAND4_X1  g081(.A1(new_n466), .A2(G126), .A3(G2105), .A4(new_n472), .ZN(new_n507));
  OR2_X1    g082(.A1(G102), .A2(G2105), .ZN(new_n508));
  XOR2_X1   g083(.A(KEYINPUT74), .B(G114), .Z(new_n509));
  OAI211_X1 g084(.A(G2104), .B(new_n508), .C1(new_n509), .C2(new_n467), .ZN(new_n510));
  AND2_X1   g085(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  AND2_X1   g086(.A1(new_n467), .A2(G138), .ZN(new_n512));
  NAND4_X1  g087(.A1(new_n472), .A2(new_n486), .A3(new_n487), .A4(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(KEYINPUT4), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT4), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n515), .A2(new_n467), .A3(G138), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n480), .A2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n514), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g094(.A(KEYINPUT75), .B1(new_n511), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n507), .A2(new_n510), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n517), .B1(new_n513), .B2(KEYINPUT4), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT75), .ZN(new_n523));
  NOR3_X1   g098(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n520), .A2(new_n524), .ZN(G164));
  INV_X1    g100(.A(G651), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT76), .ZN(new_n527));
  INV_X1    g102(.A(G543), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n527), .B1(new_n528), .B2(KEYINPUT5), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT5), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n530), .A2(KEYINPUT76), .A3(G543), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n529), .A2(new_n531), .B1(KEYINPUT5), .B2(new_n528), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G62), .ZN(new_n533));
  NAND2_X1  g108(.A1(G75), .A2(G543), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n526), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(new_n535), .ZN(new_n536));
  XNOR2_X1  g111(.A(KEYINPUT6), .B(G651), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n532), .A2(G88), .A3(new_n537), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n537), .A2(G50), .A3(G543), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(new_n540), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n536), .A2(new_n541), .A3(KEYINPUT77), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT77), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n543), .B1(new_n535), .B2(new_n540), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n542), .A2(new_n544), .ZN(G166));
  AND2_X1   g120(.A1(G63), .A2(G651), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n532), .A2(new_n546), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT78), .ZN(new_n548));
  AND2_X1   g123(.A1(new_n537), .A2(G543), .ZN(new_n549));
  XOR2_X1   g124(.A(KEYINPUT79), .B(G51), .Z(new_n550));
  NAND3_X1  g125(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(KEYINPUT7), .ZN(new_n552));
  OR2_X1    g127(.A1(new_n551), .A2(KEYINPUT7), .ZN(new_n553));
  AOI22_X1  g128(.A1(new_n549), .A2(new_n550), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n532), .A2(G89), .A3(new_n537), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  OAI21_X1  g131(.A(KEYINPUT80), .B1(new_n548), .B2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT78), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n547), .B(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT80), .ZN(new_n560));
  NAND4_X1  g135(.A1(new_n559), .A2(new_n560), .A3(new_n555), .A4(new_n554), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n557), .A2(new_n561), .ZN(G168));
  AOI22_X1  g137(.A1(new_n532), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n563));
  OR2_X1    g138(.A1(new_n563), .A2(new_n526), .ZN(new_n564));
  XOR2_X1   g139(.A(KEYINPUT81), .B(G52), .Z(new_n565));
  NAND2_X1  g140(.A1(new_n549), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n532), .A2(G90), .A3(new_n537), .ZN(new_n567));
  AND3_X1   g142(.A1(new_n566), .A2(KEYINPUT82), .A3(new_n567), .ZN(new_n568));
  AOI21_X1  g143(.A(KEYINPUT82), .B1(new_n566), .B2(new_n567), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n564), .B1(new_n568), .B2(new_n569), .ZN(G301));
  INV_X1    g145(.A(G301), .ZN(G171));
  AOI22_X1  g146(.A1(new_n532), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n572), .A2(new_n526), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n532), .A2(new_n537), .ZN(new_n574));
  INV_X1    g149(.A(G81), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n537), .A2(G543), .ZN(new_n576));
  XNOR2_X1  g151(.A(KEYINPUT83), .B(G43), .ZN(new_n577));
  OAI22_X1  g152(.A1(new_n574), .A2(new_n575), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NOR2_X1   g153(.A1(new_n573), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n579), .A2(G860), .ZN(G153));
  NAND4_X1  g155(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g156(.A1(G1), .A2(G3), .ZN(new_n582));
  XNOR2_X1  g157(.A(new_n582), .B(KEYINPUT8), .ZN(new_n583));
  NAND4_X1  g158(.A1(G319), .A2(G483), .A3(G661), .A4(new_n583), .ZN(G188));
  INV_X1    g159(.A(G53), .ZN(new_n585));
  OR3_X1    g160(.A1(new_n576), .A2(KEYINPUT9), .A3(new_n585), .ZN(new_n586));
  OAI21_X1  g161(.A(KEYINPUT9), .B1(new_n576), .B2(new_n585), .ZN(new_n587));
  INV_X1    g162(.A(new_n574), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n586), .A2(new_n587), .B1(new_n588), .B2(G91), .ZN(new_n589));
  XOR2_X1   g164(.A(KEYINPUT84), .B(G65), .Z(new_n590));
  AOI22_X1  g165(.A1(new_n532), .A2(new_n590), .B1(G78), .B2(G543), .ZN(new_n591));
  OR2_X1    g166(.A1(new_n591), .A2(new_n526), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n589), .A2(new_n592), .ZN(G299));
  INV_X1    g168(.A(G168), .ZN(G286));
  INV_X1    g169(.A(G166), .ZN(G303));
  OAI21_X1  g170(.A(G651), .B1(new_n532), .B2(G74), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n549), .A2(G49), .ZN(new_n597));
  INV_X1    g172(.A(G87), .ZN(new_n598));
  OAI211_X1 g173(.A(new_n596), .B(new_n597), .C1(new_n598), .C2(new_n574), .ZN(G288));
  AOI22_X1  g174(.A1(new_n532), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n600), .A2(new_n526), .ZN(new_n601));
  INV_X1    g176(.A(G86), .ZN(new_n602));
  INV_X1    g177(.A(G48), .ZN(new_n603));
  OAI22_X1  g178(.A1(new_n574), .A2(new_n602), .B1(new_n603), .B2(new_n576), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(new_n605), .ZN(G305));
  AOI22_X1  g181(.A1(new_n532), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n607), .A2(new_n526), .ZN(new_n608));
  INV_X1    g183(.A(G85), .ZN(new_n609));
  INV_X1    g184(.A(G47), .ZN(new_n610));
  OAI22_X1  g185(.A1(new_n574), .A2(new_n609), .B1(new_n610), .B2(new_n576), .ZN(new_n611));
  OR2_X1    g186(.A1(new_n608), .A2(new_n611), .ZN(G290));
  NAND2_X1  g187(.A1(G301), .A2(G868), .ZN(new_n613));
  AND3_X1   g188(.A1(new_n532), .A2(G92), .A3(new_n537), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT10), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n532), .A2(G66), .ZN(new_n616));
  INV_X1    g191(.A(G79), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n617), .B2(new_n528), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n549), .A2(KEYINPUT85), .ZN(new_n619));
  INV_X1    g194(.A(G54), .ZN(new_n620));
  INV_X1    g195(.A(KEYINPUT85), .ZN(new_n621));
  AOI21_X1  g196(.A(new_n620), .B1(new_n576), .B2(new_n621), .ZN(new_n622));
  AOI22_X1  g197(.A1(new_n618), .A2(G651), .B1(new_n619), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n615), .A2(new_n623), .ZN(new_n624));
  INV_X1    g199(.A(new_n624), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n613), .B1(new_n625), .B2(G868), .ZN(G284));
  OAI21_X1  g201(.A(new_n613), .B1(new_n625), .B2(G868), .ZN(G321));
  NOR2_X1   g202(.A1(G299), .A2(G868), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n628), .B1(G168), .B2(G868), .ZN(G297));
  AOI21_X1  g204(.A(new_n628), .B1(G168), .B2(G868), .ZN(G280));
  INV_X1    g205(.A(G559), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n625), .B1(new_n631), .B2(G860), .ZN(G148));
  INV_X1    g207(.A(new_n579), .ZN(new_n633));
  INV_X1    g208(.A(G868), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NOR2_X1   g210(.A1(new_n624), .A2(G559), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n635), .B1(new_n636), .B2(new_n634), .ZN(G323));
  XNOR2_X1  g212(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g213(.A1(new_n493), .A2(G123), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n498), .A2(G135), .ZN(new_n640));
  OR2_X1    g215(.A1(G99), .A2(G2105), .ZN(new_n641));
  OAI211_X1 g216(.A(new_n641), .B(G2104), .C1(G111), .C2(new_n467), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n639), .A2(new_n640), .A3(new_n642), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n643), .A2(G2096), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n643), .A2(G2096), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n467), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(KEYINPUT12), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT13), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(G2100), .Z(new_n649));
  NAND3_X1  g224(.A1(new_n644), .A2(new_n645), .A3(new_n649), .ZN(G156));
  INV_X1    g225(.A(G14), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2427), .B(G2438), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(G2430), .ZN(new_n653));
  XNOR2_X1  g228(.A(KEYINPUT15), .B(G2435), .ZN(new_n654));
  OR2_X1    g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n653), .A2(new_n654), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n655), .A2(KEYINPUT14), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2451), .B(G2454), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT16), .ZN(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2443), .B(G2446), .ZN(new_n662));
  NAND4_X1  g237(.A1(new_n655), .A2(KEYINPUT14), .A3(new_n659), .A4(new_n656), .ZN(new_n663));
  AND3_X1   g238(.A1(new_n661), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n662), .B1(new_n661), .B2(new_n663), .ZN(new_n665));
  OR2_X1    g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1341), .B(G1348), .ZN(new_n667));
  AOI21_X1  g242(.A(new_n651), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NOR4_X1   g243(.A1(new_n664), .A2(new_n665), .A3(KEYINPUT86), .A4(new_n667), .ZN(new_n669));
  INV_X1    g244(.A(KEYINPUT86), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n664), .A2(new_n665), .ZN(new_n671));
  INV_X1    g246(.A(new_n667), .ZN(new_n672));
  AOI21_X1  g247(.A(new_n670), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  OAI21_X1  g248(.A(new_n668), .B1(new_n669), .B2(new_n673), .ZN(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(G401));
  XNOR2_X1  g250(.A(G2084), .B(G2090), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT87), .ZN(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G2067), .B(G2678), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(G2072), .B(G2078), .Z(new_n681));
  NAND2_X1  g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n678), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n681), .B(KEYINPUT17), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n684), .A2(new_n680), .ZN(new_n685));
  OR3_X1    g260(.A1(new_n683), .A2(new_n685), .A3(KEYINPUT88), .ZN(new_n686));
  OAI21_X1  g261(.A(KEYINPUT88), .B1(new_n683), .B2(new_n685), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n684), .A2(new_n677), .A3(new_n680), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT89), .ZN(new_n690));
  NOR3_X1   g265(.A1(new_n678), .A2(new_n680), .A3(new_n681), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT18), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n688), .A2(new_n690), .A3(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(G2096), .B(G2100), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  NAND4_X1  g271(.A1(new_n688), .A2(new_n692), .A3(new_n690), .A4(new_n694), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n696), .A2(new_n697), .ZN(G227));
  XNOR2_X1  g273(.A(G1981), .B(G1986), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1971), .B(G1976), .ZN(new_n701));
  INV_X1    g276(.A(KEYINPUT19), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  XOR2_X1   g278(.A(G1956), .B(G2474), .Z(new_n704));
  XOR2_X1   g279(.A(G1961), .B(G1966), .Z(new_n705));
  AND2_X1   g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n703), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT20), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n704), .A2(new_n705), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n703), .A2(new_n709), .ZN(new_n710));
  OR3_X1    g285(.A1(new_n703), .A2(new_n706), .A3(new_n709), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n708), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(KEYINPUT20), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n707), .B(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n711), .A2(new_n710), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(new_n713), .ZN(new_n720));
  XOR2_X1   g295(.A(G1991), .B(G1996), .Z(new_n721));
  INV_X1    g296(.A(new_n721), .ZN(new_n722));
  AND3_X1   g297(.A1(new_n715), .A2(new_n720), .A3(new_n722), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n722), .B1(new_n715), .B2(new_n720), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n700), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n712), .A2(new_n714), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n719), .A2(new_n713), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n721), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n715), .A2(new_n720), .A3(new_n722), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n728), .A2(new_n699), .A3(new_n729), .ZN(new_n730));
  AND2_X1   g305(.A1(new_n725), .A2(new_n730), .ZN(G229));
  OR2_X1    g306(.A1(G29), .A2(G35), .ZN(new_n732));
  INV_X1    g307(.A(G29), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n732), .B1(new_n505), .B2(new_n733), .ZN(new_n734));
  XNOR2_X1  g309(.A(KEYINPUT29), .B(G2090), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(new_n735), .ZN(new_n737));
  OAI211_X1 g312(.A(new_n732), .B(new_n737), .C1(new_n505), .C2(new_n733), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  AND2_X1   g314(.A1(new_n733), .A2(G33), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n498), .A2(G139), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n467), .A2(G103), .A3(G2104), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT93), .ZN(new_n743));
  OR2_X1    g318(.A1(new_n743), .A2(KEYINPUT25), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n743), .A2(KEYINPUT25), .ZN(new_n745));
  NAND2_X1  g320(.A1(G115), .A2(G2104), .ZN(new_n746));
  INV_X1    g321(.A(G127), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n746), .B1(new_n480), .B2(new_n747), .ZN(new_n748));
  AOI22_X1  g323(.A1(new_n744), .A2(new_n745), .B1(G2105), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n741), .A2(new_n749), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n740), .B1(new_n750), .B2(G29), .ZN(new_n751));
  INV_X1    g326(.A(KEYINPUT94), .ZN(new_n752));
  OR2_X1    g327(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n751), .A2(new_n752), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n442), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n733), .A2(G27), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(G164), .B2(new_n733), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n757), .A2(new_n443), .ZN(new_n758));
  OR2_X1    g333(.A1(new_n757), .A2(new_n443), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n755), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(G16), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n761), .A2(G5), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G171), .B2(new_n761), .ZN(new_n763));
  INV_X1    g338(.A(G1961), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  AND3_X1   g340(.A1(new_n739), .A2(new_n760), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(G286), .A2(G16), .ZN(new_n767));
  INV_X1    g342(.A(G21), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n767), .B1(G16), .B2(new_n768), .ZN(new_n769));
  XNOR2_X1  g344(.A(KEYINPUT98), .B(G1966), .ZN(new_n770));
  INV_X1    g345(.A(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n643), .A2(new_n733), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT99), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n761), .A2(G4), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(new_n625), .B2(new_n761), .ZN(new_n776));
  INV_X1    g351(.A(G1348), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  OAI211_X1 g353(.A(new_n767), .B(new_n770), .C1(G16), .C2(new_n768), .ZN(new_n779));
  AND4_X1   g354(.A1(new_n772), .A2(new_n774), .A3(new_n778), .A4(new_n779), .ZN(new_n780));
  NAND3_X1  g355(.A1(new_n753), .A2(new_n442), .A3(new_n754), .ZN(new_n781));
  AND2_X1   g356(.A1(KEYINPUT24), .A2(G34), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n733), .B1(KEYINPUT24), .B2(G34), .ZN(new_n783));
  OAI22_X1  g358(.A1(G160), .A2(new_n733), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n784), .A2(G2084), .ZN(new_n785));
  AND2_X1   g360(.A1(new_n784), .A2(G2084), .ZN(new_n786));
  INV_X1    g361(.A(G1341), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n579), .A2(G16), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G16), .B2(G19), .ZN(new_n789));
  AOI211_X1 g364(.A(new_n785), .B(new_n786), .C1(new_n787), .C2(new_n789), .ZN(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT100), .B(KEYINPUT23), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n761), .A2(G20), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(G299), .B2(G16), .ZN(new_n794));
  INV_X1    g369(.A(G1956), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  INV_X1    g371(.A(G28), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n797), .A2(KEYINPUT30), .ZN(new_n798));
  AOI21_X1  g373(.A(G29), .B1(new_n797), .B2(KEYINPUT30), .ZN(new_n799));
  OR2_X1    g374(.A1(KEYINPUT31), .A2(G11), .ZN(new_n800));
  NAND2_X1  g375(.A1(KEYINPUT31), .A2(G11), .ZN(new_n801));
  AOI22_X1  g376(.A1(new_n798), .A2(new_n799), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(new_n789), .B2(new_n787), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n796), .A2(new_n803), .ZN(new_n804));
  AND3_X1   g379(.A1(new_n781), .A2(new_n790), .A3(new_n804), .ZN(new_n805));
  NAND3_X1  g380(.A1(new_n489), .A2(G129), .A3(new_n492), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n495), .A2(G141), .A3(new_n497), .ZN(new_n807));
  XNOR2_X1  g382(.A(KEYINPUT96), .B(KEYINPUT26), .ZN(new_n808));
  NAND3_X1  g383(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n474), .A2(G105), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n811), .A2(KEYINPUT95), .ZN(new_n812));
  OR2_X1    g387(.A1(new_n811), .A2(KEYINPUT95), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n810), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n806), .A2(new_n807), .A3(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(KEYINPUT97), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND4_X1  g392(.A1(new_n806), .A2(new_n807), .A3(KEYINPUT97), .A4(new_n814), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  MUX2_X1   g394(.A(G32), .B(new_n819), .S(G29), .Z(new_n820));
  XNOR2_X1  g395(.A(KEYINPUT27), .B(G1996), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  AND3_X1   g397(.A1(new_n780), .A2(new_n805), .A3(new_n822), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n489), .A2(G128), .A3(new_n492), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n495), .A2(G140), .A3(new_n497), .ZN(new_n825));
  OR2_X1    g400(.A1(G104), .A2(G2105), .ZN(new_n826));
  OAI211_X1 g401(.A(new_n826), .B(G2104), .C1(G116), .C2(new_n467), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n824), .A2(new_n825), .A3(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT92), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND4_X1  g405(.A1(new_n824), .A2(new_n825), .A3(KEYINPUT92), .A4(new_n827), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(G26), .ZN(new_n833));
  OAI21_X1  g408(.A(KEYINPUT28), .B1(new_n833), .B2(G29), .ZN(new_n834));
  OR3_X1    g409(.A1(new_n833), .A2(KEYINPUT28), .A3(G29), .ZN(new_n835));
  AOI22_X1  g410(.A1(new_n832), .A2(G29), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(G2067), .ZN(new_n837));
  NAND4_X1  g412(.A1(new_n766), .A2(new_n823), .A3(KEYINPUT101), .A4(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT101), .ZN(new_n839));
  NAND4_X1  g414(.A1(new_n739), .A2(new_n760), .A3(new_n837), .A4(new_n765), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n780), .A2(new_n805), .A3(new_n822), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n839), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n838), .A2(new_n842), .ZN(new_n843));
  NOR2_X1   g418(.A1(G6), .A2(G16), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n844), .B1(new_n605), .B2(G16), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT32), .ZN(new_n846));
  OR2_X1    g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n845), .A2(new_n846), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(G1981), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT34), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n761), .A2(G22), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n852), .B1(G166), .B2(new_n761), .ZN(new_n853));
  OR2_X1    g428(.A1(new_n853), .A2(G1971), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(G1971), .ZN(new_n855));
  MUX2_X1   g430(.A(G23), .B(G288), .S(G16), .Z(new_n856));
  XNOR2_X1  g431(.A(KEYINPUT33), .B(G1976), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n856), .B(new_n857), .ZN(new_n858));
  AND3_X1   g433(.A1(new_n854), .A2(new_n855), .A3(new_n858), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n850), .A2(new_n851), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n733), .A2(G25), .ZN(new_n861));
  XOR2_X1   g436(.A(new_n861), .B(KEYINPUT90), .Z(new_n862));
  NAND3_X1  g437(.A1(new_n489), .A2(G119), .A3(new_n492), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n495), .A2(G131), .A3(new_n497), .ZN(new_n864));
  OR2_X1    g439(.A1(G95), .A2(G2105), .ZN(new_n865));
  OAI211_X1 g440(.A(new_n865), .B(G2104), .C1(G107), .C2(new_n467), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n863), .A2(new_n864), .A3(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT91), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND4_X1  g444(.A1(new_n863), .A2(new_n864), .A3(KEYINPUT91), .A4(new_n866), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n862), .B1(new_n871), .B2(G29), .ZN(new_n872));
  XOR2_X1   g447(.A(KEYINPUT35), .B(G1991), .Z(new_n873));
  AND2_X1   g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n872), .A2(new_n873), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n761), .A2(G24), .ZN(new_n876));
  INV_X1    g451(.A(G290), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n876), .B1(new_n877), .B2(new_n761), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(G1986), .ZN(new_n879));
  NOR3_X1   g454(.A1(new_n874), .A2(new_n875), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n860), .A2(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n851), .B1(new_n850), .B2(new_n859), .ZN(new_n882));
  OR3_X1    g457(.A1(new_n881), .A2(KEYINPUT36), .A3(new_n882), .ZN(new_n883));
  OAI21_X1  g458(.A(KEYINPUT36), .B1(new_n881), .B2(new_n882), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  AND2_X1   g460(.A1(new_n843), .A2(new_n885), .ZN(G311));
  INV_X1    g461(.A(KEYINPUT102), .ZN(new_n887));
  AND3_X1   g462(.A1(new_n843), .A2(new_n887), .A3(new_n885), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n887), .B1(new_n843), .B2(new_n885), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n888), .A2(new_n889), .ZN(G150));
  NAND2_X1  g465(.A1(new_n625), .A2(G559), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(KEYINPUT38), .ZN(new_n892));
  AOI22_X1  g467(.A1(new_n532), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n893), .A2(new_n526), .ZN(new_n894));
  XNOR2_X1  g469(.A(KEYINPUT103), .B(G93), .ZN(new_n895));
  INV_X1    g470(.A(G55), .ZN(new_n896));
  OAI22_X1  g471(.A1(new_n574), .A2(new_n895), .B1(new_n896), .B2(new_n576), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n894), .A2(new_n897), .ZN(new_n898));
  XOR2_X1   g473(.A(new_n579), .B(new_n898), .Z(new_n899));
  XNOR2_X1  g474(.A(new_n892), .B(new_n899), .ZN(new_n900));
  OR2_X1    g475(.A1(new_n900), .A2(KEYINPUT39), .ZN(new_n901));
  INV_X1    g476(.A(G860), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n900), .A2(KEYINPUT39), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n898), .A2(new_n902), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n905), .B(KEYINPUT37), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n904), .A2(new_n906), .ZN(G145));
  AND3_X1   g482(.A1(new_n869), .A2(KEYINPUT104), .A3(new_n870), .ZN(new_n908));
  AOI21_X1  g483(.A(KEYINPUT104), .B1(new_n869), .B2(new_n870), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n647), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT104), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n871), .A2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n647), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n869), .A2(KEYINPUT104), .A3(new_n870), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n910), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n832), .A2(new_n750), .ZN(new_n917));
  NAND4_X1  g492(.A1(new_n830), .A2(new_n741), .A3(new_n749), .A4(new_n831), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n916), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n498), .A2(G142), .ZN(new_n922));
  OR2_X1    g497(.A1(G106), .A2(G2105), .ZN(new_n923));
  OAI211_X1 g498(.A(new_n923), .B(G2104), .C1(G118), .C2(new_n467), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n925), .B1(G130), .B2(new_n493), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n521), .A2(new_n522), .ZN(new_n927));
  AND3_X1   g502(.A1(new_n817), .A2(new_n927), .A3(new_n818), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n927), .B1(new_n817), .B2(new_n818), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n926), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  OR3_X1    g505(.A1(new_n928), .A2(new_n926), .A3(new_n929), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n910), .A2(new_n915), .A3(new_n919), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n921), .A2(new_n930), .A3(new_n931), .A4(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n931), .A2(new_n930), .ZN(new_n934));
  AND3_X1   g509(.A1(new_n910), .A2(new_n915), .A3(new_n919), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n919), .B1(new_n910), .B2(new_n915), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n934), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n933), .A2(new_n937), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n643), .B(G160), .ZN(new_n939));
  XOR2_X1   g514(.A(new_n505), .B(new_n939), .Z(new_n940));
  AOI21_X1  g515(.A(G37), .B1(new_n938), .B2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n940), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n942), .A2(new_n933), .A3(new_n937), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n944), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g520(.A1(new_n625), .A2(new_n631), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n899), .A2(new_n946), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n579), .B(new_n898), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(new_n636), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n624), .A2(G299), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n615), .A2(new_n592), .A3(new_n589), .A4(new_n623), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n947), .A2(new_n949), .A3(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT105), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n954), .B(new_n955), .ZN(new_n956));
  XNOR2_X1  g531(.A(new_n952), .B(KEYINPUT41), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n947), .A2(new_n949), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n957), .A2(new_n958), .A3(KEYINPUT106), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n957), .A2(new_n958), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT106), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n956), .A2(new_n959), .A3(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(KEYINPUT42), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT42), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n956), .A2(new_n962), .A3(new_n965), .A4(new_n959), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  XOR2_X1   g542(.A(G288), .B(KEYINPUT107), .Z(new_n968));
  AND2_X1   g543(.A1(new_n968), .A2(new_n605), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n968), .A2(new_n605), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(G166), .A2(new_n877), .ZN(new_n972));
  NAND2_X1  g547(.A1(G303), .A2(G290), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n971), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n972), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n975), .B1(new_n969), .B2(new_n970), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n634), .B1(new_n967), .B2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(new_n977), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n964), .A2(new_n966), .A3(new_n979), .ZN(new_n980));
  AND3_X1   g555(.A1(new_n978), .A2(KEYINPUT108), .A3(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT108), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n982), .B1(new_n898), .B2(G868), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n983), .B1(new_n978), .B2(new_n980), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n981), .A2(new_n984), .ZN(G295));
  NOR2_X1   g560(.A1(new_n981), .A2(new_n984), .ZN(G331));
  INV_X1    g561(.A(KEYINPUT109), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n566), .A2(new_n567), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT82), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n566), .A2(KEYINPUT82), .A3(new_n567), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n987), .B1(new_n992), .B2(new_n564), .ZN(new_n993));
  OAI211_X1 g568(.A(new_n564), .B(new_n987), .C1(new_n568), .C2(new_n569), .ZN(new_n994));
  INV_X1    g569(.A(new_n994), .ZN(new_n995));
  OAI21_X1  g570(.A(G168), .B1(new_n993), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(G301), .A2(KEYINPUT109), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n997), .A2(new_n561), .A3(new_n557), .A4(new_n994), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n948), .B1(new_n996), .B2(new_n998), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n999), .A2(new_n952), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n996), .A2(new_n948), .A3(new_n998), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(KEYINPUT110), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT110), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n996), .A2(new_n998), .A3(new_n1003), .A4(new_n948), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1000), .A2(new_n1002), .A3(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(new_n1001), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n957), .B1(new_n1006), .B2(new_n999), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1005), .A2(new_n977), .A3(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(G37), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n977), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1011));
  OAI21_X1  g586(.A(KEYINPUT43), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n996), .A2(new_n998), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(new_n899), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1002), .A2(new_n1014), .A3(new_n1004), .ZN(new_n1015));
  AOI22_X1  g590(.A1(new_n1015), .A2(new_n957), .B1(new_n1001), .B2(new_n1000), .ZN(new_n1016));
  OAI211_X1 g591(.A(new_n1008), .B(new_n1009), .C1(new_n1016), .C2(new_n977), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1012), .B1(KEYINPUT43), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT43), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1019), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1020), .B1(new_n1019), .B2(new_n1017), .ZN(new_n1021));
  MUX2_X1   g596(.A(new_n1018), .B(new_n1021), .S(KEYINPUT44), .Z(G397));
  INV_X1    g597(.A(KEYINPUT62), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT45), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n511), .A2(new_n519), .A3(KEYINPUT75), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n523), .B1(new_n521), .B2(new_n522), .ZN(new_n1026));
  AOI211_X1 g601(.A(new_n1024), .B(G1384), .C1(new_n1025), .C2(new_n1026), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n483), .A2(new_n473), .A3(G40), .A4(new_n475), .ZN(new_n1028));
  INV_X1    g603(.A(G1384), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1029), .B1(new_n521), .B2(new_n522), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1028), .B1(new_n1030), .B2(new_n1024), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1031), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n770), .B1(new_n1027), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT50), .ZN(new_n1034));
  OAI211_X1 g609(.A(new_n1034), .B(new_n1029), .C1(new_n521), .C2(new_n522), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1028), .A2(G2084), .ZN(new_n1036));
  AOI21_X1  g611(.A(G1384), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1037));
  OAI211_X1 g612(.A(new_n1035), .B(new_n1036), .C1(new_n1037), .C2(new_n1034), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1033), .A2(G168), .A3(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(G8), .ZN(new_n1040));
  AOI21_X1  g615(.A(G168), .B1(new_n1033), .B2(new_n1038), .ZN(new_n1041));
  OAI21_X1  g616(.A(KEYINPUT51), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT123), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT51), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1039), .A2(new_n1044), .A3(G8), .ZN(new_n1045));
  AND3_X1   g620(.A1(new_n1042), .A2(new_n1043), .A3(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1043), .B1(new_n1042), .B2(new_n1045), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1023), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(G8), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1035), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1029), .B1(new_n520), .B2(new_n524), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1050), .B1(new_n1051), .B2(KEYINPUT50), .ZN(new_n1052));
  OAI211_X1 g627(.A(KEYINPUT45), .B(new_n1029), .C1(new_n520), .C2(new_n524), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(new_n1031), .ZN(new_n1054));
  AOI22_X1  g629(.A1(new_n1052), .A2(new_n1036), .B1(new_n1054), .B2(new_n770), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1049), .B1(new_n1055), .B2(G168), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1041), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1044), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1045), .ZN(new_n1059));
  OAI21_X1  g634(.A(KEYINPUT123), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1042), .A2(new_n1043), .A3(new_n1045), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1060), .A2(KEYINPUT62), .A3(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1051), .A2(KEYINPUT50), .ZN(new_n1063));
  INV_X1    g638(.A(G2090), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1028), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1063), .A2(new_n1064), .A3(new_n1065), .A4(new_n1035), .ZN(new_n1066));
  AOI21_X1  g641(.A(G1384), .B1(new_n511), .B2(new_n519), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1028), .B1(new_n1067), .B2(KEYINPUT45), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1068), .B1(new_n1037), .B2(KEYINPUT45), .ZN(new_n1069));
  INV_X1    g644(.A(G1971), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1049), .B1(new_n1066), .B2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n542), .A2(G8), .A3(new_n544), .ZN(new_n1073));
  XNOR2_X1  g648(.A(KEYINPUT114), .B(KEYINPUT55), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n542), .A2(new_n544), .A3(G8), .A4(new_n1074), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(KEYINPUT115), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT115), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1076), .A2(new_n1080), .A3(new_n1077), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1072), .A2(new_n1082), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1030), .A2(new_n1028), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1084), .A2(new_n1049), .ZN(new_n1085));
  INV_X1    g660(.A(G1976), .ZN(new_n1086));
  AOI21_X1  g661(.A(KEYINPUT52), .B1(G288), .B2(new_n1086), .ZN(new_n1087));
  OAI211_X1 g662(.A(new_n1085), .B(new_n1087), .C1(new_n1086), .C2(G288), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1067), .A2(new_n1065), .ZN(new_n1089));
  OAI211_X1 g664(.A(new_n1089), .B(G8), .C1(new_n1086), .C2(G288), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(KEYINPUT52), .ZN(new_n1091));
  NOR3_X1   g666(.A1(new_n601), .A2(new_n604), .A3(G1981), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1092), .ZN(new_n1093));
  OAI21_X1  g668(.A(G1981), .B1(new_n601), .B2(new_n604), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1093), .A2(KEYINPUT49), .A3(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT49), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1094), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1096), .B1(new_n1097), .B2(new_n1092), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1095), .A2(new_n1098), .A3(new_n1085), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1088), .A2(new_n1091), .A3(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1100), .ZN(new_n1101));
  AOI211_X1 g676(.A(KEYINPUT50), .B(G1384), .C1(new_n1025), .C2(new_n1026), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1028), .B1(new_n1030), .B2(KEYINPUT50), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(KEYINPUT116), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1105));
  OAI211_X1 g680(.A(new_n1034), .B(new_n1029), .C1(new_n520), .C2(new_n524), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT116), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1106), .A2(new_n1107), .A3(new_n1103), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1105), .A2(new_n1064), .A3(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1049), .B1(new_n1109), .B2(new_n1071), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1078), .ZN(new_n1111));
  OAI211_X1 g686(.A(new_n1083), .B(new_n1101), .C1(new_n1110), .C2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT53), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1113), .B1(new_n1069), .B2(G2078), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1113), .A2(G2078), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1053), .A2(new_n1031), .A3(new_n1115), .ZN(new_n1116));
  OAI211_X1 g691(.A(new_n1065), .B(new_n1035), .C1(new_n1037), .C2(new_n1034), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(new_n764), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1114), .A2(new_n1116), .A3(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(G171), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1112), .A2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1048), .A2(new_n1062), .A3(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1051), .A2(new_n1024), .ZN(new_n1123));
  AOI21_X1  g698(.A(G1971), .B1(new_n1123), .B2(new_n1068), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1106), .A2(new_n1103), .ZN(new_n1125));
  AOI21_X1  g700(.A(G2090), .B1(new_n1125), .B2(KEYINPUT116), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1124), .B1(new_n1126), .B2(new_n1108), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1078), .B1(new_n1127), .B2(new_n1049), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1100), .B1(new_n1072), .B2(new_n1082), .ZN(new_n1129));
  NOR3_X1   g704(.A1(new_n1055), .A2(new_n1049), .A3(G286), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1128), .A2(new_n1129), .A3(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(KEYINPUT117), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT63), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT117), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1128), .A2(new_n1129), .A3(new_n1134), .A4(new_n1130), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1132), .A2(new_n1133), .A3(new_n1135), .ZN(new_n1136));
  AND2_X1   g711(.A1(new_n1130), .A2(KEYINPUT63), .ZN(new_n1137));
  AND2_X1   g712(.A1(new_n1072), .A2(KEYINPUT118), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1078), .B1(new_n1072), .B2(KEYINPUT118), .ZN(new_n1139));
  OAI211_X1 g714(.A(new_n1137), .B(new_n1129), .C1(new_n1138), .C2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1136), .A2(new_n1140), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1067), .A2(KEYINPUT45), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n483), .A2(G40), .A3(new_n1115), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT125), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1144), .B1(new_n1145), .B2(new_n476), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1030), .A2(new_n1024), .ZN(new_n1147));
  INV_X1    g722(.A(new_n476), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1148), .A2(KEYINPUT125), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n1143), .A2(new_n1146), .A3(new_n1147), .A4(new_n1149), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1114), .A2(new_n1118), .A3(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1151), .A2(G171), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1114), .A2(G301), .A3(new_n1118), .A4(new_n1116), .ZN(new_n1153));
  AND3_X1   g728(.A1(new_n1152), .A2(KEYINPUT54), .A3(new_n1153), .ZN(new_n1154));
  XOR2_X1   g729(.A(KEYINPUT124), .B(KEYINPUT54), .Z(new_n1155));
  NAND4_X1  g730(.A1(new_n1114), .A2(G301), .A3(new_n1118), .A4(new_n1150), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1155), .B1(new_n1120), .B2(new_n1156), .ZN(new_n1157));
  NOR3_X1   g732(.A1(new_n1154), .A2(new_n1112), .A3(new_n1157), .ZN(new_n1158));
  XNOR2_X1  g733(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n1159));
  XNOR2_X1  g734(.A(G299), .B(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(new_n1160), .ZN(new_n1161));
  XNOR2_X1  g736(.A(KEYINPUT56), .B(G2072), .ZN(new_n1162));
  OAI211_X1 g737(.A(new_n1068), .B(new_n1162), .C1(new_n1037), .C2(KEYINPUT45), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1163), .ZN(new_n1164));
  AOI21_X1  g739(.A(G1956), .B1(new_n1106), .B2(new_n1103), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1161), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1125), .A2(new_n795), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1168), .A2(new_n1160), .A3(new_n1163), .ZN(new_n1169));
  AND2_X1   g744(.A1(new_n1169), .A2(new_n625), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1117), .A2(new_n777), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT120), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1172), .B1(new_n1089), .B2(G2067), .ZN(new_n1173));
  INV_X1    g748(.A(G2067), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1084), .A2(KEYINPUT120), .A3(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1173), .A2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1171), .A2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1167), .B1(new_n1170), .B2(new_n1177), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT60), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1177), .A2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1171), .A2(new_n1176), .A3(KEYINPUT60), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1180), .A2(new_n625), .A3(new_n1181), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT122), .ZN(new_n1183));
  AND3_X1   g758(.A1(new_n1166), .A2(new_n1183), .A3(new_n1169), .ZN(new_n1184));
  XNOR2_X1  g759(.A(KEYINPUT121), .B(KEYINPUT61), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1185), .B1(new_n1166), .B2(new_n1183), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1182), .B1(new_n1184), .B2(new_n1186), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1166), .A2(KEYINPUT61), .A3(new_n1169), .ZN(new_n1188));
  NAND4_X1  g763(.A1(new_n1171), .A2(KEYINPUT60), .A3(new_n624), .A4(new_n1176), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT59), .ZN(new_n1190));
  INV_X1    g765(.A(G1996), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1123), .A2(new_n1191), .A3(new_n1068), .ZN(new_n1192));
  XOR2_X1   g767(.A(KEYINPUT58), .B(G1341), .Z(new_n1193));
  NAND2_X1  g768(.A1(new_n1089), .A2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1192), .A2(new_n1194), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1190), .B1(new_n1195), .B2(new_n579), .ZN(new_n1196));
  AOI211_X1 g771(.A(KEYINPUT59), .B(new_n633), .C1(new_n1192), .C2(new_n1194), .ZN(new_n1197));
  OAI211_X1 g772(.A(new_n1188), .B(new_n1189), .C1(new_n1196), .C2(new_n1197), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n1178), .B1(new_n1187), .B2(new_n1198), .ZN(new_n1199));
  NAND3_X1  g774(.A1(new_n1142), .A2(new_n1158), .A3(new_n1199), .ZN(new_n1200));
  NOR2_X1   g775(.A1(new_n1083), .A2(new_n1100), .ZN(new_n1201));
  INV_X1    g776(.A(new_n1099), .ZN(new_n1202));
  OR2_X1    g777(.A1(G288), .A2(G1976), .ZN(new_n1203));
  OAI21_X1  g778(.A(new_n1093), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g779(.A(new_n1201), .B1(new_n1204), .B2(new_n1085), .ZN(new_n1205));
  NAND4_X1  g780(.A1(new_n1122), .A2(new_n1141), .A3(new_n1200), .A4(new_n1205), .ZN(new_n1206));
  NOR2_X1   g781(.A1(new_n1147), .A2(new_n1028), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1207), .A2(new_n1191), .ZN(new_n1208));
  XOR2_X1   g783(.A(new_n1208), .B(KEYINPUT111), .Z(new_n1209));
  NOR2_X1   g784(.A1(new_n1209), .A2(new_n819), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n832), .A2(G2067), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n819), .A2(G1996), .ZN(new_n1212));
  NAND3_X1  g787(.A1(new_n830), .A2(new_n1174), .A3(new_n831), .ZN(new_n1213));
  NAND3_X1  g788(.A1(new_n1211), .A2(new_n1212), .A3(new_n1213), .ZN(new_n1214));
  AOI21_X1  g789(.A(new_n1210), .B1(new_n1207), .B2(new_n1214), .ZN(new_n1215));
  INV_X1    g790(.A(new_n1207), .ZN(new_n1216));
  XNOR2_X1  g791(.A(new_n871), .B(new_n873), .ZN(new_n1217));
  INV_X1    g792(.A(KEYINPUT112), .ZN(new_n1218));
  AOI21_X1  g793(.A(new_n1216), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  OAI21_X1  g794(.A(new_n1219), .B1(new_n1218), .B2(new_n1217), .ZN(new_n1220));
  XOR2_X1   g795(.A(G290), .B(G1986), .Z(new_n1221));
  OAI211_X1 g796(.A(new_n1215), .B(new_n1220), .C1(new_n1216), .C2(new_n1221), .ZN(new_n1222));
  XNOR2_X1  g797(.A(new_n1222), .B(KEYINPUT113), .ZN(new_n1223));
  NAND2_X1  g798(.A1(new_n1206), .A2(new_n1223), .ZN(new_n1224));
  XNOR2_X1  g799(.A(new_n1209), .B(KEYINPUT46), .ZN(new_n1225));
  NAND2_X1  g800(.A1(new_n1211), .A2(new_n1213), .ZN(new_n1226));
  OAI21_X1  g801(.A(new_n1207), .B1(new_n1226), .B2(new_n819), .ZN(new_n1227));
  NAND2_X1  g802(.A1(new_n1225), .A2(new_n1227), .ZN(new_n1228));
  XOR2_X1   g803(.A(new_n1228), .B(KEYINPUT47), .Z(new_n1229));
  NAND4_X1  g804(.A1(new_n1215), .A2(new_n873), .A3(new_n869), .A4(new_n870), .ZN(new_n1230));
  AOI21_X1  g805(.A(new_n1216), .B1(new_n1230), .B2(new_n1213), .ZN(new_n1231));
  NOR3_X1   g806(.A1(new_n1216), .A2(G1986), .A3(G290), .ZN(new_n1232));
  XOR2_X1   g807(.A(new_n1232), .B(KEYINPUT48), .Z(new_n1233));
  AND3_X1   g808(.A1(new_n1215), .A2(new_n1220), .A3(new_n1233), .ZN(new_n1234));
  NOR3_X1   g809(.A1(new_n1229), .A2(new_n1231), .A3(new_n1234), .ZN(new_n1235));
  NAND2_X1  g810(.A1(new_n1224), .A2(new_n1235), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g811(.A1(new_n696), .A2(G319), .A3(new_n697), .ZN(new_n1238));
  AOI21_X1  g812(.A(new_n1238), .B1(new_n725), .B2(new_n730), .ZN(new_n1239));
  INV_X1    g813(.A(KEYINPUT126), .ZN(new_n1240));
  AND3_X1   g814(.A1(new_n1239), .A2(new_n1240), .A3(new_n674), .ZN(new_n1241));
  AOI21_X1  g815(.A(new_n1240), .B1(new_n1239), .B2(new_n674), .ZN(new_n1242));
  NOR2_X1   g816(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  AOI21_X1  g817(.A(new_n1243), .B1(new_n941), .B2(new_n943), .ZN(new_n1244));
  INV_X1    g818(.A(KEYINPUT127), .ZN(new_n1245));
  AND3_X1   g819(.A1(new_n1244), .A2(new_n1245), .A3(new_n1018), .ZN(new_n1246));
  AOI21_X1  g820(.A(new_n1245), .B1(new_n1244), .B2(new_n1018), .ZN(new_n1247));
  NOR2_X1   g821(.A1(new_n1246), .A2(new_n1247), .ZN(G308));
  NAND2_X1  g822(.A1(new_n1244), .A2(new_n1018), .ZN(new_n1249));
  NAND2_X1  g823(.A1(new_n1249), .A2(KEYINPUT127), .ZN(new_n1250));
  NAND3_X1  g824(.A1(new_n1244), .A2(new_n1245), .A3(new_n1018), .ZN(new_n1251));
  NAND2_X1  g825(.A1(new_n1250), .A2(new_n1251), .ZN(G225));
endmodule


