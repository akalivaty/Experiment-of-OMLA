//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 1 0 1 0 0 1 0 1 1 0 1 1 0 1 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 1 1 0 0 0 1 1 1 0 1 1 1 0 0 0 1 1 1 1 1 0 0 1 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:47 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n785, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n806, new_n807, new_n808, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n919,
    new_n920, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993;
  INV_X1    g000(.A(G221), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT9), .B(G234), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G902), .ZN(new_n190));
  AOI21_X1  g004(.A(new_n187), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G146), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G143), .ZN(new_n193));
  INV_X1    g007(.A(G143), .ZN(new_n194));
  AND3_X1   g008(.A1(new_n194), .A2(KEYINPUT64), .A3(G146), .ZN(new_n195));
  AOI21_X1  g009(.A(KEYINPUT64), .B1(new_n194), .B2(G146), .ZN(new_n196));
  OAI211_X1 g010(.A(G128), .B(new_n193), .C1(new_n195), .C2(new_n196), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n194), .A2(G146), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT64), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n199), .B1(new_n192), .B2(G143), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n194), .A2(KEYINPUT64), .A3(G146), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n198), .B1(new_n200), .B2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G128), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n203), .B1(new_n193), .B2(KEYINPUT1), .ZN(new_n204));
  OAI22_X1  g018(.A1(new_n197), .A2(KEYINPUT1), .B1(new_n202), .B2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G104), .ZN(new_n206));
  OAI21_X1  g020(.A(KEYINPUT3), .B1(new_n206), .B2(G107), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT3), .ZN(new_n208));
  INV_X1    g022(.A(G107), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n208), .A2(new_n209), .A3(G104), .ZN(new_n210));
  INV_X1    g024(.A(G101), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n206), .A2(G107), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n207), .A2(new_n210), .A3(new_n211), .A4(new_n212), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n206), .A2(G107), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n209), .A2(G104), .ZN(new_n215));
  OAI21_X1  g029(.A(G101), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n213), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n205), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(KEYINPUT76), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT76), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n205), .A2(new_n221), .A3(new_n218), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT1), .ZN(new_n224));
  OAI21_X1  g038(.A(G128), .B1(new_n198), .B2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT67), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n194), .A2(G146), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n193), .A2(new_n227), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n225), .A2(new_n226), .A3(new_n228), .ZN(new_n229));
  XNOR2_X1  g043(.A(G143), .B(G146), .ZN(new_n230));
  OAI21_X1  g044(.A(KEYINPUT67), .B1(new_n204), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n202), .A2(new_n224), .A3(G128), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n232), .A2(new_n233), .A3(new_n217), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n223), .A2(new_n234), .ZN(new_n235));
  OR2_X1    g049(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n236));
  INV_X1    g050(.A(G137), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(G134), .ZN(new_n238));
  NAND2_X1  g052(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n236), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  OR2_X1    g054(.A1(KEYINPUT66), .A2(G137), .ZN(new_n241));
  NAND2_X1  g055(.A1(KEYINPUT66), .A2(G137), .ZN(new_n242));
  AND2_X1   g056(.A1(KEYINPUT11), .A2(G134), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n241), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(G134), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(G137), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n240), .A2(new_n244), .A3(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(G131), .ZN(new_n248));
  INV_X1    g062(.A(G131), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n240), .A2(new_n244), .A3(new_n249), .A4(new_n246), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  OR2_X1    g065(.A1(KEYINPUT78), .A2(KEYINPUT12), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n235), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(new_n251), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n254), .B1(new_n223), .B2(new_n234), .ZN(new_n255));
  XOR2_X1   g069(.A(KEYINPUT78), .B(KEYINPUT12), .Z(new_n256));
  OAI21_X1  g070(.A(new_n253), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n213), .A2(KEYINPUT4), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n207), .A2(new_n210), .A3(new_n212), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G101), .ZN(new_n260));
  XNOR2_X1  g074(.A(new_n258), .B(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT0), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n262), .B1(new_n228), .B2(new_n203), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(new_n197), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n262), .B1(new_n230), .B2(new_n203), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n261), .A2(new_n266), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n226), .B1(new_n225), .B2(new_n228), .ZN(new_n268));
  NOR3_X1   g082(.A1(new_n204), .A2(new_n230), .A3(KEYINPUT67), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n233), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n270), .A2(KEYINPUT10), .A3(new_n218), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n267), .A2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT77), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT10), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n274), .B1(new_n223), .B2(new_n275), .ZN(new_n276));
  AND3_X1   g090(.A1(new_n205), .A2(new_n221), .A3(new_n218), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n221), .B1(new_n205), .B2(new_n218), .ZN(new_n278));
  OAI211_X1 g092(.A(new_n274), .B(new_n275), .C1(new_n277), .C2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  OAI211_X1 g094(.A(new_n254), .B(new_n273), .C1(new_n276), .C2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n257), .A2(new_n281), .ZN(new_n282));
  XNOR2_X1  g096(.A(G110), .B(G140), .ZN(new_n283));
  INV_X1    g097(.A(G953), .ZN(new_n284));
  AND2_X1   g098(.A1(new_n284), .A2(G227), .ZN(new_n285));
  XNOR2_X1  g099(.A(new_n283), .B(new_n285), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n275), .B1(new_n277), .B2(new_n278), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(KEYINPUT77), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n272), .B1(new_n288), .B2(new_n279), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n286), .B1(new_n289), .B2(new_n254), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n273), .B1(new_n276), .B2(new_n280), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(new_n251), .ZN(new_n292));
  AOI22_X1  g106(.A1(new_n282), .A2(new_n286), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  OAI21_X1  g107(.A(G469), .B1(new_n293), .B2(G902), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT79), .ZN(new_n295));
  INV_X1    g109(.A(G469), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n289), .A2(new_n254), .ZN(new_n297));
  AOI211_X1 g111(.A(new_n251), .B(new_n272), .C1(new_n288), .C2(new_n279), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n286), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n290), .A2(new_n257), .ZN(new_n300));
  AOI21_X1  g114(.A(G902), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  AOI22_X1  g115(.A1(new_n294), .A2(new_n295), .B1(new_n296), .B2(new_n301), .ZN(new_n302));
  OAI211_X1 g116(.A(KEYINPUT79), .B(G469), .C1(new_n293), .C2(G902), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n191), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NOR2_X1   g118(.A1(G475), .A2(G902), .ZN(new_n305));
  XNOR2_X1  g119(.A(G113), .B(G122), .ZN(new_n306));
  XNOR2_X1  g120(.A(new_n306), .B(new_n206), .ZN(new_n307));
  INV_X1    g121(.A(G140), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(G125), .ZN(new_n309));
  INV_X1    g123(.A(G125), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(G140), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  OR2_X1    g126(.A1(new_n312), .A2(KEYINPUT87), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(KEYINPUT87), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n313), .A2(KEYINPUT19), .A3(new_n314), .ZN(new_n315));
  OR2_X1    g129(.A1(new_n312), .A2(KEYINPUT19), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n315), .A2(new_n192), .A3(new_n316), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n309), .A2(KEYINPUT16), .ZN(new_n318));
  INV_X1    g132(.A(new_n312), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n318), .B1(new_n319), .B2(KEYINPUT16), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(G146), .ZN(new_n321));
  NOR2_X1   g135(.A1(G237), .A2(G953), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n322), .A2(G143), .A3(G214), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  AOI21_X1  g138(.A(G143), .B1(new_n322), .B2(G214), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(new_n249), .ZN(new_n327));
  INV_X1    g141(.A(new_n325), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(new_n323), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(G131), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n327), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n317), .A2(new_n321), .A3(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n313), .A2(G146), .A3(new_n314), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n319), .A2(new_n192), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT88), .ZN(new_n336));
  NAND2_X1  g150(.A1(KEYINPUT18), .A2(G131), .ZN(new_n337));
  NOR3_X1   g151(.A1(new_n329), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  AOI22_X1  g152(.A1(new_n326), .A2(KEYINPUT88), .B1(KEYINPUT18), .B2(G131), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n335), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n307), .B1(new_n332), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(KEYINPUT89), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT16), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n312), .A2(new_n343), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n192), .B1(new_n344), .B2(new_n318), .ZN(new_n345));
  AND2_X1   g159(.A1(new_n321), .A2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT17), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n327), .A2(new_n330), .A3(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n329), .A2(KEYINPUT17), .A3(G131), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n346), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n350), .A2(new_n307), .A3(new_n340), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n342), .A2(new_n351), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n341), .A2(KEYINPUT89), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n305), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(KEYINPUT20), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT20), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n356), .B(new_n305), .C1(new_n352), .C2(new_n353), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n350), .A2(new_n340), .ZN(new_n358));
  INV_X1    g172(.A(new_n307), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(new_n351), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(new_n190), .ZN(new_n362));
  AOI22_X1  g176(.A1(new_n355), .A2(new_n357), .B1(G475), .B2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(G217), .ZN(new_n365));
  NOR3_X1   g179(.A1(new_n188), .A2(new_n365), .A3(G953), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT69), .ZN(new_n367));
  INV_X1    g181(.A(G116), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(KEYINPUT69), .A2(G116), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n369), .A2(G122), .A3(new_n370), .ZN(new_n371));
  AND2_X1   g185(.A1(new_n371), .A2(KEYINPUT14), .ZN(new_n372));
  OAI21_X1  g186(.A(KEYINPUT90), .B1(new_n368), .B2(G122), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT90), .ZN(new_n374));
  INV_X1    g188(.A(G122), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n374), .A2(new_n375), .A3(G116), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n373), .A2(new_n376), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n377), .B1(new_n371), .B2(KEYINPUT14), .ZN(new_n378));
  OAI21_X1  g192(.A(G107), .B1(new_n372), .B2(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n377), .A2(new_n371), .A3(new_n209), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n203), .A2(G143), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n194), .A2(G128), .ZN(new_n382));
  NOR3_X1   g196(.A1(new_n381), .A2(new_n382), .A3(G134), .ZN(new_n383));
  INV_X1    g197(.A(new_n382), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n194), .A2(G128), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n245), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  OAI211_X1 g200(.A(new_n379), .B(new_n380), .C1(new_n383), .C2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(new_n383), .ZN(new_n388));
  INV_X1    g202(.A(new_n380), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n209), .B1(new_n377), .B2(new_n371), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n388), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT13), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n392), .B1(new_n203), .B2(G143), .ZN(new_n393));
  OAI21_X1  g207(.A(KEYINPUT91), .B1(new_n393), .B2(new_n381), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT91), .ZN(new_n395));
  OAI211_X1 g209(.A(new_n395), .B(new_n385), .C1(new_n382), .C2(new_n392), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n381), .A2(KEYINPUT13), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n394), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(G134), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT92), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n398), .A2(KEYINPUT92), .A3(G134), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n391), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n387), .B1(new_n403), .B2(KEYINPUT93), .ZN(new_n404));
  INV_X1    g218(.A(new_n391), .ZN(new_n405));
  INV_X1    g219(.A(new_n402), .ZN(new_n406));
  AOI21_X1  g220(.A(KEYINPUT92), .B1(new_n398), .B2(G134), .ZN(new_n407));
  OAI211_X1 g221(.A(new_n405), .B(KEYINPUT93), .C1(new_n406), .C2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n366), .B1(new_n404), .B2(new_n409), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n405), .B1(new_n406), .B2(new_n407), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT93), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(new_n366), .ZN(new_n414));
  NAND4_X1  g228(.A1(new_n413), .A2(new_n408), .A3(new_n387), .A4(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n410), .A2(new_n190), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(KEYINPUT94), .ZN(new_n417));
  INV_X1    g231(.A(G478), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n418), .A2(KEYINPUT15), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT94), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n410), .A2(new_n420), .A3(new_n415), .A4(new_n190), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n417), .A2(new_n419), .A3(new_n421), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n422), .B1(new_n416), .B2(new_n419), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n364), .A2(new_n423), .ZN(new_n424));
  AND2_X1   g238(.A1(new_n304), .A2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(G119), .ZN(new_n426));
  OR3_X1    g240(.A1(new_n426), .A2(KEYINPUT75), .A3(G128), .ZN(new_n427));
  OAI21_X1  g241(.A(KEYINPUT75), .B1(new_n426), .B2(G128), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n426), .A2(G128), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n427), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  XNOR2_X1  g244(.A(KEYINPUT24), .B(G110), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n203), .A2(KEYINPUT23), .A3(G119), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n426), .A2(G128), .ZN(new_n434));
  OAI211_X1 g248(.A(new_n429), .B(new_n433), .C1(new_n434), .C2(KEYINPUT23), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n432), .B1(G110), .B2(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n436), .A2(new_n321), .A3(new_n334), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n435), .A2(G110), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n438), .B1(new_n430), .B2(new_n431), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n437), .B1(new_n346), .B2(new_n439), .ZN(new_n440));
  XNOR2_X1  g254(.A(KEYINPUT22), .B(G137), .ZN(new_n441));
  AND3_X1   g255(.A1(new_n284), .A2(G221), .A3(G234), .ZN(new_n442));
  XOR2_X1   g256(.A(new_n441), .B(new_n442), .Z(new_n443));
  XNOR2_X1  g257(.A(new_n440), .B(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(new_n190), .ZN(new_n445));
  XOR2_X1   g259(.A(new_n445), .B(KEYINPUT25), .Z(new_n446));
  AOI21_X1  g260(.A(new_n365), .B1(G234), .B2(new_n190), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n447), .A2(G902), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n444), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT2), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n452), .A2(G113), .ZN(new_n453));
  INV_X1    g267(.A(G113), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n454), .A2(KEYINPUT2), .ZN(new_n455));
  OAI21_X1  g269(.A(KEYINPUT68), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n454), .A2(KEYINPUT2), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n452), .A2(G113), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT68), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n457), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n456), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n369), .A2(G119), .A3(new_n370), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT70), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND4_X1  g278(.A1(new_n369), .A2(KEYINPUT70), .A3(G119), .A4(new_n370), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n368), .A2(G119), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n461), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n467), .B1(new_n457), .B2(new_n458), .ZN(new_n470));
  AND2_X1   g284(.A1(KEYINPUT69), .A2(G116), .ZN(new_n471));
  NOR2_X1   g285(.A1(KEYINPUT69), .A2(G116), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  AOI21_X1  g287(.A(KEYINPUT70), .B1(new_n473), .B2(G119), .ZN(new_n474));
  INV_X1    g288(.A(new_n465), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n470), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(KEYINPUT71), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT71), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n466), .A2(new_n478), .A3(new_n470), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n469), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT72), .ZN(new_n481));
  AOI21_X1  g295(.A(G134), .B1(new_n241), .B2(new_n242), .ZN(new_n482));
  INV_X1    g296(.A(new_n238), .ZN(new_n483));
  OAI21_X1  g297(.A(G131), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(new_n250), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n485), .B1(new_n233), .B2(new_n232), .ZN(new_n486));
  AOI22_X1  g300(.A1(new_n250), .A2(new_n248), .B1(new_n264), .B2(new_n265), .ZN(new_n487));
  OAI211_X1 g301(.A(new_n481), .B(KEYINPUT30), .C1(new_n486), .C2(new_n487), .ZN(new_n488));
  AND2_X1   g302(.A1(new_n484), .A2(new_n250), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n270), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n251), .A2(new_n266), .ZN(new_n491));
  OR2_X1    g305(.A1(new_n481), .A2(KEYINPUT30), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n481), .A2(KEYINPUT30), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n490), .A2(new_n491), .A3(new_n492), .A4(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n480), .B1(new_n488), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n322), .A2(G210), .ZN(new_n496));
  XOR2_X1   g310(.A(new_n496), .B(KEYINPUT27), .Z(new_n497));
  XNOR2_X1  g311(.A(KEYINPUT26), .B(G101), .ZN(new_n498));
  XNOR2_X1  g312(.A(new_n497), .B(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n477), .A2(new_n479), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n468), .B1(new_n474), .B2(new_n475), .ZN(new_n501));
  INV_X1    g315(.A(new_n461), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n500), .A2(new_n490), .A3(new_n491), .A4(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  NOR3_X1   g319(.A1(new_n495), .A2(new_n499), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(G902), .B1(new_n506), .B2(KEYINPUT31), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n488), .A2(new_n494), .ZN(new_n508));
  AND3_X1   g322(.A1(new_n466), .A2(new_n478), .A3(new_n470), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n478), .B1(new_n466), .B2(new_n470), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n503), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(new_n499), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n512), .A2(new_n513), .A3(new_n504), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT28), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n490), .A2(new_n491), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(new_n511), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n515), .B1(new_n517), .B2(new_n504), .ZN(new_n518));
  AND2_X1   g332(.A1(new_n504), .A2(new_n515), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n499), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT31), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n514), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(G472), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n507), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT32), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND4_X1  g340(.A1(new_n507), .A2(new_n522), .A3(KEYINPUT32), .A4(new_n523), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n526), .A2(KEYINPUT74), .A3(new_n527), .ZN(new_n528));
  AND2_X1   g342(.A1(new_n507), .A2(new_n522), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT74), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n529), .A2(new_n530), .A3(KEYINPUT32), .A4(new_n523), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  NOR3_X1   g346(.A1(new_n518), .A2(new_n519), .A3(new_n499), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n533), .A2(KEYINPUT29), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT73), .ZN(new_n535));
  OAI211_X1 g349(.A(new_n535), .B(new_n499), .C1(new_n495), .C2(new_n505), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n495), .A2(new_n505), .ZN(new_n537));
  OAI21_X1  g351(.A(KEYINPUT73), .B1(new_n537), .B2(new_n513), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n534), .A2(new_n536), .A3(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(G902), .B1(new_n533), .B2(KEYINPUT29), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(G472), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n451), .B1(new_n532), .B2(new_n542), .ZN(new_n543));
  OAI21_X1  g357(.A(G214), .B1(G237), .B2(G902), .ZN(new_n544));
  OAI21_X1  g358(.A(G210), .B1(G237), .B2(G902), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT6), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n546), .A2(KEYINPUT83), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  XNOR2_X1  g362(.A(G110), .B(G122), .ZN(new_n549));
  XOR2_X1   g363(.A(new_n549), .B(KEYINPUT82), .Z(new_n550));
  OAI211_X1 g364(.A(KEYINPUT5), .B(new_n468), .C1(new_n474), .C2(new_n475), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT5), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n454), .B1(new_n467), .B2(new_n552), .ZN(new_n553));
  AOI221_X4 g367(.A(new_n217), .B1(new_n551), .B2(new_n553), .C1(new_n477), .C2(new_n479), .ZN(new_n554));
  XOR2_X1   g368(.A(new_n258), .B(new_n260), .Z(new_n555));
  OAI21_X1  g369(.A(KEYINPUT80), .B1(new_n480), .B2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT80), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n511), .A2(new_n557), .A3(new_n261), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n554), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT81), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n550), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  AOI211_X1 g375(.A(KEYINPUT81), .B(new_n554), .C1(new_n558), .C2(new_n556), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n548), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(new_n554), .ZN(new_n564));
  NOR3_X1   g378(.A1(new_n480), .A2(new_n555), .A3(KEYINPUT80), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n557), .B1(new_n511), .B2(new_n261), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n564), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(KEYINPUT81), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n559), .A2(new_n560), .ZN(new_n569));
  NAND4_X1  g383(.A1(new_n568), .A2(new_n569), .A3(new_n547), .A4(new_n550), .ZN(new_n570));
  AND2_X1   g384(.A1(new_n559), .A2(new_n549), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(KEYINPUT6), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n563), .A2(new_n570), .A3(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(G125), .B1(new_n232), .B2(new_n233), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n310), .B1(new_n264), .B2(new_n265), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n284), .A2(G224), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n576), .B(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n573), .A2(new_n579), .ZN(new_n580));
  OAI211_X1 g394(.A(KEYINPUT7), .B(new_n577), .C1(new_n574), .C2(new_n575), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT86), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT85), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT7), .ZN(new_n584));
  AOI22_X1  g398(.A1(new_n583), .A2(new_n584), .B1(new_n284), .B2(G224), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n585), .B1(new_n583), .B2(new_n584), .ZN(new_n586));
  AOI22_X1  g400(.A1(new_n581), .A2(new_n582), .B1(new_n576), .B2(new_n586), .ZN(new_n587));
  OR2_X1    g401(.A1(new_n581), .A2(new_n582), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n551), .A2(new_n553), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n218), .B1(new_n500), .B2(new_n589), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n217), .B1(new_n477), .B2(new_n479), .ZN(new_n591));
  OR2_X1    g405(.A1(new_n551), .A2(KEYINPUT84), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n551), .A2(KEYINPUT84), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n592), .A2(new_n553), .A3(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n590), .B1(new_n591), .B2(new_n594), .ZN(new_n595));
  XOR2_X1   g409(.A(new_n549), .B(KEYINPUT8), .Z(new_n596));
  OAI211_X1 g410(.A(new_n587), .B(new_n588), .C1(new_n595), .C2(new_n596), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n190), .B1(new_n571), .B2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n545), .B1(new_n580), .B2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n545), .ZN(new_n601));
  AOI211_X1 g415(.A(new_n598), .B(new_n601), .C1(new_n573), .C2(new_n579), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n544), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(G952), .ZN(new_n604));
  AOI211_X1 g418(.A(G953), .B(new_n604), .C1(G234), .C2(G237), .ZN(new_n605));
  AOI211_X1 g419(.A(new_n190), .B(new_n284), .C1(G234), .C2(G237), .ZN(new_n606));
  XNOR2_X1  g420(.A(KEYINPUT21), .B(G898), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n605), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n603), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n425), .A2(new_n543), .A3(new_n609), .ZN(new_n610));
  XNOR2_X1  g424(.A(KEYINPUT95), .B(G101), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(KEYINPUT96), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n610), .B(new_n612), .ZN(G3));
  INV_X1    g427(.A(new_n304), .ZN(new_n614));
  OR2_X1    g428(.A1(new_n529), .A2(new_n523), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(new_n524), .ZN(new_n616));
  NOR3_X1   g430(.A1(new_n614), .A2(new_n451), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n603), .A2(KEYINPUT97), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT97), .ZN(new_n619));
  OAI211_X1 g433(.A(new_n619), .B(new_n544), .C1(new_n600), .C2(new_n602), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n608), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n417), .A2(new_n418), .A3(new_n421), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT100), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n417), .A2(KEYINPUT100), .A3(new_n418), .A4(new_n421), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n414), .A2(KEYINPUT98), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n627), .B1(new_n404), .B2(new_n409), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n413), .A2(new_n408), .A3(new_n387), .A4(new_n626), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n628), .A2(KEYINPUT33), .A3(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT99), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n628), .A2(KEYINPUT99), .A3(new_n629), .A4(KEYINPUT33), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT33), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n410), .A2(new_n634), .A3(new_n415), .ZN(new_n635));
  AND3_X1   g449(.A1(new_n632), .A2(new_n633), .A3(new_n635), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n418), .A2(G902), .ZN(new_n637));
  AOI22_X1  g451(.A1(new_n624), .A2(new_n625), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n638), .A2(new_n363), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n617), .A2(new_n621), .A3(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(G104), .ZN(new_n641));
  XNOR2_X1  g455(.A(KEYINPUT101), .B(KEYINPUT34), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G6));
  NAND3_X1  g457(.A1(new_n362), .A2(KEYINPUT103), .A3(G475), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT103), .ZN(new_n645));
  AOI21_X1  g459(.A(G902), .B1(new_n360), .B2(new_n351), .ZN(new_n646));
  INV_X1    g460(.A(G475), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n645), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n644), .A2(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(new_n357), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n355), .B1(new_n650), .B2(KEYINPUT102), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT102), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n354), .A2(new_n652), .A3(KEYINPUT20), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n649), .B1(new_n651), .B2(new_n653), .ZN(new_n654));
  AND2_X1   g468(.A1(new_n654), .A2(new_n423), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n617), .A2(new_n621), .A3(new_n655), .ZN(new_n656));
  XOR2_X1   g470(.A(KEYINPUT35), .B(G107), .Z(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(G9));
  INV_X1    g472(.A(new_n443), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n659), .A2(KEYINPUT36), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n440), .B(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(new_n449), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n448), .A2(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n664), .A2(new_n616), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n425), .A2(new_n609), .A3(new_n665), .ZN(new_n666));
  XOR2_X1   g480(.A(KEYINPUT37), .B(G110), .Z(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G12));
  NAND2_X1  g482(.A1(new_n532), .A2(new_n542), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n304), .A2(new_n669), .A3(new_n663), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n670), .B1(new_n618), .B2(new_n620), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT104), .ZN(new_n672));
  INV_X1    g486(.A(G900), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n605), .B1(new_n606), .B2(new_n673), .ZN(new_n674));
  AOI211_X1 g488(.A(new_n674), .B(new_n649), .C1(new_n651), .C2(new_n653), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n672), .B1(new_n675), .B2(new_n423), .ZN(new_n676));
  INV_X1    g490(.A(new_n674), .ZN(new_n677));
  AND4_X1   g491(.A1(new_n672), .A2(new_n654), .A3(new_n423), .A4(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n671), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(KEYINPUT105), .B(G128), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(G30));
  XOR2_X1   g496(.A(new_n674), .B(KEYINPUT39), .Z(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n614), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(KEYINPUT40), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n600), .A2(new_n602), .ZN(new_n687));
  XNOR2_X1  g501(.A(KEYINPUT106), .B(KEYINPUT38), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n537), .A2(new_n499), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n517), .A2(new_n499), .A3(new_n504), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n190), .ZN(new_n692));
  OAI21_X1  g506(.A(G472), .B1(new_n690), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n532), .A2(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(new_n544), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n364), .A2(new_n423), .ZN(new_n697));
  NOR4_X1   g511(.A1(new_n695), .A2(new_n696), .A3(new_n663), .A4(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n686), .A2(new_n689), .A3(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(KEYINPUT107), .B(G143), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n699), .B(new_n700), .ZN(G45));
  INV_X1    g515(.A(KEYINPUT108), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n702), .B1(new_n639), .B2(new_n677), .ZN(new_n703));
  NOR4_X1   g517(.A1(new_n638), .A2(KEYINPUT108), .A3(new_n363), .A4(new_n674), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n671), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G146), .ZN(G48));
  NAND2_X1  g521(.A1(new_n299), .A2(new_n300), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(new_n190), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(G469), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n708), .A2(new_n296), .A3(new_n190), .ZN(new_n711));
  AND2_X1   g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(new_n191), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  AND2_X1   g529(.A1(new_n715), .A2(new_n543), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n716), .A2(new_n621), .A3(new_n639), .ZN(new_n717));
  XNOR2_X1  g531(.A(KEYINPUT41), .B(G113), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(KEYINPUT109), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n717), .B(new_n719), .ZN(G15));
  NAND3_X1  g534(.A1(new_n716), .A2(new_n621), .A3(new_n655), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G116), .ZN(G18));
  AOI21_X1  g536(.A(new_n664), .B1(new_n532), .B2(new_n542), .ZN(new_n723));
  INV_X1    g537(.A(new_n608), .ZN(new_n724));
  AND3_X1   g538(.A1(new_n723), .A2(new_n724), .A3(new_n424), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT110), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n618), .A2(new_n620), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n726), .B1(new_n727), .B2(new_n715), .ZN(new_n728));
  AOI211_X1 g542(.A(KEYINPUT110), .B(new_n714), .C1(new_n618), .C2(new_n620), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n725), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT111), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  OAI211_X1 g546(.A(KEYINPUT111), .B(new_n725), .C1(new_n728), .C2(new_n729), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G119), .ZN(G21));
  AOI21_X1  g549(.A(new_n697), .B1(new_n618), .B2(new_n620), .ZN(new_n736));
  OR2_X1    g550(.A1(new_n524), .A2(KEYINPUT112), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n524), .A2(KEYINPUT112), .ZN(new_n738));
  AND3_X1   g552(.A1(new_n615), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(new_n451), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(new_n741), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n736), .A2(new_n724), .A3(new_n715), .A4(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G122), .ZN(G24));
  AND2_X1   g558(.A1(new_n739), .A2(new_n663), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n624), .A2(new_n625), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n636), .A2(new_n637), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(new_n364), .ZN(new_n749));
  OAI21_X1  g563(.A(KEYINPUT108), .B1(new_n749), .B2(new_n674), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n639), .A2(new_n702), .A3(new_n677), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n745), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(new_n752), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n753), .B1(new_n728), .B2(new_n729), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G125), .ZN(G27));
  INV_X1    g569(.A(KEYINPUT42), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT113), .ZN(new_n757));
  AND3_X1   g571(.A1(new_n294), .A2(new_n711), .A3(new_n757), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n757), .B1(new_n294), .B2(new_n711), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n713), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(new_n600), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n580), .A2(new_n599), .A3(new_n545), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n761), .A2(new_n544), .A3(new_n762), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n542), .A2(new_n527), .A3(new_n526), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n764), .A2(new_n740), .ZN(new_n765));
  NOR3_X1   g579(.A1(new_n760), .A2(new_n763), .A3(new_n765), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n756), .B1(new_n766), .B2(new_n705), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n750), .A2(new_n756), .A3(new_n751), .ZN(new_n768));
  INV_X1    g582(.A(new_n759), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n294), .A2(new_n711), .A3(new_n757), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n191), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NOR3_X1   g585(.A1(new_n600), .A2(new_n602), .A3(new_n696), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n771), .A2(new_n543), .A3(new_n772), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n768), .A2(new_n773), .ZN(new_n774));
  OAI21_X1  g588(.A(KEYINPUT114), .B1(new_n767), .B2(new_n774), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n771), .A2(new_n740), .A3(new_n772), .A4(new_n764), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n750), .A2(new_n751), .ZN(new_n777));
  OAI21_X1  g591(.A(KEYINPUT42), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n760), .A2(new_n763), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n705), .A2(new_n779), .A3(new_n756), .A4(new_n543), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT114), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n778), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  AND2_X1   g596(.A1(new_n775), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G131), .ZN(G33));
  NAND4_X1  g598(.A1(new_n679), .A2(new_n772), .A3(new_n771), .A4(new_n543), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(G134), .ZN(G36));
  NOR2_X1   g600(.A1(new_n638), .A2(new_n364), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(KEYINPUT43), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n788), .A2(new_n616), .A3(new_n663), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT44), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n763), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n293), .A2(KEYINPUT45), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n792), .A2(new_n296), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n293), .A2(KEYINPUT45), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(G469), .A2(G902), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT46), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(new_n711), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n797), .A2(new_n798), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n713), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n802), .A2(new_n684), .ZN(new_n803));
  OAI211_X1 g617(.A(new_n791), .B(new_n803), .C1(new_n790), .C2(new_n789), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(G137), .ZN(G39));
  XNOR2_X1  g619(.A(new_n802), .B(KEYINPUT47), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n772), .A2(new_n542), .A3(new_n532), .A4(new_n451), .ZN(new_n807));
  NOR3_X1   g621(.A1(new_n806), .A2(new_n777), .A3(new_n807), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(new_n308), .ZN(G42));
  NOR3_X1   g623(.A1(new_n689), .A2(new_n544), .A3(new_n714), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT116), .ZN(new_n811));
  OR2_X1    g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  AND2_X1   g626(.A1(new_n788), .A2(new_n605), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n813), .A2(new_n742), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n810), .A2(new_n811), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n812), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT50), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n816), .B(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(new_n712), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n806), .B1(new_n713), .B2(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n820), .A2(new_n772), .A3(new_n814), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n818), .A2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(new_n822), .ZN(new_n823));
  AND3_X1   g637(.A1(new_n813), .A2(new_n715), .A3(new_n772), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n695), .A2(new_n740), .A3(new_n605), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n825), .A2(new_n714), .A3(new_n763), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n748), .A2(new_n364), .ZN(new_n827));
  AOI22_X1  g641(.A1(new_n824), .A2(new_n745), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  AOI21_X1  g642(.A(KEYINPUT51), .B1(new_n823), .B2(new_n828), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n765), .B1(KEYINPUT118), .B2(KEYINPUT48), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n824), .A2(new_n830), .ZN(new_n831));
  NOR2_X1   g645(.A1(KEYINPUT118), .A2(KEYINPUT48), .ZN(new_n832));
  OR2_X1    g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n831), .A2(new_n832), .ZN(new_n834));
  AOI211_X1 g648(.A(new_n604), .B(G953), .C1(new_n826), .C2(new_n639), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n833), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  OR2_X1    g650(.A1(new_n728), .A2(new_n729), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n836), .B1(new_n837), .B2(new_n814), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT117), .ZN(new_n839));
  OR2_X1    g653(.A1(new_n828), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n828), .A2(new_n839), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n840), .A2(KEYINPUT51), .A3(new_n841), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n838), .B1(new_n822), .B2(new_n842), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n829), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n664), .A2(new_n677), .ZN(new_n845));
  NOR3_X1   g659(.A1(new_n695), .A2(new_n760), .A3(new_n845), .ZN(new_n846));
  AOI22_X1  g660(.A1(new_n671), .A2(new_n705), .B1(new_n736), .B2(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n754), .A2(new_n680), .A3(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT52), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n754), .A2(new_n847), .A3(KEYINPUT52), .A4(new_n680), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(new_n779), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n854), .A2(new_n752), .ZN(new_n855));
  INV_X1    g669(.A(new_n675), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n856), .A2(new_n423), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n723), .A2(new_n857), .A3(new_n304), .A4(new_n772), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n785), .A2(new_n858), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n855), .A2(new_n859), .ZN(new_n860));
  AND3_X1   g674(.A1(new_n775), .A2(new_n782), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n423), .A2(new_n363), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n749), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n617), .A2(new_n609), .A3(new_n863), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n743), .A2(new_n864), .A3(new_n610), .A4(new_n666), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n717), .A2(new_n721), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n861), .A2(new_n734), .A3(new_n867), .ZN(new_n868));
  OAI21_X1  g682(.A(KEYINPUT53), .B1(new_n853), .B2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT115), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n852), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n850), .A2(KEYINPUT115), .A3(new_n851), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  AND3_X1   g687(.A1(new_n861), .A2(new_n734), .A3(new_n867), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT53), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  OAI211_X1 g690(.A(new_n869), .B(KEYINPUT54), .C1(new_n873), .C2(new_n876), .ZN(new_n877));
  AND3_X1   g691(.A1(new_n850), .A2(KEYINPUT115), .A3(new_n851), .ZN(new_n878));
  AOI21_X1  g692(.A(KEYINPUT115), .B1(new_n850), .B2(new_n851), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n778), .A2(new_n780), .A3(KEYINPUT53), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n880), .A2(new_n855), .A3(new_n859), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n734), .A2(new_n867), .A3(new_n881), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n878), .A2(new_n879), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g697(.A(KEYINPUT53), .B1(new_n874), .B2(new_n852), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT54), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n844), .A2(new_n877), .A3(new_n887), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n888), .B1(G952), .B2(G953), .ZN(new_n889));
  OR2_X1    g703(.A1(new_n819), .A2(KEYINPUT49), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n819), .A2(KEYINPUT49), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n451), .A2(new_n696), .A3(new_n191), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n890), .A2(new_n787), .A3(new_n891), .A4(new_n892), .ZN(new_n893));
  OR2_X1    g707(.A1(new_n893), .A2(new_n694), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n889), .B1(new_n689), .B2(new_n894), .ZN(G75));
  NOR2_X1   g709(.A1(new_n284), .A2(G952), .ZN(new_n896));
  INV_X1    g710(.A(new_n896), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n885), .A2(new_n190), .ZN(new_n898));
  AOI21_X1  g712(.A(KEYINPUT56), .B1(new_n898), .B2(G210), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n573), .B(new_n578), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n900), .B(KEYINPUT55), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n897), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n902), .B1(new_n901), .B2(new_n899), .ZN(G51));
  INV_X1    g717(.A(new_n882), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n871), .A2(new_n872), .A3(new_n904), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n875), .B1(new_n853), .B2(new_n868), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(KEYINPUT54), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n887), .A2(KEYINPUT120), .A3(new_n908), .ZN(new_n909));
  OR3_X1    g723(.A1(new_n885), .A2(KEYINPUT120), .A3(new_n886), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n796), .B(KEYINPUT119), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n911), .B(KEYINPUT57), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n909), .A2(new_n910), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(new_n708), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n898), .A2(new_n794), .A3(new_n793), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n896), .B1(new_n914), .B2(new_n915), .ZN(G54));
  NAND3_X1  g730(.A1(new_n898), .A2(KEYINPUT58), .A3(G475), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n352), .A2(new_n353), .ZN(new_n918));
  AND2_X1   g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n917), .A2(new_n918), .ZN(new_n920));
  NOR3_X1   g734(.A1(new_n919), .A2(new_n920), .A3(new_n896), .ZN(G60));
  NAND2_X1  g735(.A1(G478), .A2(G902), .ZN(new_n922));
  XOR2_X1   g736(.A(new_n922), .B(KEYINPUT59), .Z(new_n923));
  AOI21_X1  g737(.A(new_n923), .B1(new_n887), .B2(new_n877), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n897), .B1(new_n924), .B2(new_n636), .ZN(new_n925));
  INV_X1    g739(.A(new_n636), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n926), .A2(new_n923), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n909), .A2(new_n910), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(KEYINPUT121), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT121), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n909), .A2(new_n910), .A3(new_n930), .A4(new_n927), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n925), .B1(new_n929), .B2(new_n931), .ZN(G63));
  NAND2_X1  g746(.A1(G217), .A2(G902), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(KEYINPUT60), .ZN(new_n934));
  INV_X1    g748(.A(new_n934), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n935), .B1(new_n883), .B2(new_n884), .ZN(new_n936));
  INV_X1    g750(.A(new_n444), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  OAI211_X1 g752(.A(new_n661), .B(new_n935), .C1(new_n883), .C2(new_n884), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n938), .A2(KEYINPUT61), .A3(new_n897), .A4(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(KEYINPUT122), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT122), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n907), .A2(new_n942), .A3(new_n661), .A4(new_n935), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n941), .A2(new_n938), .A3(new_n897), .A4(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT123), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT61), .ZN(new_n946));
  AND3_X1   g760(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n945), .B1(new_n944), .B2(new_n946), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n940), .B1(new_n947), .B2(new_n948), .ZN(G66));
  INV_X1    g763(.A(G224), .ZN(new_n950));
  OAI21_X1  g764(.A(G953), .B1(new_n607), .B2(new_n950), .ZN(new_n951));
  AND2_X1   g765(.A1(new_n734), .A2(new_n867), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n951), .B1(new_n952), .B2(G953), .ZN(new_n953));
  INV_X1    g767(.A(new_n573), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n954), .B1(G898), .B2(new_n284), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n953), .B(new_n955), .ZN(G69));
  AND3_X1   g770(.A1(new_n754), .A2(new_n680), .A3(new_n706), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n957), .A2(new_n804), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n958), .B(KEYINPUT125), .Z(new_n959));
  INV_X1    g773(.A(new_n785), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n808), .A2(new_n960), .ZN(new_n961));
  NAND4_X1  g775(.A1(new_n803), .A2(new_n740), .A3(new_n736), .A4(new_n764), .ZN(new_n962));
  AND3_X1   g776(.A1(new_n961), .A2(new_n783), .A3(new_n962), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n959), .A2(new_n284), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n315), .A2(new_n316), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n508), .B(new_n965), .Z(new_n966));
  OAI211_X1 g780(.A(new_n964), .B(new_n966), .C1(new_n673), .C2(new_n284), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n957), .A2(new_n699), .ZN(new_n968));
  OR2_X1    g782(.A1(new_n968), .A2(KEYINPUT62), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n968), .A2(KEYINPUT62), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n685), .A2(new_n543), .A3(new_n772), .A4(new_n863), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n804), .A2(new_n971), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n808), .A2(new_n972), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n969), .A2(new_n970), .A3(new_n973), .ZN(new_n974));
  OR2_X1    g788(.A1(new_n974), .A2(KEYINPUT124), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n974), .A2(KEYINPUT124), .ZN(new_n976));
  AOI21_X1  g790(.A(G953), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n967), .B1(new_n977), .B2(new_n966), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n284), .B1(G227), .B2(G900), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n978), .B(new_n979), .ZN(G72));
  NAND3_X1  g794(.A1(new_n959), .A2(new_n952), .A3(new_n963), .ZN(new_n981));
  XNOR2_X1  g795(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n523), .A2(new_n190), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n982), .B(new_n983), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n984), .B(KEYINPUT127), .Z(new_n985));
  NAND2_X1  g799(.A1(new_n981), .A2(new_n985), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n986), .A2(new_n499), .A3(new_n537), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n869), .B1(new_n873), .B2(new_n876), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n538), .A2(new_n536), .A3(new_n514), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n989), .A2(new_n984), .ZN(new_n990));
  OAI211_X1 g804(.A(new_n987), .B(new_n897), .C1(new_n988), .C2(new_n990), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n975), .A2(new_n952), .A3(new_n976), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n992), .A2(new_n985), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n991), .B1(new_n690), .B2(new_n993), .ZN(G57));
endmodule


