//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 0 0 1 1 0 1 0 1 0 1 0 1 0 0 1 0 1 1 1 0 1 0 0 1 1 1 1 1 1 0 1 1 1 1 0 1 1 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:56 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n683, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n730, new_n731,
    new_n732, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n901, new_n902, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  XOR2_X1   g001(.A(new_n187), .B(KEYINPUT79), .Z(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  OAI21_X1  g003(.A(G210), .B1(G237), .B2(G902), .ZN(new_n190));
  INV_X1    g004(.A(G119), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G116), .ZN(new_n192));
  INV_X1    g006(.A(G116), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G119), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n192), .A2(new_n194), .A3(KEYINPUT5), .ZN(new_n195));
  OAI211_X1 g009(.A(new_n195), .B(G113), .C1(KEYINPUT5), .C2(new_n192), .ZN(new_n196));
  INV_X1    g010(.A(G113), .ZN(new_n197));
  AND2_X1   g011(.A1(new_n197), .A2(KEYINPUT2), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n197), .A2(KEYINPUT2), .ZN(new_n199));
  OAI211_X1 g013(.A(new_n192), .B(new_n194), .C1(new_n198), .C2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G104), .ZN(new_n201));
  OAI21_X1  g015(.A(KEYINPUT3), .B1(new_n201), .B2(G107), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT3), .ZN(new_n203));
  INV_X1    g017(.A(G107), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n203), .A2(new_n204), .A3(G104), .ZN(new_n205));
  INV_X1    g019(.A(G101), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n201), .A2(G107), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n202), .A2(new_n205), .A3(new_n206), .A4(new_n207), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n201), .A2(G107), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n204), .A2(G104), .ZN(new_n210));
  OAI21_X1  g024(.A(G101), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n196), .A2(new_n200), .A3(new_n208), .A4(new_n211), .ZN(new_n212));
  XNOR2_X1  g026(.A(G110), .B(G122), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n202), .A2(new_n205), .A3(new_n207), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G101), .ZN(new_n215));
  AND3_X1   g029(.A1(new_n215), .A2(KEYINPUT4), .A3(new_n208), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n192), .A2(new_n194), .ZN(new_n217));
  XNOR2_X1  g031(.A(KEYINPUT2), .B(G113), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n200), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT4), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n214), .A2(new_n221), .A3(G101), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  OAI211_X1 g037(.A(new_n212), .B(new_n213), .C1(new_n216), .C2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(KEYINPUT6), .ZN(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n212), .B1(new_n216), .B2(new_n223), .ZN(new_n227));
  XNOR2_X1  g041(.A(new_n213), .B(KEYINPUT80), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(KEYINPUT81), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT81), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n227), .A2(new_n231), .A3(new_n228), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n226), .A2(new_n230), .A3(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT6), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n227), .A2(new_n234), .A3(new_n228), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(KEYINPUT82), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT82), .ZN(new_n237));
  NAND4_X1  g051(.A1(new_n227), .A2(new_n237), .A3(new_n234), .A4(new_n228), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(G146), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G143), .ZN(new_n241));
  INV_X1    g055(.A(G143), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G146), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n241), .A2(new_n243), .A3(KEYINPUT0), .A4(G128), .ZN(new_n244));
  XNOR2_X1  g058(.A(G143), .B(G146), .ZN(new_n245));
  XNOR2_X1  g059(.A(KEYINPUT0), .B(G128), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n244), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(G125), .ZN(new_n248));
  XNOR2_X1  g062(.A(KEYINPUT66), .B(G128), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT1), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n250), .B1(G143), .B2(new_n240), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n242), .A2(G146), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n240), .A2(G143), .ZN(new_n253));
  OAI22_X1  g067(.A1(new_n249), .A2(new_n251), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(G128), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n255), .A2(KEYINPUT1), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n256), .A2(new_n241), .A3(new_n243), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n254), .A2(new_n257), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n248), .B1(new_n258), .B2(G125), .ZN(new_n259));
  INV_X1    g073(.A(G224), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n260), .A2(G953), .ZN(new_n261));
  XNOR2_X1  g075(.A(new_n259), .B(new_n261), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n233), .A2(new_n239), .A3(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT83), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n233), .A2(new_n239), .A3(new_n262), .A4(KEYINPUT83), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  OAI21_X1  g081(.A(KEYINPUT7), .B1(new_n260), .B2(G953), .ZN(new_n268));
  XOR2_X1   g082(.A(new_n259), .B(new_n268), .Z(new_n269));
  NAND2_X1  g083(.A1(new_n196), .A2(new_n200), .ZN(new_n270));
  AND2_X1   g084(.A1(new_n208), .A2(new_n211), .ZN(new_n271));
  XNOR2_X1  g085(.A(new_n270), .B(new_n271), .ZN(new_n272));
  XOR2_X1   g086(.A(new_n213), .B(KEYINPUT8), .Z(new_n273));
  OAI211_X1 g087(.A(new_n269), .B(new_n224), .C1(new_n272), .C2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(G902), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n190), .B1(new_n267), .B2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n190), .ZN(new_n279));
  AOI211_X1 g093(.A(new_n279), .B(new_n276), .C1(new_n265), .C2(new_n266), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n189), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT84), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  OAI211_X1 g097(.A(KEYINPUT84), .B(new_n189), .C1(new_n278), .C2(new_n280), .ZN(new_n284));
  XNOR2_X1  g098(.A(KEYINPUT9), .B(G234), .ZN(new_n285));
  OAI21_X1  g099(.A(G221), .B1(new_n285), .B2(G902), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(G469), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n288), .A2(new_n275), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT10), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n257), .A2(KEYINPUT76), .ZN(new_n291));
  OAI22_X1  g105(.A1(new_n251), .A2(new_n255), .B1(new_n252), .B2(new_n253), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT76), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n245), .A2(new_n293), .A3(new_n256), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n291), .A2(new_n292), .A3(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT77), .ZN(new_n296));
  AND3_X1   g110(.A1(new_n295), .A2(new_n271), .A3(new_n296), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n296), .B1(new_n295), .B2(new_n271), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n290), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(new_n247), .ZN(new_n300));
  AND2_X1   g114(.A1(new_n300), .A2(new_n222), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n215), .A2(KEYINPUT4), .A3(new_n208), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n290), .B1(new_n254), .B2(new_n257), .ZN(new_n303));
  AOI22_X1  g117(.A1(new_n301), .A2(new_n302), .B1(new_n271), .B2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(G134), .ZN(new_n305));
  OAI21_X1  g119(.A(KEYINPUT11), .B1(new_n305), .B2(G137), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT11), .ZN(new_n307));
  INV_X1    g121(.A(G137), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n307), .A2(new_n308), .A3(G134), .ZN(new_n309));
  AND2_X1   g123(.A1(new_n306), .A2(new_n309), .ZN(new_n310));
  OAI21_X1  g124(.A(KEYINPUT64), .B1(new_n308), .B2(G134), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT64), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n312), .A2(new_n305), .A3(G137), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  OAI21_X1  g128(.A(G131), .B1(new_n310), .B2(new_n314), .ZN(new_n315));
  AND2_X1   g129(.A1(new_n311), .A2(new_n313), .ZN(new_n316));
  INV_X1    g130(.A(G131), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n306), .A2(new_n309), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n316), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n315), .A2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n299), .A2(new_n304), .A3(new_n321), .ZN(new_n322));
  OAI22_X1  g136(.A1(new_n297), .A2(new_n298), .B1(new_n258), .B2(new_n271), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n323), .A2(KEYINPUT12), .A3(new_n320), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  AOI21_X1  g139(.A(KEYINPUT12), .B1(new_n323), .B2(new_n320), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n322), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  XNOR2_X1  g141(.A(G110), .B(G140), .ZN(new_n328));
  XNOR2_X1  g142(.A(new_n328), .B(KEYINPUT75), .ZN(new_n329));
  INV_X1    g143(.A(G953), .ZN(new_n330));
  AND2_X1   g144(.A1(new_n330), .A2(G227), .ZN(new_n331));
  XNOR2_X1  g145(.A(new_n329), .B(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT78), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n295), .A2(new_n271), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(KEYINPUT77), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n295), .A2(new_n271), .A3(new_n296), .ZN(new_n337));
  AOI21_X1  g151(.A(KEYINPUT10), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n303), .A2(new_n271), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n300), .A2(new_n222), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n339), .B1(new_n340), .B2(new_n216), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n334), .B1(new_n338), .B2(new_n341), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n299), .A2(new_n304), .A3(KEYINPUT78), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n342), .A2(new_n320), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n322), .A2(new_n332), .ZN(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  AOI22_X1  g160(.A1(new_n327), .A2(new_n333), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n289), .B1(new_n347), .B2(G469), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n332), .B1(new_n344), .B2(new_n322), .ZN(new_n349));
  INV_X1    g163(.A(new_n326), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n345), .B1(new_n350), .B2(new_n324), .ZN(new_n351));
  OAI211_X1 g165(.A(new_n288), .B(new_n275), .C1(new_n349), .C2(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n287), .B1(new_n348), .B2(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n283), .A2(new_n284), .A3(new_n353), .ZN(new_n354));
  XNOR2_X1  g168(.A(KEYINPUT85), .B(KEYINPUT20), .ZN(new_n355));
  INV_X1    g169(.A(G237), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n356), .A2(new_n330), .A3(G214), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(new_n242), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n356), .A2(new_n330), .A3(G143), .A4(G214), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT18), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n361), .B1(new_n362), .B2(new_n317), .ZN(new_n363));
  INV_X1    g177(.A(G140), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(G125), .ZN(new_n365));
  INV_X1    g179(.A(G125), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(G140), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  XNOR2_X1  g182(.A(new_n368), .B(G146), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n360), .A2(KEYINPUT18), .A3(G131), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n363), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  XNOR2_X1  g185(.A(G113), .B(G122), .ZN(new_n372));
  XNOR2_X1  g186(.A(new_n372), .B(new_n201), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n360), .A2(G131), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(KEYINPUT17), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT71), .ZN(new_n377));
  NAND4_X1  g191(.A1(new_n365), .A2(new_n367), .A3(new_n377), .A4(KEYINPUT16), .ZN(new_n378));
  AND3_X1   g192(.A1(new_n365), .A2(new_n367), .A3(KEYINPUT16), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT16), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n380), .A2(new_n364), .A3(G125), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(KEYINPUT71), .ZN(new_n382));
  OAI211_X1 g196(.A(new_n240), .B(new_n378), .C1(new_n379), .C2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT72), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  OAI211_X1 g199(.A(KEYINPUT71), .B(new_n381), .C1(new_n368), .C2(new_n380), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n240), .B1(new_n386), .B2(new_n378), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  AOI211_X1 g202(.A(new_n384), .B(new_n240), .C1(new_n386), .C2(new_n378), .ZN(new_n389));
  OAI211_X1 g203(.A(KEYINPUT88), .B(new_n376), .C1(new_n388), .C2(new_n389), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n361), .A2(KEYINPUT86), .A3(new_n317), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT86), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n392), .B1(new_n360), .B2(G131), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n391), .A2(new_n374), .A3(new_n393), .ZN(new_n394));
  OR2_X1    g208(.A1(new_n394), .A2(KEYINPUT17), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n390), .A2(new_n395), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n378), .B1(new_n379), .B2(new_n382), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(G146), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n398), .A2(new_n384), .A3(new_n383), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n385), .A2(new_n387), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(KEYINPUT88), .B1(new_n401), .B2(new_n376), .ZN(new_n402));
  OAI211_X1 g216(.A(new_n371), .B(new_n373), .C1(new_n396), .C2(new_n402), .ZN(new_n403));
  XOR2_X1   g217(.A(new_n368), .B(KEYINPUT19), .Z(new_n404));
  AOI21_X1  g218(.A(new_n387), .B1(new_n240), .B2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT87), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n405), .B1(new_n406), .B2(new_n394), .ZN(new_n407));
  AND2_X1   g221(.A1(new_n394), .A2(new_n406), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n371), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(new_n373), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n403), .A2(new_n411), .ZN(new_n412));
  NOR2_X1   g226(.A1(G475), .A2(G902), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n355), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n413), .ZN(new_n415));
  AOI211_X1 g229(.A(KEYINPUT20), .B(new_n415), .C1(new_n403), .C2(new_n411), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n371), .B1(new_n396), .B2(new_n402), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(new_n410), .ZN(new_n418));
  AOI21_X1  g232(.A(G902), .B1(new_n418), .B2(new_n403), .ZN(new_n419));
  INV_X1    g233(.A(G475), .ZN(new_n420));
  OAI22_X1  g234(.A1(new_n414), .A2(new_n416), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(KEYINPUT89), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT89), .ZN(new_n423));
  OAI221_X1 g237(.A(new_n423), .B1(new_n419), .B2(new_n420), .C1(new_n414), .C2(new_n416), .ZN(new_n424));
  OR2_X1    g238(.A1(new_n193), .A2(G122), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n204), .B1(new_n425), .B2(KEYINPUT14), .ZN(new_n426));
  XOR2_X1   g240(.A(G116), .B(G122), .Z(new_n427));
  XNOR2_X1  g241(.A(new_n426), .B(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n249), .A2(G143), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n242), .A2(G128), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n429), .A2(new_n305), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n429), .A2(new_n430), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(G134), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n428), .B1(new_n431), .B2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT13), .ZN(new_n435));
  AOI22_X1  g249(.A1(new_n249), .A2(G143), .B1(new_n435), .B2(new_n430), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT90), .ZN(new_n437));
  OAI211_X1 g251(.A(new_n436), .B(new_n437), .C1(new_n435), .C2(new_n430), .ZN(new_n438));
  OAI211_X1 g252(.A(new_n438), .B(G134), .C1(new_n437), .C2(new_n436), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n427), .B(G107), .ZN(new_n440));
  AND2_X1   g254(.A1(new_n440), .A2(new_n431), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n434), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(G217), .ZN(new_n443));
  NOR3_X1   g257(.A1(new_n285), .A2(new_n443), .A3(G953), .ZN(new_n444));
  OR2_X1    g258(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n442), .A2(new_n444), .ZN(new_n446));
  AOI21_X1  g260(.A(G902), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(G478), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n448), .A2(KEYINPUT15), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  AND2_X1   g264(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n447), .A2(new_n450), .ZN(new_n452));
  AOI211_X1 g266(.A(new_n275), .B(new_n330), .C1(G234), .C2(G237), .ZN(new_n453));
  XNOR2_X1  g267(.A(KEYINPUT21), .B(G898), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  OR2_X1    g269(.A1(KEYINPUT91), .A2(G952), .ZN(new_n456));
  NAND2_X1  g270(.A1(KEYINPUT91), .A2(G952), .ZN(new_n457));
  AOI21_X1  g271(.A(G953), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(G234), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n458), .B1(new_n459), .B2(new_n356), .ZN(new_n460));
  AND2_X1   g274(.A1(new_n455), .A2(new_n460), .ZN(new_n461));
  NOR3_X1   g275(.A1(new_n451), .A2(new_n452), .A3(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n422), .A2(new_n424), .A3(new_n462), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n354), .A2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(new_n368), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n387), .B1(new_n240), .B2(new_n465), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n255), .A2(G119), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n467), .B1(new_n249), .B2(G119), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  XNOR2_X1  g283(.A(KEYINPUT24), .B(G110), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n469), .A2(KEYINPUT73), .A3(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n249), .A2(KEYINPUT23), .A3(G119), .ZN(new_n472));
  AOI21_X1  g286(.A(KEYINPUT23), .B1(new_n255), .B2(G119), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n473), .A2(new_n467), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n471), .B1(G110), .B2(new_n475), .ZN(new_n476));
  AOI21_X1  g290(.A(KEYINPUT73), .B1(new_n469), .B2(new_n470), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n466), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(new_n470), .ZN(new_n479));
  AOI22_X1  g293(.A1(new_n475), .A2(G110), .B1(new_n468), .B2(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n399), .A2(new_n400), .A3(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n330), .A2(G221), .A3(G234), .ZN(new_n482));
  XNOR2_X1  g296(.A(new_n482), .B(KEYINPUT74), .ZN(new_n483));
  XNOR2_X1  g297(.A(KEYINPUT22), .B(G137), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n483), .B(new_n484), .ZN(new_n485));
  AND3_X1   g299(.A1(new_n478), .A2(new_n481), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n485), .B1(new_n478), .B2(new_n481), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n275), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT25), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n488), .B(new_n489), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n443), .B1(G234), .B2(new_n275), .ZN(new_n491));
  OR2_X1    g305(.A1(new_n486), .A2(new_n487), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n491), .A2(G902), .ZN(new_n493));
  AOI22_X1  g307(.A1(new_n490), .A2(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  NOR2_X1   g309(.A1(G472), .A2(G902), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  OAI21_X1  g311(.A(KEYINPUT65), .B1(new_n308), .B2(G134), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n498), .B1(new_n305), .B2(G137), .ZN(new_n499));
  NOR3_X1   g313(.A1(new_n308), .A2(KEYINPUT65), .A3(G134), .ZN(new_n500));
  OAI21_X1  g314(.A(G131), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n258), .A2(new_n501), .A3(new_n319), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  NOR3_X1   g317(.A1(new_n310), .A2(G131), .A3(new_n314), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n317), .B1(new_n316), .B2(new_n318), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n300), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(KEYINPUT67), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT67), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n320), .A2(new_n508), .A3(new_n300), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n503), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n220), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n356), .A2(new_n330), .A3(G210), .ZN(new_n513));
  XOR2_X1   g327(.A(new_n513), .B(KEYINPUT27), .Z(new_n514));
  XNOR2_X1  g328(.A(KEYINPUT26), .B(G101), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n514), .B(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT30), .ZN(new_n518));
  AND3_X1   g332(.A1(new_n506), .A2(new_n502), .A3(new_n518), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n508), .B1(new_n320), .B2(new_n300), .ZN(new_n520));
  AOI211_X1 g334(.A(KEYINPUT67), .B(new_n247), .C1(new_n315), .C2(new_n319), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n502), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n519), .B1(new_n522), .B2(KEYINPUT30), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n512), .B(new_n517), .C1(new_n523), .C2(new_n511), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(KEYINPUT68), .ZN(new_n525));
  INV_X1    g339(.A(new_n519), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n526), .B1(new_n510), .B2(new_n518), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(new_n220), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT68), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n528), .A2(new_n529), .A3(new_n512), .A4(new_n517), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n525), .A2(new_n530), .A3(KEYINPUT31), .ZN(new_n531));
  AND2_X1   g345(.A1(new_n506), .A2(new_n502), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n532), .A2(new_n511), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT28), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n532), .A2(new_n511), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n510), .A2(KEYINPUT28), .A3(new_n511), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n517), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n524), .ZN(new_n539));
  XOR2_X1   g353(.A(KEYINPUT69), .B(KEYINPUT31), .Z(new_n540));
  AOI21_X1  g354(.A(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n497), .B1(new_n531), .B2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT32), .ZN(new_n543));
  XNOR2_X1  g357(.A(new_n542), .B(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n522), .A2(new_n220), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n534), .B1(new_n512), .B2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT70), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n535), .A2(new_n534), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(KEYINPUT70), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n548), .B1(new_n546), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n551), .A2(KEYINPUT29), .A3(new_n517), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n528), .A2(new_n512), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(new_n516), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT29), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n536), .A2(new_n517), .A3(new_n537), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n552), .A2(new_n275), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(G472), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n495), .B1(new_n544), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n464), .A2(new_n560), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n561), .B(G101), .ZN(G3));
  AND2_X1   g376(.A1(new_n353), .A2(new_n494), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n531), .A2(new_n541), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(new_n275), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n542), .B1(new_n565), .B2(G472), .ZN(new_n566));
  AND2_X1   g380(.A1(new_n563), .A2(new_n566), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n567), .B(KEYINPUT92), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n445), .A2(new_n446), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT93), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n445), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n569), .A2(new_n571), .A3(KEYINPUT33), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT33), .ZN(new_n573));
  OAI211_X1 g387(.A(new_n445), .B(new_n446), .C1(new_n570), .C2(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n572), .A2(G478), .A3(new_n574), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n448), .A2(new_n275), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n576), .B1(new_n447), .B2(new_n448), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n578), .B1(new_n422), .B2(new_n424), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n281), .A2(new_n461), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n568), .A2(new_n581), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n582), .B(KEYINPUT94), .ZN(new_n583));
  XOR2_X1   g397(.A(KEYINPUT34), .B(G104), .Z(new_n584));
  XNOR2_X1  g398(.A(new_n583), .B(new_n584), .ZN(G6));
  NOR2_X1   g399(.A1(new_n451), .A2(new_n452), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n394), .A2(KEYINPUT17), .ZN(new_n588));
  AOI22_X1  g402(.A1(new_n399), .A2(new_n400), .B1(KEYINPUT17), .B2(new_n375), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n588), .B1(new_n589), .B2(KEYINPUT88), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n401), .A2(new_n376), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT88), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n373), .B1(new_n594), .B2(new_n371), .ZN(new_n595));
  INV_X1    g409(.A(new_n403), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n275), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n355), .ZN(new_n598));
  AOI211_X1 g412(.A(new_n415), .B(new_n598), .C1(new_n403), .C2(new_n411), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT95), .ZN(new_n600));
  AOI22_X1  g414(.A1(G475), .A2(new_n597), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n412), .A2(new_n413), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(new_n598), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n412), .A2(new_n413), .A3(new_n355), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n603), .A2(KEYINPUT95), .A3(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n587), .A2(new_n601), .A3(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT96), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n607), .A2(new_n580), .A3(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n228), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n302), .A2(new_n220), .A3(new_n222), .ZN(new_n611));
  AOI211_X1 g425(.A(KEYINPUT81), .B(new_n610), .C1(new_n611), .C2(new_n212), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n612), .A2(new_n225), .ZN(new_n613));
  AOI22_X1  g427(.A1(new_n613), .A2(new_n230), .B1(new_n236), .B2(new_n238), .ZN(new_n614));
  AOI21_X1  g428(.A(KEYINPUT83), .B1(new_n614), .B2(new_n262), .ZN(new_n615));
  INV_X1    g429(.A(new_n266), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n277), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(new_n279), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n267), .A2(new_n190), .A3(new_n277), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n461), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n620), .A2(new_n621), .A3(new_n189), .ZN(new_n622));
  OAI21_X1  g436(.A(KEYINPUT96), .B1(new_n622), .B2(new_n606), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n568), .B1(new_n609), .B2(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(KEYINPUT35), .B(G107), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n624), .B(new_n625), .ZN(G9));
  NAND2_X1  g440(.A1(new_n490), .A2(new_n491), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n478), .A2(new_n481), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n485), .A2(KEYINPUT36), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(new_n493), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n627), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n566), .A2(new_n632), .ZN(new_n633));
  NOR3_X1   g447(.A1(new_n354), .A2(new_n633), .A3(new_n463), .ZN(new_n634));
  XNOR2_X1  g448(.A(KEYINPUT37), .B(G110), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G12));
  NOR2_X1   g450(.A1(new_n542), .A2(new_n543), .ZN(new_n637));
  AOI211_X1 g451(.A(KEYINPUT32), .B(new_n497), .C1(new_n531), .C2(new_n541), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n559), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n188), .B1(new_n618), .B2(new_n619), .ZN(new_n640));
  AND4_X1   g454(.A1(new_n639), .A2(new_n640), .A3(new_n353), .A4(new_n632), .ZN(new_n641));
  INV_X1    g455(.A(new_n453), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n460), .B1(new_n642), .B2(G900), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(KEYINPUT97), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n587), .A2(new_n601), .A3(new_n605), .A4(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n641), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(G128), .ZN(G30));
  NAND2_X1  g463(.A1(new_n422), .A2(new_n424), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NOR4_X1   g465(.A1(new_n651), .A2(new_n586), .A3(new_n188), .A4(new_n632), .ZN(new_n652));
  XOR2_X1   g466(.A(new_n644), .B(KEYINPUT39), .Z(new_n653));
  NAND2_X1  g467(.A1(new_n353), .A2(new_n653), .ZN(new_n654));
  XOR2_X1   g468(.A(new_n654), .B(KEYINPUT40), .Z(new_n655));
  INV_X1    g469(.A(G472), .ZN(new_n656));
  AND2_X1   g470(.A1(new_n525), .A2(new_n530), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n512), .A2(new_n545), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(new_n516), .ZN(new_n659));
  AOI21_X1  g473(.A(G902), .B1(new_n657), .B2(new_n659), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n544), .B1(new_n656), .B2(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(KEYINPUT98), .B(KEYINPUT38), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n620), .B(new_n662), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n652), .A2(new_n655), .A3(new_n661), .A4(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(G143), .ZN(G45));
  INV_X1    g479(.A(new_n578), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n650), .A2(new_n666), .A3(new_n645), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT99), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n579), .A2(KEYINPUT99), .A3(new_n645), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n641), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G146), .ZN(G48));
  NAND2_X1  g486(.A1(new_n352), .A2(new_n286), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n275), .B1(new_n349), .B2(new_n351), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT100), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n288), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  OAI211_X1 g490(.A(KEYINPUT100), .B(new_n275), .C1(new_n349), .C2(new_n351), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n673), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n639), .A2(new_n494), .A3(new_n678), .ZN(new_n679));
  OR2_X1    g493(.A1(new_n679), .A2(new_n581), .ZN(new_n680));
  XNOR2_X1  g494(.A(KEYINPUT41), .B(G113), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(G15));
  AOI21_X1  g496(.A(new_n679), .B1(new_n609), .B2(new_n623), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(new_n193), .ZN(G18));
  NAND2_X1  g498(.A1(new_n674), .A2(new_n675), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n685), .A2(G469), .A3(new_n677), .ZN(new_n686));
  INV_X1    g500(.A(new_n673), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT101), .ZN(new_n689));
  NOR3_X1   g503(.A1(new_n688), .A2(new_n281), .A3(new_n689), .ZN(new_n690));
  AOI21_X1  g504(.A(KEYINPUT101), .B1(new_n640), .B2(new_n678), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  AND3_X1   g506(.A1(new_n422), .A2(new_n424), .A3(new_n462), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n639), .A2(new_n693), .A3(new_n632), .ZN(new_n694));
  OAI21_X1  g508(.A(KEYINPUT102), .B1(new_n692), .B2(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(new_n632), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n696), .B1(new_n544), .B2(new_n559), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n689), .B1(new_n688), .B2(new_n281), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n640), .A2(new_n678), .A3(KEYINPUT101), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT102), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n697), .A2(new_n700), .A3(new_n701), .A4(new_n693), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n695), .A2(new_n702), .ZN(new_n703));
  XOR2_X1   g517(.A(KEYINPUT103), .B(G119), .Z(new_n704));
  XNOR2_X1  g518(.A(new_n703), .B(new_n704), .ZN(G21));
  NAND2_X1  g519(.A1(new_n539), .A2(new_n540), .ZN(new_n706));
  OAI211_X1 g520(.A(new_n531), .B(new_n706), .C1(new_n517), .C2(new_n551), .ZN(new_n707));
  AOI22_X1  g521(.A1(new_n565), .A2(G472), .B1(new_n707), .B2(new_n496), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n708), .A2(new_n494), .A3(new_n650), .A4(new_n587), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n678), .A2(new_n640), .A3(new_n621), .ZN(new_n710));
  OR2_X1    g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G122), .ZN(G24));
  NAND2_X1  g526(.A1(new_n565), .A2(G472), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n707), .A2(new_n496), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n713), .A2(new_n632), .A3(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(new_n715), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n669), .A2(new_n700), .A3(new_n670), .A4(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G125), .ZN(G27));
  INV_X1    g532(.A(KEYINPUT42), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n669), .A2(new_n670), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n278), .A2(new_n280), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n721), .A2(new_n189), .A3(new_n353), .ZN(new_n722));
  INV_X1    g536(.A(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n723), .A2(new_n639), .A3(new_n494), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n719), .B1(new_n720), .B2(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(new_n724), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n726), .A2(KEYINPUT42), .A3(new_n669), .A4(new_n670), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G131), .ZN(G33));
  INV_X1    g543(.A(KEYINPUT104), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n646), .B(new_n730), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n731), .A2(new_n560), .A3(new_n723), .ZN(new_n732));
  XOR2_X1   g546(.A(KEYINPUT105), .B(G134), .Z(new_n733));
  XNOR2_X1  g547(.A(new_n732), .B(new_n733), .ZN(G36));
  NAND2_X1  g548(.A1(new_n651), .A2(new_n666), .ZN(new_n735));
  OR2_X1    g549(.A1(new_n735), .A2(KEYINPUT43), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(KEYINPUT43), .ZN(new_n737));
  AND2_X1   g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n566), .A2(new_n696), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT44), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n721), .A2(new_n189), .ZN(new_n743));
  INV_X1    g557(.A(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n738), .A2(KEYINPUT44), .A3(new_n739), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n742), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT106), .ZN(new_n747));
  AND2_X1   g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  OR2_X1    g562(.A1(new_n347), .A2(KEYINPUT45), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n347), .A2(KEYINPUT45), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n749), .A2(G469), .A3(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(new_n289), .ZN(new_n752));
  AOI21_X1  g566(.A(KEYINPUT46), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(new_n352), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n751), .A2(KEYINPUT46), .A3(new_n752), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n287), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(new_n653), .ZN(new_n758));
  INV_X1    g572(.A(new_n758), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n759), .B1(new_n746), .B2(new_n747), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n748), .A2(new_n760), .ZN(new_n761));
  XOR2_X1   g575(.A(KEYINPUT107), .B(G137), .Z(new_n762));
  XNOR2_X1  g576(.A(new_n761), .B(new_n762), .ZN(G39));
  OR4_X1    g577(.A1(new_n639), .A2(new_n720), .A3(new_n494), .A4(new_n743), .ZN(new_n764));
  XOR2_X1   g578(.A(new_n757), .B(KEYINPUT47), .Z(new_n765));
  NOR2_X1   g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(new_n364), .ZN(G42));
  NOR4_X1   g581(.A1(new_n663), .A2(new_n495), .A3(new_n188), .A4(new_n287), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n686), .A2(new_n352), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n735), .B1(KEYINPUT49), .B2(new_n769), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n637), .A2(new_n638), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n660), .A2(new_n656), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  OR2_X1    g587(.A1(new_n769), .A2(KEYINPUT49), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n768), .A2(new_n770), .A3(new_n773), .A4(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT51), .ZN(new_n776));
  INV_X1    g590(.A(new_n460), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n743), .A2(new_n688), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n773), .A2(new_n494), .A3(new_n777), .A4(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(KEYINPUT114), .ZN(new_n780));
  NOR3_X1   g594(.A1(new_n780), .A2(new_n650), .A3(new_n666), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n736), .A2(new_n777), .A3(new_n737), .A4(new_n778), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n782), .A2(new_n715), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT115), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n776), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  XOR2_X1   g600(.A(KEYINPUT112), .B(KEYINPUT50), .Z(new_n787));
  AND2_X1   g601(.A1(new_n708), .A2(new_n494), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n736), .A2(new_n777), .A3(new_n788), .A4(new_n737), .ZN(new_n789));
  OR3_X1    g603(.A1(new_n663), .A2(new_n189), .A3(new_n688), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n787), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(KEYINPUT113), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n789), .A2(new_n790), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(KEYINPUT50), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT113), .ZN(new_n795));
  OAI211_X1 g609(.A(new_n795), .B(new_n787), .C1(new_n789), .C2(new_n790), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n792), .A2(new_n794), .A3(new_n796), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n765), .B1(new_n286), .B2(new_n769), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n789), .A2(new_n743), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  OAI21_X1  g614(.A(KEYINPUT115), .B1(new_n781), .B2(new_n783), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n786), .A2(new_n797), .A3(new_n800), .A4(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(new_n579), .ZN(new_n803));
  OAI221_X1 g617(.A(new_n458), .B1(new_n692), .B2(new_n789), .C1(new_n780), .C2(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n639), .A2(new_n494), .ZN(new_n805));
  NOR3_X1   g619(.A1(new_n782), .A2(KEYINPUT48), .A3(new_n805), .ZN(new_n806));
  XOR2_X1   g620(.A(new_n806), .B(KEYINPUT116), .Z(new_n807));
  OAI21_X1  g621(.A(KEYINPUT48), .B1(new_n782), .B2(new_n805), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(KEYINPUT117), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n804), .B1(new_n807), .B2(new_n809), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n784), .A2(new_n797), .A3(new_n800), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(new_n776), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n802), .A2(new_n810), .A3(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT54), .ZN(new_n814));
  AND2_X1   g628(.A1(new_n695), .A2(new_n702), .ZN(new_n815));
  INV_X1    g629(.A(new_n679), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n609), .A2(new_n623), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n818), .A2(new_n680), .A3(new_n711), .ZN(new_n819));
  OAI21_X1  g633(.A(KEYINPUT108), .B1(new_n815), .B2(new_n819), .ZN(new_n820));
  OAI22_X1  g634(.A1(new_n679), .A2(new_n581), .B1(new_n709), .B2(new_n710), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n683), .A2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT108), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n822), .A2(new_n703), .A3(new_n823), .ZN(new_n824));
  AND2_X1   g638(.A1(new_n820), .A2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(new_n353), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n696), .A2(KEYINPUT111), .A3(new_n645), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT111), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n828), .B1(new_n632), .B2(new_n644), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n826), .B1(new_n827), .B2(new_n829), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n651), .A2(new_n586), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n830), .A2(new_n661), .A3(new_n831), .A4(new_n640), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n671), .A2(new_n648), .A3(new_n717), .A4(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT52), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n833), .B(new_n834), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n715), .A2(new_n722), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n669), .A2(new_n836), .A3(new_n670), .ZN(new_n837));
  AND4_X1   g651(.A1(new_n586), .A2(new_n601), .A3(new_n605), .A4(new_n645), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n697), .A2(new_n723), .A3(new_n838), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n732), .A2(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n728), .A2(new_n837), .A3(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n563), .A2(new_n566), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n579), .A2(new_n283), .A3(new_n621), .A4(new_n284), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n842), .B1(new_n843), .B2(KEYINPUT109), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n283), .A2(new_n284), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT109), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n845), .A2(new_n846), .A3(new_n621), .A4(new_n579), .ZN(new_n847));
  AOI22_X1  g661(.A1(new_n844), .A2(new_n847), .B1(new_n560), .B2(new_n464), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n651), .A2(new_n563), .A3(new_n566), .A4(new_n587), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n283), .A2(new_n621), .A3(new_n284), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  OAI21_X1  g665(.A(KEYINPUT110), .B1(new_n851), .B2(new_n634), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n650), .A2(new_n586), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n567), .A2(new_n845), .A3(new_n621), .A4(new_n853), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n566), .A2(new_n632), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n845), .A2(new_n855), .A3(new_n693), .A4(new_n353), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT110), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n854), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n848), .A2(new_n852), .A3(new_n858), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n841), .A2(new_n859), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n648), .A2(new_n717), .ZN(new_n861));
  OR2_X1    g675(.A1(new_n861), .A2(new_n834), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT53), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n825), .A2(new_n835), .A3(new_n860), .A4(new_n864), .ZN(new_n865));
  AND3_X1   g679(.A1(new_n848), .A2(new_n852), .A3(new_n858), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n732), .A2(new_n839), .A3(new_n837), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n867), .B1(new_n725), .B2(new_n727), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n820), .A2(new_n866), .A3(new_n868), .A4(new_n824), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n833), .B(KEYINPUT52), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n863), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n814), .B1(new_n865), .B2(new_n871), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n815), .A2(new_n819), .A3(new_n863), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n835), .A2(new_n860), .A3(new_n862), .A4(new_n873), .ZN(new_n874));
  AND3_X1   g688(.A1(new_n871), .A2(new_n814), .A3(new_n874), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n813), .A2(new_n872), .A3(new_n875), .ZN(new_n876));
  NOR2_X1   g690(.A1(G952), .A2(G953), .ZN(new_n877));
  XOR2_X1   g691(.A(new_n877), .B(KEYINPUT118), .Z(new_n878));
  OAI21_X1  g692(.A(new_n775), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(KEYINPUT119), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT119), .ZN(new_n881));
  OAI211_X1 g695(.A(new_n881), .B(new_n775), .C1(new_n876), .C2(new_n878), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n880), .A2(new_n882), .ZN(G75));
  NOR2_X1   g697(.A1(new_n330), .A2(G952), .ZN(new_n884));
  INV_X1    g698(.A(new_n884), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n275), .B1(new_n871), .B2(new_n874), .ZN(new_n886));
  AOI21_X1  g700(.A(KEYINPUT56), .B1(new_n886), .B2(G210), .ZN(new_n887));
  XOR2_X1   g701(.A(new_n614), .B(KEYINPUT120), .Z(new_n888));
  XNOR2_X1  g702(.A(new_n888), .B(KEYINPUT55), .ZN(new_n889));
  XOR2_X1   g703(.A(new_n889), .B(KEYINPUT121), .Z(new_n890));
  XNOR2_X1  g704(.A(new_n890), .B(new_n262), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n885), .B1(new_n887), .B2(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n892), .B1(new_n887), .B2(new_n891), .ZN(G51));
  AOI21_X1  g707(.A(new_n814), .B1(new_n871), .B2(new_n874), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n875), .A2(new_n894), .ZN(new_n895));
  XOR2_X1   g709(.A(new_n289), .B(KEYINPUT57), .Z(new_n896));
  OAI22_X1  g710(.A1(new_n895), .A2(new_n896), .B1(new_n349), .B2(new_n351), .ZN(new_n897));
  INV_X1    g711(.A(new_n751), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n886), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n884), .B1(new_n897), .B2(new_n899), .ZN(G54));
  AND3_X1   g714(.A1(new_n886), .A2(KEYINPUT58), .A3(G475), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n885), .B1(new_n901), .B2(new_n412), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n902), .B1(new_n412), .B2(new_n901), .ZN(G60));
  INV_X1    g717(.A(KEYINPUT122), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n572), .A2(new_n574), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n576), .B(KEYINPUT59), .Z(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n871), .A2(new_n874), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(KEYINPUT54), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n871), .A2(new_n874), .A3(new_n814), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n907), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n904), .B1(new_n911), .B2(new_n884), .ZN(new_n912));
  OAI211_X1 g726(.A(KEYINPUT122), .B(new_n885), .C1(new_n895), .C2(new_n907), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n906), .B1(new_n875), .B2(new_n872), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n914), .A2(new_n574), .A3(new_n572), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n912), .A2(new_n913), .A3(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT123), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n912), .A2(new_n913), .A3(new_n915), .A4(KEYINPUT123), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n918), .A2(new_n919), .ZN(G63));
  NAND2_X1  g734(.A1(G217), .A2(G902), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(KEYINPUT60), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n922), .B1(new_n871), .B2(new_n874), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n885), .B1(new_n923), .B2(new_n492), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n924), .B1(new_n630), .B2(new_n923), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n925), .B(KEYINPUT61), .ZN(G66));
  OAI21_X1  g740(.A(G953), .B1(new_n454), .B2(new_n260), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n927), .B(KEYINPUT124), .Z(new_n928));
  AND2_X1   g742(.A1(new_n825), .A2(new_n866), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n928), .B1(new_n929), .B2(G953), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n888), .B1(G898), .B2(new_n330), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n930), .B(new_n931), .ZN(G69));
  NAND3_X1  g746(.A1(new_n560), .A2(new_n640), .A3(new_n831), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n732), .B1(new_n758), .B2(new_n933), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n766), .A2(new_n934), .ZN(new_n935));
  AND2_X1   g749(.A1(new_n861), .A2(new_n671), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n935), .A2(new_n728), .A3(new_n936), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n761), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(new_n330), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n523), .B(KEYINPUT125), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(new_n404), .ZN(new_n941));
  NAND2_X1  g755(.A1(G900), .A2(G953), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n939), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  OR2_X1    g757(.A1(new_n748), .A2(new_n760), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n936), .A2(new_n664), .ZN(new_n945));
  OR2_X1    g759(.A1(new_n945), .A2(KEYINPUT62), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n945), .A2(KEYINPUT62), .ZN(new_n947));
  INV_X1    g761(.A(new_n766), .ZN(new_n948));
  OAI211_X1 g762(.A(new_n726), .B(new_n653), .C1(new_n579), .C2(new_n853), .ZN(new_n949));
  AND3_X1   g763(.A1(new_n947), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n944), .A2(KEYINPUT126), .A3(new_n946), .A4(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT126), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n946), .A2(new_n948), .A3(new_n947), .A4(new_n949), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n952), .B1(new_n953), .B2(new_n761), .ZN(new_n954));
  AOI21_X1  g768(.A(G953), .B1(new_n951), .B2(new_n954), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n943), .B1(new_n955), .B2(new_n941), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n330), .B1(G227), .B2(G900), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(new_n957), .ZN(new_n959));
  OAI211_X1 g773(.A(new_n943), .B(new_n959), .C1(new_n955), .C2(new_n941), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n958), .A2(new_n960), .ZN(G72));
  NAND2_X1  g775(.A1(new_n553), .A2(new_n517), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n951), .A2(new_n954), .A3(new_n929), .ZN(new_n963));
  NAND2_X1  g777(.A1(G472), .A2(G902), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n964), .B(KEYINPUT63), .Z(new_n965));
  XOR2_X1   g779(.A(new_n965), .B(KEYINPUT127), .Z(new_n966));
  AOI21_X1  g780(.A(new_n962), .B1(new_n963), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n657), .A2(new_n554), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n968), .A2(new_n965), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n969), .B1(new_n865), .B2(new_n871), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n528), .A2(new_n512), .A3(new_n516), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n938), .A2(new_n929), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n971), .B1(new_n972), .B2(new_n966), .ZN(new_n973));
  NOR4_X1   g787(.A1(new_n967), .A2(new_n970), .A3(new_n884), .A4(new_n973), .ZN(G57));
endmodule


