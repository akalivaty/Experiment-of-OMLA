

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805;

  XNOR2_X1 U379 ( .A(n421), .B(n490), .ZN(n464) );
  XNOR2_X1 U380 ( .A(n623), .B(n622), .ZN(n736) );
  NAND2_X1 U381 ( .A1(n764), .A2(KEYINPUT79), .ZN(n378) );
  XOR2_X1 U382 ( .A(n619), .B(KEYINPUT75), .Z(n356) );
  NOR2_X1 U383 ( .A1(n726), .A2(n724), .ZN(n642) );
  OR2_X1 U384 ( .A1(n711), .A2(G902), .ZN(n443) );
  XNOR2_X1 U385 ( .A(G104), .B(G110), .ZN(n511) );
  INV_X1 U386 ( .A(KEYINPUT64), .ZN(n376) );
  NOR2_X1 U387 ( .A1(n767), .A2(n768), .ZN(n468) );
  OR2_X1 U388 ( .A1(n697), .A2(n689), .ZN(n358) );
  NOR2_X1 U389 ( .A1(n424), .A2(n730), .ZN(n423) );
  XNOR2_X1 U390 ( .A(n364), .B(n363), .ZN(n362) );
  OR2_X1 U391 ( .A1(n715), .A2(n727), .ZN(n644) );
  NAND2_X1 U392 ( .A1(n457), .A2(n454), .ZN(n804) );
  XNOR2_X1 U393 ( .A(n646), .B(KEYINPUT104), .ZN(n596) );
  XNOR2_X1 U394 ( .A(n372), .B(n371), .ZN(n743) );
  NAND2_X1 U395 ( .A1(n456), .A2(n455), .ZN(n454) );
  AND2_X1 U396 ( .A1(n459), .A2(n458), .ZN(n457) );
  AND2_X1 U397 ( .A1(n504), .A2(n606), .ZN(n730) );
  NAND2_X1 U398 ( .A1(n374), .A2(n373), .ZN(n372) );
  XNOR2_X1 U399 ( .A(n741), .B(KEYINPUT113), .ZN(n374) );
  NOR2_X1 U400 ( .A1(n671), .A2(n435), .ZN(n505) );
  INV_X1 U401 ( .A(n742), .ZN(n373) );
  XNOR2_X1 U402 ( .A(n359), .B(KEYINPUT112), .ZN(n739) );
  OR2_X1 U403 ( .A1(n360), .A2(n738), .ZN(n359) );
  OR2_X1 U404 ( .A1(n645), .A2(n662), .ZN(n436) );
  XNOR2_X1 U405 ( .A(n361), .B(KEYINPUT49), .ZN(n360) );
  NAND2_X1 U406 ( .A1(n736), .A2(n737), .ZN(n361) );
  XNOR2_X1 U407 ( .A(n569), .B(n568), .ZN(n601) );
  XNOR2_X1 U408 ( .A(n583), .B(n439), .ZN(n599) );
  OR2_X1 U409 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U410 ( .A(n429), .B(n541), .ZN(n542) );
  XNOR2_X1 U411 ( .A(n369), .B(n368), .ZN(n429) );
  AND2_X1 U412 ( .A1(n695), .A2(n690), .ZN(n691) );
  AND2_X1 U413 ( .A1(n479), .A2(KEYINPUT84), .ZN(n620) );
  XNOR2_X1 U414 ( .A(n511), .B(G107), .ZN(n420) );
  XNOR2_X1 U415 ( .A(n370), .B(KEYINPUT24), .ZN(n369) );
  INV_X1 U416 ( .A(KEYINPUT44), .ZN(n379) );
  INV_X1 U417 ( .A(KEYINPUT84), .ZN(n380) );
  XNOR2_X1 U418 ( .A(KEYINPUT114), .B(KEYINPUT51), .ZN(n371) );
  XNOR2_X1 U419 ( .A(G128), .B(G119), .ZN(n368) );
  INV_X1 U420 ( .A(KEYINPUT117), .ZN(n363) );
  INV_X1 U421 ( .A(KEYINPUT23), .ZN(n370) );
  XNOR2_X1 U422 ( .A(G101), .B(KEYINPUT67), .ZN(n405) );
  NAND2_X1 U423 ( .A1(n357), .A2(n696), .ZN(n375) );
  NAND2_X1 U424 ( .A1(n358), .A2(n691), .ZN(n357) );
  NAND2_X1 U425 ( .A1(n362), .A2(n763), .ZN(n768) );
  NAND2_X1 U426 ( .A1(n366), .A2(n365), .ZN(n364) );
  INV_X1 U427 ( .A(n760), .ZN(n365) );
  XNOR2_X1 U428 ( .A(n759), .B(n367), .ZN(n366) );
  INV_X1 U429 ( .A(KEYINPUT52), .ZN(n367) );
  NAND2_X1 U430 ( .A1(n375), .A2(n378), .ZN(n377) );
  XNOR2_X2 U431 ( .A(n377), .B(n376), .ZN(n701) );
  OR2_X2 U432 ( .A1(n697), .A2(n792), .ZN(n764) );
  OR2_X2 U433 ( .A1(n381), .A2(n379), .ZN(n649) );
  NAND2_X1 U434 ( .A1(n381), .A2(n380), .ZN(n476) );
  NAND2_X1 U435 ( .A1(n381), .A2(n620), .ZN(n630) );
  XNOR2_X1 U436 ( .A(n381), .B(G122), .ZN(G24) );
  XNOR2_X2 U437 ( .A(n480), .B(n356), .ZN(n381) );
  INV_X1 U438 ( .A(n382), .ZN(n383) );
  INV_X1 U439 ( .A(G143), .ZN(n382) );
  XNOR2_X1 U440 ( .A(n791), .B(G146), .ZN(n384) );
  BUF_X1 U441 ( .A(n567), .Z(n385) );
  XNOR2_X1 U442 ( .A(n791), .B(G146), .ZN(n555) );
  XNOR2_X2 U443 ( .A(n567), .B(n387), .ZN(n791) );
  INV_X1 U444 ( .A(G902), .ZN(n522) );
  NAND2_X1 U445 ( .A1(n596), .A2(n478), .ZN(n477) );
  NAND2_X1 U446 ( .A1(n803), .A2(n479), .ZN(n475) );
  AND2_X1 U447 ( .A1(n595), .A2(n479), .ZN(n478) );
  INV_X1 U448 ( .A(KEYINPUT0), .ZN(n416) );
  NAND2_X1 U449 ( .A1(n450), .A2(n434), .ZN(n422) );
  XNOR2_X1 U450 ( .A(n562), .B(n561), .ZN(n563) );
  INV_X1 U451 ( .A(KEYINPUT7), .ZN(n561) );
  XOR2_X1 U452 ( .A(G122), .B(KEYINPUT9), .Z(n562) );
  INV_X1 U453 ( .A(G134), .ZN(n526) );
  INV_X1 U454 ( .A(KEYINPUT87), .ZN(n486) );
  INV_X1 U455 ( .A(G237), .ZN(n521) );
  NOR2_X1 U456 ( .A1(n712), .A2(n388), .ZN(n430) );
  XNOR2_X1 U457 ( .A(n492), .B(G146), .ZN(n536) );
  INV_X1 U458 ( .A(G125), .ZN(n492) );
  XNOR2_X1 U459 ( .A(n584), .B(n440), .ZN(n439) );
  INV_X1 U460 ( .A(G475), .ZN(n440) );
  XNOR2_X1 U461 ( .A(n545), .B(KEYINPUT25), .ZN(n506) );
  XNOR2_X1 U462 ( .A(n738), .B(KEYINPUT6), .ZN(n645) );
  XNOR2_X1 U463 ( .A(n488), .B(n515), .ZN(n531) );
  XNOR2_X1 U464 ( .A(n406), .B(n405), .ZN(n488) );
  XNOR2_X1 U465 ( .A(KEYINPUT3), .B(G119), .ZN(n406) );
  XOR2_X1 U466 ( .A(G137), .B(G140), .Z(n556) );
  XNOR2_X1 U467 ( .A(n472), .B(KEYINPUT91), .ZN(n471) );
  INV_X1 U468 ( .A(G101), .ZN(n472) );
  INV_X1 U469 ( .A(KEYINPUT39), .ZN(n659) );
  INV_X1 U470 ( .A(KEYINPUT90), .ZN(n415) );
  XNOR2_X1 U471 ( .A(n407), .B(n394), .ZN(n621) );
  AND2_X1 U472 ( .A1(n441), .A2(n645), .ZN(n411) );
  NAND2_X1 U473 ( .A1(n495), .A2(n783), .ZN(n494) );
  INV_X1 U474 ( .A(n500), .ZN(n495) );
  XNOR2_X1 U475 ( .A(KEYINPUT86), .B(KEYINPUT15), .ZN(n520) );
  NAND2_X1 U476 ( .A1(G234), .A2(G237), .ZN(n546) );
  XNOR2_X1 U477 ( .A(G137), .B(KEYINPUT94), .ZN(n527) );
  INV_X1 U478 ( .A(n732), .ZN(n444) );
  INV_X1 U479 ( .A(KEYINPUT48), .ZN(n490) );
  NAND2_X1 U480 ( .A1(n423), .A2(n422), .ZN(n421) );
  XNOR2_X1 U481 ( .A(n566), .B(n431), .ZN(n782) );
  XNOR2_X1 U482 ( .A(n564), .B(n563), .ZN(n566) );
  XNOR2_X1 U483 ( .A(G116), .B(G107), .ZN(n565) );
  NOR2_X1 U484 ( .A1(G953), .A2(G237), .ZN(n570) );
  XNOR2_X1 U485 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U486 ( .A(n518), .B(n486), .ZN(n485) );
  XNOR2_X1 U487 ( .A(n413), .B(n414), .ZN(n612) );
  INV_X1 U488 ( .A(KEYINPUT71), .ZN(n414) );
  INV_X1 U489 ( .A(KEYINPUT30), .ZN(n462) );
  INV_X1 U490 ( .A(KEYINPUT19), .ZN(n425) );
  XNOR2_X1 U491 ( .A(n540), .B(n539), .ZN(n541) );
  INV_X1 U492 ( .A(G110), .ZN(n539) );
  XNOR2_X1 U493 ( .A(KEYINPUT93), .B(KEYINPUT92), .ZN(n540) );
  XNOR2_X1 U494 ( .A(n580), .B(n491), .ZN(n790) );
  INV_X1 U495 ( .A(n556), .ZN(n491) );
  XOR2_X1 U496 ( .A(G140), .B(G104), .Z(n578) );
  XNOR2_X1 U497 ( .A(n536), .B(n535), .ZN(n580) );
  INV_X1 U498 ( .A(KEYINPUT10), .ZN(n535) );
  XNOR2_X1 U499 ( .A(n409), .B(n408), .ZN(n666) );
  INV_X1 U500 ( .A(KEYINPUT28), .ZN(n408) );
  NOR2_X1 U501 ( .A1(n751), .A2(n749), .ZN(n667) );
  NOR2_X1 U502 ( .A1(n661), .A2(n460), .ZN(n455) );
  XNOR2_X1 U503 ( .A(n436), .B(KEYINPUT106), .ZN(n604) );
  XNOR2_X1 U504 ( .A(KEYINPUT68), .B(KEYINPUT34), .ZN(n615) );
  BUF_X1 U505 ( .A(n670), .Z(n435) );
  AND2_X1 U506 ( .A1(n621), .A2(n441), .ZN(n646) );
  XNOR2_X1 U507 ( .A(n531), .B(n487), .ZN(n608) );
  XNOR2_X1 U508 ( .A(n420), .B(n514), .ZN(n487) );
  INV_X1 U509 ( .A(G122), .ZN(n512) );
  XNOR2_X1 U510 ( .A(n473), .B(n470), .ZN(n469) );
  XNOR2_X1 U511 ( .A(n510), .B(n471), .ZN(n470) );
  NAND2_X1 U512 ( .A1(n435), .A2(n446), .ZN(n445) );
  XNOR2_X1 U513 ( .A(n448), .B(n447), .ZN(n446) );
  INV_X1 U514 ( .A(KEYINPUT43), .ZN(n447) );
  NOR2_X1 U515 ( .A1(n671), .A2(n606), .ZN(n448) );
  INV_X1 U516 ( .A(KEYINPUT100), .ZN(n438) );
  NOR2_X1 U517 ( .A1(n640), .A2(n639), .ZN(n724) );
  OR2_X1 U518 ( .A1(n634), .A2(n426), .ZN(n635) );
  NAND2_X1 U519 ( .A1(n663), .A2(n427), .ZN(n426) );
  INV_X1 U520 ( .A(n733), .ZN(n427) );
  AND2_X1 U521 ( .A1(n648), .A2(n647), .ZN(n712) );
  XNOR2_X1 U522 ( .A(n412), .B(KEYINPUT83), .ZN(n648) );
  NAND2_X1 U523 ( .A1(n498), .A2(n497), .ZN(n496) );
  NAND2_X1 U524 ( .A1(n494), .A2(n502), .ZN(n493) );
  INV_X1 U525 ( .A(KEYINPUT53), .ZN(n465) );
  AND2_X1 U526 ( .A1(n453), .A2(n669), .ZN(n386) );
  XOR2_X1 U527 ( .A(G131), .B(KEYINPUT4), .Z(n387) );
  AND2_X1 U528 ( .A1(n644), .A2(n643), .ZN(n388) );
  XOR2_X1 U529 ( .A(n593), .B(n592), .Z(n389) );
  OR2_X1 U530 ( .A1(n590), .A2(n589), .ZN(n390) );
  AND2_X1 U531 ( .A1(n445), .A2(n444), .ZN(n391) );
  AND2_X1 U532 ( .A1(n430), .A2(n649), .ZN(n392) );
  AND2_X1 U533 ( .A1(n391), .A2(n688), .ZN(n393) );
  XNOR2_X1 U534 ( .A(KEYINPUT69), .B(KEYINPUT22), .ZN(n394) );
  XOR2_X1 U535 ( .A(n711), .B(KEYINPUT62), .Z(n395) );
  INV_X1 U536 ( .A(KEYINPUT44), .ZN(n479) );
  INV_X1 U537 ( .A(n783), .ZN(n503) );
  XOR2_X1 U538 ( .A(KEYINPUT63), .B(KEYINPUT85), .Z(n396) );
  AND2_X1 U539 ( .A1(n707), .A2(G953), .ZN(n789) );
  INV_X1 U540 ( .A(n789), .ZN(n502) );
  XNOR2_X1 U541 ( .A(n433), .B(n790), .ZN(n787) );
  OR2_X2 U542 ( .A1(n787), .A2(G902), .ZN(n507) );
  NOR2_X1 U543 ( .A1(n701), .A2(n766), .ZN(n397) );
  NOR2_X2 U544 ( .A1(n701), .A2(n766), .ZN(n781) );
  XNOR2_X1 U545 ( .A(G131), .B(n383), .ZN(n577) );
  BUF_X1 U546 ( .A(n636), .Z(n398) );
  AND2_X1 U547 ( .A1(n454), .A2(n453), .ZN(n449) );
  XNOR2_X1 U548 ( .A(n542), .B(n538), .ZN(n433) );
  XNOR2_X1 U549 ( .A(n557), .B(G469), .ZN(n636) );
  NOR2_X1 U550 ( .A1(G902), .A2(n769), .ZN(n557) );
  XNOR2_X1 U551 ( .A(n555), .B(n469), .ZN(n769) );
  NAND2_X1 U552 ( .A1(n608), .A2(n484), .ZN(n401) );
  NAND2_X1 U553 ( .A1(n399), .A2(n400), .ZN(n402) );
  NAND2_X1 U554 ( .A1(n401), .A2(n402), .ZN(n704) );
  INV_X1 U555 ( .A(n608), .ZN(n399) );
  INV_X1 U556 ( .A(n484), .ZN(n400) );
  BUF_X1 U557 ( .A(n673), .Z(n403) );
  NOR2_X1 U558 ( .A1(n708), .A2(n789), .ZN(n710) );
  NOR2_X1 U559 ( .A1(n779), .A2(n789), .ZN(n780) );
  XNOR2_X1 U560 ( .A(n419), .B(n395), .ZN(n418) );
  NAND2_X1 U561 ( .A1(n397), .A2(G472), .ZN(n419) );
  BUF_X1 U562 ( .A(n697), .Z(n404) );
  XNOR2_X1 U563 ( .A(n432), .B(n650), .ZN(n697) );
  BUF_X1 U564 ( .A(n734), .Z(n441) );
  NAND2_X1 U565 ( .A1(n637), .A2(n389), .ZN(n407) );
  XNOR2_X2 U566 ( .A(n591), .B(n416), .ZN(n637) );
  INV_X1 U567 ( .A(n738), .ZN(n663) );
  NAND2_X1 U568 ( .A1(n410), .A2(n738), .ZN(n409) );
  XNOR2_X2 U569 ( .A(n443), .B(G472), .ZN(n738) );
  INV_X1 U570 ( .A(n662), .ZN(n410) );
  NAND2_X1 U571 ( .A1(n621), .A2(n411), .ZN(n412) );
  NOR2_X2 U572 ( .A1(n734), .A2(n733), .ZN(n413) );
  XNOR2_X1 U573 ( .A(n636), .B(n598), .ZN(n734) );
  XNOR2_X1 U574 ( .A(n637), .B(n415), .ZN(n634) );
  XNOR2_X1 U575 ( .A(n417), .B(n396), .ZN(G57) );
  NAND2_X1 U576 ( .A1(n418), .A2(n502), .ZN(n417) );
  XNOR2_X1 U577 ( .A(n420), .B(n556), .ZN(n473) );
  AND2_X1 U578 ( .A1(n612), .A2(n738), .ZN(n742) );
  INV_X1 U579 ( .A(n684), .ZN(n424) );
  NAND2_X1 U580 ( .A1(n673), .A2(n390), .ZN(n591) );
  XNOR2_X1 U581 ( .A(n489), .B(n425), .ZN(n673) );
  NOR2_X1 U582 ( .A1(n672), .A2(n761), .ZN(n668) );
  NOR2_X2 U583 ( .A1(n744), .A2(n634), .ZN(n616) );
  NAND2_X1 U584 ( .A1(n428), .A2(n392), .ZN(n432) );
  NAND2_X1 U585 ( .A1(n633), .A2(n632), .ZN(n428) );
  XNOR2_X1 U586 ( .A(n385), .B(n565), .ZN(n431) );
  INV_X1 U587 ( .A(n669), .ZN(n461) );
  XNOR2_X1 U588 ( .A(n463), .B(n462), .ZN(n509) );
  NOR2_X2 U589 ( .A1(n670), .A2(n587), .ZN(n489) );
  NAND2_X1 U590 ( .A1(n738), .A2(n745), .ZN(n463) );
  NAND2_X1 U591 ( .A1(n452), .A2(n386), .ZN(n434) );
  NOR2_X1 U592 ( .A1(n679), .A2(n437), .ZN(n681) );
  NOR2_X1 U593 ( .A1(n678), .A2(KEYINPUT47), .ZN(n437) );
  XNOR2_X2 U594 ( .A(n641), .B(n438), .ZN(n726) );
  NAND2_X1 U595 ( .A1(n477), .A2(n475), .ZN(n474) );
  XNOR2_X2 U596 ( .A(n442), .B(n526), .ZN(n567) );
  XNOR2_X1 U597 ( .A(n442), .B(n536), .ZN(n482) );
  XNOR2_X2 U598 ( .A(n519), .B(G128), .ZN(n442) );
  INV_X1 U599 ( .A(n445), .ZN(n687) );
  NAND2_X1 U600 ( .A1(n449), .A2(n457), .ZN(n451) );
  INV_X1 U601 ( .A(n804), .ZN(n452) );
  NAND2_X1 U602 ( .A1(n451), .A2(n461), .ZN(n450) );
  INV_X1 U603 ( .A(n802), .ZN(n453) );
  INV_X1 U604 ( .A(n685), .ZN(n456) );
  NAND2_X1 U605 ( .A1(n661), .A2(n460), .ZN(n458) );
  NAND2_X1 U606 ( .A1(n685), .A2(n460), .ZN(n459) );
  INV_X1 U607 ( .A(KEYINPUT40), .ZN(n460) );
  NAND2_X1 U608 ( .A1(n464), .A2(n393), .ZN(n689) );
  NAND2_X1 U609 ( .A1(n464), .A2(n391), .ZN(n792) );
  XNOR2_X1 U610 ( .A(n466), .B(n465), .ZN(G75) );
  NAND2_X1 U611 ( .A1(n467), .A2(n793), .ZN(n466) );
  XNOR2_X1 U612 ( .A(n468), .B(KEYINPUT118), .ZN(n467) );
  NAND2_X1 U613 ( .A1(n476), .A2(n474), .ZN(n632) );
  NOR2_X1 U614 ( .A1(n803), .A2(n629), .ZN(n631) );
  AND2_X1 U615 ( .A1(n596), .A2(n595), .ZN(n629) );
  NAND2_X1 U616 ( .A1(n618), .A2(n617), .ZN(n480) );
  XNOR2_X1 U617 ( .A(n481), .B(n485), .ZN(n483) );
  XNOR2_X1 U618 ( .A(n517), .B(n516), .ZN(n481) );
  XNOR2_X2 U619 ( .A(n525), .B(n524), .ZN(n670) );
  INV_X1 U620 ( .A(n701), .ZN(n501) );
  NOR2_X2 U621 ( .A1(n496), .A2(n493), .ZN(n784) );
  NAND2_X1 U622 ( .A1(n701), .A2(n783), .ZN(n497) );
  NAND2_X1 U623 ( .A1(n499), .A2(n501), .ZN(n498) );
  AND2_X1 U624 ( .A1(n500), .A2(n503), .ZN(n499) );
  NOR2_X2 U625 ( .A1(n766), .A2(n569), .ZN(n500) );
  XNOR2_X1 U626 ( .A(n505), .B(KEYINPUT36), .ZN(n504) );
  NAND2_X1 U627 ( .A1(n605), .A2(n745), .ZN(n671) );
  XNOR2_X2 U628 ( .A(n507), .B(n506), .ZN(n623) );
  XNOR2_X1 U629 ( .A(n614), .B(n613), .ZN(n744) );
  NAND2_X1 U630 ( .A1(n612), .A2(n611), .ZN(n614) );
  BUF_X1 U631 ( .A(n397), .Z(n785) );
  XNOR2_X2 U632 ( .A(n660), .B(n659), .ZN(n685) );
  XNOR2_X2 U633 ( .A(n700), .B(n699), .ZN(n766) );
  AND2_X1 U634 ( .A1(n558), .A2(n664), .ZN(n508) );
  AND2_X1 U635 ( .A1(G227), .A2(n793), .ZN(n510) );
  XNOR2_X1 U636 ( .A(KEYINPUT70), .B(KEYINPUT16), .ZN(n513) );
  XNOR2_X1 U637 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U638 ( .A(G116), .B(G113), .ZN(n515) );
  XOR2_X1 U639 ( .A(KEYINPUT74), .B(KEYINPUT18), .Z(n517) );
  XNOR2_X1 U640 ( .A(KEYINPUT4), .B(KEYINPUT17), .ZN(n516) );
  INV_X2 U641 ( .A(G953), .ZN(n793) );
  NAND2_X1 U642 ( .A1(G224), .A2(n793), .ZN(n518) );
  INV_X2 U643 ( .A(G143), .ZN(n519) );
  XNOR2_X1 U644 ( .A(n520), .B(n522), .ZN(n695) );
  INV_X1 U645 ( .A(n695), .ZN(n543) );
  NAND2_X1 U646 ( .A1(n704), .A2(n543), .ZN(n525) );
  NAND2_X1 U647 ( .A1(n522), .A2(n521), .ZN(n534) );
  NAND2_X1 U648 ( .A1(n534), .A2(G210), .ZN(n523) );
  XNOR2_X1 U649 ( .A(n523), .B(KEYINPUT88), .ZN(n524) );
  INV_X1 U650 ( .A(n435), .ZN(n586) );
  XOR2_X1 U651 ( .A(KEYINPUT95), .B(KEYINPUT5), .Z(n528) );
  XNOR2_X1 U652 ( .A(n528), .B(n527), .ZN(n530) );
  NAND2_X1 U653 ( .A1(n570), .A2(G210), .ZN(n529) );
  XNOR2_X1 U654 ( .A(n530), .B(n529), .ZN(n532) );
  XNOR2_X1 U655 ( .A(n531), .B(n532), .ZN(n533) );
  XNOR2_X1 U656 ( .A(n384), .B(n533), .ZN(n711) );
  NAND2_X1 U657 ( .A1(n534), .A2(G214), .ZN(n745) );
  NAND2_X1 U658 ( .A1(G234), .A2(n793), .ZN(n537) );
  XOR2_X1 U659 ( .A(n537), .B(KEYINPUT8), .Z(n560) );
  AND2_X1 U660 ( .A1(G221), .A2(n560), .ZN(n538) );
  NAND2_X1 U661 ( .A1(G234), .A2(n543), .ZN(n544) );
  XNOR2_X1 U662 ( .A(n544), .B(KEYINPUT20), .ZN(n551) );
  NAND2_X1 U663 ( .A1(n551), .A2(G217), .ZN(n545) );
  XNOR2_X1 U664 ( .A(n546), .B(KEYINPUT14), .ZN(n547) );
  NAND2_X1 U665 ( .A1(G952), .A2(n547), .ZN(n760) );
  NOR2_X1 U666 ( .A1(n760), .A2(G953), .ZN(n589) );
  NAND2_X1 U667 ( .A1(n547), .A2(G902), .ZN(n548) );
  XNOR2_X1 U668 ( .A(n548), .B(KEYINPUT89), .ZN(n588) );
  NAND2_X1 U669 ( .A1(G953), .A2(n588), .ZN(n549) );
  NOR2_X1 U670 ( .A1(G900), .A2(n549), .ZN(n550) );
  NOR2_X1 U671 ( .A1(n589), .A2(n550), .ZN(n553) );
  NAND2_X1 U672 ( .A1(n551), .A2(G221), .ZN(n552) );
  XNOR2_X1 U673 ( .A(n552), .B(KEYINPUT21), .ZN(n737) );
  NOR2_X1 U674 ( .A1(n553), .A2(n737), .ZN(n602) );
  INV_X1 U675 ( .A(n602), .ZN(n554) );
  NOR2_X1 U676 ( .A1(n623), .A2(n554), .ZN(n558) );
  INV_X1 U677 ( .A(n398), .ZN(n664) );
  NAND2_X1 U678 ( .A1(n509), .A2(n508), .ZN(n559) );
  XNOR2_X1 U679 ( .A(n559), .B(KEYINPUT73), .ZN(n658) );
  INV_X1 U680 ( .A(G478), .ZN(n569) );
  NAND2_X1 U681 ( .A1(G217), .A2(n560), .ZN(n564) );
  OR2_X1 U682 ( .A1(G902), .A2(n782), .ZN(n568) );
  XNOR2_X1 U683 ( .A(KEYINPUT13), .B(KEYINPUT98), .ZN(n584) );
  XOR2_X1 U684 ( .A(KEYINPUT97), .B(KEYINPUT12), .Z(n572) );
  NAND2_X1 U685 ( .A1(G214), .A2(n570), .ZN(n571) );
  XNOR2_X1 U686 ( .A(n572), .B(n571), .ZN(n576) );
  XOR2_X1 U687 ( .A(KEYINPUT11), .B(KEYINPUT96), .Z(n574) );
  XNOR2_X1 U688 ( .A(G113), .B(G122), .ZN(n573) );
  XNOR2_X1 U689 ( .A(n574), .B(n573), .ZN(n575) );
  XOR2_X1 U690 ( .A(n576), .B(n575), .Z(n582) );
  XNOR2_X1 U691 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U692 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U693 ( .A(n581), .B(n582), .ZN(n776) );
  NOR2_X1 U694 ( .A1(n776), .A2(G902), .ZN(n583) );
  NOR2_X1 U695 ( .A1(n601), .A2(n599), .ZN(n617) );
  AND2_X1 U696 ( .A1(n658), .A2(n617), .ZN(n585) );
  NAND2_X1 U697 ( .A1(n586), .A2(n585), .ZN(n676) );
  XNOR2_X1 U698 ( .A(n676), .B(n383), .ZN(G45) );
  INV_X1 U699 ( .A(n745), .ZN(n587) );
  NOR2_X1 U700 ( .A1(G898), .A2(n793), .ZN(n607) );
  AND2_X1 U701 ( .A1(n588), .A2(n607), .ZN(n590) );
  NAND2_X1 U702 ( .A1(n599), .A2(n601), .ZN(n749) );
  NOR2_X1 U703 ( .A1(n749), .A2(n737), .ZN(n593) );
  INV_X1 U704 ( .A(KEYINPUT102), .ZN(n592) );
  INV_X1 U705 ( .A(KEYINPUT65), .ZN(n594) );
  XNOR2_X1 U706 ( .A(n594), .B(KEYINPUT1), .ZN(n598) );
  AND2_X1 U707 ( .A1(n623), .A2(n663), .ZN(n595) );
  XNOR2_X1 U708 ( .A(G110), .B(KEYINPUT109), .ZN(n597) );
  XNOR2_X1 U709 ( .A(n629), .B(n597), .ZN(G12) );
  XOR2_X1 U710 ( .A(n398), .B(n598), .Z(n606) );
  INV_X1 U711 ( .A(KEYINPUT99), .ZN(n600) );
  XNOR2_X1 U712 ( .A(n600), .B(n599), .ZN(n640) );
  INV_X1 U713 ( .A(n601), .ZN(n639) );
  INV_X1 U714 ( .A(n724), .ZN(n661) );
  XNOR2_X1 U715 ( .A(n602), .B(KEYINPUT66), .ZN(n603) );
  NAND2_X1 U716 ( .A1(n603), .A2(n623), .ZN(n662) );
  NOR2_X1 U717 ( .A1(n661), .A2(n604), .ZN(n605) );
  XOR2_X1 U718 ( .A(n687), .B(G140), .Z(G42) );
  NOR2_X1 U719 ( .A1(n608), .A2(n607), .ZN(n657) );
  INV_X1 U720 ( .A(n623), .ZN(n610) );
  INV_X1 U721 ( .A(n737), .ZN(n609) );
  NAND2_X1 U722 ( .A1(n610), .A2(n609), .ZN(n733) );
  INV_X1 U723 ( .A(n645), .ZN(n611) );
  XNOR2_X1 U724 ( .A(KEYINPUT105), .B(KEYINPUT33), .ZN(n613) );
  XNOR2_X1 U725 ( .A(n616), .B(n615), .ZN(n618) );
  XNOR2_X1 U726 ( .A(KEYINPUT81), .B(KEYINPUT35), .ZN(n619) );
  INV_X1 U727 ( .A(KEYINPUT103), .ZN(n622) );
  NAND2_X1 U728 ( .A1(n736), .A2(n645), .ZN(n624) );
  NOR2_X1 U729 ( .A1(n441), .A2(n624), .ZN(n625) );
  XNOR2_X1 U730 ( .A(KEYINPUT76), .B(n625), .ZN(n626) );
  NAND2_X1 U731 ( .A1(n621), .A2(n626), .ZN(n628) );
  INV_X1 U732 ( .A(KEYINPUT32), .ZN(n627) );
  XNOR2_X1 U733 ( .A(n628), .B(n627), .ZN(n803) );
  NAND2_X1 U734 ( .A1(n630), .A2(n631), .ZN(n633) );
  NOR2_X1 U735 ( .A1(n398), .A2(n635), .ZN(n715) );
  NAND2_X1 U736 ( .A1(n742), .A2(n637), .ZN(n638) );
  XNOR2_X1 U737 ( .A(n638), .B(KEYINPUT31), .ZN(n727) );
  NAND2_X1 U738 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X2 U739 ( .A(n642), .B(KEYINPUT101), .ZN(n750) );
  XNOR2_X1 U740 ( .A(KEYINPUT78), .B(n750), .ZN(n643) );
  INV_X1 U741 ( .A(n736), .ZN(n647) );
  INV_X1 U742 ( .A(KEYINPUT45), .ZN(n650) );
  NOR2_X1 U743 ( .A1(n404), .A2(G953), .ZN(n655) );
  NAND2_X1 U744 ( .A1(G953), .A2(G224), .ZN(n651) );
  XNOR2_X1 U745 ( .A(KEYINPUT61), .B(n651), .ZN(n652) );
  NAND2_X1 U746 ( .A1(n652), .A2(G898), .ZN(n653) );
  XOR2_X1 U747 ( .A(KEYINPUT124), .B(n653), .Z(n654) );
  NOR2_X1 U748 ( .A1(n655), .A2(n654), .ZN(n656) );
  XOR2_X1 U749 ( .A(n657), .B(n656), .Z(G69) );
  XNOR2_X1 U750 ( .A(n670), .B(KEYINPUT38), .ZN(n746) );
  NAND2_X1 U751 ( .A1(n658), .A2(n746), .ZN(n660) );
  XOR2_X1 U752 ( .A(n664), .B(KEYINPUT107), .Z(n665) );
  NAND2_X1 U753 ( .A1(n666), .A2(n665), .ZN(n672) );
  NAND2_X1 U754 ( .A1(n746), .A2(n745), .ZN(n751) );
  XNOR2_X1 U755 ( .A(n667), .B(KEYINPUT41), .ZN(n761) );
  XNOR2_X1 U756 ( .A(n668), .B(KEYINPUT42), .ZN(n802) );
  XNOR2_X1 U757 ( .A(KEYINPUT46), .B(KEYINPUT82), .ZN(n669) );
  INV_X1 U758 ( .A(n672), .ZN(n674) );
  NAND2_X1 U759 ( .A1(n674), .A2(n403), .ZN(n680) );
  INV_X1 U760 ( .A(n680), .ZN(n722) );
  NAND2_X1 U761 ( .A1(n750), .A2(n722), .ZN(n675) );
  NAND2_X1 U762 ( .A1(n675), .A2(KEYINPUT47), .ZN(n677) );
  NAND2_X1 U763 ( .A1(n677), .A2(n676), .ZN(n683) );
  NOR2_X1 U764 ( .A1(KEYINPUT78), .A2(n750), .ZN(n679) );
  NAND2_X1 U765 ( .A1(n750), .A2(KEYINPUT78), .ZN(n678) );
  NOR2_X1 U766 ( .A1(n681), .A2(n680), .ZN(n682) );
  NOR2_X1 U767 ( .A1(n683), .A2(n682), .ZN(n684) );
  INV_X1 U768 ( .A(n726), .ZN(n686) );
  NOR2_X1 U769 ( .A1(n686), .A2(n685), .ZN(n732) );
  INV_X1 U770 ( .A(KEYINPUT79), .ZN(n688) );
  NAND2_X1 U771 ( .A1(KEYINPUT2), .A2(KEYINPUT80), .ZN(n690) );
  INV_X1 U772 ( .A(KEYINPUT2), .ZN(n692) );
  NOR2_X1 U773 ( .A1(KEYINPUT80), .A2(n692), .ZN(n693) );
  OR2_X1 U774 ( .A1(n693), .A2(KEYINPUT79), .ZN(n694) );
  INV_X1 U775 ( .A(n764), .ZN(n698) );
  NAND2_X1 U776 ( .A1(n698), .A2(KEYINPUT2), .ZN(n700) );
  INV_X1 U777 ( .A(KEYINPUT72), .ZN(n699) );
  NAND2_X1 U778 ( .A1(n781), .A2(G210), .ZN(n706) );
  XOR2_X1 U779 ( .A(KEYINPUT77), .B(KEYINPUT54), .Z(n702) );
  XNOR2_X1 U780 ( .A(n702), .B(KEYINPUT55), .ZN(n703) );
  XNOR2_X1 U781 ( .A(n704), .B(n703), .ZN(n705) );
  XNOR2_X1 U782 ( .A(n706), .B(n705), .ZN(n708) );
  INV_X1 U783 ( .A(G952), .ZN(n707) );
  XOR2_X1 U784 ( .A(KEYINPUT119), .B(KEYINPUT56), .Z(n709) );
  XNOR2_X1 U785 ( .A(n710), .B(n709), .ZN(G51) );
  XOR2_X1 U786 ( .A(n712), .B(G101), .Z(G3) );
  NAND2_X1 U787 ( .A1(n715), .A2(n724), .ZN(n713) );
  XNOR2_X1 U788 ( .A(n713), .B(KEYINPUT108), .ZN(n714) );
  XNOR2_X1 U789 ( .A(G104), .B(n714), .ZN(G6) );
  XOR2_X1 U790 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n717) );
  NAND2_X1 U791 ( .A1(n715), .A2(n726), .ZN(n716) );
  XNOR2_X1 U792 ( .A(n717), .B(n716), .ZN(n718) );
  XNOR2_X1 U793 ( .A(G107), .B(n718), .ZN(G9) );
  XOR2_X1 U794 ( .A(KEYINPUT29), .B(KEYINPUT110), .Z(n720) );
  NAND2_X1 U795 ( .A1(n722), .A2(n726), .ZN(n719) );
  XNOR2_X1 U796 ( .A(n720), .B(n719), .ZN(n721) );
  XNOR2_X1 U797 ( .A(G128), .B(n721), .ZN(G30) );
  NAND2_X1 U798 ( .A1(n722), .A2(n724), .ZN(n723) );
  XNOR2_X1 U799 ( .A(n723), .B(G146), .ZN(G48) );
  NAND2_X1 U800 ( .A1(n727), .A2(n724), .ZN(n725) );
  XNOR2_X1 U801 ( .A(n725), .B(G113), .ZN(G15) );
  XOR2_X1 U802 ( .A(G116), .B(KEYINPUT111), .Z(n729) );
  NAND2_X1 U803 ( .A1(n727), .A2(n726), .ZN(n728) );
  XNOR2_X1 U804 ( .A(n729), .B(n728), .ZN(G18) );
  XNOR2_X1 U805 ( .A(n730), .B(G125), .ZN(n731) );
  XNOR2_X1 U806 ( .A(n731), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U807 ( .A(G134), .B(n732), .Z(G36) );
  NAND2_X1 U808 ( .A1(n441), .A2(n733), .ZN(n735) );
  XOR2_X1 U809 ( .A(KEYINPUT50), .B(n735), .Z(n740) );
  NOR2_X1 U810 ( .A1(n740), .A2(n739), .ZN(n741) );
  NOR2_X1 U811 ( .A1(n761), .A2(n743), .ZN(n758) );
  BUF_X1 U812 ( .A(n744), .Z(n762) );
  NOR2_X1 U813 ( .A1(n746), .A2(n745), .ZN(n747) );
  XOR2_X1 U814 ( .A(KEYINPUT115), .B(n747), .Z(n748) );
  NOR2_X1 U815 ( .A1(n749), .A2(n748), .ZN(n754) );
  INV_X1 U816 ( .A(n750), .ZN(n752) );
  NOR2_X1 U817 ( .A1(n752), .A2(n751), .ZN(n753) );
  NOR2_X1 U818 ( .A1(n754), .A2(n753), .ZN(n755) );
  NOR2_X1 U819 ( .A1(n762), .A2(n755), .ZN(n756) );
  XNOR2_X1 U820 ( .A(n756), .B(KEYINPUT116), .ZN(n757) );
  NOR2_X1 U821 ( .A1(n758), .A2(n757), .ZN(n759) );
  OR2_X1 U822 ( .A1(n762), .A2(n761), .ZN(n763) );
  NOR2_X1 U823 ( .A1(n698), .A2(KEYINPUT2), .ZN(n765) );
  NOR2_X1 U824 ( .A1(n766), .A2(n765), .ZN(n767) );
  NAND2_X1 U825 ( .A1(n785), .A2(G469), .ZN(n774) );
  XOR2_X1 U826 ( .A(KEYINPUT58), .B(KEYINPUT57), .Z(n771) );
  XNOR2_X1 U827 ( .A(KEYINPUT121), .B(KEYINPUT120), .ZN(n770) );
  XNOR2_X1 U828 ( .A(n771), .B(n770), .ZN(n772) );
  XOR2_X1 U829 ( .A(n769), .B(n772), .Z(n773) );
  XNOR2_X1 U830 ( .A(n774), .B(n773), .ZN(n775) );
  NOR2_X1 U831 ( .A1(n789), .A2(n775), .ZN(G54) );
  NAND2_X1 U832 ( .A1(n781), .A2(G475), .ZN(n778) );
  XOR2_X1 U833 ( .A(n776), .B(KEYINPUT59), .Z(n777) );
  XNOR2_X1 U834 ( .A(n778), .B(n777), .ZN(n779) );
  XNOR2_X1 U835 ( .A(n780), .B(KEYINPUT60), .ZN(G60) );
  XNOR2_X1 U836 ( .A(n782), .B(KEYINPUT122), .ZN(n783) );
  XOR2_X1 U837 ( .A(KEYINPUT123), .B(n784), .Z(G63) );
  NAND2_X1 U838 ( .A1(n785), .A2(G217), .ZN(n786) );
  XNOR2_X1 U839 ( .A(n787), .B(n786), .ZN(n788) );
  NOR2_X1 U840 ( .A1(n789), .A2(n788), .ZN(G66) );
  XOR2_X1 U841 ( .A(n791), .B(n790), .Z(n795) );
  XOR2_X1 U842 ( .A(n792), .B(n795), .Z(n794) );
  NAND2_X1 U843 ( .A1(n794), .A2(n793), .ZN(n800) );
  XNOR2_X1 U844 ( .A(n795), .B(G227), .ZN(n796) );
  XNOR2_X1 U845 ( .A(n796), .B(KEYINPUT125), .ZN(n797) );
  NAND2_X1 U846 ( .A1(n797), .A2(G900), .ZN(n798) );
  NAND2_X1 U847 ( .A1(G953), .A2(n798), .ZN(n799) );
  NAND2_X1 U848 ( .A1(n800), .A2(n799), .ZN(G72) );
  XOR2_X1 U849 ( .A(G137), .B(KEYINPUT126), .Z(n801) );
  XNOR2_X1 U850 ( .A(n802), .B(n801), .ZN(G39) );
  XOR2_X1 U851 ( .A(G119), .B(n803), .Z(G21) );
  XNOR2_X1 U852 ( .A(G131), .B(KEYINPUT127), .ZN(n805) );
  XNOR2_X1 U853 ( .A(n805), .B(n804), .ZN(G33) );
endmodule

