//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 1 0 0 0 0 1 1 1 1 0 1 0 1 1 1 1 0 1 1 1 0 0 0 0 0 0 1 1 0 0 0 1 1 0 1 1 0 0 0 1 0 0 0 0 1 1 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:13 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n233, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1286, new_n1287, new_n1288, new_n1289, new_n1291,
    new_n1292, new_n1293, new_n1294, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355, new_n1356, new_n1357, new_n1358, new_n1359,
    new_n1360, new_n1361, new_n1362, new_n1363, new_n1364, new_n1365,
    new_n1366, new_n1367, new_n1368, new_n1369;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  NOR2_X1   g0001(.A1(G97), .A2(G107), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n203), .A2(G87), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT64), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  AND2_X1   g0009(.A1(new_n209), .A2(KEYINPUT65), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(KEYINPUT65), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G68), .A2(G238), .B1(G107), .B2(G264), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G50), .A2(G226), .B1(G87), .B2(G250), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n206), .B1(new_n214), .B2(new_n217), .ZN(new_n218));
  XNOR2_X1  g0018(.A(new_n218), .B(KEYINPUT1), .ZN(new_n219));
  OAI21_X1  g0019(.A(G50), .B1(G58), .B2(G68), .ZN(new_n220));
  INV_X1    g0020(.A(G20), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G13), .ZN(new_n222));
  NOR3_X1   g0022(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  NOR4_X1   g0023(.A1(new_n210), .A2(new_n211), .A3(new_n219), .A4(new_n223), .ZN(G361));
  XNOR2_X1  g0024(.A(G238), .B(G244), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(G232), .ZN(new_n226));
  XNOR2_X1  g0026(.A(KEYINPUT2), .B(G226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XOR2_X1   g0028(.A(G264), .B(G270), .Z(new_n229));
  XNOR2_X1  g0029(.A(G250), .B(G257), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n228), .B(new_n231), .ZN(G358));
  XOR2_X1   g0032(.A(G87), .B(G97), .Z(new_n233));
  XOR2_X1   g0033(.A(G107), .B(G116), .Z(new_n234));
  XOR2_X1   g0034(.A(new_n233), .B(new_n234), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT66), .ZN(new_n236));
  XOR2_X1   g0036(.A(G58), .B(G77), .Z(new_n237));
  XNOR2_X1  g0037(.A(G50), .B(G68), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G351));
  INV_X1    g0040(.A(G1698), .ZN(new_n241));
  AND2_X1   g0041(.A1(KEYINPUT3), .A2(G33), .ZN(new_n242));
  NOR2_X1   g0042(.A1(KEYINPUT3), .A2(G33), .ZN(new_n243));
  OAI211_X1 g0043(.A(G222), .B(new_n241), .C1(new_n242), .C2(new_n243), .ZN(new_n244));
  OAI211_X1 g0044(.A(G223), .B(G1698), .C1(new_n242), .C2(new_n243), .ZN(new_n245));
  INV_X1    g0045(.A(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(KEYINPUT3), .B(G33), .ZN(new_n247));
  OAI211_X1 g0047(.A(new_n244), .B(new_n245), .C1(new_n246), .C2(new_n247), .ZN(new_n248));
  AND2_X1   g0048(.A1(G33), .A2(G41), .ZN(new_n249));
  NOR2_X1   g0049(.A1(new_n249), .A2(new_n222), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  OAI21_X1  g0051(.A(G274), .B1(new_n249), .B2(new_n222), .ZN(new_n252));
  INV_X1    g0052(.A(G1), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n253), .B1(G41), .B2(G45), .ZN(new_n254));
  OAI21_X1  g0054(.A(KEYINPUT67), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G274), .ZN(new_n256));
  AND2_X1   g0056(.A1(G1), .A2(G13), .ZN(new_n257));
  NAND2_X1  g0057(.A1(G33), .A2(G41), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n256), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT67), .ZN(new_n260));
  INV_X1    g0060(.A(G41), .ZN(new_n261));
  INV_X1    g0061(.A(G45), .ZN(new_n262));
  AOI21_X1  g0062(.A(G1), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n259), .A2(new_n260), .A3(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n255), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n258), .A2(G1), .A3(G13), .ZN(new_n266));
  AND3_X1   g0066(.A1(new_n266), .A2(KEYINPUT68), .A3(new_n254), .ZN(new_n267));
  AOI21_X1  g0067(.A(KEYINPUT68), .B1(new_n266), .B2(new_n254), .ZN(new_n268));
  OAI21_X1  g0068(.A(G226), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n251), .A2(new_n265), .A3(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT69), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND4_X1  g0072(.A1(new_n251), .A2(KEYINPUT69), .A3(new_n265), .A4(new_n269), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G179), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(new_n222), .ZN(new_n278));
  XNOR2_X1  g0078(.A(KEYINPUT8), .B(G58), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n221), .A2(G33), .ZN(new_n280));
  INV_X1    g0080(.A(G150), .ZN(new_n281));
  NOR2_X1   g0081(.A1(G20), .A2(G33), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  OAI22_X1  g0083(.A1(new_n279), .A2(new_n280), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  NOR2_X1   g0084(.A1(G58), .A2(G68), .ZN(new_n285));
  INV_X1    g0085(.A(G50), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n221), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n278), .B1(new_n284), .B2(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n253), .A2(G13), .A3(G20), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT70), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND4_X1  g0091(.A1(new_n253), .A2(KEYINPUT70), .A3(G13), .A4(G20), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(new_n286), .ZN(new_n295));
  INV_X1    g0095(.A(new_n278), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n253), .A2(G20), .ZN(new_n297));
  NAND4_X1  g0097(.A1(new_n293), .A2(G50), .A3(new_n296), .A4(new_n297), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n288), .A2(new_n295), .A3(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G169), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n272), .A2(new_n300), .A3(new_n273), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n276), .A2(new_n299), .A3(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n272), .A2(G200), .A3(new_n273), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n299), .A2(KEYINPUT9), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT9), .ZN(new_n306));
  NAND4_X1  g0106(.A1(new_n288), .A2(new_n295), .A3(new_n306), .A4(new_n298), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  AND2_X1   g0108(.A1(new_n304), .A2(new_n308), .ZN(new_n309));
  AOI21_X1  g0109(.A(KEYINPUT71), .B1(new_n274), .B2(G190), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT71), .ZN(new_n311));
  INV_X1    g0111(.A(G190), .ZN(new_n312));
  AOI211_X1 g0112(.A(new_n311), .B(new_n312), .C1(new_n272), .C2(new_n273), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n309), .B1(new_n310), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(KEYINPUT10), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT10), .ZN(new_n316));
  OAI211_X1 g0116(.A(new_n309), .B(new_n316), .C1(new_n310), .C2(new_n313), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n303), .B1(new_n315), .B2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(G68), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n294), .A2(new_n319), .ZN(new_n320));
  XNOR2_X1  g0120(.A(new_n320), .B(KEYINPUT12), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n283), .A2(new_n286), .ZN(new_n322));
  OAI22_X1  g0122(.A1(new_n280), .A2(new_n246), .B1(new_n221), .B2(G68), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n278), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  XNOR2_X1  g0124(.A(new_n324), .B(KEYINPUT11), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n294), .A2(new_n278), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n326), .A2(G68), .A3(new_n297), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n321), .A2(new_n325), .A3(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  OAI21_X1  g0129(.A(G238), .B1(new_n267), .B2(new_n268), .ZN(new_n330));
  NAND2_X1  g0130(.A1(G33), .A2(G97), .ZN(new_n331));
  INV_X1    g0131(.A(G232), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(G1698), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n333), .B1(G226), .B2(G1698), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n242), .A2(new_n243), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n331), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(new_n250), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n330), .A2(new_n265), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(KEYINPUT13), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT13), .ZN(new_n340));
  NAND4_X1  g0140(.A1(new_n265), .A2(new_n330), .A3(new_n337), .A4(new_n340), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n339), .A2(G179), .A3(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT72), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n339), .A2(new_n344), .A3(new_n341), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n338), .A2(KEYINPUT72), .A3(KEYINPUT13), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n345), .A2(G169), .A3(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n343), .B1(new_n347), .B2(KEYINPUT14), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT14), .ZN(new_n349));
  NAND4_X1  g0149(.A1(new_n345), .A2(new_n349), .A3(G169), .A4(new_n346), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n329), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n339), .A2(G190), .A3(new_n341), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n329), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n345), .A2(G200), .A3(new_n346), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT73), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND4_X1  g0156(.A1(new_n345), .A2(KEYINPUT73), .A3(G200), .A4(new_n346), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n353), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n351), .A2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(G58), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(KEYINPUT8), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT8), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(G58), .ZN(new_n363));
  AOI22_X1  g0163(.A1(new_n361), .A2(new_n363), .B1(new_n253), .B2(G20), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n293), .A2(new_n296), .A3(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n291), .A2(new_n279), .A3(new_n292), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT75), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n365), .A2(KEYINPUT75), .A3(new_n366), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT16), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT3), .ZN(new_n373));
  INV_X1    g0173(.A(G33), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(KEYINPUT3), .A2(G33), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n375), .A2(new_n221), .A3(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT7), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND4_X1  g0179(.A1(new_n375), .A2(KEYINPUT7), .A3(new_n221), .A4(new_n376), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n319), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n360), .A2(new_n319), .ZN(new_n382));
  OAI21_X1  g0182(.A(G20), .B1(new_n382), .B2(new_n285), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n282), .A2(G159), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n372), .B1(new_n381), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(new_n278), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n383), .A2(KEYINPUT16), .A3(new_n384), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n380), .A2(KEYINPUT74), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT74), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n335), .A2(new_n390), .A3(KEYINPUT7), .A4(new_n221), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n389), .A2(new_n391), .A3(new_n379), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n388), .B1(new_n392), .B2(G68), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n371), .B1(new_n387), .B2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT76), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n250), .A2(new_n263), .ZN(new_n396));
  AOI22_X1  g0196(.A1(new_n255), .A2(new_n264), .B1(new_n396), .B2(G232), .ZN(new_n397));
  OAI211_X1 g0197(.A(G223), .B(new_n241), .C1(new_n242), .C2(new_n243), .ZN(new_n398));
  OAI211_X1 g0198(.A(G226), .B(G1698), .C1(new_n242), .C2(new_n243), .ZN(new_n399));
  NAND2_X1  g0199(.A1(G33), .A2(G87), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n398), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(new_n250), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n397), .A2(G179), .A3(new_n402), .ZN(new_n403));
  AND2_X1   g0203(.A1(new_n397), .A2(new_n402), .ZN(new_n404));
  OAI211_X1 g0204(.A(new_n395), .B(new_n403), .C1(new_n404), .C2(new_n300), .ZN(new_n405));
  AND3_X1   g0205(.A1(new_n397), .A2(G179), .A3(new_n402), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n300), .B1(new_n397), .B2(new_n402), .ZN(new_n407));
  OAI21_X1  g0207(.A(KEYINPUT76), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n394), .A2(new_n405), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(KEYINPUT18), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT18), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n394), .A2(new_n405), .A3(new_n408), .A4(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT17), .ZN(new_n414));
  AND3_X1   g0214(.A1(new_n397), .A2(new_n312), .A3(new_n402), .ZN(new_n415));
  AOI21_X1  g0215(.A(G200), .B1(new_n397), .B2(new_n402), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  OAI21_X1  g0217(.A(KEYINPUT77), .B1(new_n394), .B2(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n397), .A2(new_n312), .A3(new_n402), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n419), .B1(new_n404), .B2(G200), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n392), .A2(G68), .ZN(new_n421));
  INV_X1    g0221(.A(new_n388), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n423), .A2(new_n278), .A3(new_n386), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT77), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n420), .A2(new_n424), .A3(new_n425), .A4(new_n371), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n414), .B1(new_n418), .B2(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(KEYINPUT7), .B1(new_n335), .B2(new_n221), .ZN(new_n428));
  INV_X1    g0228(.A(new_n380), .ZN(new_n429));
  OAI21_X1  g0229(.A(G68), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(new_n385), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n296), .B1(new_n432), .B2(new_n372), .ZN(new_n433));
  AOI22_X1  g0233(.A1(new_n433), .A2(new_n423), .B1(new_n369), .B2(new_n370), .ZN(new_n434));
  AOI21_X1  g0234(.A(KEYINPUT17), .B1(new_n434), .B2(new_n420), .ZN(new_n435));
  NOR3_X1   g0235(.A1(new_n413), .A2(new_n427), .A3(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n279), .ZN(new_n437));
  AOI22_X1  g0237(.A1(new_n437), .A2(new_n282), .B1(G20), .B2(G77), .ZN(new_n438));
  XNOR2_X1  g0238(.A(KEYINPUT15), .B(G87), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n438), .B1(new_n280), .B2(new_n439), .ZN(new_n440));
  AOI22_X1  g0240(.A1(new_n440), .A2(new_n278), .B1(new_n246), .B2(new_n294), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n326), .A2(G77), .A3(new_n297), .ZN(new_n442));
  AND2_X1   g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n247), .A2(G232), .A3(new_n241), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n247), .A2(G238), .A3(G1698), .ZN(new_n445));
  INV_X1    g0245(.A(G107), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n444), .B(new_n445), .C1(new_n446), .C2(new_n247), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(new_n250), .ZN(new_n448));
  OAI21_X1  g0248(.A(G244), .B1(new_n267), .B2(new_n268), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n448), .A2(new_n265), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(G200), .ZN(new_n451));
  OAI211_X1 g0251(.A(new_n443), .B(new_n451), .C1(new_n312), .C2(new_n450), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n450), .A2(new_n300), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n441), .A2(new_n442), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n453), .B(new_n454), .C1(G179), .C2(new_n450), .ZN(new_n455));
  AND2_X1   g0255(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n318), .A2(new_n359), .A3(new_n436), .A4(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(KEYINPUT78), .ZN(new_n458));
  INV_X1    g0258(.A(new_n413), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n418), .A2(new_n426), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n435), .B1(new_n460), .B2(KEYINPUT17), .ZN(new_n461));
  AND3_X1   g0261(.A1(new_n459), .A2(new_n461), .A3(new_n456), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT78), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n462), .A2(new_n463), .A3(new_n359), .A4(new_n318), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n458), .A2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(G97), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n293), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n253), .A2(G33), .ZN(new_n468));
  AND3_X1   g0268(.A1(new_n293), .A2(new_n296), .A3(new_n468), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n467), .B1(new_n469), .B2(new_n466), .ZN(new_n470));
  OAI21_X1  g0270(.A(G107), .B1(new_n428), .B2(new_n429), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT6), .ZN(new_n472));
  AND2_X1   g0272(.A1(G97), .A2(G107), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n472), .B1(new_n473), .B2(new_n202), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n446), .A2(KEYINPUT6), .A3(G97), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  AOI22_X1  g0276(.A1(new_n476), .A2(G20), .B1(G77), .B2(new_n282), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n296), .B1(new_n471), .B2(new_n477), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n478), .A2(KEYINPUT79), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT79), .ZN(new_n480));
  AOI211_X1 g0280(.A(new_n480), .B(new_n296), .C1(new_n471), .C2(new_n477), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n470), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT80), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT5), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n483), .B1(new_n484), .B2(G41), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n261), .A2(KEYINPUT80), .A3(KEYINPUT5), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n262), .A2(G1), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n484), .A2(G41), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n485), .A2(new_n486), .A3(new_n487), .A4(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n489), .A2(G257), .A3(new_n266), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n253), .B(G45), .C1(new_n261), .C2(KEYINPUT5), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n492), .A2(new_n259), .A3(new_n486), .A4(new_n485), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  OAI211_X1 g0294(.A(G244), .B(new_n241), .C1(new_n242), .C2(new_n243), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT4), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(G33), .A2(G283), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(G250), .A2(G1698), .ZN(new_n500));
  NAND2_X1  g0300(.A1(KEYINPUT4), .A2(G244), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n500), .B1(new_n501), .B2(G1698), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n499), .B1(new_n247), .B2(new_n502), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n266), .B1(new_n497), .B2(new_n503), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n494), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(new_n275), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n300), .B1(new_n494), .B2(new_n504), .ZN(new_n507));
  AND2_X1   g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n482), .A2(new_n508), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n221), .B(G87), .C1(new_n242), .C2(new_n243), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT83), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n511), .A2(KEYINPUT22), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n247), .A2(new_n221), .A3(G87), .A4(new_n512), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n511), .A2(KEYINPUT22), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT23), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n518), .B1(new_n221), .B2(G107), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n446), .A2(KEYINPUT23), .A3(G20), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(G33), .A2(G116), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n521), .B1(G20), .B2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n517), .A2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT84), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT24), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n525), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(new_n516), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n529), .B1(new_n510), .B2(new_n513), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n523), .B1(new_n530), .B2(new_n515), .ZN(new_n531));
  OAI21_X1  g0331(.A(KEYINPUT24), .B1(new_n531), .B2(KEYINPUT84), .ZN(new_n532));
  AND3_X1   g0332(.A1(new_n517), .A2(KEYINPUT84), .A3(new_n524), .ZN(new_n533));
  OAI211_X1 g0333(.A(new_n278), .B(new_n528), .C1(new_n532), .C2(new_n533), .ZN(new_n534));
  XOR2_X1   g0334(.A(KEYINPUT85), .B(KEYINPUT25), .Z(new_n535));
  NAND3_X1  g0335(.A1(new_n294), .A2(new_n446), .A3(new_n535), .ZN(new_n536));
  OAI211_X1 g0336(.A(KEYINPUT85), .B(KEYINPUT25), .C1(new_n293), .C2(G107), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n538), .B1(G107), .B2(new_n469), .ZN(new_n539));
  OAI211_X1 g0339(.A(G257), .B(G1698), .C1(new_n242), .C2(new_n243), .ZN(new_n540));
  OAI211_X1 g0340(.A(G250), .B(new_n241), .C1(new_n242), .C2(new_n243), .ZN(new_n541));
  NAND2_X1  g0341(.A1(G33), .A2(G294), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(new_n250), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n489), .A2(G264), .A3(new_n266), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n544), .A2(new_n493), .A3(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(G200), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n548), .B1(G190), .B2(new_n546), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n534), .A2(new_n539), .A3(new_n549), .ZN(new_n550));
  OAI211_X1 g0350(.A(G244), .B(G1698), .C1(new_n242), .C2(new_n243), .ZN(new_n551));
  OAI211_X1 g0351(.A(G238), .B(new_n241), .C1(new_n242), .C2(new_n243), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n551), .A2(new_n552), .A3(new_n522), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(new_n250), .ZN(new_n554));
  INV_X1    g0354(.A(G250), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n555), .B1(new_n262), .B2(G1), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n253), .A2(new_n256), .A3(G45), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n266), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(KEYINPUT81), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT81), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n266), .A2(new_n556), .A3(new_n557), .A4(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n554), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(G200), .ZN(new_n564));
  AOI22_X1  g0364(.A1(new_n250), .A2(new_n553), .B1(new_n559), .B2(new_n561), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(G190), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n247), .A2(new_n221), .A3(G68), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT19), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n221), .B1(new_n331), .B2(new_n568), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n569), .B1(G87), .B2(new_n203), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n221), .A2(G33), .A3(G97), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT82), .ZN(new_n572));
  AND3_X1   g0372(.A1(new_n571), .A2(new_n572), .A3(new_n568), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n572), .B1(new_n571), .B2(new_n568), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n567), .B(new_n570), .C1(new_n573), .C2(new_n574), .ZN(new_n575));
  AOI22_X1  g0375(.A1(new_n575), .A2(new_n278), .B1(new_n294), .B2(new_n439), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n469), .A2(G87), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n564), .A2(new_n566), .A3(new_n576), .A4(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n575), .A2(new_n278), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n294), .A2(new_n439), .ZN(new_n580));
  INV_X1    g0380(.A(new_n439), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n293), .A2(new_n296), .A3(new_n581), .A4(new_n468), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n579), .A2(new_n580), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n563), .A2(new_n300), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n565), .A2(new_n275), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  AND2_X1   g0386(.A1(new_n578), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n476), .A2(G20), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n282), .A2(G77), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n446), .B1(new_n379), .B2(new_n380), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n278), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n480), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n478), .A2(KEYINPUT79), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  AND2_X1   g0395(.A1(new_n490), .A2(new_n493), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n497), .A2(new_n503), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n250), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n596), .A2(new_n598), .A3(new_n312), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n599), .B1(new_n505), .B2(G200), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n595), .A2(new_n470), .A3(new_n600), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n509), .A2(new_n550), .A3(new_n587), .A4(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n534), .A2(new_n539), .ZN(new_n603));
  AOI21_X1  g0403(.A(KEYINPUT80), .B1(new_n261), .B2(KEYINPUT5), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n491), .A2(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n250), .B1(new_n605), .B2(new_n486), .ZN(new_n606));
  AOI22_X1  g0406(.A1(new_n606), .A2(G264), .B1(new_n543), .B2(new_n250), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT86), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n607), .A2(new_n608), .A3(G179), .A4(new_n493), .ZN(new_n609));
  AOI21_X1  g0409(.A(KEYINPUT86), .B1(new_n546), .B2(G169), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n546), .A2(new_n275), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n609), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n603), .A2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT21), .ZN(new_n614));
  OAI211_X1 g0414(.A(G264), .B(G1698), .C1(new_n242), .C2(new_n243), .ZN(new_n615));
  OAI211_X1 g0415(.A(G257), .B(new_n241), .C1(new_n242), .C2(new_n243), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n375), .A2(G303), .A3(new_n376), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n615), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  AND2_X1   g0418(.A1(new_n618), .A2(new_n250), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n489), .A2(G270), .A3(new_n266), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(new_n493), .ZN(new_n621));
  OAI21_X1  g0421(.A(G169), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n293), .A2(G116), .A3(new_n296), .A4(new_n468), .ZN(new_n623));
  INV_X1    g0423(.A(G116), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n291), .A2(new_n624), .A3(new_n292), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  AOI22_X1  g0426(.A1(new_n277), .A2(new_n222), .B1(G20), .B2(new_n624), .ZN(new_n627));
  OAI211_X1 g0427(.A(new_n498), .B(new_n221), .C1(G33), .C2(new_n466), .ZN(new_n628));
  AND3_X1   g0428(.A1(new_n627), .A2(KEYINPUT20), .A3(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(KEYINPUT20), .B1(new_n627), .B2(new_n628), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n626), .A2(new_n631), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n614), .B1(new_n622), .B2(new_n632), .ZN(new_n633));
  OAI211_X1 g0433(.A(new_n623), .B(new_n625), .C1(new_n630), .C2(new_n629), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n618), .A2(new_n250), .ZN(new_n635));
  INV_X1    g0435(.A(new_n621), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n634), .A2(G179), .A3(new_n635), .A4(new_n636), .ZN(new_n637));
  OAI21_X1  g0437(.A(G200), .B1(new_n619), .B2(new_n621), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n635), .A2(G190), .A3(new_n493), .A4(new_n620), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n638), .A2(new_n632), .A3(new_n639), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n635), .A2(new_n493), .A3(new_n620), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n634), .A2(new_n641), .A3(KEYINPUT21), .A4(G169), .ZN(new_n642));
  AND4_X1   g0442(.A1(new_n633), .A2(new_n637), .A3(new_n640), .A4(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n613), .A2(new_n643), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n602), .A2(new_n644), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n465), .A2(new_n645), .ZN(G372));
  OAI21_X1  g0446(.A(new_n506), .B1(new_n505), .B2(G169), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n647), .B1(new_n595), .B2(new_n470), .ZN(new_n648));
  XOR2_X1   g0448(.A(KEYINPUT88), .B(KEYINPUT26), .Z(new_n649));
  NAND3_X1  g0449(.A1(new_n648), .A2(new_n587), .A3(new_n649), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n482), .A2(new_n508), .A3(new_n586), .A4(new_n578), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(KEYINPUT26), .ZN(new_n652));
  XNOR2_X1  g0452(.A(new_n586), .B(KEYINPUT87), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n650), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n633), .A2(new_n637), .A3(new_n642), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n655), .B1(new_n603), .B2(new_n612), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n602), .A2(new_n656), .ZN(new_n657));
  OR2_X1    g0457(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n465), .A2(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n403), .B1(new_n404), .B2(new_n300), .ZN(new_n660));
  AND3_X1   g0460(.A1(new_n394), .A2(new_n411), .A3(new_n660), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n411), .B1(new_n394), .B2(new_n660), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n347), .A2(KEYINPUT14), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n665), .A2(new_n350), .A3(new_n342), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(new_n328), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n667), .B1(new_n358), .B2(new_n455), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n664), .B1(new_n668), .B2(new_n461), .ZN(new_n669));
  AND2_X1   g0469(.A1(new_n314), .A2(KEYINPUT10), .ZN(new_n670));
  INV_X1    g0470(.A(new_n317), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n302), .B1(new_n669), .B2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n659), .A2(new_n674), .ZN(G369));
  AND2_X1   g0475(.A1(new_n603), .A2(new_n612), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n253), .A2(new_n221), .A3(G13), .ZN(new_n677));
  OR2_X1    g0477(.A1(new_n677), .A2(KEYINPUT27), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(KEYINPUT27), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n678), .A2(G213), .A3(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(G343), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n603), .A2(new_n682), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n676), .B1(new_n550), .B2(new_n683), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n613), .A2(new_n682), .ZN(new_n685));
  OAI21_X1  g0485(.A(KEYINPUT89), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n683), .A2(new_n550), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(new_n613), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT89), .ZN(new_n689));
  INV_X1    g0489(.A(new_n682), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n676), .A2(new_n690), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n688), .A2(new_n689), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n655), .A2(new_n690), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n686), .A2(new_n692), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(new_n691), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n686), .A2(new_n692), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n632), .A2(new_n690), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n655), .A2(new_n698), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n633), .A2(new_n640), .A3(new_n637), .A4(new_n642), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n699), .B1(new_n700), .B2(new_n698), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(G330), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n697), .A2(new_n702), .ZN(new_n703));
  OR2_X1    g0503(.A1(new_n696), .A2(new_n703), .ZN(G399));
  INV_X1    g0504(.A(new_n207), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(G41), .ZN(new_n706));
  INV_X1    g0506(.A(G87), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n202), .A2(new_n707), .A3(new_n624), .ZN(new_n708));
  NOR3_X1   g0508(.A1(new_n706), .A2(new_n253), .A3(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n220), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n709), .B1(new_n710), .B2(new_n706), .ZN(new_n711));
  XOR2_X1   g0511(.A(new_n711), .B(KEYINPUT28), .Z(new_n712));
  INV_X1    g0512(.A(KEYINPUT29), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n658), .A2(new_n713), .A3(new_n690), .ZN(new_n714));
  INV_X1    g0514(.A(new_n649), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n651), .A2(new_n715), .ZN(new_n716));
  OAI211_X1 g0516(.A(new_n716), .B(new_n653), .C1(KEYINPUT26), .C2(new_n651), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n717), .A2(new_n657), .ZN(new_n718));
  OAI21_X1  g0518(.A(KEYINPUT29), .B1(new_n718), .B2(new_n682), .ZN(new_n719));
  AND3_X1   g0519(.A1(new_n509), .A2(new_n601), .A3(new_n587), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n700), .B1(new_n603), .B2(new_n612), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n720), .A2(new_n721), .A3(new_n550), .A4(new_n690), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT30), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n607), .A2(new_n565), .A3(new_n596), .A4(new_n598), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n635), .A2(G179), .A3(new_n493), .A4(new_n620), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n723), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(KEYINPUT91), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n641), .A2(new_n275), .A3(new_n563), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(KEYINPUT90), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT90), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n641), .A2(new_n563), .A3(new_n730), .A4(new_n275), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n505), .B1(new_n493), .B2(new_n607), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n729), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  OR3_X1    g0533(.A1(new_n724), .A2(new_n723), .A3(new_n725), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT91), .ZN(new_n735));
  OAI211_X1 g0535(.A(new_n735), .B(new_n723), .C1(new_n724), .C2(new_n725), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n727), .A2(new_n733), .A3(new_n734), .A4(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(new_n682), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT31), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n733), .A2(new_n734), .A3(new_n726), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n741), .A2(KEYINPUT31), .A3(new_n682), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n722), .A2(new_n740), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(G330), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n714), .A2(new_n719), .A3(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n712), .B1(new_n746), .B2(G1), .ZN(G364));
  INV_X1    g0547(.A(new_n702), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n221), .A2(G13), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n253), .B1(new_n750), .B2(G45), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n706), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n748), .A2(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n754), .B1(G330), .B2(new_n701), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n207), .A2(G355), .A3(new_n247), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n756), .B1(G116), .B2(new_n207), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n207), .A2(new_n335), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n758), .B1(new_n262), .B2(new_n710), .ZN(new_n759));
  OR2_X1    g0559(.A1(new_n239), .A2(new_n262), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n757), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(G13), .A2(G33), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(G20), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n222), .B1(G20), .B2(new_n300), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n753), .B1(new_n761), .B2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n221), .A2(new_n275), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n769), .A2(new_n312), .A3(G200), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  XNOR2_X1  g0571(.A(KEYINPUT33), .B(G317), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n769), .A2(G190), .A3(new_n547), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  AOI22_X1  g0574(.A1(new_n771), .A2(new_n772), .B1(new_n774), .B2(G322), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  OR2_X1    g0576(.A1(new_n776), .A2(KEYINPUT94), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n769), .A2(G190), .A3(G200), .ZN(new_n778));
  INV_X1    g0578(.A(KEYINPUT92), .ZN(new_n779));
  AND2_X1   g0579(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n778), .A2(new_n779), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n221), .A2(G179), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n784), .A2(G190), .A3(G200), .ZN(new_n785));
  XOR2_X1   g0585(.A(new_n785), .B(KEYINPUT93), .Z(new_n786));
  AOI22_X1  g0586(.A1(new_n783), .A2(G326), .B1(G303), .B2(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(G190), .A2(G200), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n769), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(G311), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n335), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NOR3_X1   g0591(.A1(new_n312), .A2(G179), .A3(G200), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(new_n221), .ZN(new_n793));
  INV_X1    g0593(.A(G294), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n784), .A2(new_n312), .A3(G200), .ZN(new_n795));
  INV_X1    g0595(.A(G283), .ZN(new_n796));
  OAI22_X1  g0596(.A1(new_n793), .A2(new_n794), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n784), .A2(new_n788), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  AOI211_X1 g0599(.A(new_n791), .B(new_n797), .C1(G329), .C2(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n776), .A2(KEYINPUT94), .ZN(new_n801));
  NAND4_X1  g0601(.A1(new_n777), .A2(new_n787), .A3(new_n800), .A4(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n782), .A2(new_n286), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n793), .A2(new_n466), .ZN(new_n804));
  OAI22_X1  g0604(.A1(new_n770), .A2(new_n319), .B1(new_n785), .B2(new_n707), .ZN(new_n805));
  INV_X1    g0605(.A(new_n795), .ZN(new_n806));
  AOI211_X1 g0606(.A(new_n804), .B(new_n805), .C1(G107), .C2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(G159), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n798), .A2(new_n808), .ZN(new_n809));
  XNOR2_X1  g0609(.A(new_n809), .B(KEYINPUT32), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n247), .B1(new_n773), .B2(new_n360), .ZN(new_n811));
  INV_X1    g0611(.A(new_n789), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n811), .B1(G77), .B2(new_n812), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n807), .A2(new_n810), .A3(new_n813), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n802), .B1(new_n803), .B2(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n768), .B1(new_n815), .B2(new_n765), .ZN(new_n816));
  XNOR2_X1  g0616(.A(new_n764), .B(KEYINPUT95), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n816), .B1(new_n701), .B2(new_n817), .ZN(new_n818));
  AND2_X1   g0618(.A1(new_n755), .A2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(G396));
  NOR2_X1   g0620(.A1(new_n765), .A2(new_n762), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n786), .ZN(new_n823));
  INV_X1    g0623(.A(G303), .ZN(new_n824));
  OAI22_X1  g0624(.A1(new_n823), .A2(new_n446), .B1(new_n824), .B2(new_n782), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n247), .B1(new_n799), .B2(G311), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n826), .B1(new_n624), .B2(new_n789), .C1(new_n794), .C2(new_n773), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n804), .B1(G283), .B2(new_n771), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n828), .B1(new_n707), .B2(new_n795), .ZN(new_n829));
  NOR3_X1   g0629(.A1(new_n825), .A2(new_n827), .A3(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n823), .A2(new_n286), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n335), .B1(new_n799), .B2(G132), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n832), .B1(new_n360), .B2(new_n793), .C1(new_n319), .C2(new_n795), .ZN(new_n833));
  AOI22_X1  g0633(.A1(new_n774), .A2(G143), .B1(new_n812), .B2(G159), .ZN(new_n834));
  AOI22_X1  g0634(.A1(new_n783), .A2(G137), .B1(G150), .B2(new_n771), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n836), .A2(KEYINPUT96), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n836), .A2(KEYINPUT96), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n834), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT34), .ZN(new_n841));
  AOI211_X1 g0641(.A(new_n831), .B(new_n833), .C1(new_n840), .C2(new_n841), .ZN(new_n842));
  OR2_X1    g0642(.A1(new_n840), .A2(new_n841), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n830), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n765), .ZN(new_n845));
  OAI221_X1 g0645(.A(new_n753), .B1(G77), .B2(new_n822), .C1(new_n844), .C2(new_n845), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n455), .A2(new_n682), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n452), .B1(new_n443), .B2(new_n690), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n847), .B1(new_n848), .B2(new_n455), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n846), .B1(new_n762), .B2(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n849), .B1(new_n658), .B2(new_n690), .ZN(new_n852));
  OAI211_X1 g0652(.A(new_n690), .B(new_n849), .C1(new_n654), .C2(new_n657), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  OR2_X1    g0654(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  OR2_X1    g0655(.A1(new_n855), .A2(new_n744), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n753), .B1(new_n855), .B2(new_n744), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n851), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(G384));
  NOR3_X1   g0659(.A1(new_n222), .A2(new_n221), .A3(new_n624), .ZN(new_n860));
  XNOR2_X1  g0660(.A(new_n476), .B(KEYINPUT97), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT35), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n860), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n863), .B1(new_n862), .B2(new_n861), .ZN(new_n864));
  XOR2_X1   g0664(.A(KEYINPUT98), .B(KEYINPUT36), .Z(new_n865));
  XNOR2_X1  g0665(.A(new_n864), .B(new_n865), .ZN(new_n866));
  NOR3_X1   g0666(.A1(new_n382), .A2(new_n220), .A3(new_n246), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT99), .ZN(new_n868));
  OR2_X1    g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  AOI22_X1  g0669(.A1(new_n867), .A2(new_n868), .B1(new_n286), .B2(G68), .ZN(new_n870));
  AOI211_X1 g0670(.A(new_n253), .B(G13), .C1(new_n869), .C2(new_n870), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n866), .A2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT38), .ZN(new_n873));
  INV_X1    g0673(.A(new_n680), .ZN(new_n874));
  AOI21_X1  g0674(.A(KEYINPUT37), .B1(new_n394), .B2(new_n874), .ZN(new_n875));
  NAND4_X1  g0675(.A1(new_n418), .A2(new_n875), .A3(new_n409), .A4(new_n426), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n367), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n423), .A2(new_n278), .ZN(new_n879));
  AOI21_X1  g0679(.A(KEYINPUT16), .B1(new_n421), .B2(new_n431), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n878), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(new_n660), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n882), .A2(new_n418), .A3(new_n426), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT100), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND4_X1  g0685(.A1(new_n882), .A2(new_n418), .A3(KEYINPUT100), .A4(new_n426), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n881), .A2(new_n874), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n877), .B1(new_n888), .B2(KEYINPUT37), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n887), .B1(new_n459), .B2(new_n461), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n873), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n459), .A2(new_n461), .ZN(new_n892));
  INV_X1    g0692(.A(new_n887), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT37), .ZN(new_n895));
  AND2_X1   g0695(.A1(new_n886), .A2(new_n887), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n895), .B1(new_n896), .B2(new_n885), .ZN(new_n897));
  OAI211_X1 g0697(.A(KEYINPUT38), .B(new_n894), .C1(new_n897), .C2(new_n877), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n891), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n329), .A2(new_n690), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(new_n358), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n901), .B1(new_n902), .B2(new_n667), .ZN(new_n903));
  NOR3_X1   g0703(.A1(new_n351), .A2(new_n358), .A3(new_n900), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n849), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n737), .A2(KEYINPUT31), .A3(new_n682), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n722), .A2(new_n740), .A3(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT104), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND4_X1  g0709(.A1(new_n722), .A2(new_n740), .A3(KEYINPUT104), .A4(new_n906), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n905), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(KEYINPUT40), .B1(new_n899), .B2(new_n911), .ZN(new_n912));
  XOR2_X1   g0712(.A(KEYINPUT102), .B(KEYINPUT38), .Z(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n425), .B1(new_n434), .B2(new_n420), .ZN(new_n915));
  NOR3_X1   g0715(.A1(new_n394), .A2(new_n417), .A3(KEYINPUT77), .ZN(new_n916));
  OAI21_X1  g0716(.A(KEYINPUT17), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(new_n435), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n917), .A2(new_n918), .A3(new_n663), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n394), .A2(new_n874), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n394), .A2(new_n660), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n923), .B(new_n920), .C1(new_n394), .C2(new_n417), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(KEYINPUT37), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(new_n876), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n914), .B1(new_n922), .B2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n898), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n902), .A2(new_n667), .A3(new_n901), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n900), .B1(new_n351), .B2(new_n358), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n850), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(KEYINPUT31), .B1(new_n737), .B2(new_n682), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n933), .B1(new_n645), .B2(new_n690), .ZN(new_n934));
  AOI21_X1  g0734(.A(KEYINPUT104), .B1(new_n934), .B2(new_n906), .ZN(new_n935));
  INV_X1    g0735(.A(new_n910), .ZN(new_n936));
  OAI211_X1 g0736(.A(KEYINPUT40), .B(new_n932), .C1(new_n935), .C2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n912), .B1(new_n929), .B2(new_n938), .ZN(new_n939));
  AOI22_X1  g0739(.A1(new_n458), .A2(new_n464), .B1(new_n909), .B2(new_n910), .ZN(new_n940));
  AND2_X1   g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n939), .A2(new_n940), .ZN(new_n942));
  INV_X1    g0742(.A(G330), .ZN(new_n943));
  NOR3_X1   g0743(.A1(new_n941), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT39), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n929), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n351), .A2(new_n690), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT101), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n947), .B(new_n948), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n891), .A2(new_n898), .A3(KEYINPUT39), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n946), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(new_n847), .ZN(new_n952));
  AOI22_X1  g0752(.A1(new_n853), .A2(new_n952), .B1(new_n930), .B2(new_n931), .ZN(new_n953));
  AOI22_X1  g0753(.A1(new_n899), .A2(new_n953), .B1(new_n664), .B2(new_n680), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n951), .A2(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n714), .A2(new_n719), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n673), .B1(new_n465), .B2(new_n957), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n958), .B(KEYINPUT103), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n956), .B(new_n959), .ZN(new_n960));
  OAI22_X1  g0760(.A1(new_n944), .A2(new_n960), .B1(new_n253), .B2(new_n750), .ZN(new_n961));
  AND2_X1   g0761(.A1(new_n944), .A2(new_n960), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n872), .B1(new_n961), .B2(new_n962), .ZN(G367));
  NAND2_X1  g0763(.A1(new_n576), .A2(new_n577), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n964), .A2(new_n682), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n653), .A2(new_n965), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n966), .B1(new_n587), .B2(new_n965), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT43), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  OR2_X1    g0769(.A1(new_n967), .A2(new_n968), .ZN(new_n970));
  INV_X1    g0770(.A(new_n695), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n482), .A2(new_n682), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n509), .A2(new_n972), .A3(new_n601), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n648), .A2(new_n682), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n971), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(KEYINPUT42), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n509), .B1(new_n973), .B2(new_n613), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n978), .A2(new_n690), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n976), .A2(KEYINPUT42), .ZN(new_n981));
  OAI211_X1 g0781(.A(new_n969), .B(new_n970), .C1(new_n980), .C2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(new_n703), .ZN(new_n983));
  INV_X1    g0783(.A(new_n975), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(new_n981), .ZN(new_n986));
  AOI22_X1  g0786(.A1(new_n976), .A2(KEYINPUT42), .B1(new_n690), .B2(new_n978), .ZN(new_n987));
  NAND4_X1  g0787(.A1(new_n986), .A2(new_n987), .A3(new_n968), .A4(new_n967), .ZN(new_n988));
  AND3_X1   g0788(.A1(new_n982), .A2(new_n985), .A3(new_n988), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n985), .B1(new_n982), .B2(new_n988), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  XNOR2_X1  g0791(.A(KEYINPUT105), .B(KEYINPUT41), .ZN(new_n992));
  XOR2_X1   g0792(.A(new_n706), .B(new_n992), .Z(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  AOI21_X1  g0794(.A(KEYINPUT44), .B1(new_n696), .B2(new_n984), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT44), .ZN(new_n996));
  AOI211_X1 g0796(.A(new_n996), .B(new_n975), .C1(new_n695), .C2(new_n691), .ZN(new_n997));
  OR2_X1    g0797(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n695), .A2(new_n691), .A3(new_n975), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT45), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n999), .B(new_n1000), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n998), .A2(new_n983), .A3(new_n1001), .ZN(new_n1002));
  AND2_X1   g0802(.A1(new_n999), .A2(new_n1000), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n999), .A2(new_n1000), .ZN(new_n1004));
  OAI22_X1  g0804(.A1(new_n1003), .A2(new_n1004), .B1(new_n995), .B2(new_n997), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1005), .A2(new_n703), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n697), .A2(new_n693), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n702), .B1(new_n1007), .B2(KEYINPUT106), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n694), .B1(new_n686), .B2(new_n692), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT106), .ZN(new_n1010));
  NOR3_X1   g0810(.A1(new_n1009), .A2(new_n1010), .A3(new_n748), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n695), .B1(new_n1008), .B2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1007), .A2(KEYINPUT106), .A3(new_n702), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n748), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1013), .A2(new_n971), .A3(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n745), .B1(new_n1012), .B2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1002), .A2(new_n1006), .A3(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n994), .B1(new_n1017), .B2(new_n746), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n991), .B1(new_n1018), .B2(new_n752), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n766), .B1(new_n207), .B2(new_n439), .C1(new_n758), .C2(new_n231), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n783), .A2(G311), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n793), .A2(new_n446), .B1(new_n795), .B2(new_n466), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1022), .B1(G294), .B2(new_n771), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n786), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n785), .ZN(new_n1025));
  AOI21_X1  g0825(.A(KEYINPUT46), .B1(new_n1025), .B2(G116), .ZN(new_n1026));
  INV_X1    g0826(.A(G317), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n773), .A2(new_n824), .B1(new_n798), .B2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n335), .B1(new_n789), .B2(new_n796), .ZN(new_n1029));
  NOR3_X1   g0829(.A1(new_n1026), .A2(new_n1028), .A3(new_n1029), .ZN(new_n1030));
  NAND4_X1  g0830(.A1(new_n1021), .A2(new_n1023), .A3(new_n1024), .A4(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(G137), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n247), .B1(new_n798), .B2(new_n1032), .C1(new_n286), .C2(new_n789), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n806), .A2(G77), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1034), .B1(new_n808), .B2(new_n770), .ZN(new_n1035));
  AOI211_X1 g0835(.A(new_n1033), .B(new_n1035), .C1(G58), .C2(new_n1025), .ZN(new_n1036));
  INV_X1    g0836(.A(G143), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1036), .B1(new_n1037), .B2(new_n782), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n793), .A2(new_n319), .B1(new_n773), .B2(new_n281), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1039), .B(KEYINPUT107), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1031), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1041));
  XOR2_X1   g0841(.A(new_n1041), .B(KEYINPUT47), .Z(new_n1042));
  OAI211_X1 g0842(.A(new_n753), .B(new_n1020), .C1(new_n1042), .C2(new_n845), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n817), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1043), .B1(new_n1044), .B2(new_n967), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT108), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1019), .A2(new_n1046), .ZN(G387));
  NAND2_X1  g0847(.A1(new_n1012), .A2(new_n1015), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1048), .A2(new_n746), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1012), .A2(new_n745), .A3(new_n1015), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1049), .A2(new_n706), .A3(new_n1050), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n789), .A2(new_n319), .B1(new_n798), .B2(new_n281), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n335), .B(new_n1052), .C1(G50), .C2(new_n774), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n793), .A2(new_n439), .B1(new_n785), .B2(new_n246), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n770), .A2(new_n279), .B1(new_n795), .B2(new_n466), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n1053), .B(new_n1056), .C1(new_n808), .C2(new_n782), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1057), .B(KEYINPUT110), .ZN(new_n1058));
  INV_X1    g0858(.A(G322), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n782), .A2(new_n1059), .B1(new_n790), .B2(new_n770), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT111), .ZN(new_n1061));
  OR2_X1    g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n774), .A2(G317), .B1(new_n812), .B2(G303), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1062), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT48), .ZN(new_n1066));
  OR2_X1    g0866(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n793), .A2(new_n796), .B1(new_n785), .B2(new_n794), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1068), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1067), .A2(KEYINPUT49), .A3(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n247), .B1(new_n799), .B2(G326), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n1070), .B(new_n1071), .C1(new_n624), .C2(new_n795), .ZN(new_n1072));
  AOI21_X1  g0872(.A(KEYINPUT49), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1058), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n765), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n753), .ZN(new_n1076));
  NOR3_X1   g0876(.A1(new_n228), .A2(new_n262), .A3(new_n247), .ZN(new_n1077));
  XOR2_X1   g0877(.A(KEYINPUT109), .B(KEYINPUT50), .Z(new_n1078));
  INV_X1    g0878(.A(new_n1078), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1079), .B1(new_n279), .B2(G50), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n437), .A2(new_n286), .A3(new_n1078), .ZN(new_n1081));
  AOI21_X1  g0881(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1080), .A2(new_n1081), .A3(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n708), .B1(new_n1083), .B2(new_n335), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n207), .B1(new_n1077), .B2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n767), .B1(new_n705), .B2(G107), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1076), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1075), .A2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1088), .B1(new_n697), .B2(new_n1044), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1089), .B1(new_n1048), .B2(new_n752), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1051), .A2(new_n1090), .ZN(G393));
  INV_X1    g0891(.A(KEYINPUT112), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1002), .A2(new_n1006), .A3(new_n1092), .ZN(new_n1093));
  NAND4_X1  g0893(.A1(new_n998), .A2(KEYINPUT112), .A3(new_n983), .A4(new_n1001), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1093), .A2(new_n1049), .A3(new_n1094), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1095), .A2(new_n706), .A3(new_n1017), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n235), .A2(new_n758), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n766), .B1(new_n207), .B2(new_n466), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n753), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  NOR3_X1   g0899(.A1(new_n975), .A2(G20), .A3(new_n763), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n782), .A2(new_n1027), .B1(new_n790), .B2(new_n773), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(new_n1101), .B(KEYINPUT52), .ZN(new_n1102));
  OAI221_X1 g0902(.A(new_n335), .B1(new_n798), .B2(new_n1059), .C1(new_n794), .C2(new_n789), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n770), .A2(new_n824), .B1(new_n795), .B2(new_n446), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n793), .A2(new_n624), .B1(new_n785), .B2(new_n796), .ZN(new_n1105));
  NOR3_X1   g0905(.A1(new_n1103), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n782), .A2(new_n281), .B1(new_n808), .B2(new_n773), .ZN(new_n1107));
  XNOR2_X1  g0907(.A(new_n1107), .B(KEYINPUT51), .ZN(new_n1108));
  OAI221_X1 g0908(.A(new_n247), .B1(new_n798), .B2(new_n1037), .C1(new_n279), .C2(new_n789), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n770), .A2(new_n286), .B1(new_n795), .B2(new_n707), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n793), .A2(new_n246), .B1(new_n785), .B2(new_n319), .ZN(new_n1111));
  NOR3_X1   g0911(.A1(new_n1109), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n1102), .A2(new_n1106), .B1(new_n1108), .B2(new_n1112), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(new_n1113), .B(KEYINPUT113), .ZN(new_n1114));
  AOI211_X1 g0914(.A(new_n1099), .B(new_n1100), .C1(new_n765), .C2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1115), .B1(new_n1116), .B2(new_n752), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1096), .A2(new_n1117), .ZN(G390));
  AOI21_X1  g0918(.A(new_n943), .B1(new_n909), .B2(new_n910), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(new_n932), .ZN(new_n1120));
  INV_X1    g0920(.A(KEYINPUT114), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1121), .B1(new_n953), .B2(new_n949), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(new_n947), .B(KEYINPUT101), .ZN(new_n1123));
  AND2_X1   g0923(.A1(new_n853), .A2(new_n952), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n903), .A2(new_n904), .ZN(new_n1125));
  OAI211_X1 g0925(.A(KEYINPUT114), .B(new_n1123), .C1(new_n1124), .C2(new_n1125), .ZN(new_n1126));
  AND3_X1   g0926(.A1(new_n891), .A2(KEYINPUT39), .A3(new_n898), .ZN(new_n1127));
  AOI21_X1  g0927(.A(KEYINPUT39), .B1(new_n898), .B2(new_n928), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n1122), .B(new_n1126), .C1(new_n1127), .C2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n848), .A2(new_n455), .ZN(new_n1130));
  OAI211_X1 g0930(.A(new_n690), .B(new_n1130), .C1(new_n717), .C2(new_n657), .ZN(new_n1131));
  AND2_X1   g0931(.A1(new_n1131), .A2(new_n952), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1123), .B1(new_n1132), .B2(new_n1125), .ZN(new_n1133));
  AND2_X1   g0933(.A1(new_n883), .A2(new_n884), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n886), .A2(new_n887), .ZN(new_n1135));
  OAI21_X1  g0935(.A(KEYINPUT37), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n890), .B1(new_n1136), .B2(new_n876), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n927), .B1(new_n1137), .B2(KEYINPUT38), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n1133), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1120), .B1(new_n1129), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1125), .ZN(new_n1143));
  NAND4_X1  g0943(.A1(new_n1143), .A2(G330), .A3(new_n743), .A4(new_n849), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1129), .A2(new_n1140), .A3(new_n1144), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n849), .B1(new_n1119), .B2(KEYINPUT116), .ZN(new_n1146));
  INV_X1    g0946(.A(KEYINPUT116), .ZN(new_n1147));
  AOI211_X1 g0947(.A(new_n1147), .B(new_n943), .C1(new_n909), .C2(new_n910), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1125), .B1(new_n1146), .B2(new_n1148), .ZN(new_n1149));
  AND2_X1   g0949(.A1(new_n1144), .A2(new_n1132), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1125), .B1(new_n744), .B2(new_n850), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1124), .B1(new_n1120), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1151), .A2(new_n1154), .ZN(new_n1155));
  AND3_X1   g0955(.A1(new_n465), .A2(KEYINPUT115), .A3(new_n1119), .ZN(new_n1156));
  AOI21_X1  g0956(.A(KEYINPUT115), .B1(new_n465), .B2(new_n1119), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n958), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n1142), .A2(new_n1145), .A3(new_n1155), .A4(new_n1159), .ZN(new_n1160));
  AND3_X1   g0960(.A1(new_n1129), .A2(new_n1140), .A3(new_n1144), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1153), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1162));
  OAI22_X1  g0962(.A1(new_n1161), .A2(new_n1141), .B1(new_n1162), .B2(new_n1158), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1160), .A2(new_n706), .A3(new_n1163), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n1161), .A2(new_n1141), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n946), .A2(new_n950), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1166), .A2(new_n762), .ZN(new_n1167));
  INV_X1    g0967(.A(KEYINPUT119), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n753), .B1(new_n437), .B2(new_n822), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n785), .A2(new_n281), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(new_n1170), .B(KEYINPUT53), .ZN(new_n1171));
  INV_X1    g0971(.A(G128), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1171), .B1(new_n782), .B2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n335), .B1(new_n774), .B2(G132), .ZN(new_n1174));
  INV_X1    g0974(.A(G125), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(KEYINPUT54), .B(G143), .ZN(new_n1176));
  OAI221_X1 g0976(.A(new_n1174), .B1(new_n1175), .B2(new_n798), .C1(new_n789), .C2(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n793), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n1178), .A2(G159), .B1(new_n806), .B2(G50), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1179), .B1(new_n1032), .B2(new_n770), .ZN(new_n1180));
  NOR3_X1   g0980(.A1(new_n1173), .A2(new_n1177), .A3(new_n1180), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(new_n771), .A2(G107), .B1(new_n812), .B2(G97), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1182), .B1(new_n782), .B2(new_n796), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(new_n1183), .B(KEYINPUT117), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n335), .B1(new_n798), .B2(new_n794), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(G116), .B2(new_n774), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n1178), .A2(G77), .B1(new_n806), .B2(G68), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1188), .B1(G87), .B2(new_n786), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1181), .B1(new_n1184), .B2(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n1191), .A2(KEYINPUT118), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n845), .B1(new_n1191), .B2(KEYINPUT118), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1169), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1167), .A2(new_n1168), .A3(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1167), .A2(new_n1195), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1197), .A2(KEYINPUT119), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(new_n1165), .A2(new_n752), .B1(new_n1196), .B2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1164), .A2(new_n1199), .ZN(G378));
  NAND2_X1  g1000(.A1(new_n299), .A2(new_n874), .ZN(new_n1201));
  AND2_X1   g1001(.A1(new_n318), .A2(new_n1201), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n318), .A2(new_n1201), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1204), .ZN(new_n1205));
  OR3_X1    g1005(.A1(new_n1202), .A2(new_n1203), .A3(new_n1205), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1205), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(new_n1209));
  OAI21_X1  g1009(.A(G330), .B1(new_n937), .B2(new_n1138), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n899), .A2(new_n911), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT40), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1209), .B1(new_n1211), .B2(new_n1214), .ZN(new_n1215));
  NOR3_X1   g1015(.A1(new_n912), .A2(new_n1210), .A3(new_n1208), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n956), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1211), .A2(new_n1214), .A3(new_n1209), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1208), .B1(new_n912), .B2(new_n1210), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1218), .A2(new_n955), .A3(new_n1219), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1217), .A2(KEYINPUT122), .A3(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n955), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT122), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1221), .A2(new_n752), .A3(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1209), .A2(new_n762), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n753), .B1(G50), .B2(new_n822), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n774), .A2(G128), .B1(new_n812), .B2(G137), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1228), .B1(new_n785), .B2(new_n1176), .ZN(new_n1229));
  OAI22_X1  g1029(.A1(new_n782), .A2(new_n1175), .B1(new_n281), .B2(new_n793), .ZN(new_n1230));
  XNOR2_X1  g1030(.A(new_n1230), .B(KEYINPUT121), .ZN(new_n1231));
  AOI211_X1 g1031(.A(new_n1229), .B(new_n1231), .C1(G132), .C2(new_n771), .ZN(new_n1232));
  XNOR2_X1  g1032(.A(new_n1232), .B(KEYINPUT59), .ZN(new_n1233));
  AOI211_X1 g1033(.A(G33), .B(G41), .C1(new_n799), .C2(G124), .ZN(new_n1234));
  OAI211_X1 g1034(.A(new_n1233), .B(new_n1234), .C1(new_n808), .C2(new_n795), .ZN(new_n1235));
  OAI211_X1 g1035(.A(new_n261), .B(new_n335), .C1(new_n785), .C2(new_n246), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(new_n783), .A2(G116), .B1(new_n1236), .B2(KEYINPUT120), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1237), .B1(KEYINPUT120), .B2(new_n1236), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n581), .A2(new_n812), .B1(new_n799), .B2(G283), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1239), .B1(new_n446), .B2(new_n773), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n806), .A2(G58), .ZN(new_n1241));
  OAI221_X1 g1041(.A(new_n1241), .B1(new_n466), .B2(new_n770), .C1(new_n319), .C2(new_n793), .ZN(new_n1242));
  NOR3_X1   g1042(.A1(new_n1238), .A2(new_n1240), .A3(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1243), .A2(KEYINPUT58), .ZN(new_n1244));
  AOI21_X1  g1044(.A(G50), .B1(new_n374), .B2(new_n261), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1245), .B1(new_n247), .B2(G41), .ZN(new_n1246));
  OR2_X1    g1046(.A1(new_n1243), .A2(KEYINPUT58), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n1235), .A2(new_n1244), .A3(new_n1246), .A4(new_n1247), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1227), .B1(new_n1248), .B2(new_n765), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1226), .A2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1225), .A2(new_n1250), .ZN(new_n1251));
  AND2_X1   g1051(.A1(new_n1126), .A2(new_n1122), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1139), .B1(new_n1252), .B2(new_n1166), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1145), .B1(new_n1253), .B2(new_n1120), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1159), .B1(new_n1254), .B2(new_n1162), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1255), .A2(new_n1221), .A3(new_n1224), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT57), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n706), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1257), .B1(new_n1217), .B2(new_n1220), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1259), .B1(new_n1260), .B2(new_n1255), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1251), .B1(new_n1258), .B2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(G375));
  NAND2_X1  g1063(.A1(new_n1125), .A2(new_n762), .ZN(new_n1264));
  XOR2_X1   g1064(.A(new_n1264), .B(KEYINPUT123), .Z(new_n1265));
  AOI22_X1  g1065(.A1(new_n786), .A2(G97), .B1(G303), .B2(new_n799), .ZN(new_n1266));
  XNOR2_X1  g1066(.A(new_n1266), .B(KEYINPUT124), .ZN(new_n1267));
  OAI221_X1 g1067(.A(new_n335), .B1(new_n789), .B2(new_n446), .C1(new_n796), .C2(new_n773), .ZN(new_n1268));
  OAI221_X1 g1068(.A(new_n1034), .B1(new_n624), .B2(new_n770), .C1(new_n439), .C2(new_n793), .ZN(new_n1269));
  AOI211_X1 g1069(.A(new_n1268), .B(new_n1269), .C1(G294), .C2(new_n783), .ZN(new_n1270));
  OAI221_X1 g1070(.A(new_n1241), .B1(new_n770), .B2(new_n1176), .C1(new_n286), .C2(new_n793), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n247), .B1(new_n773), .B2(new_n1032), .ZN(new_n1272));
  OAI22_X1  g1072(.A1(new_n789), .A2(new_n281), .B1(new_n798), .B2(new_n1172), .ZN(new_n1273));
  NOR3_X1   g1073(.A1(new_n1271), .A2(new_n1272), .A3(new_n1273), .ZN(new_n1274));
  AOI22_X1  g1074(.A1(new_n783), .A2(G132), .B1(G159), .B2(new_n786), .ZN(new_n1275));
  AOI22_X1  g1075(.A1(new_n1267), .A2(new_n1270), .B1(new_n1274), .B2(new_n1275), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1276), .A2(new_n845), .ZN(new_n1277));
  AOI211_X1 g1077(.A(new_n1076), .B(new_n1277), .C1(new_n319), .C2(new_n821), .ZN(new_n1278));
  AOI22_X1  g1078(.A1(new_n1155), .A2(new_n752), .B1(new_n1265), .B2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1162), .A2(new_n1158), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1281), .A2(new_n994), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1162), .A2(new_n1158), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1280), .B1(new_n1282), .B2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1284), .ZN(G381));
  AND2_X1   g1085(.A1(new_n1096), .A2(new_n1117), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1051), .A2(new_n819), .A3(new_n1090), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1287), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1286), .A2(new_n858), .A3(new_n1284), .A4(new_n1288), .ZN(new_n1289));
  OR4_X1    g1089(.A1(G387), .A2(G375), .A3(G378), .A4(new_n1289), .ZN(G407));
  INV_X1    g1090(.A(G378), .ZN(new_n1291));
  INV_X1    g1091(.A(G213), .ZN(new_n1292));
  NOR2_X1   g1092(.A1(new_n1292), .A2(G343), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1262), .A2(new_n1291), .A3(new_n1293), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(G407), .A2(G213), .A3(new_n1294), .ZN(G409));
  INV_X1    g1095(.A(KEYINPUT61), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1286), .A2(G387), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(G390), .A2(new_n1046), .A3(new_n1019), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n819), .B1(new_n1051), .B2(new_n1090), .ZN(new_n1299));
  OAI21_X1  g1099(.A(KEYINPUT126), .B1(new_n1288), .B2(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1299), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT126), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1301), .A2(new_n1302), .A3(new_n1287), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1300), .A2(new_n1303), .ZN(new_n1304));
  AND3_X1   g1104(.A1(new_n1297), .A2(new_n1298), .A3(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1300), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1306), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1296), .B1(new_n1305), .B2(new_n1307), .ZN(new_n1308));
  NAND4_X1  g1108(.A1(new_n1151), .A2(KEYINPUT60), .A3(new_n1158), .A4(new_n1154), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1309), .A2(new_n706), .ZN(new_n1310));
  OAI21_X1  g1110(.A(KEYINPUT60), .B1(new_n1162), .B2(new_n1158), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1310), .B1(new_n1283), .B2(new_n1311), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n858), .B1(new_n1312), .B2(new_n1280), .ZN(new_n1313));
  AND2_X1   g1113(.A1(new_n1311), .A2(new_n1283), .ZN(new_n1314));
  OAI211_X1 g1114(.A(G384), .B(new_n1279), .C1(new_n1314), .C2(new_n1310), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1293), .A2(G2897), .ZN(new_n1316));
  AND3_X1   g1116(.A1(new_n1313), .A2(new_n1315), .A3(new_n1316), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1316), .B1(new_n1313), .B2(new_n1315), .ZN(new_n1318));
  NOR2_X1   g1118(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1319));
  NAND4_X1  g1119(.A1(new_n1255), .A2(new_n1221), .A3(new_n993), .A4(new_n1224), .ZN(new_n1320));
  AND3_X1   g1120(.A1(new_n1218), .A2(new_n955), .A3(new_n1219), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n752), .B1(new_n1321), .B2(new_n1222), .ZN(new_n1322));
  AND2_X1   g1122(.A1(new_n1322), .A2(new_n1250), .ZN(new_n1323));
  AOI21_X1  g1123(.A(G378), .B1(new_n1320), .B2(new_n1323), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1324), .B1(new_n1262), .B2(G378), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1319), .B1(new_n1325), .B2(new_n1293), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1308), .B1(new_n1326), .B2(KEYINPUT125), .ZN(new_n1327));
  INV_X1    g1127(.A(KEYINPUT125), .ZN(new_n1328));
  OAI211_X1 g1128(.A(new_n1319), .B(new_n1328), .C1(new_n1325), .C2(new_n1293), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1258), .A2(new_n1261), .ZN(new_n1330));
  INV_X1    g1130(.A(new_n1251), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1330), .A2(G378), .A3(new_n1331), .ZN(new_n1332));
  INV_X1    g1132(.A(new_n1324), .ZN(new_n1333));
  AOI21_X1  g1133(.A(new_n1293), .B1(new_n1332), .B2(new_n1333), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1313), .A2(new_n1315), .ZN(new_n1335));
  INV_X1    g1135(.A(new_n1335), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1334), .A2(new_n1336), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT63), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1337), .A2(new_n1338), .ZN(new_n1339));
  NAND3_X1  g1139(.A1(new_n1334), .A2(KEYINPUT63), .A3(new_n1336), .ZN(new_n1340));
  NAND4_X1  g1140(.A1(new_n1327), .A2(new_n1329), .A3(new_n1339), .A4(new_n1340), .ZN(new_n1341));
  NOR2_X1   g1141(.A1(new_n1305), .A2(new_n1307), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1332), .A2(new_n1333), .ZN(new_n1343));
  INV_X1    g1143(.A(KEYINPUT62), .ZN(new_n1344));
  INV_X1    g1144(.A(new_n1293), .ZN(new_n1345));
  NAND4_X1  g1145(.A1(new_n1343), .A2(new_n1344), .A3(new_n1345), .A4(new_n1336), .ZN(new_n1346));
  NAND3_X1  g1146(.A1(new_n1346), .A2(new_n1326), .A3(new_n1296), .ZN(new_n1347));
  AOI21_X1  g1147(.A(new_n1344), .B1(new_n1334), .B2(new_n1336), .ZN(new_n1348));
  OAI21_X1  g1148(.A(new_n1342), .B1(new_n1347), .B2(new_n1348), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1341), .A2(new_n1349), .ZN(G405));
  INV_X1    g1150(.A(new_n1342), .ZN(new_n1351));
  INV_X1    g1151(.A(KEYINPUT127), .ZN(new_n1352));
  AND3_X1   g1152(.A1(new_n1330), .A2(G378), .A3(new_n1331), .ZN(new_n1353));
  AOI21_X1  g1153(.A(G378), .B1(new_n1330), .B2(new_n1331), .ZN(new_n1354));
  OAI21_X1  g1154(.A(new_n1352), .B1(new_n1353), .B2(new_n1354), .ZN(new_n1355));
  AOI21_X1  g1155(.A(new_n1158), .B1(new_n1165), .B2(new_n1281), .ZN(new_n1356));
  OAI21_X1  g1156(.A(KEYINPUT57), .B1(new_n1321), .B2(new_n1222), .ZN(new_n1357));
  OAI21_X1  g1157(.A(new_n706), .B1(new_n1356), .B2(new_n1357), .ZN(new_n1358));
  AOI21_X1  g1158(.A(new_n1358), .B1(new_n1257), .B2(new_n1256), .ZN(new_n1359));
  OAI21_X1  g1159(.A(new_n1291), .B1(new_n1359), .B2(new_n1251), .ZN(new_n1360));
  NAND3_X1  g1160(.A1(new_n1360), .A2(KEYINPUT127), .A3(new_n1332), .ZN(new_n1361));
  AND3_X1   g1161(.A1(new_n1355), .A2(new_n1361), .A3(new_n1335), .ZN(new_n1362));
  AOI21_X1  g1162(.A(new_n1335), .B1(new_n1355), .B2(new_n1361), .ZN(new_n1363));
  OAI21_X1  g1163(.A(new_n1351), .B1(new_n1362), .B2(new_n1363), .ZN(new_n1364));
  NOR3_X1   g1164(.A1(new_n1353), .A2(new_n1354), .A3(new_n1352), .ZN(new_n1365));
  AOI21_X1  g1165(.A(KEYINPUT127), .B1(new_n1360), .B2(new_n1332), .ZN(new_n1366));
  OAI21_X1  g1166(.A(new_n1336), .B1(new_n1365), .B2(new_n1366), .ZN(new_n1367));
  NAND3_X1  g1167(.A1(new_n1355), .A2(new_n1361), .A3(new_n1335), .ZN(new_n1368));
  NAND3_X1  g1168(.A1(new_n1367), .A2(new_n1342), .A3(new_n1368), .ZN(new_n1369));
  NAND2_X1  g1169(.A1(new_n1364), .A2(new_n1369), .ZN(G402));
endmodule


