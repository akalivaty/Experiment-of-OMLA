//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 1 0 0 1 0 1 0 0 1 1 1 1 1 0 0 1 1 1 0 1 0 1 1 1 0 0 0 1 0 1 1 1 0 1 1 1 0 0 1 1 1 1 0 1 1 1 1 1 1 1 1 1 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:19 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1284, new_n1285,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(new_n207), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  OAI21_X1  g0015(.A(G50), .B1(G58), .B2(G68), .ZN(new_n216));
  XOR2_X1   g0016(.A(new_n216), .B(KEYINPUT64), .Z(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n218));
  XOR2_X1   g0018(.A(new_n218), .B(KEYINPUT65), .Z(new_n219));
  AOI22_X1  g0019(.A1(G77), .A2(G244), .B1(G87), .B2(G250), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G68), .A2(G238), .B1(G107), .B2(G264), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n222));
  NAND3_X1  g0022(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n209), .B1(new_n219), .B2(new_n223), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n212), .B1(new_n215), .B2(new_n217), .C1(new_n224), .C2(KEYINPUT1), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n225), .B1(KEYINPUT1), .B2(new_n224), .ZN(G361));
  XNOR2_X1  g0026(.A(G238), .B(G244), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT2), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(G226), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(G232), .ZN(new_n230));
  XOR2_X1   g0030(.A(G250), .B(G257), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT66), .ZN(new_n232));
  XOR2_X1   g0032(.A(G264), .B(G270), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n230), .B(new_n234), .ZN(G358));
  XOR2_X1   g0035(.A(G68), .B(G77), .Z(new_n236));
  XNOR2_X1  g0036(.A(G50), .B(G58), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XNOR2_X1  g0039(.A(G107), .B(G116), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G351));
  NOR2_X1   g0042(.A1(G20), .A2(G33), .ZN(new_n243));
  AOI22_X1  g0043(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(KEYINPUT8), .B(G58), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n207), .A2(G33), .ZN(new_n246));
  OAI21_X1  g0046(.A(new_n244), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NAND3_X1  g0047(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(new_n213), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(G13), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n251), .A2(G1), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(G20), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(new_n202), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n249), .B1(new_n206), .B2(G20), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n254), .B1(new_n255), .B2(new_n202), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n250), .A2(new_n256), .ZN(new_n257));
  XNOR2_X1  g0057(.A(new_n257), .B(KEYINPUT9), .ZN(new_n258));
  NAND2_X1  g0058(.A1(G33), .A2(G41), .ZN(new_n259));
  NAND4_X1  g0059(.A1(new_n259), .A2(KEYINPUT68), .A3(G1), .A4(G13), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  AND2_X1   g0061(.A1(G1), .A2(G13), .ZN(new_n262));
  AOI21_X1  g0062(.A(KEYINPUT68), .B1(new_n262), .B2(new_n259), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  AND2_X1   g0064(.A1(KEYINPUT67), .A2(G41), .ZN(new_n265));
  NOR2_X1   g0065(.A1(KEYINPUT67), .A2(G41), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G45), .ZN(new_n268));
  AOI21_X1  g0068(.A(G1), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n264), .A2(new_n269), .A3(G274), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n264), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G226), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n270), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  XNOR2_X1  g0075(.A(KEYINPUT3), .B(G33), .ZN(new_n276));
  INV_X1    g0076(.A(G1698), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n276), .A2(G222), .A3(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G77), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n276), .A2(G1698), .ZN(new_n280));
  INV_X1    g0080(.A(G223), .ZN(new_n281));
  OAI221_X1 g0081(.A(new_n278), .B1(new_n279), .B2(new_n276), .C1(new_n280), .C2(new_n281), .ZN(new_n282));
  AND2_X1   g0082(.A1(G33), .A2(G41), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n283), .A2(new_n213), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n275), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(G200), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n275), .A2(G190), .A3(new_n285), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n258), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(KEYINPUT10), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT10), .ZN(new_n291));
  NAND4_X1  g0091(.A1(new_n258), .A2(new_n287), .A3(new_n291), .A4(new_n288), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G179), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n286), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G169), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n296), .B1(new_n275), .B2(new_n285), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n257), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n293), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G68), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n252), .A2(G20), .A3(new_n301), .ZN(new_n302));
  XOR2_X1   g0102(.A(new_n302), .B(KEYINPUT12), .Z(new_n303));
  AOI21_X1  g0103(.A(new_n303), .B1(G68), .B2(new_n255), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  AOI22_X1  g0105(.A1(new_n243), .A2(G50), .B1(G20), .B2(new_n301), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n306), .B1(new_n279), .B2(new_n246), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(new_n249), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT11), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n308), .A2(new_n309), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  NOR3_X1   g0112(.A1(new_n305), .A2(new_n310), .A3(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT13), .ZN(new_n315));
  INV_X1    g0115(.A(G238), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n270), .B1(new_n272), .B2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(G33), .A2(G97), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n276), .A2(G226), .A3(new_n277), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n276), .A2(G232), .A3(G1698), .ZN(new_n321));
  OAI211_X1 g0121(.A(new_n319), .B(new_n320), .C1(new_n321), .C2(KEYINPUT70), .ZN(new_n322));
  AND2_X1   g0122(.A1(new_n321), .A2(KEYINPUT70), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n284), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n315), .B1(new_n318), .B2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n318), .A2(new_n315), .A3(new_n324), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n296), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT14), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n326), .A2(G179), .A3(new_n327), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n332), .B1(new_n328), .B2(new_n329), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n314), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(G200), .ZN(new_n335));
  INV_X1    g0135(.A(new_n327), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n335), .B1(new_n336), .B2(new_n325), .ZN(new_n337));
  INV_X1    g0137(.A(G190), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n326), .A2(new_n338), .A3(new_n327), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n314), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n276), .A2(G232), .A3(new_n277), .ZN(new_n342));
  INV_X1    g0142(.A(G107), .ZN(new_n343));
  OAI221_X1 g0143(.A(new_n342), .B1(new_n343), .B2(new_n276), .C1(new_n280), .C2(new_n316), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(new_n284), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n264), .A2(G244), .A3(new_n271), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n345), .A2(new_n270), .A3(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(G179), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n347), .A2(G169), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n245), .ZN(new_n352));
  AND2_X1   g0152(.A1(new_n243), .A2(KEYINPUT69), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n243), .A2(KEYINPUT69), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n352), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  XNOR2_X1  g0155(.A(KEYINPUT15), .B(G87), .ZN(new_n356));
  OAI221_X1 g0156(.A(new_n355), .B1(new_n207), .B2(new_n279), .C1(new_n246), .C2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(new_n249), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n253), .A2(G77), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n359), .B1(G77), .B2(new_n255), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n351), .A2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n348), .A2(new_n338), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n347), .A2(new_n335), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n361), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n363), .A2(new_n366), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n300), .A2(new_n334), .A3(new_n341), .A4(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT16), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT7), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n370), .B1(new_n276), .B2(G20), .ZN(new_n371));
  INV_X1    g0171(.A(G33), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n372), .A2(KEYINPUT3), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT3), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n374), .A2(G33), .ZN(new_n375));
  OAI211_X1 g0175(.A(KEYINPUT7), .B(new_n207), .C1(new_n373), .C2(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n301), .B1(new_n371), .B2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(G58), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n378), .A2(new_n301), .ZN(new_n379));
  OAI21_X1  g0179(.A(G20), .B1(new_n379), .B2(new_n201), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n243), .A2(G159), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n369), .B1(new_n377), .B2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT72), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  OAI21_X1  g0185(.A(KEYINPUT71), .B1(new_n372), .B2(KEYINPUT3), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT71), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n387), .A2(new_n374), .A3(G33), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n372), .A2(KEYINPUT3), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n386), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(new_n207), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(KEYINPUT7), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n390), .A2(new_n370), .A3(new_n207), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n392), .A2(G68), .A3(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n382), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n394), .A2(KEYINPUT16), .A3(new_n395), .ZN(new_n396));
  OAI211_X1 g0196(.A(KEYINPUT72), .B(new_n369), .C1(new_n377), .C2(new_n382), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n385), .A2(new_n396), .A3(new_n249), .A4(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n253), .A2(new_n245), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n399), .B1(new_n255), .B2(new_n245), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(G226), .A2(G1698), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n402), .B1(new_n281), .B2(G1698), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n403), .A2(new_n386), .A3(new_n388), .A4(new_n389), .ZN(new_n404));
  NAND2_X1  g0204(.A1(G33), .A2(G87), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(new_n284), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT68), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n408), .B1(new_n283), .B2(new_n213), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n409), .A2(G232), .A3(new_n260), .A4(new_n271), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n407), .A2(new_n270), .A3(new_n294), .A4(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n409), .A2(G274), .A3(new_n260), .ZN(new_n412));
  OR2_X1    g0212(.A1(KEYINPUT67), .A2(G41), .ZN(new_n413));
  NAND2_X1  g0213(.A1(KEYINPUT67), .A2(G41), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n413), .A2(new_n268), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(new_n206), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n410), .B1(new_n412), .B2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(new_n284), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n418), .B1(new_n404), .B2(new_n405), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n296), .B1(new_n417), .B2(new_n419), .ZN(new_n420));
  AND2_X1   g0220(.A1(new_n411), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n401), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(KEYINPUT18), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n411), .A2(new_n420), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n424), .B1(new_n398), .B2(new_n400), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT18), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n407), .A2(new_n270), .A3(G190), .A4(new_n410), .ZN(new_n428));
  OAI21_X1  g0228(.A(G200), .B1(new_n417), .B2(new_n419), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT73), .ZN(new_n430));
  AND3_X1   g0230(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n430), .B1(new_n428), .B2(new_n429), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n398), .B(new_n400), .C1(new_n431), .C2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT17), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(new_n432), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n438), .A2(KEYINPUT17), .A3(new_n398), .A4(new_n400), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n423), .A2(new_n427), .A3(new_n435), .A4(new_n439), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n368), .A2(new_n440), .ZN(new_n441));
  AND2_X1   g0241(.A1(new_n248), .A2(new_n213), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n206), .A2(G33), .ZN(new_n443));
  AND3_X1   g0243(.A1(new_n442), .A2(new_n253), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(G97), .ZN(new_n445));
  INV_X1    g0245(.A(new_n253), .ZN(new_n446));
  INV_X1    g0246(.A(G97), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n445), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n343), .A2(KEYINPUT6), .A3(G97), .ZN(new_n450));
  XOR2_X1   g0250(.A(G97), .B(G107), .Z(new_n451));
  OAI21_X1  g0251(.A(new_n450), .B1(new_n451), .B2(KEYINPUT6), .ZN(new_n452));
  AOI22_X1  g0252(.A1(new_n452), .A2(G20), .B1(G77), .B2(new_n243), .ZN(new_n453));
  AND2_X1   g0253(.A1(new_n371), .A2(new_n376), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n453), .B1(new_n454), .B2(new_n343), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n449), .B1(new_n455), .B2(new_n249), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n276), .A2(G250), .A3(G1698), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT4), .ZN(new_n458));
  INV_X1    g0258(.A(G244), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n276), .A2(new_n277), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(G33), .A2(G283), .ZN(new_n462));
  AND3_X1   g0262(.A1(new_n457), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n459), .A2(G1698), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n386), .A2(new_n388), .A3(new_n389), .A4(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT74), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n458), .B1(new_n465), .B2(new_n466), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n463), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(new_n284), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n268), .A2(G1), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT5), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n413), .A2(new_n474), .A3(new_n414), .ZN(new_n475));
  NAND2_X1  g0275(.A1(KEYINPUT5), .A2(G41), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n473), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NOR3_X1   g0277(.A1(new_n477), .A2(new_n263), .A3(new_n261), .ZN(new_n478));
  AND3_X1   g0278(.A1(new_n409), .A2(G274), .A3(new_n260), .ZN(new_n479));
  AOI22_X1  g0279(.A1(new_n478), .A2(G257), .B1(new_n479), .B2(new_n477), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n471), .A2(new_n480), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n456), .B1(new_n481), .B2(new_n338), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n457), .A2(new_n461), .A3(new_n462), .ZN(new_n483));
  AND4_X1   g0283(.A1(new_n388), .A2(new_n386), .A3(new_n389), .A4(new_n464), .ZN(new_n484));
  AOI21_X1  g0284(.A(KEYINPUT4), .B1(new_n484), .B2(KEYINPUT74), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n483), .B1(new_n485), .B2(new_n467), .ZN(new_n486));
  OAI21_X1  g0286(.A(KEYINPUT75), .B1(new_n486), .B2(new_n418), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT75), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n470), .A2(new_n488), .A3(new_n284), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n487), .A2(new_n480), .A3(new_n489), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n482), .B1(G200), .B2(new_n490), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n487), .A2(new_n294), .A3(new_n480), .A4(new_n489), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n481), .A2(new_n296), .ZN(new_n493));
  INV_X1    g0293(.A(new_n456), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n492), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT76), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n492), .A2(new_n493), .A3(KEYINPUT76), .A4(new_n494), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n491), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT79), .ZN(new_n500));
  NAND2_X1  g0300(.A1(KEYINPUT77), .A2(G116), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  NOR2_X1   g0302(.A1(KEYINPUT77), .A2(G116), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  AOI22_X1  g0304(.A1(new_n444), .A2(G116), .B1(new_n446), .B2(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(new_n503), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n207), .B1(new_n506), .B2(new_n501), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n372), .A2(G97), .ZN(new_n508));
  AOI21_X1  g0308(.A(G20), .B1(new_n508), .B2(new_n462), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n249), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT20), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n462), .B1(new_n447), .B2(G33), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(new_n207), .ZN(new_n514));
  OAI21_X1  g0314(.A(G20), .B1(new_n502), .B2(new_n503), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AOI21_X1  g0316(.A(KEYINPUT20), .B1(new_n516), .B2(new_n249), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n505), .B1(new_n512), .B2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n475), .A2(new_n476), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n472), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n521), .A2(G270), .A3(new_n264), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n479), .A2(new_n477), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n277), .A2(G257), .ZN(new_n524));
  NAND2_X1  g0324(.A1(G264), .A2(G1698), .ZN(new_n525));
  AND2_X1   g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(G303), .ZN(new_n527));
  OAI22_X1  g0327(.A1(new_n390), .A2(new_n526), .B1(new_n527), .B2(new_n276), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n284), .ZN(new_n529));
  AND3_X1   g0329(.A1(new_n522), .A2(new_n523), .A3(new_n529), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n500), .B(new_n519), .C1(new_n530), .C2(new_n335), .ZN(new_n531));
  AOI22_X1  g0331(.A1(new_n284), .A2(new_n528), .B1(new_n479), .B2(new_n477), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n335), .B1(new_n532), .B2(new_n522), .ZN(new_n533));
  OAI21_X1  g0333(.A(KEYINPUT79), .B1(new_n533), .B2(new_n518), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n522), .A2(new_n523), .A3(new_n529), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n535), .A2(new_n338), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n531), .A2(new_n534), .A3(KEYINPUT80), .A4(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n530), .A2(G179), .A3(new_n518), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n518), .A2(new_n535), .A3(KEYINPUT21), .A4(G169), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n510), .A2(new_n511), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n516), .A2(KEYINPUT20), .A3(new_n249), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n296), .B1(new_n544), .B2(new_n505), .ZN(new_n545));
  AOI21_X1  g0345(.A(KEYINPUT21), .B1(new_n545), .B2(new_n535), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n541), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n538), .A2(new_n547), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n533), .A2(new_n518), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n536), .B1(new_n549), .B2(new_n500), .ZN(new_n550));
  AOI21_X1  g0350(.A(KEYINPUT80), .B1(new_n550), .B2(new_n534), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n521), .A2(G264), .A3(new_n264), .ZN(new_n553));
  NAND2_X1  g0353(.A1(G33), .A2(G294), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n277), .A2(G250), .ZN(new_n555));
  NAND2_X1  g0355(.A1(G257), .A2(G1698), .ZN(new_n556));
  AND2_X1   g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n554), .B1(new_n390), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(new_n284), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n553), .A2(new_n523), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n335), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(KEYINPUT83), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT83), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n560), .A2(new_n563), .A3(new_n335), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n559), .A2(KEYINPUT82), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT82), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n558), .A2(new_n566), .A3(new_n284), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n565), .A2(new_n523), .A3(new_n567), .A4(new_n553), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n562), .B(new_n564), .C1(G190), .C2(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(new_n252), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT25), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n343), .A2(G20), .ZN(new_n572));
  NOR3_X1   g0372(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(KEYINPUT81), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT81), .ZN(new_n575));
  INV_X1    g0375(.A(new_n572), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n252), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n575), .B1(new_n577), .B2(new_n571), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n574), .B1(new_n573), .B2(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(new_n444), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n579), .B1(new_n343), .B2(new_n580), .ZN(new_n581));
  XNOR2_X1  g0381(.A(new_n572), .B(KEYINPUT23), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n504), .A2(new_n372), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n582), .B1(new_n207), .B2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(new_n390), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n585), .A2(KEYINPUT22), .A3(new_n207), .A4(G87), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT22), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n374), .A2(G33), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n389), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n207), .A2(G87), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n587), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n584), .A2(new_n586), .A3(KEYINPUT24), .A4(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n249), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT24), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n584), .A2(new_n591), .ZN(new_n596));
  INV_X1    g0396(.A(new_n586), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n595), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n581), .B1(new_n594), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n569), .A2(new_n599), .ZN(new_n600));
  MUX2_X1   g0400(.A(new_n316), .B(new_n459), .S(G1698), .Z(new_n601));
  NOR2_X1   g0401(.A1(new_n390), .A2(new_n601), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n284), .B1(new_n602), .B2(new_n583), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n472), .A2(G274), .ZN(new_n604));
  INV_X1    g0404(.A(G250), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n604), .B1(new_n472), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n264), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n603), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n296), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n585), .A2(new_n207), .A3(G68), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT19), .ZN(new_n611));
  INV_X1    g0411(.A(G87), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n612), .A2(new_n447), .A3(new_n343), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n319), .A2(new_n207), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n611), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NOR3_X1   g0415(.A1(new_n319), .A2(KEYINPUT19), .A3(G20), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n610), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  AOI22_X1  g0417(.A1(new_n617), .A2(new_n249), .B1(new_n446), .B2(new_n356), .ZN(new_n618));
  INV_X1    g0418(.A(new_n356), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n444), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g0420(.A(new_n620), .B(KEYINPUT78), .ZN(new_n621));
  INV_X1    g0421(.A(new_n608), .ZN(new_n622));
  AOI22_X1  g0422(.A1(new_n618), .A2(new_n621), .B1(new_n294), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n444), .A2(G87), .ZN(new_n624));
  AND2_X1   g0424(.A1(new_n618), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n335), .B1(new_n603), .B2(new_n607), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n626), .B1(new_n622), .B2(G190), .ZN(new_n627));
  AOI22_X1  g0427(.A1(new_n609), .A2(new_n623), .B1(new_n625), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n568), .A2(G169), .ZN(new_n629));
  OR2_X1    g0429(.A1(new_n560), .A2(new_n294), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AND3_X1   g0431(.A1(new_n598), .A2(new_n249), .A3(new_n592), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n631), .B1(new_n632), .B2(new_n581), .ZN(new_n633));
  AND3_X1   g0433(.A1(new_n600), .A2(new_n628), .A3(new_n633), .ZN(new_n634));
  AND4_X1   g0434(.A1(new_n441), .A2(new_n499), .A3(new_n552), .A4(new_n634), .ZN(G372));
  INV_X1    g0435(.A(new_n298), .ZN(new_n636));
  XNOR2_X1  g0436(.A(new_n425), .B(KEYINPUT18), .ZN(new_n637));
  OR2_X1    g0437(.A1(new_n331), .A2(new_n333), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n362), .A2(KEYINPUT86), .ZN(new_n639));
  OR2_X1    g0439(.A1(new_n362), .A2(KEYINPUT86), .ZN(new_n640));
  AOI22_X1  g0440(.A1(new_n638), .A2(new_n314), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  AND2_X1   g0441(.A1(new_n435), .A2(new_n439), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(new_n341), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n637), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n636), .B1(new_n644), .B2(new_n293), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n497), .A2(new_n498), .A3(new_n628), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(KEYINPUT26), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n608), .A2(KEYINPUT84), .A3(new_n296), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT84), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n609), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n623), .A2(new_n648), .A3(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n647), .A2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  AOI22_X1  g0453(.A1(new_n633), .A2(new_n547), .B1(new_n569), .B2(new_n599), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n499), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n492), .A2(new_n493), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT85), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n492), .A2(new_n493), .A3(KEYINPUT85), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n456), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT26), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  AND2_X1   g0462(.A1(new_n655), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n625), .A2(new_n627), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n653), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(new_n441), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n645), .A2(new_n667), .ZN(G369));
  INV_X1    g0468(.A(new_n547), .ZN(new_n669));
  OR3_X1    g0469(.A1(new_n570), .A2(KEYINPUT27), .A3(G20), .ZN(new_n670));
  OAI21_X1  g0470(.A(KEYINPUT27), .B1(new_n570), .B2(G20), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n670), .A2(G213), .A3(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(G343), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n518), .A2(new_n674), .ZN(new_n675));
  MUX2_X1   g0475(.A(new_n669), .B(new_n552), .S(new_n675), .Z(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(G330), .ZN(new_n677));
  INV_X1    g0477(.A(new_n674), .ZN(new_n678));
  OAI211_X1 g0478(.A(new_n600), .B(new_n633), .C1(new_n599), .C2(new_n678), .ZN(new_n679));
  OR2_X1    g0479(.A1(new_n633), .A2(new_n678), .ZN(new_n680));
  AND2_X1   g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n677), .A2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n654), .A2(new_n678), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(new_n684), .ZN(G399));
  NAND2_X1  g0485(.A1(new_n210), .A2(new_n267), .ZN(new_n686));
  NOR4_X1   g0486(.A1(G87), .A2(G97), .A3(G107), .A4(G116), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n686), .A2(G1), .A3(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n688), .B1(new_n216), .B2(new_n686), .ZN(new_n689));
  XNOR2_X1  g0489(.A(new_n689), .B(KEYINPUT28), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT90), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT29), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n497), .A2(new_n498), .ZN(new_n693));
  INV_X1    g0493(.A(new_n491), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n693), .A2(new_n654), .A3(new_n694), .A4(new_n664), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(new_n651), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n665), .A2(new_n661), .ZN(new_n697));
  AOI22_X1  g0497(.A1(new_n661), .A2(new_n646), .B1(new_n660), .B2(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n678), .B1(new_n696), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(KEYINPUT89), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT89), .ZN(new_n701));
  OAI211_X1 g0501(.A(new_n701), .B(new_n678), .C1(new_n696), .C2(new_n698), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n692), .B1(new_n700), .B2(new_n702), .ZN(new_n703));
  AOI21_X1  g0503(.A(KEYINPUT29), .B1(new_n666), .B2(new_n678), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  AOI21_X1  g0505(.A(G179), .B1(new_n603), .B2(new_n607), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT87), .ZN(new_n707));
  AND3_X1   g0507(.A1(new_n706), .A2(new_n535), .A3(new_n707), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n707), .B1(new_n706), .B2(new_n535), .ZN(new_n709));
  OAI211_X1 g0509(.A(new_n490), .B(new_n560), .C1(new_n708), .C2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT30), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n553), .A2(new_n559), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n530), .A2(new_n713), .A3(new_n622), .A4(G179), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n711), .B1(new_n714), .B2(new_n481), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n532), .A2(G179), .A3(new_n522), .ZN(new_n716));
  NOR3_X1   g0516(.A1(new_n716), .A2(new_n712), .A3(new_n608), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n717), .A2(KEYINPUT30), .A3(new_n471), .A4(new_n480), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n710), .A2(new_n715), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(KEYINPUT88), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT88), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n710), .A2(new_n721), .A3(new_n715), .A4(new_n718), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n678), .B1(new_n720), .B2(new_n722), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n499), .A2(new_n634), .A3(new_n552), .A4(new_n678), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n723), .B1(new_n724), .B2(KEYINPUT31), .ZN(new_n725));
  AND3_X1   g0525(.A1(new_n719), .A2(KEYINPUT31), .A3(new_n674), .ZN(new_n726));
  OR2_X1    g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(G330), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n691), .B1(new_n705), .B2(new_n729), .ZN(new_n730));
  OAI211_X1 g0530(.A(KEYINPUT90), .B(new_n728), .C1(new_n703), .C2(new_n704), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n690), .B1(new_n732), .B2(G1), .ZN(G364));
  NOR2_X1   g0533(.A1(new_n251), .A2(G20), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(G45), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n686), .A2(G1), .A3(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n677), .A2(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n676), .A2(G330), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(G13), .A2(G33), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n741), .A2(G20), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  OR2_X1    g0543(.A1(new_n676), .A2(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n213), .B1(G20), .B2(new_n296), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n742), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n210), .A2(new_n276), .ZN(new_n747));
  INV_X1    g0547(.A(G355), .ZN(new_n748));
  OAI22_X1  g0548(.A1(new_n747), .A2(new_n748), .B1(G116), .B2(new_n210), .ZN(new_n749));
  XNOR2_X1  g0549(.A(new_n749), .B(KEYINPUT92), .ZN(new_n750));
  AND2_X1   g0550(.A1(new_n210), .A2(new_n390), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n238), .A2(G45), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n217), .A2(new_n268), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n752), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n746), .B1(new_n750), .B2(new_n755), .ZN(new_n756));
  XOR2_X1   g0556(.A(new_n736), .B(KEYINPUT91), .Z(new_n757));
  NAND2_X1  g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n207), .A2(new_n338), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n294), .A2(G200), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(G322), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n589), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n207), .A2(G190), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n760), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(G179), .A2(G200), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n764), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  AOI22_X1  g0569(.A1(G311), .A2(new_n766), .B1(new_n769), .B2(G329), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n759), .A2(new_n294), .A3(G200), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n770), .B1(new_n527), .B2(new_n771), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n207), .B1(new_n767), .B2(G190), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  AOI211_X1 g0574(.A(new_n763), .B(new_n772), .C1(G294), .C2(new_n774), .ZN(new_n775));
  NOR3_X1   g0575(.A1(new_n207), .A2(new_n294), .A3(new_n335), .ZN(new_n776));
  XNOR2_X1  g0576(.A(new_n776), .B(KEYINPUT93), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(new_n338), .ZN(new_n778));
  XOR2_X1   g0578(.A(KEYINPUT96), .B(G326), .Z(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n777), .A2(G190), .ZN(new_n781));
  XNOR2_X1  g0581(.A(KEYINPUT33), .B(G317), .ZN(new_n782));
  AOI22_X1  g0582(.A1(new_n778), .A2(new_n780), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(G283), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n764), .A2(new_n294), .A3(G200), .ZN(new_n785));
  XNOR2_X1  g0585(.A(new_n785), .B(KEYINPUT95), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  OAI211_X1 g0587(.A(new_n775), .B(new_n783), .C1(new_n784), .C2(new_n787), .ZN(new_n788));
  XOR2_X1   g0588(.A(new_n788), .B(KEYINPUT97), .Z(new_n789));
  OAI22_X1  g0589(.A1(new_n761), .A2(new_n378), .B1(new_n765), .B2(new_n279), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n790), .B1(new_n778), .B2(G50), .ZN(new_n791));
  XNOR2_X1  g0591(.A(new_n791), .B(KEYINPUT94), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n787), .A2(new_n343), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n769), .A2(G159), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n795), .B(KEYINPUT32), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n773), .A2(new_n447), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n276), .B1(new_n771), .B2(new_n612), .ZN(new_n798));
  NOR3_X1   g0598(.A1(new_n796), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n781), .ZN(new_n800));
  OAI211_X1 g0600(.A(new_n794), .B(new_n799), .C1(new_n301), .C2(new_n800), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n789), .B1(new_n792), .B2(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n758), .B1(new_n802), .B2(new_n745), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n739), .B1(new_n744), .B2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(G396));
  INV_X1    g0605(.A(new_n757), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n745), .A2(new_n740), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n806), .B1(new_n279), .B2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n761), .ZN(new_n809));
  AOI22_X1  g0609(.A1(G143), .A2(new_n809), .B1(new_n766), .B2(G159), .ZN(new_n810));
  INV_X1    g0610(.A(new_n778), .ZN(new_n811));
  INV_X1    g0611(.A(G137), .ZN(new_n812));
  INV_X1    g0612(.A(G150), .ZN(new_n813));
  OAI221_X1 g0613(.A(new_n810), .B1(new_n811), .B2(new_n812), .C1(new_n813), .C2(new_n800), .ZN(new_n814));
  XNOR2_X1  g0614(.A(new_n814), .B(KEYINPUT34), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n786), .A2(G68), .ZN(new_n816));
  INV_X1    g0616(.A(new_n771), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n817), .A2(G50), .B1(new_n774), .B2(G58), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(G132), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n585), .B1(new_n820), .B2(new_n768), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n819), .B1(KEYINPUT98), .B2(new_n821), .ZN(new_n822));
  OAI211_X1 g0622(.A(new_n815), .B(new_n822), .C1(KEYINPUT98), .C2(new_n821), .ZN(new_n823));
  AOI22_X1  g0623(.A1(G283), .A2(new_n781), .B1(new_n778), .B2(G303), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n786), .A2(G87), .ZN(new_n825));
  INV_X1    g0625(.A(G294), .ZN(new_n826));
  OAI22_X1  g0626(.A1(new_n504), .A2(new_n765), .B1(new_n761), .B2(new_n826), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n827), .B1(G311), .B2(new_n769), .ZN(new_n828));
  AOI211_X1 g0628(.A(new_n276), .B(new_n797), .C1(G107), .C2(new_n817), .ZN(new_n829));
  NAND4_X1  g0629(.A1(new_n824), .A2(new_n825), .A3(new_n828), .A4(new_n829), .ZN(new_n830));
  AND2_X1   g0630(.A1(new_n823), .A2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n745), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n361), .A2(new_n674), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n640), .A2(new_n639), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n367), .A2(new_n833), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  OAI221_X1 g0637(.A(new_n808), .B1(new_n831), .B2(new_n832), .C1(new_n741), .C2(new_n837), .ZN(new_n838));
  XOR2_X1   g0638(.A(new_n838), .B(KEYINPUT99), .Z(new_n839));
  AOI21_X1  g0639(.A(new_n837), .B1(new_n666), .B2(new_n678), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n665), .B1(new_n655), .B2(new_n662), .ZN(new_n841));
  OAI211_X1 g0641(.A(new_n678), .B(new_n837), .C1(new_n841), .C2(new_n652), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n840), .A2(new_n843), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n844), .A2(new_n729), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n736), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n847), .B1(new_n844), .B2(new_n729), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n839), .B1(new_n846), .B2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(G384));
  OAI211_X1 g0650(.A(G116), .B(new_n214), .C1(new_n452), .C2(KEYINPUT35), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n851), .B1(KEYINPUT35), .B2(new_n452), .ZN(new_n852));
  XNOR2_X1  g0652(.A(new_n852), .B(KEYINPUT36), .ZN(new_n853));
  OR3_X1    g0653(.A1(new_n379), .A2(new_n216), .A3(new_n279), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n202), .A2(G68), .ZN(new_n855));
  AOI211_X1 g0655(.A(new_n206), .B(G13), .C1(new_n854), .C2(new_n855), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n853), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n837), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n724), .A2(KEYINPUT31), .ZN(new_n859));
  INV_X1    g0659(.A(new_n723), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n723), .A2(KEYINPUT31), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n858), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  OAI211_X1 g0663(.A(new_n314), .B(new_n674), .C1(new_n638), .C2(new_n340), .ZN(new_n864));
  OAI211_X1 g0664(.A(new_n334), .B(new_n341), .C1(new_n313), .C2(new_n678), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT38), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT37), .ZN(new_n868));
  INV_X1    g0668(.A(new_n672), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n401), .A2(new_n869), .ZN(new_n870));
  AND4_X1   g0670(.A1(new_n868), .A2(new_n422), .A3(new_n870), .A4(new_n433), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n396), .A2(new_n249), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n301), .B1(new_n391), .B2(KEYINPUT7), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n382), .B1(new_n873), .B2(new_n393), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n874), .A2(KEYINPUT16), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n400), .B1(new_n872), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n424), .A2(new_n672), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  AOI211_X1 g0678(.A(KEYINPUT101), .B(new_n868), .C1(new_n878), .C2(new_n433), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT101), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n431), .A2(new_n432), .ZN(new_n881));
  INV_X1    g0681(.A(new_n400), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n442), .B1(new_n874), .B2(KEYINPUT16), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n394), .A2(new_n395), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(new_n369), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n882), .B1(new_n883), .B2(new_n885), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n421), .A2(new_n869), .ZN(new_n887));
  OAI22_X1  g0687(.A1(new_n401), .A2(new_n881), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n880), .B1(new_n888), .B2(KEYINPUT37), .ZN(new_n889));
  NOR3_X1   g0689(.A1(new_n871), .A2(new_n879), .A3(new_n889), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n886), .A2(new_n672), .ZN(new_n891));
  AND2_X1   g0691(.A1(new_n440), .A2(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n867), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n888), .A2(KEYINPUT37), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(KEYINPUT101), .ZN(new_n895));
  INV_X1    g0695(.A(new_n401), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n425), .B1(new_n896), .B2(new_n438), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n897), .A2(new_n868), .A3(new_n870), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n888), .A2(new_n880), .A3(KEYINPUT37), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n895), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n440), .A2(new_n891), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n900), .A2(new_n901), .A3(KEYINPUT38), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n893), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n863), .A2(new_n866), .A3(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT40), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  AND3_X1   g0706(.A1(new_n900), .A2(new_n901), .A3(KEYINPUT38), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n440), .A2(new_n401), .A3(new_n869), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n422), .A2(new_n870), .A3(new_n433), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(KEYINPUT37), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n898), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(KEYINPUT38), .B1(new_n908), .B2(new_n911), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n907), .A2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  NAND4_X1  g0714(.A1(new_n914), .A2(new_n863), .A3(KEYINPUT40), .A4(new_n866), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n906), .A2(new_n915), .ZN(new_n916));
  AND2_X1   g0716(.A1(new_n723), .A2(KEYINPUT31), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n441), .B1(new_n725), .B2(new_n917), .ZN(new_n918));
  XOR2_X1   g0718(.A(new_n916), .B(new_n918), .Z(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(G330), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n700), .A2(new_n702), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(KEYINPUT29), .ZN(new_n922));
  INV_X1    g0722(.A(new_n704), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n922), .A2(new_n923), .A3(new_n441), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(new_n645), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n362), .A2(new_n674), .ZN(new_n926));
  XOR2_X1   g0726(.A(new_n926), .B(KEYINPUT100), .Z(new_n927));
  NAND2_X1  g0727(.A1(new_n842), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n928), .A2(new_n866), .A3(new_n903), .ZN(new_n929));
  OR2_X1    g0729(.A1(new_n637), .A2(new_n869), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n868), .B1(new_n897), .B2(new_n870), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n931), .A2(new_n871), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n870), .B1(new_n642), .B2(new_n637), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n867), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT102), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n935), .A2(KEYINPUT39), .ZN(new_n936));
  AND3_X1   g0736(.A1(new_n934), .A2(new_n902), .A3(new_n936), .ZN(new_n937));
  OAI211_X1 g0737(.A(new_n893), .B(new_n902), .C1(KEYINPUT102), .C2(new_n912), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n937), .B1(new_n938), .B2(KEYINPUT39), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n334), .A2(new_n674), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  OAI211_X1 g0741(.A(new_n929), .B(new_n930), .C1(new_n939), .C2(new_n941), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n925), .B(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n920), .A2(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n944), .B1(new_n206), .B2(new_n734), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n920), .A2(new_n943), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n857), .B1(new_n945), .B2(new_n946), .ZN(G367));
  OAI21_X1  g0747(.A(new_n746), .B1(new_n210), .B2(new_n356), .ZN(new_n948));
  INV_X1    g0748(.A(new_n234), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n948), .B1(new_n949), .B2(new_n751), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n950), .A2(new_n806), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n774), .A2(G68), .ZN(new_n952));
  OAI211_X1 g0752(.A(new_n952), .B(new_n276), .C1(new_n378), .C2(new_n771), .ZN(new_n953));
  OAI22_X1  g0753(.A1(new_n761), .A2(new_n813), .B1(new_n768), .B2(new_n812), .ZN(new_n954));
  OAI22_X1  g0754(.A1(new_n785), .A2(new_n279), .B1(new_n765), .B2(new_n202), .ZN(new_n955));
  NOR3_X1   g0755(.A1(new_n953), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(G143), .ZN(new_n957));
  INV_X1    g0757(.A(G159), .ZN(new_n958));
  OAI221_X1 g0758(.A(new_n956), .B1(new_n811), .B2(new_n957), .C1(new_n958), .C2(new_n800), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n506), .A2(new_n501), .ZN(new_n960));
  AOI21_X1  g0760(.A(KEYINPUT46), .B1(new_n817), .B2(new_n960), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n961), .B1(G107), .B2(new_n774), .ZN(new_n962));
  AND3_X1   g0762(.A1(new_n817), .A2(KEYINPUT46), .A3(G116), .ZN(new_n963));
  OAI22_X1  g0763(.A1(new_n447), .A2(new_n785), .B1(new_n761), .B2(new_n527), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  AOI22_X1  g0765(.A1(G283), .A2(new_n766), .B1(new_n769), .B2(G317), .ZN(new_n966));
  NAND4_X1  g0766(.A1(new_n962), .A2(new_n390), .A3(new_n965), .A4(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(G311), .ZN(new_n968));
  OAI22_X1  g0768(.A1(new_n826), .A2(new_n800), .B1(new_n811), .B2(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n959), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT47), .ZN(new_n971));
  AND2_X1   g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n745), .B1(new_n970), .B2(new_n971), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n625), .A2(new_n678), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n651), .B1(new_n665), .B2(new_n974), .ZN(new_n975));
  OR2_X1    g0775(.A1(new_n651), .A2(new_n974), .ZN(new_n976));
  AND2_X1   g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  OAI221_X1 g0777(.A(new_n951), .B1(new_n972), .B2(new_n973), .C1(new_n977), .C2(new_n743), .ZN(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n499), .B1(new_n456), .B2(new_n678), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n660), .A2(new_n674), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n669), .A2(new_n678), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n679), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n985), .A2(KEYINPUT42), .ZN(new_n986));
  XOR2_X1   g0786(.A(new_n986), .B(KEYINPUT103), .Z(new_n987));
  INV_X1    g0787(.A(new_n982), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n693), .B1(new_n988), .B2(new_n633), .ZN(new_n989));
  AOI22_X1  g0789(.A1(new_n989), .A2(new_n678), .B1(KEYINPUT42), .B2(new_n985), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n987), .A2(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(new_n977), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT43), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n977), .A2(KEYINPUT43), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n991), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  NAND4_X1  g0796(.A1(new_n987), .A2(new_n993), .A3(new_n992), .A4(new_n990), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n683), .A2(new_n988), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n998), .B(new_n999), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n686), .B(KEYINPUT41), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n982), .A2(new_n684), .ZN(new_n1002));
  XOR2_X1   g0802(.A(new_n1002), .B(KEYINPUT45), .Z(new_n1003));
  NOR2_X1   g0803(.A1(new_n982), .A2(new_n684), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT44), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1006), .A2(new_n682), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1003), .A2(new_n683), .A3(new_n1005), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT105), .ZN(new_n1011));
  AND2_X1   g0811(.A1(new_n681), .A2(new_n983), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n677), .A2(KEYINPUT104), .B1(new_n1012), .B2(new_n984), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n677), .A2(KEYINPUT104), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1013), .B(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n1015), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1011), .B1(new_n732), .B2(new_n1016), .ZN(new_n1017));
  AOI211_X1 g0817(.A(KEYINPUT105), .B(new_n1015), .C1(new_n730), .C2(new_n731), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1010), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1001), .B1(new_n1019), .B2(new_n732), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n735), .A2(G1), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1000), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(KEYINPUT106), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  OAI211_X1 g0824(.A(KEYINPUT106), .B(new_n1000), .C1(new_n1020), .C2(new_n1021), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n979), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  OR2_X1    g0826(.A1(new_n1026), .A2(KEYINPUT107), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1026), .A2(KEYINPUT107), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n1029), .ZN(G387));
  NAND2_X1  g0830(.A1(new_n922), .A2(new_n923), .ZN(new_n1031));
  AOI21_X1  g0831(.A(KEYINPUT90), .B1(new_n1031), .B2(new_n728), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n731), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1016), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n686), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n730), .A2(new_n731), .A3(new_n1015), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1034), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  INV_X1    g0837(.A(KEYINPUT108), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n268), .B1(new_n301), .B2(new_n279), .C1(new_n687), .C2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1039), .B1(new_n1038), .B2(new_n687), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n245), .A2(G50), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(KEYINPUT109), .B(KEYINPUT50), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1041), .B(new_n1042), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n752), .B1(new_n1040), .B2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1044), .B1(new_n230), .B2(new_n268), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n1045), .B1(G107), .B2(new_n210), .C1(new_n687), .C2(new_n747), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n806), .B1(new_n1046), .B2(new_n746), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n585), .B1(new_n356), .B2(new_n773), .ZN(new_n1048));
  XOR2_X1   g0848(.A(KEYINPUT110), .B(G150), .Z(new_n1049));
  OAI22_X1  g0849(.A1(new_n1049), .A2(new_n768), .B1(new_n761), .B2(new_n202), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n771), .A2(new_n279), .B1(new_n765), .B2(new_n301), .ZN(new_n1051));
  OR3_X1    g0851(.A1(new_n1048), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n958), .A2(new_n811), .B1(new_n800), .B2(new_n245), .ZN(new_n1053));
  AOI211_X1 g0853(.A(new_n1052), .B(new_n1053), .C1(G97), .C2(new_n786), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n504), .A2(new_n785), .B1(new_n779), .B2(new_n768), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n817), .A2(G294), .B1(new_n774), .B2(G283), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(G317), .A2(new_n809), .B1(new_n766), .B2(G303), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n1057), .B1(new_n811), .B2(new_n762), .C1(new_n968), .C2(new_n800), .ZN(new_n1058));
  INV_X1    g0858(.A(KEYINPUT48), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1056), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1060), .B1(new_n1059), .B2(new_n1058), .ZN(new_n1061));
  AOI211_X1 g0861(.A(new_n585), .B(new_n1055), .C1(new_n1061), .C2(KEYINPUT49), .ZN(new_n1062));
  OR2_X1    g0862(.A1(new_n1061), .A2(KEYINPUT49), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1054), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1047), .B1(new_n1064), .B2(new_n832), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1065), .B1(new_n681), .B2(new_n742), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(new_n1016), .B2(new_n1021), .ZN(new_n1067));
  AOI21_X1  g0867(.A(KEYINPUT111), .B1(new_n1037), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n1068), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1037), .A2(KEYINPUT111), .A3(new_n1067), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1069), .A2(new_n1070), .ZN(G393));
  AOI21_X1  g0871(.A(new_n686), .B1(new_n1034), .B2(new_n1009), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1019), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n988), .A2(new_n742), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n746), .B1(new_n447), .B2(new_n210), .C1(new_n752), .C2(new_n241), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n757), .A2(new_n1075), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT112), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n778), .A2(G317), .B1(G311), .B2(new_n809), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(new_n1078), .B(KEYINPUT52), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n781), .A2(G303), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n774), .A2(new_n960), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n765), .A2(new_n826), .B1(new_n768), .B2(new_n762), .ZN(new_n1082));
  AOI211_X1 g0882(.A(new_n276), .B(new_n1082), .C1(G283), .C2(new_n817), .ZN(new_n1083));
  NAND4_X1  g0883(.A1(new_n794), .A2(new_n1080), .A3(new_n1081), .A4(new_n1083), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n778), .A2(G150), .B1(G159), .B2(new_n809), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1085), .B(KEYINPUT51), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n817), .A2(G68), .B1(new_n766), .B2(new_n352), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1087), .B1(new_n957), .B2(new_n768), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n773), .A2(new_n279), .ZN(new_n1089));
  NOR3_X1   g0889(.A1(new_n1088), .A2(new_n390), .A3(new_n1089), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n1090), .B(new_n825), .C1(new_n202), .C2(new_n800), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n1079), .A2(new_n1084), .B1(new_n1086), .B2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1077), .B1(new_n745), .B2(new_n1092), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n1010), .A2(new_n1021), .B1(new_n1074), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1073), .A2(new_n1094), .ZN(G390));
  NAND2_X1  g0895(.A1(new_n938), .A2(KEYINPUT39), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n937), .ZN(new_n1097));
  AND2_X1   g0897(.A1(new_n864), .A2(new_n865), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1098), .B1(new_n842), .B2(new_n927), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n1096), .B(new_n1097), .C1(new_n1099), .C2(new_n940), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n646), .A2(new_n661), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n660), .A2(new_n697), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1103), .A2(new_n651), .A3(new_n695), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n701), .B1(new_n1104), .B2(new_n678), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n702), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n837), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n926), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1098), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n913), .A2(new_n940), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1100), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n863), .A2(KEYINPUT113), .A3(new_n866), .A4(G330), .ZN(new_n1113));
  INV_X1    g0913(.A(KEYINPUT113), .ZN(new_n1114));
  OAI211_X1 g0914(.A(G330), .B(new_n837), .C1(new_n725), .C2(new_n917), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1114), .B1(new_n1115), .B2(new_n1098), .ZN(new_n1116));
  AND2_X1   g0916(.A1(new_n1113), .A2(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1112), .A2(new_n1118), .ZN(new_n1119));
  OAI211_X1 g0919(.A(G330), .B(new_n837), .C1(new_n725), .C2(new_n726), .ZN(new_n1120));
  OR2_X1    g0920(.A1(new_n1120), .A2(new_n1098), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1100), .B(new_n1121), .C1(new_n1109), .C2(new_n1111), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1119), .A2(new_n1122), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n441), .B(G330), .C1(new_n725), .C2(new_n917), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(new_n1124), .B(KEYINPUT114), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1125), .A2(new_n924), .A3(new_n645), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1120), .A2(new_n1098), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1113), .A2(new_n1116), .A3(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1129), .A2(new_n928), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n926), .B1(new_n921), .B2(new_n837), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1115), .A2(new_n1098), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1131), .A2(new_n1121), .A3(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1130), .A2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1127), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1123), .A2(new_n1135), .ZN(new_n1136));
  NAND4_X1  g0936(.A1(new_n1119), .A2(new_n1127), .A3(new_n1134), .A4(new_n1122), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1136), .A2(new_n1035), .A3(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1122), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1110), .B1(new_n1131), .B2(new_n1098), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1117), .B1(new_n1140), .B2(new_n1100), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1142), .A2(new_n1021), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n939), .A2(new_n740), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n806), .B1(new_n245), .B2(new_n807), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(KEYINPUT54), .B(G143), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(new_n809), .A2(G132), .B1(new_n766), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(G125), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1148), .B1(new_n1149), .B2(new_n768), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n771), .A2(new_n1049), .ZN(new_n1151));
  INV_X1    g0951(.A(KEYINPUT53), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1153), .B1(new_n958), .B2(new_n773), .ZN(new_n1154));
  OAI221_X1 g0954(.A(new_n276), .B1(new_n202), .B2(new_n785), .C1(new_n1151), .C2(new_n1152), .ZN(new_n1155));
  NOR3_X1   g0955(.A1(new_n1150), .A2(new_n1154), .A3(new_n1155), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(G128), .A2(new_n778), .B1(new_n781), .B2(G137), .ZN(new_n1157));
  AOI211_X1 g0957(.A(new_n276), .B(new_n1089), .C1(G87), .C2(new_n817), .ZN(new_n1158));
  INV_X1    g0958(.A(G116), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n761), .A2(new_n1159), .B1(new_n765), .B2(new_n447), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1160), .B1(G294), .B2(new_n769), .ZN(new_n1161));
  AND3_X1   g0961(.A1(new_n1158), .A2(new_n816), .A3(new_n1161), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(G107), .A2(new_n781), .B1(new_n778), .B2(G283), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n1156), .A2(new_n1157), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  OAI211_X1 g0964(.A(new_n1144), .B(new_n1145), .C1(new_n832), .C2(new_n1164), .ZN(new_n1165));
  AND3_X1   g0965(.A1(new_n1143), .A2(KEYINPUT115), .A3(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(KEYINPUT115), .B1(new_n1143), .B2(new_n1165), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1138), .B1(new_n1166), .B2(new_n1167), .ZN(G378));
  INV_X1    g0968(.A(KEYINPUT119), .ZN(new_n1169));
  XOR2_X1   g0969(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n257), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1172), .A2(new_n672), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT118), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n299), .A2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n299), .A2(new_n1174), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1173), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1176), .A2(new_n1173), .A3(new_n1177), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1171), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1180), .ZN(new_n1182));
  NOR3_X1   g0982(.A1(new_n1182), .A2(new_n1178), .A3(new_n1170), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n1181), .A2(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n942), .A2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(KEYINPUT39), .ZN(new_n1187));
  AOI21_X1  g0987(.A(KEYINPUT38), .B1(new_n900), .B2(new_n901), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n907), .A2(new_n1188), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n934), .A2(new_n935), .A3(new_n902), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1187), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n940), .B1(new_n1191), .B2(new_n937), .ZN(new_n1192));
  NAND4_X1  g0992(.A1(new_n1192), .A2(new_n929), .A3(new_n1184), .A4(new_n930), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1186), .A2(new_n1193), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n906), .A2(G330), .A3(new_n915), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1194), .A2(new_n1196), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1186), .A2(new_n1195), .A3(new_n1193), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(new_n1137), .A2(new_n1127), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1169), .B1(new_n1199), .B2(KEYINPUT57), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n686), .B1(new_n1199), .B2(KEYINPUT57), .ZN(new_n1201));
  INV_X1    g1001(.A(KEYINPUT57), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1126), .B1(new_n1142), .B2(new_n1134), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1198), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1195), .B1(new_n1186), .B2(new_n1193), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  OAI211_X1 g1006(.A(KEYINPUT119), .B(new_n1202), .C1(new_n1203), .C2(new_n1206), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1200), .A2(new_n1201), .A3(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1184), .A2(new_n740), .ZN(new_n1209));
  NOR3_X1   g1009(.A1(new_n745), .A2(G50), .A3(new_n740), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(G107), .A2(new_n809), .B1(new_n769), .B2(G283), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1211), .B1(new_n356), .B2(new_n765), .ZN(new_n1212));
  OAI221_X1 g1012(.A(new_n952), .B1(new_n378), .B2(new_n785), .C1(new_n279), .C2(new_n771), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n390), .A2(new_n267), .ZN(new_n1214));
  NOR3_X1   g1014(.A1(new_n1212), .A2(new_n1213), .A3(new_n1214), .ZN(new_n1215));
  OAI221_X1 g1015(.A(new_n1215), .B1(new_n447), .B2(new_n800), .C1(new_n1159), .C2(new_n811), .ZN(new_n1216));
  XOR2_X1   g1016(.A(new_n1216), .B(KEYINPUT116), .Z(new_n1217));
  OR2_X1    g1017(.A1(new_n1217), .A2(KEYINPUT58), .ZN(new_n1218));
  OAI211_X1 g1018(.A(new_n1214), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1219));
  INV_X1    g1019(.A(G128), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n761), .A2(new_n1220), .B1(new_n765), .B2(new_n812), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n771), .A2(new_n1146), .ZN(new_n1222));
  XNOR2_X1  g1022(.A(new_n1222), .B(KEYINPUT117), .ZN(new_n1223));
  AOI211_X1 g1023(.A(new_n1221), .B(new_n1223), .C1(G150), .C2(new_n774), .ZN(new_n1224));
  OAI221_X1 g1024(.A(new_n1224), .B1(new_n1149), .B2(new_n811), .C1(new_n820), .C2(new_n800), .ZN(new_n1225));
  OR2_X1    g1025(.A1(new_n1225), .A2(KEYINPUT59), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1225), .A2(KEYINPUT59), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(G33), .A2(G41), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1228), .B1(new_n785), .B2(new_n958), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1229), .B1(G124), .B2(new_n769), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1226), .A2(new_n1227), .A3(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1217), .A2(KEYINPUT58), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n1218), .A2(new_n1219), .A3(new_n1231), .A4(new_n1232), .ZN(new_n1233));
  AOI211_X1 g1033(.A(new_n736), .B(new_n1210), .C1(new_n1233), .C2(new_n745), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1209), .A2(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1021), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1235), .B1(new_n1206), .B2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1208), .A2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT120), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1208), .A2(KEYINPUT120), .A3(new_n1238), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(G375));
  INV_X1    g1044(.A(new_n1001), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1126), .A2(new_n1130), .A3(new_n1133), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1135), .A2(new_n1245), .A3(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1098), .A2(new_n740), .ZN(new_n1248));
  XNOR2_X1  g1048(.A(new_n1248), .B(KEYINPUT121), .ZN(new_n1249));
  OAI221_X1 g1049(.A(new_n589), .B1(new_n768), .B2(new_n527), .C1(new_n356), .C2(new_n773), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(new_n817), .A2(G97), .B1(new_n766), .B2(G107), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1251), .B1(new_n784), .B2(new_n761), .ZN(new_n1252));
  AOI211_X1 g1052(.A(new_n1250), .B(new_n1252), .C1(G77), .C2(new_n786), .ZN(new_n1253));
  AOI22_X1  g1053(.A1(G294), .A2(new_n778), .B1(new_n781), .B2(new_n960), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(new_n817), .A2(G159), .B1(new_n769), .B2(G128), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1255), .B1(new_n813), .B2(new_n765), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n773), .A2(new_n202), .ZN(new_n1257));
  OAI22_X1  g1057(.A1(new_n378), .A2(new_n785), .B1(new_n761), .B2(new_n812), .ZN(new_n1258));
  NOR4_X1   g1058(.A1(new_n1256), .A2(new_n390), .A3(new_n1257), .A4(new_n1258), .ZN(new_n1259));
  AOI22_X1  g1059(.A1(G132), .A2(new_n778), .B1(new_n781), .B2(new_n1147), .ZN(new_n1260));
  AOI22_X1  g1060(.A1(new_n1253), .A2(new_n1254), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1261), .A2(new_n832), .ZN(new_n1262));
  AOI211_X1 g1062(.A(new_n806), .B(new_n1262), .C1(new_n301), .C2(new_n807), .ZN(new_n1263));
  AOI22_X1  g1063(.A1(new_n1134), .A2(new_n1021), .B1(new_n1249), .B2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1247), .A2(new_n1264), .ZN(G381));
  AND3_X1   g1065(.A1(new_n1138), .A2(new_n1143), .A3(new_n1165), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1243), .A2(KEYINPUT123), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT123), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1241), .A2(new_n1269), .A3(new_n1242), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1267), .B1(new_n1268), .B2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1070), .ZN(new_n1272));
  NOR3_X1   g1072(.A1(new_n1272), .A2(G396), .A3(new_n1068), .ZN(new_n1273));
  AOI21_X1  g1073(.A(KEYINPUT122), .B1(new_n1273), .B2(new_n849), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1069), .A2(new_n804), .A3(new_n1070), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT122), .ZN(new_n1276));
  NOR3_X1   g1076(.A1(new_n1275), .A2(new_n1276), .A3(G384), .ZN(new_n1277));
  OR2_X1    g1077(.A1(G390), .A2(G381), .ZN(new_n1278));
  OR3_X1    g1078(.A1(new_n1274), .A2(new_n1277), .A3(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1279), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1280));
  AND3_X1   g1080(.A1(new_n1271), .A2(KEYINPUT124), .A3(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(KEYINPUT124), .B1(new_n1271), .B2(new_n1280), .ZN(new_n1282));
  OR2_X1    g1082(.A1(new_n1281), .A2(new_n1282), .ZN(G407));
  INV_X1    g1083(.A(G213), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1284), .B1(new_n1271), .B2(new_n673), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1285), .B1(new_n1281), .B2(new_n1282), .ZN(G409));
  AND3_X1   g1086(.A1(new_n1073), .A2(KEYINPUT107), .A3(new_n1094), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n804), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1287), .B1(new_n1288), .B2(new_n1273), .ZN(new_n1289));
  OAI21_X1  g1089(.A(G396), .B1(new_n1272), .B2(new_n1068), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1290), .A2(new_n1275), .A3(G390), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1289), .A2(new_n1291), .ZN(new_n1292));
  AND2_X1   g1092(.A1(new_n1026), .A2(new_n1292), .ZN(new_n1293));
  NOR2_X1   g1093(.A1(new_n1026), .A2(new_n1292), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1295));
  XOR2_X1   g1095(.A(KEYINPUT127), .B(KEYINPUT62), .Z(new_n1296));
  NOR2_X1   g1096(.A1(new_n1284), .A2(G343), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1208), .A2(G378), .A3(new_n1238), .ZN(new_n1298));
  NOR3_X1   g1098(.A1(new_n1203), .A2(new_n1206), .A3(new_n1001), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1266), .B1(new_n1237), .B2(new_n1299), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1297), .B1(new_n1298), .B2(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1135), .A2(new_n1035), .ZN(new_n1302));
  OR2_X1    g1102(.A1(new_n1246), .A2(KEYINPUT60), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1246), .A2(KEYINPUT60), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1302), .B1(new_n1303), .B2(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1264), .ZN(new_n1306));
  OR3_X1    g1106(.A1(new_n1305), .A2(new_n849), .A3(new_n1306), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n849), .B1(new_n1305), .B2(new_n1306), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1309), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1296), .B1(new_n1301), .B2(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT126), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1298), .A2(new_n1300), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1297), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1312), .B1(new_n1313), .B2(new_n1314), .ZN(new_n1315));
  AOI211_X1 g1115(.A(KEYINPUT126), .B(new_n1297), .C1(new_n1298), .C2(new_n1300), .ZN(new_n1316));
  NOR2_X1   g1116(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1317));
  AND2_X1   g1117(.A1(new_n1310), .A2(KEYINPUT62), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1311), .B1(new_n1317), .B2(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1297), .A2(G2897), .ZN(new_n1320));
  OR2_X1    g1120(.A1(new_n1309), .A2(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1309), .A2(new_n1320), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1321), .A2(new_n1322), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1323), .B1(new_n1315), .B2(new_n1316), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT61), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1324), .A2(new_n1325), .ZN(new_n1326));
  OAI21_X1  g1126(.A(new_n1295), .B1(new_n1319), .B2(new_n1326), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n1325), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n1301), .B1(new_n1321), .B2(new_n1322), .ZN(new_n1329));
  NOR2_X1   g1129(.A1(new_n1328), .A2(new_n1329), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT63), .ZN(new_n1331));
  INV_X1    g1131(.A(new_n1301), .ZN(new_n1332));
  OAI21_X1  g1132(.A(new_n1331), .B1(new_n1332), .B2(new_n1309), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1333), .A2(KEYINPUT125), .ZN(new_n1334));
  NOR2_X1   g1134(.A1(new_n1309), .A2(new_n1331), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1317), .A2(new_n1335), .ZN(new_n1336));
  INV_X1    g1136(.A(KEYINPUT125), .ZN(new_n1337));
  OAI211_X1 g1137(.A(new_n1337), .B(new_n1331), .C1(new_n1332), .C2(new_n1309), .ZN(new_n1338));
  NAND4_X1  g1138(.A1(new_n1330), .A2(new_n1334), .A3(new_n1336), .A4(new_n1338), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1327), .A2(new_n1339), .ZN(G405));
  NAND2_X1  g1140(.A1(new_n1295), .A2(new_n1310), .ZN(new_n1341));
  OAI21_X1  g1141(.A(new_n1298), .B1(new_n1243), .B2(new_n1267), .ZN(new_n1342));
  OAI21_X1  g1142(.A(new_n1309), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1343));
  AND3_X1   g1143(.A1(new_n1341), .A2(new_n1342), .A3(new_n1343), .ZN(new_n1344));
  AOI21_X1  g1144(.A(new_n1342), .B1(new_n1341), .B2(new_n1343), .ZN(new_n1345));
  NOR2_X1   g1145(.A1(new_n1344), .A2(new_n1345), .ZN(G402));
endmodule


