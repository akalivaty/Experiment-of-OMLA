//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 0 0 1 0 0 1 0 1 1 1 0 0 0 1 1 1 1 1 1 0 1 1 1 0 1 0 0 1 0 1 0 0 0 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 0 1 0 0 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:24 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n594, new_n595,
    new_n596, new_n597, new_n598, new_n599, new_n601, new_n602, new_n603,
    new_n604, new_n605, new_n606, new_n607, new_n608, new_n609, new_n610,
    new_n611, new_n612, new_n613, new_n614, new_n615, new_n616, new_n617,
    new_n618, new_n619, new_n620, new_n621, new_n622, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n663,
    new_n664, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n714, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G104), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n189), .A2(G107), .ZN(new_n190));
  AND2_X1   g004(.A1(KEYINPUT81), .A2(KEYINPUT3), .ZN(new_n191));
  NOR2_X1   g005(.A1(KEYINPUT81), .A2(KEYINPUT3), .ZN(new_n192));
  OAI21_X1  g006(.A(new_n190), .B1(new_n191), .B2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G107), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n194), .A2(G104), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  OAI211_X1 g010(.A(new_n193), .B(new_n196), .C1(new_n190), .C2(new_n192), .ZN(new_n197));
  OR2_X1    g011(.A1(new_n197), .A2(G101), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(G101), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n198), .A2(KEYINPUT4), .A3(new_n199), .ZN(new_n200));
  XNOR2_X1  g014(.A(new_n200), .B(KEYINPUT82), .ZN(new_n201));
  OR2_X1    g015(.A1(new_n199), .A2(KEYINPUT4), .ZN(new_n202));
  AND2_X1   g016(.A1(KEYINPUT66), .A2(G119), .ZN(new_n203));
  NOR2_X1   g017(.A1(KEYINPUT66), .A2(G119), .ZN(new_n204));
  OAI21_X1  g018(.A(G116), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G116), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G119), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  XNOR2_X1  g022(.A(KEYINPUT2), .B(G113), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  XOR2_X1   g024(.A(KEYINPUT2), .B(G113), .Z(new_n211));
  NAND3_X1  g025(.A1(new_n211), .A2(new_n205), .A3(new_n207), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n201), .A2(new_n202), .A3(new_n213), .ZN(new_n214));
  OAI21_X1  g028(.A(G101), .B1(new_n190), .B2(new_n195), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n198), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(KEYINPUT83), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT83), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n205), .A2(KEYINPUT5), .A3(new_n207), .ZN(new_n221));
  OAI211_X1 g035(.A(new_n221), .B(G113), .C1(KEYINPUT5), .C2(new_n205), .ZN(new_n222));
  OR2_X1    g036(.A1(new_n222), .A2(KEYINPUT88), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(KEYINPUT88), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n223), .A2(new_n212), .A3(new_n224), .ZN(new_n225));
  OR2_X1    g039(.A1(new_n220), .A2(new_n225), .ZN(new_n226));
  XOR2_X1   g040(.A(G110), .B(G122), .Z(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n214), .A2(new_n226), .A3(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(KEYINPUT6), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n228), .B1(new_n214), .B2(new_n226), .ZN(new_n231));
  OR2_X1    g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(G146), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(G143), .ZN(new_n234));
  INV_X1    g048(.A(G143), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G146), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  NOR2_X1   g051(.A1(KEYINPUT0), .A2(G128), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT0), .ZN(new_n239));
  INV_X1    g053(.A(G128), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n237), .B1(new_n238), .B2(new_n241), .ZN(new_n242));
  OAI211_X1 g056(.A(new_n234), .B(new_n236), .C1(new_n239), .C2(new_n240), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G125), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n240), .A2(KEYINPUT1), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n246), .A2(new_n234), .A3(new_n236), .ZN(new_n247));
  OAI211_X1 g061(.A(new_n235), .B(G146), .C1(new_n240), .C2(KEYINPUT1), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n240), .A2(new_n233), .A3(G143), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n247), .A2(new_n248), .A3(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n245), .B1(G125), .B2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(G953), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G224), .ZN(new_n254));
  XNOR2_X1  g068(.A(new_n252), .B(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT6), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n231), .A2(new_n256), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n257), .A2(KEYINPUT89), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT89), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n259), .B1(new_n231), .B2(new_n256), .ZN(new_n260));
  OAI211_X1 g074(.A(new_n232), .B(new_n255), .C1(new_n258), .C2(new_n260), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n252), .B1(KEYINPUT7), .B2(new_n254), .ZN(new_n262));
  AND3_X1   g076(.A1(new_n252), .A2(KEYINPUT7), .A3(new_n254), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT90), .ZN(new_n264));
  OR2_X1    g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n263), .A2(new_n264), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n262), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n219), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n268), .B1(new_n216), .B2(KEYINPUT83), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n222), .A2(new_n212), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  XOR2_X1   g085(.A(new_n227), .B(KEYINPUT8), .Z(new_n272));
  OAI211_X1 g086(.A(new_n271), .B(new_n272), .C1(new_n269), .C2(new_n225), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n229), .A2(new_n267), .A3(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(G902), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(KEYINPUT91), .ZN(new_n277));
  OR2_X1    g091(.A1(new_n276), .A2(KEYINPUT91), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n261), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(G210), .B1(G237), .B2(G902), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  NAND4_X1  g096(.A1(new_n261), .A2(new_n277), .A3(new_n280), .A4(new_n278), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n188), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(KEYINPUT76), .A2(G125), .ZN(new_n285));
  OAI21_X1  g099(.A(KEYINPUT77), .B1(new_n285), .B2(G140), .ZN(new_n286));
  INV_X1    g100(.A(G125), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(G140), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n285), .A2(KEYINPUT77), .A3(G140), .ZN(new_n290));
  AND3_X1   g104(.A1(new_n289), .A2(KEYINPUT16), .A3(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT78), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  OR2_X1    g107(.A1(new_n287), .A2(G140), .ZN(new_n294));
  OAI21_X1  g108(.A(KEYINPUT78), .B1(new_n294), .B2(KEYINPUT16), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n293), .B1(new_n291), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(G146), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n296), .A2(G146), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NOR2_X1   g114(.A1(G237), .A2(G953), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(G214), .ZN(new_n302));
  XNOR2_X1  g116(.A(new_n302), .B(G143), .ZN(new_n303));
  INV_X1    g117(.A(G131), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(KEYINPUT17), .ZN(new_n306));
  XNOR2_X1  g120(.A(new_n303), .B(new_n304), .ZN(new_n307));
  OAI211_X1 g121(.A(new_n300), .B(new_n306), .C1(KEYINPUT17), .C2(new_n307), .ZN(new_n308));
  XNOR2_X1  g122(.A(G113), .B(G122), .ZN(new_n309));
  XNOR2_X1  g123(.A(new_n309), .B(KEYINPUT92), .ZN(new_n310));
  XNOR2_X1  g124(.A(new_n310), .B(G104), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n294), .A2(new_n233), .A3(new_n288), .ZN(new_n312));
  XNOR2_X1  g126(.A(new_n312), .B(KEYINPUT79), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n289), .A2(new_n290), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n314), .B1(new_n233), .B2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT18), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n303), .B1(new_n318), .B2(new_n304), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n305), .A2(KEYINPUT18), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n317), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n308), .A2(new_n311), .A3(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT19), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n294), .A2(new_n323), .A3(new_n288), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n324), .B1(new_n316), .B2(new_n323), .ZN(new_n325));
  OAI211_X1 g139(.A(new_n297), .B(new_n307), .C1(G146), .C2(new_n325), .ZN(new_n326));
  AND2_X1   g140(.A1(new_n326), .A2(new_n321), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n322), .B1(new_n311), .B2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(G475), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n328), .A2(new_n329), .A3(new_n275), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT20), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(new_n322), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n311), .B1(new_n308), .B2(new_n321), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n275), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(G475), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n328), .A2(KEYINPUT20), .A3(new_n329), .A4(new_n275), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n332), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  OR2_X1    g152(.A1(KEYINPUT64), .A2(G134), .ZN(new_n339));
  NAND2_X1  g153(.A1(KEYINPUT64), .A2(G134), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  XNOR2_X1  g155(.A(G128), .B(G143), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n240), .A2(G143), .ZN(new_n345));
  OR2_X1    g159(.A1(new_n345), .A2(KEYINPUT13), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(KEYINPUT13), .ZN(new_n347));
  OAI211_X1 g161(.A(new_n346), .B(new_n347), .C1(G128), .C2(new_n235), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n344), .B1(new_n348), .B2(G134), .ZN(new_n349));
  XNOR2_X1  g163(.A(G116), .B(G122), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n350), .A2(new_n194), .ZN(new_n351));
  AND2_X1   g165(.A1(new_n350), .A2(new_n194), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n349), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  OAI21_X1  g167(.A(KEYINPUT14), .B1(new_n206), .B2(G122), .ZN(new_n354));
  OR2_X1    g168(.A1(new_n194), .A2(KEYINPUT14), .ZN(new_n355));
  AOI22_X1  g169(.A1(new_n351), .A2(new_n354), .B1(new_n350), .B2(new_n355), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n341), .A2(new_n342), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n356), .B1(new_n344), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n353), .A2(new_n358), .ZN(new_n359));
  XOR2_X1   g173(.A(KEYINPUT9), .B(G234), .Z(new_n360));
  NAND3_X1  g174(.A1(new_n360), .A2(G217), .A3(new_n253), .ZN(new_n361));
  XNOR2_X1  g175(.A(new_n359), .B(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(new_n275), .ZN(new_n363));
  INV_X1    g177(.A(G478), .ZN(new_n364));
  OR2_X1    g178(.A1(new_n364), .A2(KEYINPUT15), .ZN(new_n365));
  XNOR2_X1  g179(.A(new_n363), .B(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n338), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(G234), .A2(G237), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n369), .A2(G952), .A3(new_n253), .ZN(new_n370));
  XOR2_X1   g184(.A(KEYINPUT21), .B(G898), .Z(new_n371));
  NAND3_X1  g185(.A1(new_n369), .A2(G902), .A3(G953), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n370), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  AND3_X1   g187(.A1(new_n284), .A2(new_n368), .A3(new_n373), .ZN(new_n374));
  OR2_X1    g188(.A1(new_n203), .A2(new_n204), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT23), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n375), .B1(new_n376), .B2(G128), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n240), .A2(KEYINPUT23), .A3(G119), .ZN(new_n378));
  OAI211_X1 g192(.A(new_n377), .B(new_n378), .C1(KEYINPUT23), .C2(new_n240), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(G110), .ZN(new_n380));
  MUX2_X1   g194(.A(G119), .B(new_n375), .S(G128), .Z(new_n381));
  XOR2_X1   g195(.A(KEYINPUT24), .B(G110), .Z(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  OAI221_X1 g197(.A(new_n380), .B1(new_n381), .B2(new_n383), .C1(new_n298), .C2(new_n299), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n381), .A2(new_n383), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n385), .B1(new_n379), .B2(G110), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n297), .A2(new_n314), .A3(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n253), .A2(G221), .A3(G234), .ZN(new_n388));
  XNOR2_X1  g202(.A(new_n388), .B(KEYINPUT80), .ZN(new_n389));
  XNOR2_X1  g203(.A(new_n389), .B(KEYINPUT22), .ZN(new_n390));
  XNOR2_X1  g204(.A(new_n390), .B(G137), .ZN(new_n391));
  AND3_X1   g205(.A1(new_n384), .A2(new_n387), .A3(new_n391), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n391), .B1(new_n384), .B2(new_n387), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  OAI21_X1  g208(.A(KEYINPUT25), .B1(new_n394), .B2(G902), .ZN(new_n395));
  INV_X1    g209(.A(G217), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n396), .B1(G234), .B2(new_n275), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(KEYINPUT75), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT25), .ZN(new_n399));
  OAI211_X1 g213(.A(new_n399), .B(new_n275), .C1(new_n392), .C2(new_n393), .ZN(new_n400));
  OR2_X1    g214(.A1(new_n397), .A2(KEYINPUT75), .ZN(new_n401));
  NAND4_X1  g215(.A1(new_n395), .A2(new_n398), .A3(new_n400), .A4(new_n401), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n397), .A2(G902), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n403), .B1(new_n392), .B2(new_n393), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT74), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT30), .ZN(new_n408));
  OR2_X1    g222(.A1(new_n408), .A2(KEYINPUT65), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(KEYINPUT65), .ZN(new_n410));
  INV_X1    g224(.A(G137), .ZN(new_n411));
  AOI22_X1  g225(.A1(new_n339), .A2(new_n340), .B1(KEYINPUT11), .B2(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n411), .A2(KEYINPUT11), .A3(G134), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT11), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(G137), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  OAI21_X1  g230(.A(G131), .B1(new_n412), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n411), .A2(KEYINPUT11), .ZN(new_n418));
  AND2_X1   g232(.A1(KEYINPUT64), .A2(G134), .ZN(new_n419));
  NOR2_X1   g233(.A1(KEYINPUT64), .A2(G134), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n418), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND4_X1  g235(.A1(new_n421), .A2(new_n304), .A3(new_n413), .A4(new_n415), .ZN(new_n422));
  AOI22_X1  g236(.A1(new_n417), .A2(new_n422), .B1(new_n242), .B2(new_n243), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n411), .B1(new_n419), .B2(new_n420), .ZN(new_n424));
  NAND2_X1  g238(.A1(G134), .A2(G137), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n424), .A2(G131), .A3(new_n425), .ZN(new_n426));
  AND3_X1   g240(.A1(new_n422), .A2(new_n250), .A3(new_n426), .ZN(new_n427));
  OAI211_X1 g241(.A(new_n409), .B(new_n410), .C1(new_n423), .C2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n422), .ZN(new_n429));
  AND2_X1   g243(.A1(new_n413), .A2(new_n415), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n304), .B1(new_n430), .B2(new_n421), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n244), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n422), .A2(new_n250), .A3(new_n426), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n432), .A2(KEYINPUT65), .A3(new_n408), .A4(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n428), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(new_n213), .ZN(new_n436));
  INV_X1    g250(.A(G210), .ZN(new_n437));
  NOR3_X1   g251(.A1(new_n437), .A2(G237), .A3(G953), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n438), .B(KEYINPUT27), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n439), .B(KEYINPUT26), .ZN(new_n440));
  INV_X1    g254(.A(G101), .ZN(new_n441));
  XNOR2_X1  g255(.A(new_n440), .B(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n212), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n211), .B1(new_n205), .B2(new_n207), .ZN(new_n444));
  OAI21_X1  g258(.A(KEYINPUT67), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT67), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n210), .A2(new_n446), .A3(new_n212), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n432), .A2(new_n445), .A3(new_n447), .A4(new_n433), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n436), .A2(new_n442), .A3(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT31), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND4_X1  g265(.A1(new_n436), .A2(KEYINPUT31), .A3(new_n442), .A4(new_n448), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n213), .B1(new_n423), .B2(new_n427), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT68), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  OAI211_X1 g270(.A(KEYINPUT68), .B(new_n213), .C1(new_n423), .C2(new_n427), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n456), .A2(new_n448), .A3(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT69), .ZN(new_n459));
  AND3_X1   g273(.A1(new_n458), .A2(new_n459), .A3(KEYINPUT28), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n459), .B1(new_n458), .B2(KEYINPUT28), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT28), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n448), .A2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  NOR3_X1   g278(.A1(new_n460), .A2(new_n461), .A3(new_n464), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n453), .B1(new_n465), .B2(new_n442), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(KEYINPUT70), .ZN(new_n467));
  NOR2_X1   g281(.A1(G472), .A2(G902), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n443), .A2(new_n444), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n469), .B1(new_n432), .B2(new_n433), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n448), .B1(new_n470), .B2(KEYINPUT68), .ZN(new_n471));
  INV_X1    g285(.A(new_n457), .ZN(new_n472));
  OAI21_X1  g286(.A(KEYINPUT28), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(KEYINPUT69), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n458), .A2(new_n459), .A3(KEYINPUT28), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n474), .A2(new_n463), .A3(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(new_n442), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT70), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n478), .A2(new_n479), .A3(new_n453), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n467), .A2(new_n468), .A3(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT32), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n481), .A2(KEYINPUT71), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT71), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n467), .A2(new_n485), .A3(new_n468), .A4(new_n480), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n483), .B1(new_n487), .B2(new_n482), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n474), .A2(new_n442), .A3(new_n463), .A4(new_n475), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n436), .A2(new_n448), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(new_n477), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT29), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n489), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(KEYINPUT72), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n463), .A2(KEYINPUT73), .ZN(new_n495));
  AND2_X1   g309(.A1(new_n463), .A2(KEYINPUT73), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n432), .A2(new_n433), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n445), .A2(new_n447), .ZN(new_n498));
  XNOR2_X1  g312(.A(new_n497), .B(new_n498), .ZN(new_n499));
  AOI211_X1 g313(.A(new_n495), .B(new_n496), .C1(KEYINPUT28), .C2(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n500), .A2(KEYINPUT29), .A3(new_n442), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT72), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n489), .A2(new_n491), .A3(new_n502), .A4(new_n492), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n494), .A2(new_n501), .A3(new_n275), .A4(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(G472), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n407), .B1(new_n488), .B2(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(KEYINPUT32), .B1(new_n484), .B2(new_n486), .ZN(new_n507));
  INV_X1    g321(.A(new_n505), .ZN(new_n508));
  NOR4_X1   g322(.A1(new_n507), .A2(KEYINPUT74), .A3(new_n508), .A4(new_n483), .ZN(new_n509));
  OAI211_X1 g323(.A(new_n374), .B(new_n406), .C1(new_n506), .C2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n360), .ZN(new_n511));
  OAI21_X1  g325(.A(G221), .B1(new_n511), .B2(G902), .ZN(new_n512));
  INV_X1    g326(.A(G469), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n201), .A2(new_n244), .A3(new_n202), .ZN(new_n514));
  INV_X1    g328(.A(new_n247), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n248), .A2(new_n249), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n516), .B(KEYINPUT84), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n269), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT10), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n269), .A2(KEYINPUT10), .A3(new_n250), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n417), .A2(new_n422), .ZN(new_n522));
  XOR2_X1   g336(.A(new_n522), .B(KEYINPUT85), .Z(new_n523));
  NAND4_X1  g337(.A1(new_n514), .A2(new_n520), .A3(new_n521), .A4(new_n523), .ZN(new_n524));
  AND3_X1   g338(.A1(new_n514), .A2(new_n520), .A3(new_n521), .ZN(new_n525));
  INV_X1    g339(.A(new_n522), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  XNOR2_X1  g341(.A(G110), .B(G140), .ZN(new_n528));
  INV_X1    g342(.A(G227), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n529), .A2(G953), .ZN(new_n530));
  XOR2_X1   g344(.A(new_n528), .B(new_n530), .Z(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n527), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n220), .A2(new_n251), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n526), .B1(new_n534), .B2(new_n518), .ZN(new_n535));
  XNOR2_X1  g349(.A(new_n535), .B(KEYINPUT12), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n531), .B1(new_n536), .B2(new_n524), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n533), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(KEYINPUT86), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT86), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n540), .B1(new_n533), .B2(new_n537), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n513), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT87), .ZN(new_n543));
  AND2_X1   g357(.A1(new_n534), .A2(new_n518), .ZN(new_n544));
  OAI21_X1  g358(.A(KEYINPUT12), .B1(new_n544), .B2(new_n526), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT12), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n535), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n545), .A2(new_n524), .A3(new_n547), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n543), .B1(new_n548), .B2(new_n532), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n536), .A2(KEYINPUT87), .A3(new_n524), .A4(new_n531), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n527), .A2(new_n532), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n552), .A2(new_n513), .A3(new_n275), .ZN(new_n553));
  NAND2_X1  g367(.A1(G469), .A2(G902), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n512), .B1(new_n542), .B2(new_n555), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n510), .A2(new_n556), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n557), .B(new_n441), .ZN(G3));
  INV_X1    g372(.A(new_n338), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n362), .B(KEYINPUT33), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n560), .A2(G478), .A3(new_n275), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n363), .A2(new_n364), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n559), .A2(new_n564), .ZN(new_n565));
  AND3_X1   g379(.A1(new_n284), .A2(new_n373), .A3(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n556), .ZN(new_n567));
  AOI221_X4 g381(.A(KEYINPUT70), .B1(new_n451), .B2(new_n452), .C1(new_n476), .C2(new_n477), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n479), .B1(new_n478), .B2(new_n453), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  OAI21_X1  g385(.A(G472), .B1(new_n571), .B2(G902), .ZN(new_n572));
  AND2_X1   g386(.A1(new_n572), .A2(new_n487), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n566), .A2(new_n567), .A3(new_n406), .A4(new_n573), .ZN(new_n574));
  XOR2_X1   g388(.A(KEYINPUT34), .B(G104), .Z(new_n575));
  XNOR2_X1  g389(.A(new_n574), .B(new_n575), .ZN(G6));
  NOR2_X1   g390(.A1(new_n338), .A2(new_n366), .ZN(new_n577));
  AND3_X1   g391(.A1(new_n284), .A2(new_n373), .A3(new_n577), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n578), .A2(new_n567), .A3(new_n406), .A4(new_n573), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n579), .B(KEYINPUT93), .ZN(new_n580));
  XOR2_X1   g394(.A(KEYINPUT35), .B(G107), .Z(new_n581));
  XNOR2_X1  g395(.A(new_n580), .B(new_n581), .ZN(G9));
  NAND2_X1  g396(.A1(new_n384), .A2(new_n387), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n583), .B(KEYINPUT94), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n391), .A2(KEYINPUT36), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT94), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n583), .B(new_n588), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n589), .A2(new_n585), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n403), .B1(new_n587), .B2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT95), .ZN(new_n592));
  AND3_X1   g406(.A1(new_n591), .A2(new_n592), .A3(new_n402), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n592), .B1(new_n591), .B2(new_n402), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND4_X1  g409(.A1(new_n374), .A2(new_n567), .A3(new_n573), .A4(new_n595), .ZN(new_n596));
  XNOR2_X1  g410(.A(KEYINPUT37), .B(G110), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n596), .B(new_n597), .ZN(new_n598));
  XNOR2_X1  g412(.A(KEYINPUT96), .B(KEYINPUT97), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n598), .B(new_n599), .ZN(G12));
  INV_X1    g414(.A(KEYINPUT100), .ZN(new_n601));
  OAI211_X1 g415(.A(new_n567), .B(new_n595), .C1(new_n506), .C2(new_n509), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n282), .A2(new_n283), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(new_n187), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n370), .B(KEYINPUT99), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(KEYINPUT98), .B(G900), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n606), .B1(new_n372), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n577), .A2(new_n608), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n604), .A2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n601), .B1(new_n602), .B2(new_n611), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n485), .B1(new_n570), .B2(new_n468), .ZN(new_n613));
  INV_X1    g427(.A(new_n486), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n482), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n570), .A2(KEYINPUT32), .A3(new_n468), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n615), .A2(new_n616), .A3(new_n505), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(KEYINPUT74), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n488), .A2(new_n407), .A3(new_n505), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n556), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n620), .A2(KEYINPUT100), .A3(new_n595), .A4(new_n610), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n612), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(G128), .ZN(G30));
  XNOR2_X1  g437(.A(new_n603), .B(KEYINPUT101), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(KEYINPUT38), .ZN(new_n625));
  XOR2_X1   g439(.A(new_n608), .B(KEYINPUT39), .Z(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n567), .A2(new_n627), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n628), .A2(KEYINPUT40), .ZN(new_n629));
  NOR4_X1   g443(.A1(new_n625), .A2(new_n188), .A3(new_n595), .A4(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n338), .A2(new_n367), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n631), .B1(new_n628), .B2(KEYINPUT40), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n490), .A2(new_n442), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n275), .B1(new_n499), .B2(new_n442), .ZN(new_n635));
  OAI21_X1  g449(.A(G472), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n488), .A2(new_n636), .ZN(new_n637));
  AND3_X1   g451(.A1(new_n630), .A2(new_n632), .A3(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(KEYINPUT102), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(new_n235), .ZN(G45));
  AND3_X1   g454(.A1(new_n338), .A2(new_n563), .A3(new_n608), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  OAI21_X1  g456(.A(KEYINPUT103), .B1(new_n604), .B2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT103), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n284), .A2(new_n644), .A3(new_n641), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n602), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(new_n233), .ZN(G48));
  INV_X1    g462(.A(KEYINPUT104), .ZN(new_n649));
  INV_X1    g463(.A(new_n553), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n513), .B1(new_n552), .B2(new_n275), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(new_n512), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  OAI211_X1 g468(.A(new_n654), .B(new_n406), .C1(new_n506), .C2(new_n509), .ZN(new_n655));
  INV_X1    g469(.A(new_n566), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n649), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n405), .B1(new_n618), .B2(new_n619), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n658), .A2(KEYINPUT104), .A3(new_n566), .A4(new_n654), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(KEYINPUT41), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(G113), .ZN(G15));
  INV_X1    g476(.A(new_n655), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n578), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(G116), .ZN(G18));
  NAND4_X1  g479(.A1(new_n595), .A2(new_n284), .A3(new_n368), .A4(new_n373), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n666), .B1(new_n619), .B2(new_n618), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(new_n654), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(G119), .ZN(G21));
  INV_X1    g483(.A(KEYINPUT108), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n631), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n338), .A2(KEYINPUT108), .A3(new_n367), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n673), .A2(new_n284), .A3(new_n373), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n453), .B1(new_n500), .B2(new_n442), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(new_n468), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(KEYINPUT105), .ZN(new_n677));
  AND2_X1   g491(.A1(new_n572), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n405), .A2(KEYINPUT106), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT106), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n680), .B1(new_n402), .B2(new_n404), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n678), .A2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT107), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n678), .A2(new_n682), .A3(KEYINPUT107), .ZN(new_n686));
  AOI211_X1 g500(.A(new_n653), .B(new_n674), .C1(new_n685), .C2(new_n686), .ZN(new_n687));
  XOR2_X1   g501(.A(new_n687), .B(G122), .Z(G24));
  AND2_X1   g502(.A1(new_n595), .A2(new_n678), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n604), .A2(new_n642), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n689), .A2(new_n690), .A3(new_n654), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G125), .ZN(G27));
  NAND2_X1  g506(.A1(new_n538), .A2(G469), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n553), .A2(new_n554), .A3(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(new_n512), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n695), .A2(new_n188), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n694), .A2(new_n282), .A3(new_n283), .A4(new_n696), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n697), .A2(new_n642), .ZN(new_n698));
  OAI211_X1 g512(.A(new_n698), .B(new_n406), .C1(new_n506), .C2(new_n509), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT109), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n658), .A2(KEYINPUT109), .A3(new_n698), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT42), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n701), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  OR2_X1    g518(.A1(new_n616), .A2(KEYINPUT110), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n616), .A2(KEYINPUT110), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n481), .A2(new_n482), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n705), .A2(new_n706), .A3(new_n505), .A4(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(new_n682), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(KEYINPUT111), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n710), .A2(KEYINPUT42), .A3(new_n698), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n704), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G131), .ZN(G33));
  NAND2_X1  g527(.A1(new_n618), .A2(new_n619), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(new_n406), .ZN(new_n715));
  OR3_X1    g529(.A1(new_n715), .A2(new_n609), .A3(new_n697), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G134), .ZN(G36));
  INV_X1    g531(.A(KEYINPUT45), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n539), .A2(new_n541), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n538), .A2(KEYINPUT45), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n719), .A2(G469), .A3(new_n720), .ZN(new_n721));
  AOI21_X1  g535(.A(KEYINPUT46), .B1(new_n721), .B2(new_n554), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n722), .A2(new_n650), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n721), .A2(KEYINPUT46), .A3(new_n554), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(new_n512), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n726), .A2(new_n626), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n603), .A2(new_n188), .ZN(new_n728));
  NOR3_X1   g542(.A1(new_n573), .A2(new_n594), .A3(new_n593), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n559), .A2(new_n563), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT43), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(new_n732), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n730), .A2(new_n731), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n729), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT44), .ZN(new_n736));
  OR2_X1    g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n735), .A2(new_n736), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n727), .A2(new_n728), .A3(new_n737), .A4(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G137), .ZN(G39));
  NAND2_X1  g554(.A1(new_n726), .A2(KEYINPUT47), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT47), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n725), .A2(new_n742), .A3(new_n512), .ZN(new_n743));
  AND2_X1   g557(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n641), .A2(new_n405), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n714), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n744), .A2(new_n728), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(KEYINPUT112), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT112), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n744), .A2(new_n749), .A3(new_n728), .A4(new_n746), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G140), .ZN(G42));
  INV_X1    g566(.A(KEYINPUT53), .ZN(new_n753));
  AOI22_X1  g567(.A1(new_n663), .A2(new_n578), .B1(new_n667), .B2(new_n654), .ZN(new_n754));
  INV_X1    g568(.A(new_n687), .ZN(new_n755));
  AND4_X1   g569(.A1(new_n596), .A2(new_n660), .A3(new_n754), .A4(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(new_n602), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n757), .A2(new_n368), .A3(new_n608), .A4(new_n728), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n698), .A2(new_n689), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(KEYINPUT113), .ZN(new_n760));
  AND3_X1   g574(.A1(new_n716), .A2(new_n758), .A3(new_n760), .ZN(new_n761));
  OAI211_X1 g575(.A(new_n574), .B(new_n579), .C1(new_n510), .C2(new_n556), .ZN(new_n762));
  INV_X1    g576(.A(new_n762), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n756), .A2(new_n712), .A3(new_n761), .A4(new_n763), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n691), .B1(new_n602), .B2(new_n646), .ZN(new_n765));
  INV_X1    g579(.A(new_n765), .ZN(new_n766));
  AND4_X1   g580(.A1(new_n402), .A2(new_n637), .A3(new_n591), .A4(new_n608), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n673), .A2(new_n284), .ZN(new_n768));
  INV_X1    g582(.A(new_n768), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n767), .A2(new_n512), .A3(new_n694), .A4(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n622), .A2(new_n766), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(KEYINPUT52), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n765), .B1(new_n612), .B2(new_n621), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT52), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n773), .A2(new_n774), .A3(new_n770), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n772), .A2(new_n775), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n753), .B1(new_n764), .B2(new_n776), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n774), .B1(new_n773), .B2(new_n770), .ZN(new_n778));
  AND4_X1   g592(.A1(new_n774), .A2(new_n622), .A3(new_n766), .A4(new_n770), .ZN(new_n779));
  OAI21_X1  g593(.A(KEYINPUT114), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT114), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n772), .A2(new_n775), .A3(new_n781), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n764), .B1(new_n780), .B2(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(new_n783), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n777), .B1(new_n784), .B2(new_n753), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(KEYINPUT54), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n685), .A2(new_n686), .ZN(new_n787));
  INV_X1    g601(.A(new_n734), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n606), .B1(new_n788), .B2(new_n732), .ZN(new_n789));
  AND2_X1   g603(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  NOR3_X1   g604(.A1(new_n650), .A2(new_n512), .A3(new_n651), .ZN(new_n791));
  OAI211_X1 g605(.A(new_n728), .B(new_n790), .C1(new_n744), .C2(new_n791), .ZN(new_n792));
  NOR3_X1   g606(.A1(new_n653), .A2(new_n188), .A3(new_n603), .ZN(new_n793));
  AND2_X1   g607(.A1(new_n789), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(new_n689), .ZN(new_n795));
  XOR2_X1   g609(.A(new_n795), .B(KEYINPUT117), .Z(new_n796));
  INV_X1    g610(.A(new_n637), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n793), .A2(new_n797), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n405), .A2(new_n370), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n798), .A2(new_n559), .A3(new_n564), .A4(new_n799), .ZN(new_n800));
  NOR2_X1   g614(.A1(KEYINPUT116), .A2(KEYINPUT50), .ZN(new_n801));
  NOR3_X1   g615(.A1(new_n653), .A2(new_n187), .A3(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n790), .A2(new_n625), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(KEYINPUT116), .A2(KEYINPUT50), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n803), .B(new_n804), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n792), .A2(new_n796), .A3(new_n800), .A4(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT51), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n710), .A2(new_n794), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(KEYINPUT48), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n787), .A2(new_n284), .A3(new_n654), .A4(new_n789), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n808), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  AND3_X1   g626(.A1(new_n798), .A2(new_n565), .A3(new_n799), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n806), .A2(new_n807), .ZN(new_n814));
  NOR3_X1   g628(.A1(new_n812), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n687), .B1(new_n657), .B2(new_n659), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n816), .A2(new_n763), .A3(new_n596), .A4(new_n754), .ZN(new_n817));
  AND2_X1   g631(.A1(new_n704), .A2(new_n711), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n716), .A2(new_n758), .A3(new_n760), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n817), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n778), .A2(new_n779), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n753), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n822), .B1(new_n783), .B2(new_n753), .ZN(new_n823));
  OAI21_X1  g637(.A(KEYINPUT115), .B1(new_n823), .B2(KEYINPUT54), .ZN(new_n824));
  AND3_X1   g638(.A1(new_n772), .A2(new_n781), .A3(new_n775), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n781), .B1(new_n772), .B2(new_n775), .ZN(new_n826));
  OAI211_X1 g640(.A(new_n753), .B(new_n820), .C1(new_n825), .C2(new_n826), .ZN(new_n827));
  OAI21_X1  g641(.A(KEYINPUT53), .B1(new_n764), .B2(new_n776), .ZN(new_n828));
  AOI21_X1  g642(.A(KEYINPUT54), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT115), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n786), .A2(new_n815), .A3(new_n824), .A4(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT118), .ZN(new_n833));
  OAI211_X1 g647(.A(G952), .B(new_n253), .C1(new_n832), .C2(new_n833), .ZN(new_n834));
  OAI21_X1  g648(.A(G953), .B1(new_n832), .B2(KEYINPUT118), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT49), .ZN(new_n836));
  AOI211_X1 g650(.A(new_n681), .B(new_n679), .C1(new_n652), .C2(new_n836), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n652), .A2(new_n836), .ZN(new_n838));
  NOR4_X1   g652(.A1(new_n838), .A2(new_n695), .A3(new_n188), .A4(new_n730), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n625), .A2(new_n797), .A3(new_n837), .A4(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n834), .A2(new_n835), .A3(new_n840), .ZN(G75));
  OAI21_X1  g655(.A(new_n232), .B1(new_n258), .B2(new_n260), .ZN(new_n842));
  XOR2_X1   g656(.A(new_n842), .B(KEYINPUT119), .Z(new_n843));
  XOR2_X1   g657(.A(new_n843), .B(KEYINPUT55), .Z(new_n844));
  XNOR2_X1  g658(.A(new_n844), .B(new_n255), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n827), .A2(G902), .A3(new_n828), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(KEYINPUT120), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT120), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n827), .A2(new_n848), .A3(G902), .A4(new_n828), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  AOI211_X1 g664(.A(KEYINPUT56), .B(new_n845), .C1(new_n850), .C2(new_n281), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n846), .A2(new_n437), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n845), .B1(new_n852), .B2(KEYINPUT56), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n253), .A2(G952), .ZN(new_n854));
  INV_X1    g668(.A(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n851), .A2(new_n856), .ZN(G51));
  XOR2_X1   g671(.A(new_n554), .B(KEYINPUT57), .Z(new_n858));
  AND3_X1   g672(.A1(new_n827), .A2(KEYINPUT54), .A3(new_n828), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n858), .B1(new_n859), .B2(new_n829), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n860), .A2(new_n552), .ZN(new_n861));
  INV_X1    g675(.A(new_n721), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n850), .A2(new_n862), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n854), .B1(new_n861), .B2(new_n863), .ZN(G54));
  AOI21_X1  g678(.A(new_n848), .B1(new_n823), .B2(G902), .ZN(new_n865));
  INV_X1    g679(.A(new_n849), .ZN(new_n866));
  OAI211_X1 g680(.A(KEYINPUT58), .B(G475), .C1(new_n865), .C2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT121), .ZN(new_n868));
  INV_X1    g682(.A(new_n328), .ZN(new_n869));
  AND3_X1   g683(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n868), .B1(new_n867), .B2(new_n869), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n850), .A2(KEYINPUT58), .A3(G475), .A4(new_n328), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n872), .A2(new_n855), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n870), .A2(new_n871), .A3(new_n873), .ZN(G60));
  XNOR2_X1  g688(.A(new_n560), .B(KEYINPUT122), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n786), .A2(new_n824), .A3(new_n831), .ZN(new_n876));
  NAND2_X1  g690(.A1(G478), .A2(G902), .ZN(new_n877));
  XNOR2_X1  g691(.A(new_n877), .B(KEYINPUT59), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n875), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  OAI211_X1 g693(.A(new_n878), .B(new_n875), .C1(new_n859), .C2(new_n829), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT123), .ZN(new_n881));
  AND3_X1   g695(.A1(new_n880), .A2(new_n881), .A3(new_n855), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n881), .B1(new_n880), .B2(new_n855), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n879), .A2(new_n882), .A3(new_n883), .ZN(G63));
  NAND2_X1  g698(.A1(G217), .A2(G902), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n885), .B(KEYINPUT60), .ZN(new_n886));
  INV_X1    g700(.A(new_n886), .ZN(new_n887));
  OAI211_X1 g701(.A(new_n823), .B(new_n887), .C1(new_n587), .C2(new_n590), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n827), .A2(new_n828), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n394), .B1(new_n889), .B2(new_n886), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n888), .A2(new_n890), .A3(KEYINPUT61), .A4(new_n855), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT125), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n891), .B(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT61), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n823), .A2(new_n887), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n854), .B1(new_n895), .B2(new_n394), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT124), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n888), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  AND3_X1   g712(.A1(new_n890), .A2(new_n897), .A3(new_n855), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n894), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n893), .A2(new_n900), .ZN(G66));
  AOI21_X1  g715(.A(new_n253), .B1(new_n371), .B2(G224), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n817), .B(KEYINPUT126), .ZN(new_n903));
  INV_X1    g717(.A(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n902), .B1(new_n904), .B2(new_n253), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n843), .B1(G898), .B2(new_n253), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(KEYINPUT127), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n905), .B(new_n907), .ZN(G69));
  XOR2_X1   g722(.A(new_n435), .B(new_n325), .Z(new_n909));
  NAND2_X1  g723(.A1(new_n529), .A2(G953), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n751), .A2(new_n712), .A3(new_n716), .ZN(new_n911));
  INV_X1    g725(.A(new_n739), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n727), .A2(new_n710), .A3(new_n769), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(new_n773), .ZN(new_n914));
  NOR3_X1   g728(.A1(new_n911), .A2(new_n912), .A3(new_n914), .ZN(new_n915));
  OAI211_X1 g729(.A(new_n909), .B(new_n910), .C1(new_n915), .C2(G953), .ZN(new_n916));
  OAI21_X1  g730(.A(G900), .B1(new_n909), .B2(G227), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(G953), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n565), .A2(new_n577), .ZN(new_n919));
  NOR4_X1   g733(.A1(new_n628), .A2(new_n188), .A3(new_n603), .A4(new_n919), .ZN(new_n920));
  AOI22_X1  g734(.A1(new_n748), .A2(new_n750), .B1(new_n658), .B2(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(new_n638), .ZN(new_n922));
  AND3_X1   g736(.A1(new_n922), .A2(KEYINPUT62), .A3(new_n773), .ZN(new_n923));
  AOI21_X1  g737(.A(KEYINPUT62), .B1(new_n922), .B2(new_n773), .ZN(new_n924));
  OAI211_X1 g738(.A(new_n739), .B(new_n921), .C1(new_n923), .C2(new_n924), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n909), .A2(G953), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n916), .A2(new_n918), .A3(new_n927), .ZN(G72));
  NAND2_X1  g742(.A1(G472), .A2(G902), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n929), .B(KEYINPUT63), .Z(new_n930));
  INV_X1    g744(.A(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n931), .B1(new_n915), .B2(new_n903), .ZN(new_n932));
  NOR3_X1   g746(.A1(new_n932), .A2(new_n442), .A3(new_n490), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n930), .B1(new_n925), .B2(new_n904), .ZN(new_n934));
  AND2_X1   g748(.A1(new_n934), .A2(new_n634), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n477), .A2(new_n448), .A3(new_n436), .ZN(new_n936));
  AND4_X1   g750(.A1(new_n633), .A2(new_n785), .A3(new_n930), .A4(new_n936), .ZN(new_n937));
  NOR4_X1   g751(.A1(new_n933), .A2(new_n935), .A3(new_n937), .A4(new_n854), .ZN(G57));
endmodule


