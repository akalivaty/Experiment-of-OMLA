//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 0 0 1 1 1 0 0 1 1 0 0 1 0 1 1 0 1 1 1 0 0 1 1 1 0 1 1 0 0 0 0 0 1 0 0 0 0 0 0 1 1 1 1 0 0 0 0 1 1 0 1 0 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:10 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n444, new_n448, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n560, new_n561, new_n563, new_n564, new_n565,
    new_n566, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n586, new_n587, new_n588, new_n589, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n625,
    new_n627, new_n628, new_n629, new_n630, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT64), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  XOR2_X1   g013(.A(KEYINPUT65), .B(G69), .Z(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  XNOR2_X1  g015(.A(KEYINPUT66), .B(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XOR2_X1   g019(.A(new_n444), .B(KEYINPUT67), .Z(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(new_n453), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n457), .A2(G2106), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OR2_X1    g034(.A1(new_n454), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  AND2_X1   g037(.A1(KEYINPUT68), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT68), .A2(G2104), .ZN(new_n464));
  OAI21_X1  g039(.A(KEYINPUT3), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT69), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  OR2_X1    g042(.A1(new_n467), .A2(KEYINPUT3), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT69), .ZN(new_n469));
  OAI211_X1 g044(.A(new_n469), .B(KEYINPUT3), .C1(new_n463), .C2(new_n464), .ZN(new_n470));
  AND3_X1   g045(.A1(new_n466), .A2(new_n468), .A3(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT70), .ZN(new_n472));
  INV_X1    g047(.A(G2105), .ZN(new_n473));
  NAND4_X1  g048(.A1(new_n471), .A2(new_n472), .A3(G137), .A4(new_n473), .ZN(new_n474));
  XNOR2_X1  g049(.A(KEYINPUT3), .B(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G125), .ZN(new_n476));
  INV_X1    g051(.A(G113), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n476), .B1(new_n477), .B2(new_n467), .ZN(new_n478));
  NOR3_X1   g053(.A1(new_n463), .A2(new_n464), .A3(G2105), .ZN(new_n479));
  AOI22_X1  g054(.A1(new_n478), .A2(G2105), .B1(new_n479), .B2(G101), .ZN(new_n480));
  NAND4_X1  g055(.A1(new_n466), .A2(new_n473), .A3(new_n468), .A4(new_n470), .ZN(new_n481));
  INV_X1    g056(.A(G137), .ZN(new_n482));
  OAI21_X1  g057(.A(KEYINPUT70), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n474), .A2(new_n480), .A3(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G160));
  NAND4_X1  g060(.A1(new_n466), .A2(G2105), .A3(new_n468), .A4(new_n470), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n481), .ZN(new_n488));
  AOI22_X1  g063(.A1(G124), .A2(new_n487), .B1(new_n488), .B2(G136), .ZN(new_n489));
  OR2_X1    g064(.A1(G100), .A2(G2105), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n490), .B(G2104), .C1(G112), .C2(new_n473), .ZN(new_n491));
  XNOR2_X1  g066(.A(new_n491), .B(KEYINPUT71), .ZN(new_n492));
  AND2_X1   g067(.A1(new_n489), .A2(new_n492), .ZN(G162));
  INV_X1    g068(.A(KEYINPUT72), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n494), .B1(new_n473), .B2(G114), .ZN(new_n495));
  INV_X1    g070(.A(G114), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n496), .A2(KEYINPUT72), .A3(G2105), .ZN(new_n497));
  OR2_X1    g072(.A1(G102), .A2(G2105), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n495), .A2(new_n497), .A3(new_n498), .A4(G2104), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(KEYINPUT73), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n496), .A2(G2105), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n467), .B1(new_n501), .B2(new_n494), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT73), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n502), .A2(new_n503), .A3(new_n498), .A4(new_n497), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n500), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(G126), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n505), .B1(new_n486), .B2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT4), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n473), .A2(G138), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n508), .B1(new_n509), .B2(KEYINPUT74), .ZN(new_n510));
  OR2_X1    g085(.A1(new_n508), .A2(KEYINPUT74), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n510), .A2(new_n475), .A3(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(new_n509), .ZN(new_n514));
  NAND4_X1  g089(.A1(new_n466), .A2(new_n468), .A3(new_n470), .A4(new_n514), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n513), .B1(new_n515), .B2(KEYINPUT4), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n507), .A2(new_n516), .ZN(G164));
  AND2_X1   g092(.A1(KEYINPUT6), .A2(G651), .ZN(new_n518));
  NOR2_X1   g093(.A1(KEYINPUT6), .A2(G651), .ZN(new_n519));
  OAI21_X1  g094(.A(G543), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G50), .ZN(new_n522));
  XOR2_X1   g097(.A(new_n522), .B(KEYINPUT75), .Z(new_n523));
  INV_X1    g098(.A(G543), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(KEYINPUT5), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT5), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G543), .ZN(new_n527));
  OAI211_X1 g102(.A(new_n525), .B(new_n527), .C1(new_n518), .C2(new_n519), .ZN(new_n528));
  INV_X1    g103(.A(new_n528), .ZN(new_n529));
  XNOR2_X1  g104(.A(KEYINPUT76), .B(G88), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n525), .A2(new_n527), .ZN(new_n532));
  INV_X1    g107(.A(new_n532), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n533), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n534));
  INV_X1    g109(.A(G651), .ZN(new_n535));
  OR2_X1    g110(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n523), .A2(new_n531), .A3(new_n536), .ZN(G303));
  INV_X1    g112(.A(G303), .ZN(G166));
  NAND2_X1  g113(.A1(G63), .A2(G651), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n518), .A2(new_n519), .ZN(new_n540));
  INV_X1    g115(.A(G89), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n542), .A2(new_n533), .B1(new_n521), .B2(G51), .ZN(new_n543));
  NAND3_X1  g118(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT7), .ZN(new_n545));
  AND2_X1   g120(.A1(new_n543), .A2(new_n545), .ZN(G168));
  AOI22_X1  g121(.A1(new_n533), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n547), .A2(new_n535), .ZN(new_n548));
  INV_X1    g123(.A(G90), .ZN(new_n549));
  INV_X1    g124(.A(G52), .ZN(new_n550));
  OAI22_X1  g125(.A1(new_n528), .A2(new_n549), .B1(new_n520), .B2(new_n550), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n548), .A2(new_n551), .ZN(G171));
  AOI22_X1  g127(.A1(new_n533), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n553), .A2(new_n535), .ZN(new_n554));
  INV_X1    g129(.A(G81), .ZN(new_n555));
  INV_X1    g130(.A(G43), .ZN(new_n556));
  OAI22_X1  g131(.A1(new_n528), .A2(new_n555), .B1(new_n520), .B2(new_n556), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G860), .ZN(G153));
  AND3_X1   g134(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G36), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT77), .ZN(G176));
  NAND2_X1  g137(.A1(G1), .A2(G3), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT79), .ZN(new_n564));
  XNOR2_X1  g139(.A(KEYINPUT78), .B(KEYINPUT8), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n564), .B(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n560), .A2(new_n566), .ZN(G188));
  NAND2_X1  g142(.A1(G78), .A2(G543), .ZN(new_n568));
  INV_X1    g143(.A(G65), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n568), .B1(new_n532), .B2(new_n569), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT80), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(G651), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n521), .A2(G53), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n573), .B(KEYINPUT9), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n529), .A2(G91), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n572), .A2(new_n574), .A3(new_n575), .ZN(G299));
  INV_X1    g151(.A(G171), .ZN(G301));
  INV_X1    g152(.A(G168), .ZN(G286));
  OAI21_X1  g153(.A(G651), .B1(new_n533), .B2(G74), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n579), .A2(KEYINPUT81), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n529), .A2(G87), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n521), .A2(G49), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT81), .ZN(new_n583));
  OAI211_X1 g158(.A(new_n583), .B(G651), .C1(new_n533), .C2(G74), .ZN(new_n584));
  NAND4_X1  g159(.A1(new_n580), .A2(new_n581), .A3(new_n582), .A4(new_n584), .ZN(G288));
  AOI22_X1  g160(.A1(new_n533), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n586), .A2(new_n535), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n533), .A2(G86), .B1(G48), .B2(G543), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n588), .A2(new_n540), .ZN(new_n589));
  OR2_X1    g164(.A1(new_n587), .A2(new_n589), .ZN(G305));
  INV_X1    g165(.A(G85), .ZN(new_n591));
  INV_X1    g166(.A(G47), .ZN(new_n592));
  OAI22_X1  g167(.A1(new_n528), .A2(new_n591), .B1(new_n520), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(G72), .A2(G543), .ZN(new_n594));
  INV_X1    g169(.A(G60), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n532), .B2(new_n595), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n593), .B1(G651), .B2(new_n596), .ZN(new_n597));
  XNOR2_X1  g172(.A(new_n597), .B(KEYINPUT82), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(G290));
  NAND2_X1  g174(.A1(G301), .A2(G868), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n529), .A2(G92), .ZN(new_n601));
  XOR2_X1   g176(.A(new_n601), .B(KEYINPUT10), .Z(new_n602));
  NAND2_X1  g177(.A1(new_n521), .A2(G54), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n525), .A2(new_n527), .A3(G66), .ZN(new_n604));
  NAND2_X1  g179(.A1(G79), .A2(G543), .ZN(new_n605));
  AND2_X1   g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n603), .B1(new_n606), .B2(new_n535), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT83), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  OAI211_X1 g184(.A(new_n603), .B(KEYINPUT83), .C1(new_n606), .C2(new_n535), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  AND3_X1   g186(.A1(new_n602), .A2(new_n611), .A3(KEYINPUT84), .ZN(new_n612));
  AOI21_X1  g187(.A(KEYINPUT84), .B1(new_n602), .B2(new_n611), .ZN(new_n613));
  NOR2_X1   g188(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n600), .B1(new_n614), .B2(G868), .ZN(G284));
  OAI21_X1  g190(.A(new_n600), .B1(new_n614), .B2(G868), .ZN(G321));
  INV_X1    g191(.A(G868), .ZN(new_n617));
  NOR2_X1   g192(.A1(G168), .A2(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(new_n618), .ZN(new_n619));
  INV_X1    g194(.A(G299), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n620), .B2(G868), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n621), .A2(KEYINPUT85), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(KEYINPUT85), .B2(new_n618), .ZN(G297));
  OAI21_X1  g198(.A(new_n622), .B1(KEYINPUT85), .B2(new_n618), .ZN(G280));
  INV_X1    g199(.A(G559), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n614), .B1(new_n625), .B2(G860), .ZN(G148));
  INV_X1    g201(.A(new_n558), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(new_n617), .ZN(new_n628));
  OR2_X1    g203(.A1(new_n612), .A2(new_n613), .ZN(new_n629));
  NOR2_X1   g204(.A1(new_n629), .A2(G559), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n628), .B1(new_n630), .B2(new_n617), .ZN(G323));
  XNOR2_X1  g206(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g207(.A1(new_n479), .A2(new_n475), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT12), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT13), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2100), .ZN(new_n636));
  INV_X1    g211(.A(G135), .ZN(new_n637));
  NOR2_X1   g212(.A1(G99), .A2(G2105), .ZN(new_n638));
  OAI21_X1  g213(.A(G2104), .B1(new_n473), .B2(G111), .ZN(new_n639));
  OAI22_X1  g214(.A1(new_n481), .A2(new_n637), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  AOI21_X1  g215(.A(new_n640), .B1(new_n487), .B2(G123), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT86), .B(G2096), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n636), .A2(new_n643), .ZN(G156));
  XNOR2_X1  g219(.A(G1341), .B(G1348), .ZN(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2427), .B(G2438), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2430), .ZN(new_n648));
  XOR2_X1   g223(.A(KEYINPUT15), .B(G2435), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n650), .A2(KEYINPUT14), .ZN(new_n651));
  XNOR2_X1  g226(.A(KEYINPUT87), .B(KEYINPUT16), .ZN(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n651), .B(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(G2451), .B(G2454), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(G2443), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(G2446), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n654), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n651), .B(new_n652), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n660), .A2(new_n657), .ZN(new_n661));
  OAI21_X1  g236(.A(new_n646), .B1(new_n659), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n660), .A2(new_n657), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n654), .A2(new_n658), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n663), .A2(new_n664), .A3(new_n645), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n662), .A2(G14), .A3(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(KEYINPUT88), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n666), .A2(new_n667), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(G401));
  XNOR2_X1  g246(.A(G2072), .B(G2078), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n672), .B(KEYINPUT17), .Z(new_n673));
  XOR2_X1   g248(.A(G2067), .B(G2678), .Z(new_n674));
  XOR2_X1   g249(.A(G2084), .B(G2090), .Z(new_n675));
  NAND3_X1  g250(.A1(new_n673), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n676), .B(KEYINPUT89), .Z(new_n677));
  NOR2_X1   g252(.A1(new_n673), .A2(new_n674), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n678), .A2(new_n675), .ZN(new_n679));
  INV_X1    g254(.A(new_n674), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n679), .B1(new_n680), .B2(new_n672), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n680), .A2(new_n672), .A3(new_n675), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n682), .B(KEYINPUT18), .Z(new_n683));
  NAND3_X1  g258(.A1(new_n677), .A2(new_n681), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(G2100), .ZN(new_n685));
  XNOR2_X1  g260(.A(KEYINPUT90), .B(G2096), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(G227));
  XNOR2_X1  g263(.A(G1961), .B(G1966), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT91), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1956), .B(G2474), .ZN(new_n691));
  OR2_X1    g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n690), .A2(new_n691), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT93), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1971), .B(G1976), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT19), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n692), .A2(new_n697), .ZN(new_n699));
  XOR2_X1   g274(.A(new_n699), .B(KEYINPUT20), .Z(new_n700));
  NOR2_X1   g275(.A1(new_n693), .A2(new_n697), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n701), .B(KEYINPUT92), .Z(new_n702));
  NAND3_X1  g277(.A1(new_n698), .A2(new_n700), .A3(new_n702), .ZN(new_n703));
  AND2_X1   g278(.A1(new_n703), .A2(KEYINPUT95), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n703), .A2(KEYINPUT95), .ZN(new_n705));
  OR3_X1    g280(.A1(new_n704), .A2(new_n705), .A3(KEYINPUT94), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n703), .B(KEYINPUT95), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n707), .A2(KEYINPUT94), .ZN(new_n708));
  XOR2_X1   g283(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n709));
  XNOR2_X1  g284(.A(G1981), .B(G1986), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  XNOR2_X1  g286(.A(G1991), .B(G1996), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  AND3_X1   g288(.A1(new_n706), .A2(new_n708), .A3(new_n713), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n713), .B1(new_n706), .B2(new_n708), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(G229));
  INV_X1    g292(.A(G16), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(G23), .ZN(new_n719));
  INV_X1    g294(.A(G288), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n719), .B1(new_n720), .B2(new_n718), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT33), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(G1976), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n718), .A2(G6), .ZN(new_n724));
  INV_X1    g299(.A(G305), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n724), .B1(new_n725), .B2(new_n718), .ZN(new_n726));
  XOR2_X1   g301(.A(KEYINPUT32), .B(G1981), .Z(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n718), .A2(G22), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(G166), .B2(new_n718), .ZN(new_n730));
  XNOR2_X1  g305(.A(KEYINPUT99), .B(G1971), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n723), .A2(new_n728), .A3(new_n732), .ZN(new_n733));
  OR2_X1    g308(.A1(new_n733), .A2(KEYINPUT34), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n718), .A2(G24), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(new_n598), .B2(new_n718), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT98), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(G1986), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n733), .A2(KEYINPUT34), .ZN(new_n739));
  NOR2_X1   g314(.A1(G25), .A2(G29), .ZN(new_n740));
  INV_X1    g315(.A(G119), .ZN(new_n741));
  INV_X1    g316(.A(G131), .ZN(new_n742));
  OAI22_X1  g317(.A1(new_n741), .A2(new_n486), .B1(new_n481), .B2(new_n742), .ZN(new_n743));
  OR2_X1    g318(.A1(G95), .A2(G2105), .ZN(new_n744));
  OAI211_X1 g319(.A(new_n744), .B(G2104), .C1(G107), .C2(new_n473), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT96), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n743), .A2(new_n746), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n740), .B1(new_n747), .B2(G29), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT97), .ZN(new_n749));
  XNOR2_X1  g324(.A(KEYINPUT35), .B(G1991), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NAND4_X1  g326(.A1(new_n734), .A2(new_n738), .A3(new_n739), .A4(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(KEYINPUT100), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  AND2_X1   g329(.A1(new_n739), .A2(new_n751), .ZN(new_n755));
  NAND4_X1  g330(.A1(new_n755), .A2(KEYINPUT100), .A3(new_n738), .A4(new_n734), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n754), .A2(new_n756), .A3(KEYINPUT36), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n614), .A2(new_n718), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(G4), .B2(new_n718), .ZN(new_n759));
  INV_X1    g334(.A(G1348), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(KEYINPUT36), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n752), .A2(new_n753), .A3(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n641), .A2(G29), .ZN(new_n764));
  INV_X1    g339(.A(KEYINPUT108), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G5), .B2(G16), .ZN(new_n766));
  OR3_X1    g341(.A1(new_n765), .A2(G5), .A3(G16), .ZN(new_n767));
  OAI211_X1 g342(.A(new_n766), .B(new_n767), .C1(G301), .C2(new_n718), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT109), .ZN(new_n769));
  INV_X1    g344(.A(G1961), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n764), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n769), .A2(new_n770), .ZN(new_n772));
  XNOR2_X1  g347(.A(KEYINPUT31), .B(G11), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n718), .A2(G19), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(new_n558), .B2(new_n718), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n775), .A2(G1341), .ZN(new_n776));
  INV_X1    g351(.A(G1966), .ZN(new_n777));
  NAND2_X1  g352(.A1(G168), .A2(G16), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G16), .B2(G21), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n776), .B1(new_n777), .B2(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(G29), .ZN(new_n781));
  XNOR2_X1  g356(.A(KEYINPUT30), .B(G28), .ZN(new_n782));
  AOI22_X1  g357(.A1(new_n775), .A2(G1341), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NAND4_X1  g358(.A1(new_n772), .A2(new_n773), .A3(new_n780), .A4(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n488), .A2(G139), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT102), .ZN(new_n786));
  AOI22_X1  g361(.A1(new_n475), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n787), .A2(new_n473), .ZN(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT101), .B(KEYINPUT25), .ZN(new_n789));
  NAND3_X1  g364(.A1(new_n473), .A2(G103), .A3(G2104), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NOR3_X1   g366(.A1(new_n786), .A2(new_n788), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n792), .A2(G29), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G29), .B2(G33), .ZN(new_n794));
  INV_X1    g369(.A(G2072), .ZN(new_n795));
  AOI211_X1 g370(.A(new_n771), .B(new_n784), .C1(new_n794), .C2(new_n795), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n779), .A2(new_n777), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT107), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n781), .A2(G26), .ZN(new_n799));
  INV_X1    g374(.A(G140), .ZN(new_n800));
  NOR2_X1   g375(.A1(G104), .A2(G2105), .ZN(new_n801));
  OAI21_X1  g376(.A(G2104), .B1(new_n473), .B2(G116), .ZN(new_n802));
  OAI22_X1  g377(.A1(new_n481), .A2(new_n800), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n803), .B1(new_n487), .B2(G128), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n799), .B1(new_n804), .B2(new_n781), .ZN(new_n805));
  MUX2_X1   g380(.A(new_n799), .B(new_n805), .S(KEYINPUT28), .Z(new_n806));
  INV_X1    g381(.A(G2067), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n718), .A2(G20), .ZN(new_n809));
  OAI211_X1 g384(.A(KEYINPUT23), .B(new_n809), .C1(new_n620), .C2(new_n718), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(KEYINPUT23), .B2(new_n809), .ZN(new_n811));
  INV_X1    g386(.A(G1956), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  NOR2_X1   g388(.A1(G164), .A2(new_n781), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n814), .B1(G27), .B2(new_n781), .ZN(new_n815));
  INV_X1    g390(.A(G2078), .ZN(new_n816));
  AND2_X1   g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n815), .A2(new_n816), .ZN(new_n818));
  NOR3_X1   g393(.A1(new_n813), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  NAND4_X1  g394(.A1(new_n796), .A2(new_n798), .A3(new_n808), .A4(new_n819), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n794), .A2(new_n795), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT104), .ZN(new_n822));
  NOR2_X1   g397(.A1(G29), .A2(G32), .ZN(new_n823));
  AOI22_X1  g398(.A1(new_n487), .A2(G129), .B1(G105), .B2(new_n479), .ZN(new_n824));
  NAND3_X1  g399(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n825), .B(KEYINPUT26), .Z(new_n826));
  NAND2_X1  g401(.A1(new_n488), .A2(G141), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n824), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(KEYINPUT105), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n823), .B1(new_n829), .B2(G29), .ZN(new_n830));
  XOR2_X1   g405(.A(KEYINPUT27), .B(G1996), .Z(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT106), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n830), .B(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n781), .A2(G35), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n834), .B1(G162), .B2(new_n781), .ZN(new_n835));
  MUX2_X1   g410(.A(new_n834), .B(new_n835), .S(KEYINPUT110), .Z(new_n836));
  XOR2_X1   g411(.A(KEYINPUT111), .B(KEYINPUT29), .Z(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(G2090), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n836), .B(new_n838), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n822), .A2(new_n833), .A3(new_n839), .ZN(new_n840));
  OR2_X1    g415(.A1(KEYINPUT24), .A2(G34), .ZN(new_n841));
  NAND2_X1  g416(.A1(KEYINPUT24), .A2(G34), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n841), .A2(new_n781), .A3(new_n842), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n843), .B1(G160), .B2(new_n781), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n844), .A2(G2084), .ZN(new_n845));
  XOR2_X1   g420(.A(new_n845), .B(KEYINPUT103), .Z(new_n846));
  OAI221_X1 g421(.A(new_n846), .B1(G2084), .B2(new_n844), .C1(new_n760), .C2(new_n759), .ZN(new_n847));
  NOR3_X1   g422(.A1(new_n820), .A2(new_n840), .A3(new_n847), .ZN(new_n848));
  NAND4_X1  g423(.A1(new_n757), .A2(new_n761), .A3(new_n763), .A4(new_n848), .ZN(G150));
  INV_X1    g424(.A(G150), .ZN(G311));
  AOI22_X1  g425(.A1(new_n533), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n851));
  OR2_X1    g426(.A1(new_n851), .A2(new_n535), .ZN(new_n852));
  INV_X1    g427(.A(G93), .ZN(new_n853));
  INV_X1    g428(.A(G55), .ZN(new_n854));
  OAI22_X1  g429(.A1(new_n528), .A2(new_n853), .B1(new_n520), .B2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT112), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n858), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n856), .A2(new_n857), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n852), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n862), .A2(new_n627), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n861), .A2(new_n558), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  XOR2_X1   g440(.A(new_n865), .B(KEYINPUT39), .Z(new_n866));
  NAND2_X1  g441(.A1(new_n614), .A2(G559), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(KEYINPUT38), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n866), .B(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(G860), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  XOR2_X1   g446(.A(new_n871), .B(KEYINPUT113), .Z(new_n872));
  NAND2_X1  g447(.A1(new_n861), .A2(G860), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(KEYINPUT114), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(KEYINPUT37), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n872), .A2(new_n875), .ZN(G145));
  NAND2_X1  g451(.A1(new_n487), .A2(G130), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n488), .A2(G142), .ZN(new_n878));
  NOR2_X1   g453(.A1(G106), .A2(G2105), .ZN(new_n879));
  OAI21_X1  g454(.A(G2104), .B1(new_n473), .B2(G118), .ZN(new_n880));
  OAI211_X1 g455(.A(new_n877), .B(new_n878), .C1(new_n879), .C2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(new_n804), .ZN(new_n882));
  INV_X1    g457(.A(new_n747), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n882), .B(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n507), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n515), .A2(KEYINPUT4), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n886), .A2(new_n512), .ZN(new_n887));
  AOI21_X1  g462(.A(KEYINPUT115), .B1(new_n885), .B2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT115), .ZN(new_n889));
  NOR3_X1   g464(.A1(new_n507), .A2(new_n516), .A3(new_n889), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(new_n634), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n884), .B(new_n892), .ZN(new_n893));
  MUX2_X1   g468(.A(new_n828), .B(new_n829), .S(new_n792), .Z(new_n894));
  OR2_X1    g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n893), .A2(new_n894), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n641), .B(new_n484), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n898), .B(G162), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(G37), .ZN(new_n901));
  INV_X1    g476(.A(new_n899), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n895), .A2(new_n902), .A3(new_n896), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n900), .A2(new_n901), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(KEYINPUT40), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT40), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n900), .A2(new_n906), .A3(new_n901), .A4(new_n903), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n905), .A2(new_n907), .ZN(G395));
  NAND2_X1  g483(.A1(new_n865), .A2(KEYINPUT116), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT116), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n863), .A2(new_n910), .A3(new_n864), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n912), .B1(G559), .B2(new_n629), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n630), .A2(new_n909), .A3(new_n911), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n602), .A2(new_n611), .ZN(new_n915));
  OR3_X1    g490(.A1(new_n620), .A2(new_n915), .A3(KEYINPUT117), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n620), .A2(new_n915), .ZN(new_n917));
  NAND3_X1  g492(.A1(G299), .A2(new_n611), .A3(new_n602), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n917), .A2(KEYINPUT117), .A3(new_n918), .ZN(new_n919));
  NAND4_X1  g494(.A1(new_n913), .A2(new_n914), .A3(new_n916), .A4(new_n919), .ZN(new_n920));
  AND2_X1   g495(.A1(new_n913), .A2(new_n914), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT41), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n917), .A2(new_n922), .A3(new_n918), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n919), .A2(new_n916), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n923), .B1(new_n924), .B2(new_n922), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n920), .B1(new_n921), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n926), .A2(KEYINPUT42), .ZN(new_n927));
  NAND2_X1  g502(.A1(G166), .A2(G288), .ZN(new_n928));
  NAND2_X1  g503(.A1(G303), .A2(new_n720), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n930), .A2(new_n725), .ZN(new_n931));
  XNOR2_X1  g506(.A(G303), .B(G288), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n932), .A2(G305), .ZN(new_n933));
  OAI21_X1  g508(.A(G290), .B1(new_n931), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n930), .A2(new_n725), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n932), .A2(G305), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n935), .A2(new_n936), .A3(new_n598), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n934), .A2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT42), .ZN(new_n939));
  OAI211_X1 g514(.A(new_n939), .B(new_n920), .C1(new_n921), .C2(new_n925), .ZN(new_n940));
  AND3_X1   g515(.A1(new_n927), .A2(new_n938), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n938), .B1(new_n927), .B2(new_n940), .ZN(new_n942));
  OAI21_X1  g517(.A(G868), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n943), .B1(G868), .B2(new_n862), .ZN(G295));
  OAI21_X1  g519(.A(new_n943), .B1(G868), .B2(new_n862), .ZN(G331));
  AOI21_X1  g520(.A(G168), .B1(G301), .B2(KEYINPUT118), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  NOR2_X1   g522(.A1(G301), .A2(KEYINPUT118), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n863), .A2(new_n864), .A3(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n949), .B1(new_n863), .B2(new_n864), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n947), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(new_n952), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n954), .A2(new_n946), .A3(new_n950), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(new_n924), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n925), .A2(new_n953), .A3(new_n955), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(new_n938), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n924), .B1(new_n956), .B2(new_n922), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n917), .A2(new_n918), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n953), .A2(new_n955), .A3(KEYINPUT41), .A4(new_n962), .ZN(new_n963));
  NAND4_X1  g538(.A1(new_n961), .A2(new_n937), .A3(new_n934), .A4(new_n963), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n960), .A2(new_n964), .A3(KEYINPUT43), .A4(new_n901), .ZN(new_n965));
  AND3_X1   g540(.A1(new_n934), .A2(new_n937), .A3(KEYINPUT119), .ZN(new_n966));
  AND3_X1   g541(.A1(new_n966), .A2(new_n957), .A3(new_n958), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n966), .B1(new_n957), .B2(new_n958), .ZN(new_n968));
  NOR3_X1   g543(.A1(new_n967), .A2(new_n968), .A3(G37), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n965), .B1(new_n969), .B2(KEYINPUT43), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(KEYINPUT44), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT43), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n960), .A2(new_n964), .A3(new_n972), .A4(new_n901), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n973), .B1(new_n969), .B2(new_n972), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT44), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n971), .A2(new_n976), .ZN(G397));
  INV_X1    g552(.A(G1384), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n978), .B1(new_n888), .B2(new_n890), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT45), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n474), .A2(G40), .A3(new_n483), .A4(new_n480), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(G1996), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n829), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n828), .A2(G1996), .ZN(new_n987));
  XNOR2_X1  g562(.A(new_n804), .B(G2067), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n986), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  OR3_X1    g564(.A1(new_n989), .A2(new_n750), .A3(new_n883), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n804), .A2(new_n807), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n984), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  XOR2_X1   g567(.A(KEYINPUT126), .B(KEYINPUT46), .Z(new_n993));
  OAI21_X1  g568(.A(new_n993), .B1(new_n984), .B2(G1996), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT126), .ZN(new_n995));
  OAI211_X1 g570(.A(new_n983), .B(new_n985), .C1(new_n995), .C2(KEYINPUT46), .ZN(new_n996));
  INV_X1    g571(.A(new_n988), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n983), .B1(new_n997), .B2(new_n828), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n994), .A2(new_n996), .A3(new_n998), .ZN(new_n999));
  XOR2_X1   g574(.A(new_n999), .B(KEYINPUT47), .Z(new_n1000));
  XNOR2_X1  g575(.A(new_n747), .B(new_n750), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  OR2_X1    g577(.A1(new_n989), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(new_n983), .ZN(new_n1004));
  NOR3_X1   g579(.A1(new_n984), .A2(G1986), .A3(G290), .ZN(new_n1005));
  XOR2_X1   g580(.A(new_n1005), .B(KEYINPUT48), .Z(new_n1006));
  AOI211_X1 g581(.A(new_n992), .B(new_n1000), .C1(new_n1004), .C2(new_n1006), .ZN(new_n1007));
  OAI211_X1 g582(.A(KEYINPUT45), .B(new_n978), .C1(new_n888), .C2(new_n890), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n978), .B1(new_n507), .B2(new_n516), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n982), .B1(new_n980), .B2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(G1971), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1009), .A2(KEYINPUT50), .ZN(new_n1012));
  INV_X1    g587(.A(new_n982), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT50), .ZN(new_n1014));
  OAI211_X1 g589(.A(new_n1014), .B(new_n978), .C1(new_n507), .C2(new_n516), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1012), .A2(new_n1013), .A3(new_n1015), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n1016), .A2(G2090), .ZN(new_n1017));
  OR2_X1    g592(.A1(new_n1011), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(G303), .A2(G8), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT55), .ZN(new_n1020));
  XNOR2_X1  g595(.A(new_n1019), .B(new_n1020), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n1018), .A2(KEYINPUT120), .A3(G8), .A4(new_n1021), .ZN(new_n1022));
  OAI211_X1 g597(.A(new_n1021), .B(G8), .C1(new_n1011), .C2(new_n1017), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT120), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1022), .A2(new_n1025), .ZN(new_n1026));
  XOR2_X1   g601(.A(G305), .B(G1981), .Z(new_n1027));
  AND2_X1   g602(.A1(new_n1027), .A2(KEYINPUT49), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n982), .A2(new_n1009), .ZN(new_n1029));
  INV_X1    g604(.A(G8), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1031), .B1(new_n1027), .B2(KEYINPUT49), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1028), .A2(new_n1032), .ZN(new_n1033));
  OR3_X1    g608(.A1(new_n1029), .A2(KEYINPUT121), .A3(new_n1030), .ZN(new_n1034));
  INV_X1    g609(.A(G1976), .ZN(new_n1035));
  NOR2_X1   g610(.A1(G288), .A2(new_n1035), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1034), .A2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1031), .A2(new_n1035), .A3(G288), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1037), .B1(new_n1039), .B2(KEYINPUT52), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT52), .ZN(new_n1041));
  OAI211_X1 g616(.A(new_n1038), .B(new_n1041), .C1(new_n1034), .C2(new_n1036), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1033), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1016), .A2(G2084), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1009), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(KEYINPUT45), .ZN(new_n1046));
  AOI21_X1  g621(.A(G1966), .B1(new_n1010), .B2(new_n1046), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1044), .A2(new_n1047), .ZN(new_n1048));
  NOR3_X1   g623(.A1(new_n1048), .A2(new_n1030), .A3(G286), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1018), .A2(G8), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1021), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1026), .A2(new_n1043), .A3(new_n1049), .A4(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(KEYINPUT63), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1043), .A2(new_n1025), .A3(new_n1022), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1035), .B1(new_n1028), .B2(new_n1032), .ZN(new_n1056));
  OAI22_X1  g631(.A1(new_n1056), .A2(G288), .B1(G1981), .B2(G305), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(new_n1031), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1054), .A2(new_n1055), .A3(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT63), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1049), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT125), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1008), .A2(new_n816), .A3(new_n1010), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT53), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1016), .A2(new_n770), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1064), .A2(G2078), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1010), .A2(new_n1046), .A3(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1065), .A2(new_n1066), .A3(new_n1068), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1062), .B1(new_n1069), .B2(G171), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1069), .A2(new_n1062), .A3(G171), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NOR2_X1   g648(.A1(G168), .A2(new_n1030), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(KEYINPUT51), .B1(new_n1075), .B2(KEYINPUT124), .ZN(new_n1076));
  AND2_X1   g651(.A1(new_n1010), .A2(new_n1046), .ZN(new_n1077));
  OAI22_X1  g652(.A1(new_n1077), .A2(G1966), .B1(G2084), .B2(new_n1016), .ZN(new_n1078));
  OAI211_X1 g653(.A(G8), .B(new_n1076), .C1(new_n1078), .C2(G286), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1076), .ZN(new_n1080));
  OAI211_X1 g655(.A(new_n1075), .B(new_n1080), .C1(new_n1048), .C2(new_n1030), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1078), .A2(G8), .A3(G286), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1079), .A2(new_n1081), .A3(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(KEYINPUT62), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT62), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1079), .A2(new_n1081), .A3(new_n1085), .A4(new_n1082), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1073), .A2(new_n1084), .A3(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT57), .ZN(new_n1088));
  XNOR2_X1  g663(.A(G299), .B(new_n1088), .ZN(new_n1089));
  XNOR2_X1  g664(.A(KEYINPUT56), .B(G2072), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1008), .A2(new_n1010), .A3(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1016), .A2(new_n812), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1089), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1091), .A2(new_n1092), .A3(new_n1089), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1016), .A2(new_n760), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1029), .A2(new_n807), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n629), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1093), .B1(new_n1094), .B2(new_n1097), .ZN(new_n1098));
  OR2_X1    g673(.A1(new_n1094), .A2(KEYINPUT61), .ZN(new_n1099));
  AND3_X1   g674(.A1(new_n1095), .A2(new_n629), .A3(new_n1096), .ZN(new_n1100));
  OAI21_X1  g675(.A(KEYINPUT60), .B1(new_n1100), .B2(new_n1097), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n629), .A2(KEYINPUT60), .ZN(new_n1102));
  AOI22_X1  g677(.A1(new_n1016), .A2(new_n760), .B1(new_n807), .B2(new_n1029), .ZN(new_n1103));
  AOI22_X1  g678(.A1(new_n1094), .A2(KEYINPUT61), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1099), .A2(new_n1101), .A3(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1008), .A2(new_n985), .A3(new_n1010), .ZN(new_n1106));
  XNOR2_X1  g681(.A(KEYINPUT122), .B(KEYINPUT58), .ZN(new_n1107));
  XNOR2_X1  g682(.A(new_n1107), .B(G1341), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1108), .B1(new_n982), .B2(new_n1009), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n627), .B1(new_n1106), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(KEYINPUT123), .A2(KEYINPUT59), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1111), .ZN(new_n1112));
  XNOR2_X1  g687(.A(new_n1110), .B(new_n1112), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1098), .B1(new_n1105), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(new_n1083), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n981), .A2(new_n1013), .A3(new_n1008), .A4(new_n1067), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1065), .A2(new_n1116), .A3(G171), .A4(new_n1066), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(KEYINPUT54), .ZN(new_n1118));
  AOI22_X1  g693(.A1(new_n1063), .A2(new_n1064), .B1(new_n770), .B2(new_n1016), .ZN(new_n1119));
  AOI21_X1  g694(.A(G171), .B1(new_n1119), .B2(new_n1068), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1121));
  AOI211_X1 g696(.A(KEYINPUT125), .B(G301), .C1(new_n1119), .C2(new_n1068), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1122), .A2(new_n1070), .ZN(new_n1123));
  AND2_X1   g698(.A1(new_n1119), .A2(new_n1116), .ZN(new_n1124));
  AOI21_X1  g699(.A(KEYINPUT54), .B1(new_n1124), .B2(G301), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1121), .B1(new_n1123), .B2(new_n1125), .ZN(new_n1126));
  OAI211_X1 g701(.A(new_n1061), .B(new_n1087), .C1(new_n1115), .C2(new_n1126), .ZN(new_n1127));
  AND3_X1   g702(.A1(new_n1026), .A2(new_n1043), .A3(new_n1052), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1059), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1003), .ZN(new_n1130));
  XNOR2_X1  g705(.A(new_n598), .B(G1986), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n984), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1007), .B1(new_n1129), .B2(new_n1132), .ZN(G329));
  assign    G231 = 1'b0;
  NAND4_X1  g708(.A1(new_n670), .A2(KEYINPUT127), .A3(G319), .A4(new_n687), .ZN(new_n1135));
  NAND2_X1  g709(.A1(new_n1135), .A2(new_n716), .ZN(new_n1136));
  AOI21_X1  g710(.A(new_n461), .B1(new_n668), .B2(new_n669), .ZN(new_n1137));
  AOI21_X1  g711(.A(KEYINPUT127), .B1(new_n1137), .B2(new_n687), .ZN(new_n1138));
  NOR2_X1   g712(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1139));
  AND3_X1   g713(.A1(new_n1139), .A2(new_n904), .A3(new_n974), .ZN(G308));
  NAND3_X1  g714(.A1(new_n1139), .A2(new_n904), .A3(new_n974), .ZN(G225));
endmodule


