

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587;

  XOR2_X1 U325 ( .A(G190GAT), .B(KEYINPUT75), .Z(n412) );
  XNOR2_X1 U326 ( .A(n424), .B(n423), .ZN(n426) );
  XNOR2_X1 U327 ( .A(n471), .B(KEYINPUT55), .ZN(n472) );
  XOR2_X1 U328 ( .A(n360), .B(n316), .Z(n537) );
  XNOR2_X1 U329 ( .A(n362), .B(n361), .ZN(n366) );
  AND2_X1 U330 ( .A1(G226GAT), .A2(G233GAT), .ZN(n293) );
  XOR2_X1 U331 ( .A(KEYINPUT33), .B(KEYINPUT32), .Z(n294) );
  XNOR2_X1 U332 ( .A(n422), .B(KEYINPUT31), .ZN(n423) );
  INV_X1 U333 ( .A(KEYINPUT48), .ZN(n463) );
  XNOR2_X1 U334 ( .A(n463), .B(KEYINPUT64), .ZN(n464) );
  XNOR2_X1 U335 ( .A(n412), .B(n293), .ZN(n357) );
  XNOR2_X1 U336 ( .A(n427), .B(n294), .ZN(n428) );
  XNOR2_X1 U337 ( .A(n427), .B(n413), .ZN(n414) );
  XNOR2_X1 U338 ( .A(n430), .B(n357), .ZN(n358) );
  XNOR2_X1 U339 ( .A(n429), .B(n428), .ZN(n433) );
  XNOR2_X1 U340 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U341 ( .A(n360), .B(n359), .ZN(n361) );
  OR2_X1 U342 ( .A1(n522), .A2(n491), .ZN(n448) );
  INV_X1 U343 ( .A(G43GAT), .ZN(n449) );
  XNOR2_X1 U344 ( .A(n448), .B(KEYINPUT38), .ZN(n507) );
  XNOR2_X1 U345 ( .A(n484), .B(KEYINPUT58), .ZN(n485) );
  XNOR2_X1 U346 ( .A(n449), .B(KEYINPUT40), .ZN(n450) );
  XNOR2_X1 U347 ( .A(n486), .B(n485), .ZN(G1351GAT) );
  XNOR2_X1 U348 ( .A(n451), .B(n450), .ZN(G1330GAT) );
  XOR2_X1 U349 ( .A(KEYINPUT19), .B(KEYINPUT85), .Z(n296) );
  XNOR2_X1 U350 ( .A(KEYINPUT17), .B(G183GAT), .ZN(n295) );
  XNOR2_X1 U351 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U352 ( .A(KEYINPUT18), .B(n297), .Z(n360) );
  XOR2_X1 U353 ( .A(G176GAT), .B(KEYINPUT86), .Z(n299) );
  XNOR2_X1 U354 ( .A(KEYINPUT20), .B(KEYINPUT83), .ZN(n298) );
  XNOR2_X1 U355 ( .A(n299), .B(n298), .ZN(n303) );
  XOR2_X1 U356 ( .A(KEYINPUT87), .B(KEYINPUT82), .Z(n301) );
  XNOR2_X1 U357 ( .A(G169GAT), .B(G15GAT), .ZN(n300) );
  XNOR2_X1 U358 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U359 ( .A(n303), .B(n302), .Z(n315) );
  XNOR2_X1 U360 ( .A(G127GAT), .B(KEYINPUT80), .ZN(n304) );
  XNOR2_X1 U361 ( .A(n304), .B(KEYINPUT81), .ZN(n305) );
  XOR2_X1 U362 ( .A(n305), .B(KEYINPUT0), .Z(n307) );
  XNOR2_X1 U363 ( .A(G113GAT), .B(G134GAT), .ZN(n306) );
  XNOR2_X1 U364 ( .A(n307), .B(n306), .ZN(n355) );
  XOR2_X1 U365 ( .A(G120GAT), .B(G71GAT), .Z(n431) );
  XOR2_X1 U366 ( .A(KEYINPUT84), .B(G190GAT), .Z(n309) );
  XNOR2_X1 U367 ( .A(G43GAT), .B(G99GAT), .ZN(n308) );
  XNOR2_X1 U368 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U369 ( .A(n431), .B(n310), .Z(n312) );
  NAND2_X1 U370 ( .A1(G227GAT), .A2(G233GAT), .ZN(n311) );
  XNOR2_X1 U371 ( .A(n312), .B(n311), .ZN(n313) );
  XNOR2_X1 U372 ( .A(n355), .B(n313), .ZN(n314) );
  XNOR2_X1 U373 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U374 ( .A(G211GAT), .B(G155GAT), .Z(n318) );
  XNOR2_X1 U375 ( .A(G183GAT), .B(G71GAT), .ZN(n317) );
  XNOR2_X1 U376 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U377 ( .A(KEYINPUT13), .B(G57GAT), .Z(n425) );
  XOR2_X1 U378 ( .A(n319), .B(n425), .Z(n321) );
  XNOR2_X1 U379 ( .A(G22GAT), .B(G78GAT), .ZN(n320) );
  XNOR2_X1 U380 ( .A(n321), .B(n320), .ZN(n326) );
  XNOR2_X1 U381 ( .A(G15GAT), .B(G1GAT), .ZN(n322) );
  XNOR2_X1 U382 ( .A(n322), .B(KEYINPUT71), .ZN(n434) );
  XOR2_X1 U383 ( .A(n434), .B(KEYINPUT12), .Z(n324) );
  NAND2_X1 U384 ( .A1(G231GAT), .A2(G233GAT), .ZN(n323) );
  XNOR2_X1 U385 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U386 ( .A(n326), .B(n325), .Z(n334) );
  XOR2_X1 U387 ( .A(KEYINPUT78), .B(G64GAT), .Z(n328) );
  XNOR2_X1 U388 ( .A(G8GAT), .B(G127GAT), .ZN(n327) );
  XNOR2_X1 U389 ( .A(n328), .B(n327), .ZN(n332) );
  XOR2_X1 U390 ( .A(KEYINPUT77), .B(KEYINPUT76), .Z(n330) );
  XNOR2_X1 U391 ( .A(KEYINPUT15), .B(KEYINPUT14), .ZN(n329) );
  XNOR2_X1 U392 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U393 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U394 ( .A(n334), .B(n333), .Z(n567) );
  XOR2_X1 U395 ( .A(KEYINPUT6), .B(G57GAT), .Z(n336) );
  XNOR2_X1 U396 ( .A(G1GAT), .B(G120GAT), .ZN(n335) );
  XNOR2_X1 U397 ( .A(n336), .B(n335), .ZN(n340) );
  XOR2_X1 U398 ( .A(G85GAT), .B(G148GAT), .Z(n338) );
  XNOR2_X1 U399 ( .A(G29GAT), .B(G141GAT), .ZN(n337) );
  XNOR2_X1 U400 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U401 ( .A(n340), .B(n339), .ZN(n353) );
  XOR2_X1 U402 ( .A(KEYINPUT4), .B(KEYINPUT95), .Z(n342) );
  XNOR2_X1 U403 ( .A(KEYINPUT94), .B(KEYINPUT93), .ZN(n341) );
  XNOR2_X1 U404 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U405 ( .A(KEYINPUT5), .B(n343), .Z(n345) );
  NAND2_X1 U406 ( .A1(G225GAT), .A2(G233GAT), .ZN(n344) );
  XNOR2_X1 U407 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U408 ( .A(n346), .B(KEYINPUT1), .Z(n351) );
  XOR2_X1 U409 ( .A(KEYINPUT90), .B(G162GAT), .Z(n348) );
  XNOR2_X1 U410 ( .A(KEYINPUT2), .B(G155GAT), .ZN(n347) );
  XNOR2_X1 U411 ( .A(n348), .B(n347), .ZN(n349) );
  XOR2_X1 U412 ( .A(KEYINPUT3), .B(n349), .Z(n380) );
  XNOR2_X1 U413 ( .A(n380), .B(KEYINPUT96), .ZN(n350) );
  XNOR2_X1 U414 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U415 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U416 ( .A(n355), .B(n354), .ZN(n523) );
  XNOR2_X1 U417 ( .A(G176GAT), .B(G92GAT), .ZN(n356) );
  XNOR2_X1 U418 ( .A(n356), .B(G64GAT), .ZN(n430) );
  XOR2_X1 U419 ( .A(n358), .B(G204GAT), .Z(n362) );
  XOR2_X1 U420 ( .A(G169GAT), .B(G8GAT), .Z(n438) );
  XNOR2_X1 U421 ( .A(G36GAT), .B(n438), .ZN(n359) );
  XOR2_X1 U422 ( .A(KEYINPUT89), .B(G218GAT), .Z(n364) );
  XNOR2_X1 U423 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n363) );
  XNOR2_X1 U424 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U425 ( .A(G197GAT), .B(n365), .ZN(n379) );
  XOR2_X1 U426 ( .A(n366), .B(n379), .Z(n525) );
  XNOR2_X1 U427 ( .A(KEYINPUT27), .B(n525), .ZN(n387) );
  NOR2_X1 U428 ( .A1(n523), .A2(n387), .ZN(n367) );
  XOR2_X1 U429 ( .A(KEYINPUT97), .B(n367), .Z(n532) );
  XOR2_X1 U430 ( .A(KEYINPUT88), .B(KEYINPUT22), .Z(n369) );
  XNOR2_X1 U431 ( .A(KEYINPUT91), .B(KEYINPUT24), .ZN(n368) );
  XNOR2_X1 U432 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U433 ( .A(n370), .B(KEYINPUT23), .Z(n372) );
  XOR2_X1 U434 ( .A(G141GAT), .B(G22GAT), .Z(n435) );
  XNOR2_X1 U435 ( .A(G50GAT), .B(n435), .ZN(n371) );
  XNOR2_X1 U436 ( .A(n372), .B(n371), .ZN(n378) );
  XOR2_X1 U437 ( .A(G78GAT), .B(G148GAT), .Z(n374) );
  XNOR2_X1 U438 ( .A(G106GAT), .B(G204GAT), .ZN(n373) );
  XNOR2_X1 U439 ( .A(n374), .B(n373), .ZN(n424) );
  XOR2_X1 U440 ( .A(KEYINPUT92), .B(n424), .Z(n376) );
  NAND2_X1 U441 ( .A1(G228GAT), .A2(G233GAT), .ZN(n375) );
  XNOR2_X1 U442 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U443 ( .A(n378), .B(n377), .Z(n382) );
  XOR2_X1 U444 ( .A(n380), .B(n379), .Z(n381) );
  XOR2_X1 U445 ( .A(n382), .B(n381), .Z(n388) );
  XNOR2_X1 U446 ( .A(n388), .B(KEYINPUT28), .ZN(n535) );
  AND2_X1 U447 ( .A1(n537), .A2(n535), .ZN(n383) );
  NAND2_X1 U448 ( .A1(n532), .A2(n383), .ZN(n384) );
  XNOR2_X1 U449 ( .A(n384), .B(KEYINPUT98), .ZN(n396) );
  INV_X1 U450 ( .A(n388), .ZN(n470) );
  NAND2_X1 U451 ( .A1(n470), .A2(n537), .ZN(n385) );
  XNOR2_X1 U452 ( .A(n385), .B(KEYINPUT99), .ZN(n386) );
  XNOR2_X1 U453 ( .A(KEYINPUT26), .B(n386), .ZN(n552) );
  INV_X1 U454 ( .A(n552), .ZN(n571) );
  OR2_X1 U455 ( .A1(n571), .A2(n387), .ZN(n393) );
  INV_X1 U456 ( .A(n537), .ZN(n474) );
  INV_X1 U457 ( .A(n525), .ZN(n466) );
  NAND2_X1 U458 ( .A1(n474), .A2(n466), .ZN(n389) );
  NAND2_X1 U459 ( .A1(n389), .A2(n388), .ZN(n390) );
  XNOR2_X1 U460 ( .A(n390), .B(KEYINPUT100), .ZN(n391) );
  XOR2_X1 U461 ( .A(KEYINPUT25), .B(n391), .Z(n392) );
  NAND2_X1 U462 ( .A1(n393), .A2(n392), .ZN(n394) );
  NAND2_X1 U463 ( .A1(n394), .A2(n523), .ZN(n395) );
  NAND2_X1 U464 ( .A1(n396), .A2(n395), .ZN(n489) );
  NAND2_X1 U465 ( .A1(n567), .A2(n489), .ZN(n397) );
  XNOR2_X1 U466 ( .A(KEYINPUT104), .B(n397), .ZN(n420) );
  XOR2_X1 U467 ( .A(G43GAT), .B(G29GAT), .Z(n399) );
  XNOR2_X1 U468 ( .A(KEYINPUT8), .B(G50GAT), .ZN(n398) );
  XNOR2_X1 U469 ( .A(n399), .B(n398), .ZN(n400) );
  XOR2_X1 U470 ( .A(n400), .B(KEYINPUT70), .Z(n402) );
  XNOR2_X1 U471 ( .A(G36GAT), .B(KEYINPUT7), .ZN(n401) );
  XNOR2_X1 U472 ( .A(n402), .B(n401), .ZN(n445) );
  XOR2_X1 U473 ( .A(KEYINPUT65), .B(KEYINPUT9), .Z(n404) );
  XNOR2_X1 U474 ( .A(G106GAT), .B(KEYINPUT67), .ZN(n403) );
  XNOR2_X1 U475 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U476 ( .A(n445), .B(n405), .ZN(n419) );
  XOR2_X1 U477 ( .A(KEYINPUT74), .B(KEYINPUT73), .Z(n407) );
  XNOR2_X1 U478 ( .A(G218GAT), .B(G92GAT), .ZN(n406) );
  XNOR2_X1 U479 ( .A(n407), .B(n406), .ZN(n411) );
  XOR2_X1 U480 ( .A(KEYINPUT66), .B(KEYINPUT11), .Z(n409) );
  XNOR2_X1 U481 ( .A(G134GAT), .B(G162GAT), .ZN(n408) );
  XNOR2_X1 U482 ( .A(n409), .B(n408), .ZN(n410) );
  XOR2_X1 U483 ( .A(n411), .B(n410), .Z(n417) );
  XOR2_X1 U484 ( .A(KEYINPUT10), .B(n412), .Z(n415) );
  XOR2_X1 U485 ( .A(G99GAT), .B(G85GAT), .Z(n427) );
  NAND2_X1 U486 ( .A1(G232GAT), .A2(G233GAT), .ZN(n413) );
  XNOR2_X1 U487 ( .A(n417), .B(n416), .ZN(n418) );
  XOR2_X1 U488 ( .A(n419), .B(n418), .Z(n547) );
  XOR2_X1 U489 ( .A(KEYINPUT36), .B(n547), .Z(n584) );
  NOR2_X1 U490 ( .A1(n420), .A2(n584), .ZN(n421) );
  XNOR2_X1 U491 ( .A(n421), .B(KEYINPUT37), .ZN(n522) );
  NAND2_X1 U492 ( .A1(G230GAT), .A2(G233GAT), .ZN(n422) );
  XNOR2_X1 U493 ( .A(n426), .B(n425), .ZN(n429) );
  XNOR2_X1 U494 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U495 ( .A(n433), .B(n432), .ZN(n576) );
  XOR2_X1 U496 ( .A(n435), .B(n434), .Z(n437) );
  NAND2_X1 U497 ( .A1(G229GAT), .A2(G233GAT), .ZN(n436) );
  XNOR2_X1 U498 ( .A(n437), .B(n436), .ZN(n439) );
  XOR2_X1 U499 ( .A(n439), .B(n438), .Z(n441) );
  XNOR2_X1 U500 ( .A(G197GAT), .B(G113GAT), .ZN(n440) );
  XNOR2_X1 U501 ( .A(n441), .B(n440), .ZN(n447) );
  XOR2_X1 U502 ( .A(KEYINPUT68), .B(KEYINPUT69), .Z(n443) );
  XNOR2_X1 U503 ( .A(KEYINPUT30), .B(KEYINPUT29), .ZN(n442) );
  XNOR2_X1 U504 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U505 ( .A(n445), .B(n444), .Z(n446) );
  XOR2_X1 U506 ( .A(n447), .B(n446), .Z(n572) );
  XOR2_X1 U507 ( .A(KEYINPUT72), .B(n572), .Z(n478) );
  INV_X1 U508 ( .A(n478), .ZN(n538) );
  NAND2_X1 U509 ( .A1(n576), .A2(n538), .ZN(n491) );
  NOR2_X1 U510 ( .A1(n537), .A2(n507), .ZN(n451) );
  XNOR2_X1 U511 ( .A(n576), .B(KEYINPUT41), .ZN(n540) );
  AND2_X1 U512 ( .A1(n572), .A2(n540), .ZN(n453) );
  XNOR2_X1 U513 ( .A(KEYINPUT46), .B(KEYINPUT112), .ZN(n452) );
  XNOR2_X1 U514 ( .A(n453), .B(n452), .ZN(n455) );
  INV_X1 U515 ( .A(n547), .ZN(n565) );
  NAND2_X1 U516 ( .A1(n567), .A2(n565), .ZN(n454) );
  OR2_X1 U517 ( .A1(n455), .A2(n454), .ZN(n456) );
  XNOR2_X1 U518 ( .A(n456), .B(KEYINPUT47), .ZN(n462) );
  NOR2_X1 U519 ( .A1(n584), .A2(n567), .ZN(n457) );
  XNOR2_X1 U520 ( .A(KEYINPUT45), .B(n457), .ZN(n458) );
  AND2_X1 U521 ( .A1(n458), .A2(n576), .ZN(n459) );
  XNOR2_X1 U522 ( .A(n459), .B(KEYINPUT113), .ZN(n460) );
  NOR2_X1 U523 ( .A1(n538), .A2(n460), .ZN(n461) );
  NOR2_X1 U524 ( .A1(n462), .A2(n461), .ZN(n465) );
  XNOR2_X1 U525 ( .A(n465), .B(n464), .ZN(n533) );
  NAND2_X1 U526 ( .A1(n466), .A2(n533), .ZN(n467) );
  XNOR2_X1 U527 ( .A(n467), .B(KEYINPUT121), .ZN(n468) );
  XNOR2_X1 U528 ( .A(n468), .B(KEYINPUT54), .ZN(n469) );
  NAND2_X1 U529 ( .A1(n469), .A2(n523), .ZN(n570) );
  NOR2_X1 U530 ( .A1(n470), .A2(n570), .ZN(n473) );
  XNOR2_X1 U531 ( .A(KEYINPUT122), .B(KEYINPUT123), .ZN(n471) );
  XNOR2_X1 U532 ( .A(n473), .B(n472), .ZN(n475) );
  AND2_X1 U533 ( .A1(n475), .A2(n474), .ZN(n477) );
  INV_X1 U534 ( .A(KEYINPUT124), .ZN(n476) );
  XNOR2_X1 U535 ( .A(n477), .B(n476), .ZN(n568) );
  NOR2_X1 U536 ( .A1(n478), .A2(n568), .ZN(n480) );
  XNOR2_X1 U537 ( .A(G169GAT), .B(KEYINPUT125), .ZN(n479) );
  XNOR2_X1 U538 ( .A(n480), .B(n479), .ZN(G1348GAT) );
  INV_X1 U539 ( .A(n540), .ZN(n555) );
  NOR2_X1 U540 ( .A1(n555), .A2(n568), .ZN(n483) );
  XNOR2_X1 U541 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n481) );
  XNOR2_X1 U542 ( .A(n481), .B(G176GAT), .ZN(n482) );
  XNOR2_X1 U543 ( .A(n483), .B(n482), .ZN(G1349GAT) );
  NOR2_X1 U544 ( .A1(n565), .A2(n568), .ZN(n486) );
  INV_X1 U545 ( .A(G190GAT), .ZN(n484) );
  INV_X1 U546 ( .A(n567), .ZN(n580) );
  NAND2_X1 U547 ( .A1(n580), .A2(n565), .ZN(n487) );
  XNOR2_X1 U548 ( .A(n487), .B(KEYINPUT79), .ZN(n488) );
  XNOR2_X1 U549 ( .A(n488), .B(KEYINPUT16), .ZN(n490) );
  NAND2_X1 U550 ( .A1(n490), .A2(n489), .ZN(n510) );
  NOR2_X1 U551 ( .A1(n510), .A2(n491), .ZN(n492) );
  XNOR2_X1 U552 ( .A(n492), .B(KEYINPUT101), .ZN(n498) );
  NOR2_X1 U553 ( .A1(n523), .A2(n498), .ZN(n493) );
  XOR2_X1 U554 ( .A(KEYINPUT34), .B(n493), .Z(n494) );
  XNOR2_X1 U555 ( .A(G1GAT), .B(n494), .ZN(G1324GAT) );
  NOR2_X1 U556 ( .A1(n525), .A2(n498), .ZN(n495) );
  XOR2_X1 U557 ( .A(G8GAT), .B(n495), .Z(G1325GAT) );
  NOR2_X1 U558 ( .A1(n537), .A2(n498), .ZN(n497) );
  XNOR2_X1 U559 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n496) );
  XNOR2_X1 U560 ( .A(n497), .B(n496), .ZN(G1326GAT) );
  NOR2_X1 U561 ( .A1(n535), .A2(n498), .ZN(n499) );
  XOR2_X1 U562 ( .A(KEYINPUT102), .B(n499), .Z(n500) );
  XNOR2_X1 U563 ( .A(G22GAT), .B(n500), .ZN(G1327GAT) );
  NOR2_X1 U564 ( .A1(n507), .A2(n523), .ZN(n503) );
  XOR2_X1 U565 ( .A(G29GAT), .B(KEYINPUT103), .Z(n501) );
  XNOR2_X1 U566 ( .A(KEYINPUT39), .B(n501), .ZN(n502) );
  XNOR2_X1 U567 ( .A(n503), .B(n502), .ZN(G1328GAT) );
  XNOR2_X1 U568 ( .A(KEYINPUT105), .B(KEYINPUT106), .ZN(n505) );
  NOR2_X1 U569 ( .A1(n525), .A2(n507), .ZN(n504) );
  XNOR2_X1 U570 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U571 ( .A(G36GAT), .B(n506), .ZN(G1329GAT) );
  XNOR2_X1 U572 ( .A(G50GAT), .B(KEYINPUT107), .ZN(n509) );
  NOR2_X1 U573 ( .A1(n535), .A2(n507), .ZN(n508) );
  XNOR2_X1 U574 ( .A(n509), .B(n508), .ZN(G1331GAT) );
  INV_X1 U575 ( .A(n572), .ZN(n553) );
  NAND2_X1 U576 ( .A1(n553), .A2(n540), .ZN(n521) );
  OR2_X1 U577 ( .A1(n521), .A2(n510), .ZN(n518) );
  NOR2_X1 U578 ( .A1(n523), .A2(n518), .ZN(n511) );
  XOR2_X1 U579 ( .A(n511), .B(KEYINPUT42), .Z(n512) );
  XNOR2_X1 U580 ( .A(G57GAT), .B(n512), .ZN(G1332GAT) );
  NOR2_X1 U581 ( .A1(n525), .A2(n518), .ZN(n514) );
  XNOR2_X1 U582 ( .A(KEYINPUT108), .B(KEYINPUT109), .ZN(n513) );
  XNOR2_X1 U583 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U584 ( .A(G64GAT), .B(n515), .ZN(G1333GAT) );
  NOR2_X1 U585 ( .A1(n537), .A2(n518), .ZN(n516) );
  XOR2_X1 U586 ( .A(KEYINPUT110), .B(n516), .Z(n517) );
  XNOR2_X1 U587 ( .A(G71GAT), .B(n517), .ZN(G1334GAT) );
  NOR2_X1 U588 ( .A1(n535), .A2(n518), .ZN(n520) );
  XNOR2_X1 U589 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n519) );
  XNOR2_X1 U590 ( .A(n520), .B(n519), .ZN(G1335GAT) );
  OR2_X1 U591 ( .A1(n522), .A2(n521), .ZN(n529) );
  NOR2_X1 U592 ( .A1(n523), .A2(n529), .ZN(n524) );
  XOR2_X1 U593 ( .A(G85GAT), .B(n524), .Z(G1336GAT) );
  NOR2_X1 U594 ( .A1(n525), .A2(n529), .ZN(n527) );
  XNOR2_X1 U595 ( .A(G92GAT), .B(KEYINPUT111), .ZN(n526) );
  XNOR2_X1 U596 ( .A(n527), .B(n526), .ZN(G1337GAT) );
  NOR2_X1 U597 ( .A1(n537), .A2(n529), .ZN(n528) );
  XOR2_X1 U598 ( .A(G99GAT), .B(n528), .Z(G1338GAT) );
  NOR2_X1 U599 ( .A1(n535), .A2(n529), .ZN(n530) );
  XOR2_X1 U600 ( .A(KEYINPUT44), .B(n530), .Z(n531) );
  XNOR2_X1 U601 ( .A(G106GAT), .B(n531), .ZN(G1339GAT) );
  NAND2_X1 U602 ( .A1(n533), .A2(n532), .ZN(n534) );
  XOR2_X1 U603 ( .A(KEYINPUT114), .B(n534), .Z(n551) );
  NAND2_X1 U604 ( .A1(n535), .A2(n551), .ZN(n536) );
  NOR2_X1 U605 ( .A1(n537), .A2(n536), .ZN(n548) );
  NAND2_X1 U606 ( .A1(n548), .A2(n538), .ZN(n539) );
  XNOR2_X1 U607 ( .A(G113GAT), .B(n539), .ZN(G1340GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT115), .B(KEYINPUT49), .Z(n542) );
  NAND2_X1 U609 ( .A1(n548), .A2(n540), .ZN(n541) );
  XNOR2_X1 U610 ( .A(n542), .B(n541), .ZN(n543) );
  XOR2_X1 U611 ( .A(G120GAT), .B(n543), .Z(G1341GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT116), .B(KEYINPUT50), .Z(n545) );
  NAND2_X1 U613 ( .A1(n548), .A2(n580), .ZN(n544) );
  XNOR2_X1 U614 ( .A(n545), .B(n544), .ZN(n546) );
  XOR2_X1 U615 ( .A(G127GAT), .B(n546), .Z(G1342GAT) );
  XOR2_X1 U616 ( .A(G134GAT), .B(KEYINPUT51), .Z(n550) );
  NAND2_X1 U617 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U618 ( .A(n550), .B(n549), .ZN(G1343GAT) );
  NAND2_X1 U619 ( .A1(n552), .A2(n551), .ZN(n564) );
  NOR2_X1 U620 ( .A1(n553), .A2(n564), .ZN(n554) );
  XOR2_X1 U621 ( .A(G141GAT), .B(n554), .Z(G1344GAT) );
  NOR2_X1 U622 ( .A1(n564), .A2(n555), .ZN(n562) );
  XOR2_X1 U623 ( .A(KEYINPUT117), .B(KEYINPUT119), .Z(n557) );
  XNOR2_X1 U624 ( .A(KEYINPUT52), .B(KEYINPUT53), .ZN(n556) );
  XNOR2_X1 U625 ( .A(n557), .B(n556), .ZN(n558) );
  XOR2_X1 U626 ( .A(n558), .B(KEYINPUT120), .Z(n560) );
  XNOR2_X1 U627 ( .A(G148GAT), .B(KEYINPUT118), .ZN(n559) );
  XNOR2_X1 U628 ( .A(n560), .B(n559), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n562), .B(n561), .ZN(G1345GAT) );
  NOR2_X1 U630 ( .A1(n567), .A2(n564), .ZN(n563) );
  XOR2_X1 U631 ( .A(G155GAT), .B(n563), .Z(G1346GAT) );
  NOR2_X1 U632 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U633 ( .A(G162GAT), .B(n566), .Z(G1347GAT) );
  NOR2_X1 U634 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U635 ( .A(G183GAT), .B(n569), .Z(G1350GAT) );
  XOR2_X1 U636 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n574) );
  NOR2_X1 U637 ( .A1(n571), .A2(n570), .ZN(n581) );
  NAND2_X1 U638 ( .A1(n581), .A2(n572), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U640 ( .A(G197GAT), .B(n575), .ZN(G1352GAT) );
  XOR2_X1 U641 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n578) );
  INV_X1 U642 ( .A(n581), .ZN(n583) );
  OR2_X1 U643 ( .A1(n583), .A2(n576), .ZN(n577) );
  XNOR2_X1 U644 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U645 ( .A(G204GAT), .B(n579), .ZN(G1353GAT) );
  NAND2_X1 U646 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n582), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U648 ( .A1(n584), .A2(n583), .ZN(n586) );
  XNOR2_X1 U649 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n585) );
  XNOR2_X1 U650 ( .A(n586), .B(n585), .ZN(n587) );
  XNOR2_X1 U651 ( .A(G218GAT), .B(n587), .ZN(G1355GAT) );
endmodule

