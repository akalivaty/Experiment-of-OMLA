//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 0 1 1 0 0 0 1 0 0 0 0 1 1 0 0 0 1 1 1 0 0 1 1 0 0 0 0 0 0 0 1 1 0 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 0 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:43 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n682,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n699, new_n701, new_n702, new_n703, new_n704, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n730, new_n731, new_n732, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n744, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n768,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n885, new_n886, new_n887, new_n889, new_n890, new_n891, new_n892,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  XOR2_X1   g001(.A(KEYINPUT9), .B(G234), .Z(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  OAI21_X1  g003(.A(G221), .B1(new_n189), .B2(G902), .ZN(new_n190));
  XOR2_X1   g004(.A(new_n190), .B(KEYINPUT75), .Z(new_n191));
  AND2_X1   g005(.A1(KEYINPUT3), .A2(G107), .ZN(new_n192));
  NOR2_X1   g006(.A1(KEYINPUT3), .A2(G107), .ZN(new_n193));
  AOI21_X1  g007(.A(new_n192), .B1(G104), .B2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT3), .ZN(new_n195));
  INV_X1    g009(.A(G107), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  AND2_X1   g011(.A1(KEYINPUT76), .A2(G104), .ZN(new_n198));
  NOR2_X1   g012(.A1(KEYINPUT76), .A2(G104), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n197), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G101), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n194), .A2(new_n200), .A3(new_n201), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n196), .B1(new_n198), .B2(new_n199), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n201), .B1(G104), .B2(G107), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n202), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT1), .ZN(new_n207));
  INV_X1    g021(.A(G146), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G143), .ZN(new_n209));
  INV_X1    g023(.A(G143), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G146), .ZN(new_n211));
  AND4_X1   g025(.A1(new_n207), .A2(new_n209), .A3(new_n211), .A4(G128), .ZN(new_n212));
  OAI21_X1  g026(.A(KEYINPUT1), .B1(new_n210), .B2(G146), .ZN(new_n213));
  AOI22_X1  g027(.A1(new_n213), .A2(G128), .B1(new_n209), .B2(new_n211), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n206), .A2(new_n215), .ZN(new_n216));
  OAI211_X1 g030(.A(new_n202), .B(new_n205), .C1(new_n212), .C2(new_n214), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(KEYINPUT65), .A2(G131), .ZN(new_n219));
  INV_X1    g033(.A(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT11), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(KEYINPUT64), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  XNOR2_X1  g037(.A(G134), .B(G137), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT64), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(KEYINPUT11), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n223), .B1(new_n224), .B2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G137), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n222), .B1(G134), .B2(new_n228), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n220), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n228), .A2(G134), .ZN(new_n231));
  INV_X1    g045(.A(G134), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(G137), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n226), .A2(new_n231), .A3(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(new_n222), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n223), .A2(new_n231), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n235), .A2(new_n219), .A3(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n230), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n218), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT12), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n218), .A2(KEYINPUT12), .A3(new_n238), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT4), .ZN(new_n244));
  OR2_X1    g058(.A1(KEYINPUT76), .A2(G104), .ZN(new_n245));
  NAND2_X1  g059(.A1(KEYINPUT76), .A2(G104), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n193), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n195), .A2(new_n196), .A3(G104), .ZN(new_n248));
  NAND2_X1  g062(.A1(KEYINPUT3), .A2(G107), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  OAI211_X1 g064(.A(new_n244), .B(G101), .C1(new_n247), .C2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT77), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n201), .B1(new_n194), .B2(new_n200), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n254), .A2(KEYINPUT77), .A3(new_n244), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n194), .A2(new_n200), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n244), .B1(new_n256), .B2(G101), .ZN(new_n257));
  AOI22_X1  g071(.A1(new_n253), .A2(new_n255), .B1(new_n257), .B2(new_n202), .ZN(new_n258));
  XNOR2_X1  g072(.A(G143), .B(G146), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n259), .A2(KEYINPUT0), .A3(G128), .ZN(new_n260));
  XNOR2_X1  g074(.A(KEYINPUT0), .B(G128), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n260), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n258), .A2(new_n263), .ZN(new_n264));
  XNOR2_X1  g078(.A(new_n217), .B(KEYINPUT10), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n264), .A2(new_n265), .A3(new_n230), .A4(new_n237), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n243), .A2(new_n266), .ZN(new_n267));
  XNOR2_X1  g081(.A(G110), .B(G140), .ZN(new_n268));
  INV_X1    g082(.A(G227), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n269), .A2(G953), .ZN(new_n270));
  XOR2_X1   g084(.A(new_n268), .B(new_n270), .Z(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n267), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n264), .A2(new_n265), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(new_n238), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n275), .A2(new_n266), .A3(new_n271), .ZN(new_n276));
  AND3_X1   g090(.A1(new_n273), .A2(G469), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n243), .A2(KEYINPUT78), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT78), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n241), .A2(new_n279), .A3(new_n242), .ZN(new_n280));
  NAND4_X1  g094(.A1(new_n278), .A2(new_n266), .A3(new_n271), .A4(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n275), .A2(new_n266), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(new_n272), .ZN(new_n283));
  AOI21_X1  g097(.A(G902), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(G469), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n277), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(G469), .A2(G902), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n191), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  OAI21_X1  g102(.A(G210), .B1(G237), .B2(G902), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT6), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT66), .ZN(new_n291));
  INV_X1    g105(.A(G119), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n291), .A2(new_n292), .A3(G116), .ZN(new_n293));
  INV_X1    g107(.A(G116), .ZN(new_n294));
  AOI21_X1  g108(.A(KEYINPUT66), .B1(new_n294), .B2(G119), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n294), .A2(G119), .ZN(new_n296));
  OAI211_X1 g110(.A(KEYINPUT5), .B(new_n293), .C1(new_n295), .C2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(G113), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT5), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n298), .B1(new_n296), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n291), .B1(new_n292), .B2(G116), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n302), .B1(new_n294), .B2(G119), .ZN(new_n303));
  XOR2_X1   g117(.A(KEYINPUT2), .B(G113), .Z(new_n304));
  NAND3_X1  g118(.A1(new_n303), .A2(new_n293), .A3(new_n304), .ZN(new_n305));
  NAND4_X1  g119(.A1(new_n301), .A2(new_n305), .A3(new_n202), .A4(new_n205), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT80), .ZN(new_n307));
  XNOR2_X1  g121(.A(new_n306), .B(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n303), .A2(new_n293), .ZN(new_n309));
  INV_X1    g123(.A(new_n304), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(new_n305), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n256), .A2(G101), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n313), .A2(KEYINPUT4), .A3(new_n202), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n251), .A2(new_n252), .ZN(new_n315));
  AOI21_X1  g129(.A(KEYINPUT77), .B1(new_n254), .B2(new_n244), .ZN(new_n316));
  OAI211_X1 g130(.A(new_n312), .B(new_n314), .C1(new_n315), .C2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT79), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n258), .A2(KEYINPUT79), .A3(new_n312), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n308), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  XOR2_X1   g135(.A(G110), .B(G122), .Z(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n290), .B1(new_n321), .B2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(new_n308), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n317), .A2(new_n318), .ZN(new_n326));
  AOI21_X1  g140(.A(KEYINPUT79), .B1(new_n258), .B2(new_n312), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n325), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(new_n322), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n324), .A2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(G125), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n215), .A2(new_n331), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n332), .B1(new_n263), .B2(new_n331), .ZN(new_n333));
  INV_X1    g147(.A(G224), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n334), .A2(G953), .ZN(new_n335));
  XNOR2_X1  g149(.A(new_n333), .B(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n328), .A2(new_n290), .A3(new_n322), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n330), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(KEYINPUT81), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT81), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n330), .A2(new_n340), .A3(new_n336), .A4(new_n337), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT7), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n333), .B1(new_n343), .B2(new_n335), .ZN(new_n344));
  OR2_X1    g158(.A1(new_n333), .A2(new_n335), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n344), .B1(new_n345), .B2(new_n343), .ZN(new_n346));
  XOR2_X1   g160(.A(new_n322), .B(KEYINPUT8), .Z(new_n347));
  AOI22_X1  g161(.A1(new_n301), .A2(new_n305), .B1(new_n202), .B2(new_n205), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT82), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(new_n306), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n348), .A2(new_n349), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n347), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n346), .B1(new_n353), .B2(KEYINPUT83), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n321), .A2(new_n323), .ZN(new_n355));
  OR2_X1    g169(.A1(new_n353), .A2(KEYINPUT83), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n354), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(G902), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n289), .B1(new_n342), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n289), .ZN(new_n362));
  AOI211_X1 g176(.A(new_n362), .B(new_n359), .C1(new_n339), .C2(new_n341), .ZN(new_n363));
  OAI211_X1 g177(.A(new_n187), .B(new_n288), .C1(new_n361), .C2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT20), .ZN(new_n366));
  INV_X1    g180(.A(G237), .ZN(new_n367));
  INV_X1    g181(.A(G953), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n367), .A2(new_n368), .A3(G143), .A4(G214), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(KEYINPUT85), .ZN(new_n370));
  NOR2_X1   g184(.A1(G237), .A2(G953), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT85), .ZN(new_n372));
  NAND4_X1  g186(.A1(new_n371), .A2(new_n372), .A3(G143), .A4(G214), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n370), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(G131), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n371), .A2(G214), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n376), .A2(KEYINPUT84), .A3(new_n210), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  AOI21_X1  g192(.A(KEYINPUT84), .B1(new_n376), .B2(new_n210), .ZN(new_n379));
  OAI211_X1 g193(.A(new_n374), .B(new_n375), .C1(new_n378), .C2(new_n379), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n374), .B1(new_n378), .B2(new_n379), .ZN(new_n381));
  OAI211_X1 g195(.A(new_n380), .B(KEYINPUT87), .C1(new_n381), .C2(KEYINPUT18), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT84), .ZN(new_n383));
  INV_X1    g197(.A(G214), .ZN(new_n384));
  NOR3_X1   g198(.A1(new_n384), .A2(G237), .A3(G953), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n383), .B1(new_n385), .B2(G143), .ZN(new_n386));
  AOI22_X1  g200(.A1(new_n386), .A2(new_n377), .B1(new_n370), .B2(new_n373), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT87), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT18), .ZN(new_n389));
  OAI211_X1 g203(.A(new_n387), .B(new_n388), .C1(new_n389), .C2(new_n375), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n382), .A2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(G140), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(G125), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n331), .A2(G140), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n395), .A2(G146), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(KEYINPUT86), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT86), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n393), .A2(new_n394), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n396), .B1(new_n400), .B2(G146), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n387), .A2(new_n375), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n401), .B1(new_n402), .B2(KEYINPUT18), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n391), .A2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT88), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n391), .A2(KEYINPUT88), .A3(new_n403), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  XNOR2_X1  g222(.A(G113), .B(G122), .ZN(new_n409));
  XOR2_X1   g223(.A(new_n409), .B(G104), .Z(new_n410));
  INV_X1    g224(.A(KEYINPUT89), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n411), .B1(new_n381), .B2(G131), .ZN(new_n412));
  NOR3_X1   g226(.A1(new_n387), .A2(KEYINPUT89), .A3(new_n375), .ZN(new_n413));
  OAI21_X1  g227(.A(KEYINPUT17), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(KEYINPUT93), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT93), .ZN(new_n416));
  OAI211_X1 g230(.A(new_n416), .B(KEYINPUT17), .C1(new_n412), .C2(new_n413), .ZN(new_n417));
  AND2_X1   g231(.A1(new_n393), .A2(new_n394), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(KEYINPUT16), .ZN(new_n419));
  OR2_X1    g233(.A1(new_n393), .A2(KEYINPUT16), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n419), .A2(G146), .A3(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  AOI21_X1  g236(.A(G146), .B1(new_n419), .B2(new_n420), .ZN(new_n423));
  OR2_X1    g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  AND2_X1   g238(.A1(new_n424), .A2(KEYINPUT92), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n424), .A2(KEYINPUT92), .ZN(new_n426));
  OAI211_X1 g240(.A(new_n415), .B(new_n417), .C1(new_n425), .C2(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n381), .A2(new_n411), .A3(G131), .ZN(new_n428));
  OAI21_X1  g242(.A(KEYINPUT89), .B1(new_n387), .B2(new_n375), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT17), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n428), .A2(new_n429), .A3(new_n430), .A4(new_n380), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n431), .B(KEYINPUT94), .ZN(new_n432));
  OAI211_X1 g246(.A(new_n408), .B(new_n410), .C1(new_n427), .C2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n400), .A2(KEYINPUT19), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT90), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n435), .B1(new_n395), .B2(KEYINPUT19), .ZN(new_n436));
  OR3_X1    g250(.A1(new_n395), .A2(new_n435), .A3(KEYINPUT19), .ZN(new_n437));
  NAND4_X1  g251(.A1(new_n434), .A2(new_n208), .A3(new_n436), .A4(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(new_n421), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(KEYINPUT91), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n428), .A2(new_n429), .A3(new_n380), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT91), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n438), .A2(new_n442), .A3(new_n421), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n440), .A2(new_n441), .A3(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(new_n407), .ZN(new_n445));
  AOI21_X1  g259(.A(KEYINPUT88), .B1(new_n391), .B2(new_n403), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n444), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(new_n410), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n433), .A2(new_n449), .ZN(new_n450));
  NOR2_X1   g264(.A1(G475), .A2(G902), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n366), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(new_n451), .ZN(new_n453));
  AOI211_X1 g267(.A(KEYINPUT20), .B(new_n453), .C1(new_n433), .C2(new_n449), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n408), .B1(new_n427), .B2(new_n432), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(new_n448), .ZN(new_n456));
  AOI21_X1  g270(.A(G902), .B1(new_n456), .B2(new_n433), .ZN(new_n457));
  INV_X1    g271(.A(G475), .ZN(new_n458));
  OAI22_X1  g272(.A1(new_n452), .A2(new_n454), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(G478), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n461), .A2(KEYINPUT15), .ZN(new_n462));
  INV_X1    g276(.A(G217), .ZN(new_n463));
  NOR3_X1   g277(.A1(new_n189), .A2(new_n463), .A3(G953), .ZN(new_n464));
  INV_X1    g278(.A(G128), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(G143), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n210), .A2(G128), .ZN(new_n467));
  AND2_X1   g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(new_n232), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT13), .ZN(new_n470));
  OAI21_X1  g284(.A(KEYINPUT96), .B1(new_n467), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n467), .A2(new_n470), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n471), .A2(new_n466), .A3(new_n472), .ZN(new_n473));
  NOR3_X1   g287(.A1(new_n467), .A2(KEYINPUT96), .A3(new_n470), .ZN(new_n474));
  OAI21_X1  g288(.A(G134), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  XNOR2_X1  g289(.A(new_n468), .B(new_n232), .ZN(new_n476));
  XNOR2_X1  g290(.A(KEYINPUT95), .B(G122), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(G116), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n478), .A2(KEYINPUT14), .A3(G107), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  AOI22_X1  g294(.A1(new_n469), .A2(new_n475), .B1(new_n476), .B2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(G122), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n478), .B1(G116), .B2(new_n482), .ZN(new_n483));
  XNOR2_X1  g297(.A(new_n483), .B(new_n196), .ZN(new_n484));
  OR2_X1    g298(.A1(new_n481), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n484), .A2(new_n476), .A3(new_n479), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n464), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n485), .A2(new_n486), .A3(new_n464), .ZN(new_n489));
  AND2_X1   g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n462), .B1(new_n490), .B2(G902), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n488), .A2(new_n489), .ZN(new_n492));
  INV_X1    g306(.A(new_n462), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n492), .A2(new_n358), .A3(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n491), .A2(KEYINPUT97), .A3(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT97), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n493), .B1(new_n492), .B2(new_n358), .ZN(new_n497));
  AOI211_X1 g311(.A(G902), .B(new_n462), .C1(new_n488), .C2(new_n489), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(G952), .ZN(new_n500));
  AOI211_X1 g314(.A(G953), .B(new_n500), .C1(G234), .C2(G237), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  AOI211_X1 g316(.A(new_n358), .B(new_n368), .C1(G234), .C2(G237), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  XOR2_X1   g318(.A(KEYINPUT21), .B(G898), .Z(new_n505));
  OAI21_X1  g319(.A(new_n502), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  AND3_X1   g320(.A1(new_n495), .A2(new_n499), .A3(new_n506), .ZN(new_n507));
  AND2_X1   g321(.A1(new_n460), .A2(new_n507), .ZN(new_n508));
  NOR2_X1   g322(.A1(G472), .A2(G902), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n367), .A2(new_n368), .A3(G210), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT68), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n510), .B(new_n511), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n512), .B(KEYINPUT67), .ZN(new_n513));
  XOR2_X1   g327(.A(KEYINPUT26), .B(G101), .Z(new_n514));
  XNOR2_X1  g328(.A(new_n514), .B(KEYINPUT27), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n513), .B(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  XNOR2_X1  g331(.A(KEYINPUT70), .B(KEYINPUT28), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  NOR3_X1   g333(.A1(new_n227), .A2(G131), .A3(new_n229), .ZN(new_n520));
  OR2_X1    g334(.A1(new_n224), .A2(new_n375), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n521), .B1(new_n212), .B2(new_n214), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n262), .B1(new_n230), .B2(new_n237), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n312), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NOR3_X1   g339(.A1(new_n227), .A2(new_n220), .A3(new_n229), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n219), .B1(new_n235), .B2(new_n236), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n263), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n312), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n235), .A2(new_n375), .A3(new_n236), .ZN(new_n530));
  OAI211_X1 g344(.A(new_n530), .B(new_n521), .C1(new_n212), .C2(new_n214), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n528), .A2(new_n529), .A3(new_n531), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n519), .B1(new_n525), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n523), .A2(new_n524), .ZN(new_n534));
  AOI21_X1  g348(.A(KEYINPUT28), .B1(new_n534), .B2(new_n529), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n517), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT71), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  OAI211_X1 g352(.A(new_n517), .B(KEYINPUT71), .C1(new_n533), .C2(new_n535), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT30), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n540), .B1(new_n523), .B2(new_n524), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n528), .A2(KEYINPUT30), .A3(new_n531), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n541), .A2(new_n542), .A3(new_n312), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT31), .ZN(new_n544));
  NAND4_X1  g358(.A1(new_n543), .A2(new_n516), .A3(new_n544), .A4(new_n532), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n538), .A2(new_n539), .A3(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n543), .A2(new_n532), .A3(new_n516), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT69), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n543), .A2(new_n516), .A3(KEYINPUT69), .A4(new_n532), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n544), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n509), .B1(new_n546), .B2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT32), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  OAI211_X1 g368(.A(KEYINPUT32), .B(new_n509), .C1(new_n546), .C2(new_n551), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n543), .A2(new_n532), .ZN(new_n556));
  AOI21_X1  g370(.A(KEYINPUT29), .B1(new_n556), .B2(new_n517), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT72), .ZN(new_n558));
  INV_X1    g372(.A(new_n533), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT28), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n532), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n559), .A2(new_n516), .A3(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n557), .A2(new_n558), .A3(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n560), .B1(new_n525), .B2(new_n532), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n564), .A2(new_n535), .ZN(new_n565));
  AND2_X1   g379(.A1(new_n516), .A2(KEYINPUT29), .ZN(new_n566));
  AOI21_X1  g380(.A(G902), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n563), .A2(new_n567), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n558), .B1(new_n557), .B2(new_n562), .ZN(new_n569));
  OAI21_X1  g383(.A(G472), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n554), .A2(new_n555), .A3(new_n570), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n463), .B1(G234), .B2(new_n358), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n292), .A2(G128), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n465), .A2(G119), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n575), .A2(KEYINPUT23), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT23), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n577), .B1(G119), .B2(new_n465), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n574), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n579), .A2(G110), .ZN(new_n580));
  XOR2_X1   g394(.A(KEYINPUT24), .B(G110), .Z(new_n581));
  AOI21_X1  g395(.A(new_n581), .B1(new_n575), .B2(new_n574), .ZN(new_n582));
  OAI221_X1 g396(.A(new_n421), .B1(G146), .B2(new_n395), .C1(new_n580), .C2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n579), .A2(G110), .ZN(new_n584));
  XNOR2_X1  g398(.A(new_n584), .B(KEYINPUT73), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n581), .A2(new_n575), .A3(new_n574), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n586), .B1(new_n422), .B2(new_n423), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n583), .B1(new_n585), .B2(new_n587), .ZN(new_n588));
  XNOR2_X1  g402(.A(KEYINPUT22), .B(G137), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n368), .A2(G221), .A3(G234), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n589), .B(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n588), .A2(new_n592), .ZN(new_n593));
  OAI211_X1 g407(.A(new_n583), .B(new_n591), .C1(new_n585), .C2(new_n587), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n593), .A2(new_n358), .A3(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT25), .ZN(new_n596));
  OR2_X1    g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n595), .A2(new_n596), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n573), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n573), .A2(new_n358), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n601), .B(KEYINPUT74), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n593), .A2(new_n602), .A3(new_n594), .ZN(new_n603));
  AND2_X1   g417(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n571), .A2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n365), .A2(new_n508), .A3(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(G101), .ZN(G3));
  OR2_X1    g422(.A1(new_n546), .A2(new_n551), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n358), .B1(new_n546), .B2(new_n551), .ZN(new_n610));
  AOI22_X1  g424(.A1(new_n609), .A2(new_n509), .B1(new_n610), .B2(G472), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n611), .A2(new_n288), .A3(new_n604), .ZN(new_n612));
  XOR2_X1   g426(.A(new_n612), .B(KEYINPUT98), .Z(new_n613));
  INV_X1    g427(.A(new_n187), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n342), .A2(new_n360), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(new_n362), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n342), .A2(new_n289), .A3(new_n360), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n614), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  AOI21_X1  g432(.A(KEYINPUT99), .B1(new_n485), .B2(new_n486), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT33), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n492), .B(new_n621), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n461), .A2(G902), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n461), .B1(new_n490), .B2(G902), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n459), .A2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n618), .A2(new_n506), .A3(new_n628), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n613), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(KEYINPUT34), .B(G104), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G6));
  INV_X1    g446(.A(KEYINPUT101), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n453), .B1(new_n433), .B2(new_n449), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(new_n366), .ZN(new_n635));
  OR2_X1    g449(.A1(new_n457), .A2(new_n458), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n495), .A2(new_n499), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n635), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  XOR2_X1   g452(.A(new_n506), .B(KEYINPUT100), .Z(new_n639));
  OAI21_X1  g453(.A(new_n633), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n639), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n460), .A2(KEYINPUT101), .A3(new_n637), .A4(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n640), .A2(new_n642), .A3(new_n618), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n613), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(KEYINPUT35), .B(G107), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G9));
  INV_X1    g460(.A(KEYINPUT102), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n592), .A2(KEYINPUT36), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n588), .B(new_n648), .ZN(new_n649));
  AND2_X1   g463(.A1(new_n649), .A2(new_n602), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n599), .A2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n611), .A2(new_n647), .A3(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n611), .ZN(new_n654));
  OAI21_X1  g468(.A(KEYINPUT102), .B1(new_n654), .B2(new_n651), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n365), .A2(new_n508), .A3(new_n653), .A4(new_n655), .ZN(new_n656));
  XOR2_X1   g470(.A(KEYINPUT37), .B(G110), .Z(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(G12));
  OAI21_X1  g472(.A(new_n502), .B1(new_n504), .B2(G900), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n635), .A2(new_n636), .A3(new_n637), .A4(new_n659), .ZN(new_n660));
  AND3_X1   g474(.A1(new_n554), .A2(new_n555), .A3(new_n570), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n365), .A2(new_n652), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G128), .ZN(G30));
  NOR2_X1   g478(.A1(new_n361), .A2(new_n363), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(KEYINPUT38), .ZN(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n516), .B1(new_n532), .B2(new_n525), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n668), .B1(new_n549), .B2(new_n550), .ZN(new_n669));
  OAI21_X1  g483(.A(G472), .B1(new_n669), .B2(G902), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n670), .A2(new_n554), .A3(new_n555), .ZN(new_n671));
  AND3_X1   g485(.A1(new_n671), .A2(new_n187), .A3(new_n651), .ZN(new_n672));
  AND2_X1   g486(.A1(new_n495), .A2(new_n499), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n460), .A2(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(new_n288), .ZN(new_n675));
  XOR2_X1   g489(.A(new_n659), .B(KEYINPUT39), .Z(new_n676));
  NOR2_X1   g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(KEYINPUT40), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n667), .A2(new_n672), .A3(new_n674), .A4(new_n678), .ZN(new_n679));
  XOR2_X1   g493(.A(KEYINPUT103), .B(G143), .Z(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(G45));
  NAND3_X1  g495(.A1(new_n459), .A2(new_n626), .A3(new_n659), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n682), .A2(new_n661), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n683), .A2(new_n618), .A3(new_n288), .A4(new_n652), .ZN(new_n684));
  XNOR2_X1  g498(.A(KEYINPUT104), .B(G146), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(G48));
  NAND2_X1  g500(.A1(new_n281), .A2(new_n283), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(new_n358), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(G469), .ZN(new_n689));
  INV_X1    g503(.A(new_n191), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n284), .A2(new_n285), .ZN(new_n691));
  AND3_X1   g505(.A1(new_n689), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n605), .A2(new_n693), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n694), .A2(new_n618), .A3(new_n506), .A4(new_n628), .ZN(new_n695));
  XNOR2_X1  g509(.A(KEYINPUT41), .B(G113), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n695), .B(new_n696), .ZN(G15));
  NAND4_X1  g511(.A1(new_n640), .A2(new_n694), .A3(new_n618), .A4(new_n642), .ZN(new_n698));
  XOR2_X1   g512(.A(KEYINPUT105), .B(G116), .Z(new_n699));
  XNOR2_X1  g513(.A(new_n698), .B(new_n699), .ZN(G18));
  OAI211_X1 g514(.A(new_n187), .B(new_n692), .C1(new_n361), .C2(new_n363), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  AND4_X1   g516(.A1(new_n460), .A2(new_n507), .A3(new_n571), .A4(new_n652), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G119), .ZN(G21));
  OAI211_X1 g519(.A(new_n187), .B(new_n641), .C1(new_n361), .C2(new_n363), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n549), .A2(new_n550), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(KEYINPUT31), .ZN(new_n709));
  NOR3_X1   g523(.A1(new_n523), .A2(new_n524), .A3(new_n312), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n529), .B1(new_n528), .B2(new_n531), .ZN(new_n711));
  OAI21_X1  g525(.A(KEYINPUT28), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT106), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n712), .A2(new_n713), .A3(new_n561), .ZN(new_n714));
  OAI21_X1  g528(.A(KEYINPUT106), .B1(new_n564), .B2(new_n535), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n714), .A2(new_n715), .A3(new_n517), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n709), .A2(KEYINPUT107), .A3(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT107), .ZN(new_n718));
  AND3_X1   g532(.A1(new_n714), .A2(new_n715), .A3(new_n517), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n718), .B1(new_n551), .B2(new_n719), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n717), .A2(new_n720), .A3(new_n545), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(new_n509), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n610), .A2(G472), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n722), .A2(new_n604), .A3(new_n723), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n692), .A2(new_n459), .A3(new_n637), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n707), .A2(new_n726), .ZN(new_n727));
  XOR2_X1   g541(.A(KEYINPUT108), .B(G122), .Z(new_n728));
  XNOR2_X1  g542(.A(new_n727), .B(new_n728), .ZN(G24));
  AND3_X1   g543(.A1(new_n722), .A2(new_n723), .A3(new_n652), .ZN(new_n730));
  INV_X1    g544(.A(new_n682), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n618), .A2(new_n730), .A3(new_n731), .A4(new_n692), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G125), .ZN(G27));
  NOR3_X1   g547(.A1(new_n361), .A2(new_n363), .A3(new_n614), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n287), .B(KEYINPUT109), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n191), .B1(new_n286), .B2(new_n735), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n734), .A2(new_n731), .A3(new_n606), .A4(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT42), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  AND4_X1   g553(.A1(new_n187), .A2(new_n616), .A3(new_n617), .A4(new_n736), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n740), .A2(KEYINPUT42), .A3(new_n606), .A4(new_n731), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G131), .ZN(G33));
  NAND3_X1  g557(.A1(new_n665), .A2(new_n187), .A3(new_n736), .ZN(new_n744));
  NOR3_X1   g558(.A1(new_n744), .A2(new_n605), .A3(new_n660), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(new_n232), .ZN(G36));
  NAND2_X1  g560(.A1(new_n460), .A2(new_n626), .ZN(new_n747));
  XOR2_X1   g561(.A(new_n747), .B(KEYINPUT43), .Z(new_n748));
  OR2_X1    g562(.A1(new_n748), .A2(KEYINPUT110), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(KEYINPUT110), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n749), .A2(new_n654), .A3(new_n652), .A4(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT44), .ZN(new_n752));
  OR2_X1    g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n751), .A2(new_n752), .ZN(new_n754));
  AOI21_X1  g568(.A(KEYINPUT45), .B1(new_n273), .B2(new_n276), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n755), .A2(new_n285), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n273), .A2(KEYINPUT45), .A3(new_n276), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  AND2_X1   g572(.A1(new_n758), .A2(new_n735), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(KEYINPUT46), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(new_n691), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n759), .A2(KEYINPUT46), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n690), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  OR2_X1    g577(.A1(new_n763), .A2(new_n676), .ZN(new_n764));
  INV_X1    g578(.A(new_n764), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n753), .A2(new_n734), .A3(new_n754), .A4(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G137), .ZN(G39));
  XNOR2_X1  g581(.A(new_n763), .B(KEYINPUT47), .ZN(new_n768));
  INV_X1    g582(.A(new_n604), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n734), .A2(new_n769), .A3(new_n661), .A4(new_n731), .ZN(new_n770));
  OR2_X1    g584(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G140), .ZN(G42));
  INV_X1    g586(.A(KEYINPUT51), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n724), .A2(new_n502), .ZN(new_n774));
  AND2_X1   g588(.A1(new_n748), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(new_n734), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT112), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n775), .A2(KEYINPUT112), .A3(new_n734), .ZN(new_n779));
  AND2_X1   g593(.A1(new_n689), .A2(new_n691), .ZN(new_n780));
  INV_X1    g594(.A(new_n780), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n768), .B1(new_n690), .B2(new_n781), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n778), .A2(new_n779), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n783), .A2(KEYINPUT113), .ZN(new_n784));
  AND3_X1   g598(.A1(new_n734), .A2(new_n501), .A3(new_n692), .ZN(new_n785));
  AND2_X1   g599(.A1(new_n748), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(new_n730), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n769), .A2(new_n671), .ZN(new_n788));
  AND2_X1   g602(.A1(new_n785), .A2(new_n788), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n789), .A2(new_n460), .A3(new_n625), .A4(new_n624), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n787), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n692), .A2(new_n614), .ZN(new_n792));
  XOR2_X1   g606(.A(new_n792), .B(KEYINPUT114), .Z(new_n793));
  NOR2_X1   g607(.A1(new_n667), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n775), .A2(KEYINPUT50), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n775), .A2(new_n794), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT50), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n791), .B1(new_n795), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n784), .A2(new_n799), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n783), .A2(KEYINPUT113), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n773), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(KEYINPUT115), .ZN(new_n803));
  INV_X1    g617(.A(new_n799), .ZN(new_n804));
  OR2_X1    g618(.A1(new_n804), .A2(KEYINPUT116), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(KEYINPUT116), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n805), .A2(KEYINPUT51), .A3(new_n783), .A4(new_n806), .ZN(new_n807));
  OAI211_X1 g621(.A(new_n635), .B(new_n636), .C1(new_n498), .C2(new_n497), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n612), .B1(new_n627), .B2(new_n808), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n707), .B1(new_n809), .B2(new_n726), .ZN(new_n810));
  AND3_X1   g624(.A1(new_n810), .A2(new_n656), .A3(new_n698), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n745), .B1(new_n739), .B2(new_n741), .ZN(new_n812));
  AND3_X1   g626(.A1(new_n607), .A2(new_n695), .A3(new_n704), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n652), .A2(new_n494), .A3(new_n491), .A4(new_n659), .ZN(new_n814));
  NOR4_X1   g628(.A1(new_n814), .A2(new_n661), .A3(new_n675), .A4(new_n459), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n722), .A2(new_n723), .A3(new_n652), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n816), .A2(new_n682), .ZN(new_n817));
  AOI22_X1  g631(.A1(new_n815), .A2(new_n734), .B1(new_n740), .B2(new_n817), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n811), .A2(new_n812), .A3(new_n813), .A4(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(new_n819), .ZN(new_n820));
  AND3_X1   g634(.A1(new_n736), .A2(new_n651), .A3(new_n659), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n618), .A2(new_n671), .A3(new_n674), .A4(new_n821), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n663), .A2(new_n684), .A3(new_n732), .A4(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n823), .A2(KEYINPUT52), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n364), .A2(new_n651), .ZN(new_n825));
  AOI22_X1  g639(.A1(new_n825), .A2(new_n662), .B1(new_n702), .B2(new_n817), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT52), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n826), .A2(new_n827), .A3(new_n684), .A4(new_n822), .ZN(new_n828));
  AND2_X1   g642(.A1(new_n824), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n820), .A2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT111), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n824), .A2(new_n828), .A3(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n831), .B1(new_n824), .B2(new_n828), .ZN(new_n834));
  NOR3_X1   g648(.A1(new_n833), .A2(new_n834), .A3(new_n819), .ZN(new_n835));
  MUX2_X1   g649(.A(new_n830), .B(new_n835), .S(KEYINPUT53), .Z(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(KEYINPUT54), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT54), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n820), .A2(KEYINPUT53), .A3(new_n829), .ZN(new_n839));
  OAI211_X1 g653(.A(new_n838), .B(new_n839), .C1(new_n835), .C2(KEYINPUT53), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n837), .A2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n775), .A2(new_n702), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n843), .A2(G952), .A3(new_n368), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT48), .ZN(new_n845));
  OAI211_X1 g659(.A(new_n786), .B(new_n606), .C1(KEYINPUT117), .C2(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(KEYINPUT117), .ZN(new_n847));
  XOR2_X1   g661(.A(new_n846), .B(new_n847), .Z(new_n848));
  AOI211_X1 g662(.A(new_n844), .B(new_n848), .C1(new_n628), .C2(new_n789), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n803), .A2(new_n807), .A3(new_n842), .A4(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n500), .A2(new_n368), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  XNOR2_X1  g666(.A(new_n780), .B(KEYINPUT49), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n853), .A2(new_n187), .A3(new_n690), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n854), .A2(new_n747), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n855), .A2(new_n666), .A3(new_n788), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n852), .A2(new_n856), .ZN(G75));
  NOR2_X1   g671(.A1(new_n834), .A2(new_n819), .ZN(new_n858));
  AOI21_X1  g672(.A(KEYINPUT53), .B1(new_n858), .B2(new_n832), .ZN(new_n859));
  AND3_X1   g673(.A1(new_n820), .A2(KEYINPUT53), .A3(new_n829), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n861), .A2(new_n358), .ZN(new_n862));
  AOI21_X1  g676(.A(KEYINPUT56), .B1(new_n862), .B2(G210), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n330), .A2(new_n337), .ZN(new_n864));
  XNOR2_X1  g678(.A(new_n864), .B(new_n336), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n865), .B(KEYINPUT55), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n863), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n863), .A2(new_n866), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n368), .A2(G952), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(G51));
  NOR3_X1   g684(.A1(new_n861), .A2(new_n358), .A3(new_n758), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT119), .ZN(new_n872));
  OAI21_X1  g686(.A(KEYINPUT54), .B1(new_n859), .B2(new_n860), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n873), .A2(new_n840), .ZN(new_n874));
  XNOR2_X1  g688(.A(KEYINPUT118), .B(KEYINPUT57), .ZN(new_n875));
  XOR2_X1   g689(.A(new_n735), .B(new_n875), .Z(new_n876));
  AOI21_X1  g690(.A(new_n872), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(new_n876), .ZN(new_n878));
  AOI211_X1 g692(.A(KEYINPUT119), .B(new_n878), .C1(new_n873), .C2(new_n840), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n687), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n871), .B1(new_n880), .B2(KEYINPUT120), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT120), .ZN(new_n882));
  OAI211_X1 g696(.A(new_n882), .B(new_n687), .C1(new_n877), .C2(new_n879), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n869), .B1(new_n881), .B2(new_n883), .ZN(G54));
  AND3_X1   g698(.A1(new_n862), .A2(KEYINPUT58), .A3(G475), .ZN(new_n885));
  AND2_X1   g699(.A1(new_n885), .A2(new_n450), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n885), .A2(new_n450), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n886), .A2(new_n887), .A3(new_n869), .ZN(G60));
  NAND2_X1  g702(.A1(G478), .A2(G902), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n889), .B(KEYINPUT59), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n622), .B1(new_n841), .B2(new_n890), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n874), .A2(new_n622), .A3(new_n890), .ZN(new_n892));
  NOR3_X1   g706(.A1(new_n891), .A2(new_n869), .A3(new_n892), .ZN(G63));
  NAND2_X1  g707(.A1(G217), .A2(G902), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n894), .B(KEYINPUT60), .ZN(new_n895));
  OR2_X1    g709(.A1(new_n861), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n593), .A2(new_n594), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n869), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  AOI21_X1  g712(.A(KEYINPUT61), .B1(new_n898), .B2(KEYINPUT121), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n861), .A2(new_n895), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(new_n649), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n899), .B(new_n902), .ZN(G66));
  INV_X1    g717(.A(new_n505), .ZN(new_n904));
  OAI21_X1  g718(.A(G953), .B1(new_n904), .B2(new_n334), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n811), .A2(new_n813), .ZN(new_n906));
  XOR2_X1   g720(.A(new_n906), .B(KEYINPUT122), .Z(new_n907));
  OAI21_X1  g721(.A(new_n905), .B1(new_n907), .B2(G953), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n864), .B1(G898), .B2(new_n368), .ZN(new_n909));
  XOR2_X1   g723(.A(new_n909), .B(KEYINPUT123), .Z(new_n910));
  XNOR2_X1  g724(.A(new_n908), .B(new_n910), .ZN(G69));
  NAND2_X1  g725(.A1(new_n541), .A2(new_n542), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n434), .A2(new_n436), .A3(new_n437), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(KEYINPUT124), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n912), .B(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(new_n269), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n368), .B1(new_n916), .B2(G900), .ZN(new_n917));
  INV_X1    g731(.A(new_n812), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n918), .A2(KEYINPUT127), .ZN(new_n919));
  OR2_X1    g733(.A1(new_n918), .A2(KEYINPUT127), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n766), .A2(new_n771), .A3(new_n919), .A4(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n826), .A2(new_n684), .ZN(new_n922));
  XOR2_X1   g736(.A(new_n922), .B(KEYINPUT125), .Z(new_n923));
  NAND4_X1  g737(.A1(new_n765), .A2(new_n618), .A3(new_n606), .A4(new_n674), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n368), .B1(new_n921), .B2(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n915), .B1(new_n269), .B2(G953), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n917), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n923), .A2(new_n679), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(KEYINPUT62), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n808), .A2(new_n627), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n931), .B(KEYINPUT126), .Z(new_n932));
  NAND4_X1  g746(.A1(new_n932), .A2(new_n606), .A3(new_n677), .A4(new_n734), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n766), .A2(new_n771), .A3(new_n933), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n930), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n915), .A2(new_n368), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n928), .B1(new_n935), .B2(new_n936), .ZN(G72));
  NAND2_X1  g751(.A1(new_n556), .A2(new_n517), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(new_n547), .ZN(new_n939));
  INV_X1    g753(.A(new_n556), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n940), .B1(new_n921), .B2(new_n925), .ZN(new_n941));
  OAI211_X1 g755(.A(new_n941), .B(new_n907), .C1(new_n935), .C2(new_n940), .ZN(new_n942));
  NAND2_X1  g756(.A1(G472), .A2(G902), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n943), .B(KEYINPUT63), .Z(new_n944));
  AOI21_X1  g758(.A(new_n939), .B1(new_n942), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n708), .A2(new_n938), .ZN(new_n946));
  AND3_X1   g760(.A1(new_n836), .A2(new_n944), .A3(new_n946), .ZN(new_n947));
  NOR3_X1   g761(.A1(new_n945), .A2(new_n869), .A3(new_n947), .ZN(G57));
endmodule


