

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764;

  XNOR2_X1 U369 ( .A(n375), .B(KEYINPUT108), .ZN(n649) );
  AND2_X1 U370 ( .A1(n403), .A2(n558), .ZN(n652) );
  OR2_X1 U371 ( .A1(n642), .A2(n629), .ZN(n541) );
  XOR2_X1 U372 ( .A(G146), .B(G125), .Z(n523) );
  XNOR2_X1 U373 ( .A(G113), .B(G143), .ZN(n455) );
  XNOR2_X2 U374 ( .A(n563), .B(KEYINPUT6), .ZN(n588) );
  XOR2_X2 U375 ( .A(n723), .B(KEYINPUT59), .Z(n724) );
  OR2_X1 U376 ( .A1(n616), .A2(n596), .ZN(n382) );
  XNOR2_X2 U377 ( .A(n402), .B(KEYINPUT0), .ZN(n616) );
  XNOR2_X2 U378 ( .A(n475), .B(n474), .ZN(n618) );
  XNOR2_X1 U379 ( .A(G119), .B(G110), .ZN(n482) );
  AND2_X2 U380 ( .A1(n676), .A2(n631), .ZN(n445) );
  XNOR2_X2 U381 ( .A(n423), .B(n586), .ZN(n613) );
  NAND2_X1 U382 ( .A1(n740), .A2(n446), .ZN(n676) );
  NOR2_X1 U383 ( .A1(n572), .A2(n404), .ZN(n430) );
  AND2_X1 U384 ( .A1(n411), .A2(n394), .ZN(n393) );
  NAND2_X1 U385 ( .A1(n381), .A2(n378), .ZN(n598) );
  AND2_X1 U386 ( .A1(n363), .A2(n760), .ZN(n394) );
  NAND2_X1 U387 ( .A1(n380), .A2(n379), .ZN(n378) );
  XNOR2_X1 U388 ( .A(n430), .B(n429), .ZN(n761) );
  AND2_X1 U389 ( .A1(n361), .A2(n351), .ZN(n363) );
  AND2_X1 U390 ( .A1(n383), .A2(n354), .ZN(n381) );
  XNOR2_X1 U391 ( .A(n431), .B(KEYINPUT42), .ZN(n764) );
  AND2_X1 U392 ( .A1(n561), .A2(n544), .ZN(n662) );
  NOR2_X1 U393 ( .A1(n595), .A2(n594), .ZN(n402) );
  OR2_X1 U394 ( .A1(n403), .A2(n558), .ZN(n473) );
  XNOR2_X1 U395 ( .A(n642), .B(n641), .ZN(n643) );
  XNOR2_X1 U396 ( .A(n433), .B(n748), .ZN(n365) );
  OR2_X1 U397 ( .A1(n634), .A2(G902), .ZN(n514) );
  XNOR2_X1 U398 ( .A(n523), .B(n450), .ZN(n483) );
  XNOR2_X1 U399 ( .A(n386), .B(KEYINPUT87), .ZN(n531) );
  AND2_X1 U400 ( .A1(n447), .A2(n445), .ZN(n349) );
  AND2_X2 U401 ( .A1(n445), .A2(n447), .ZN(n732) );
  NAND2_X1 U402 ( .A1(n444), .A2(n627), .ZN(n447) );
  NOR2_X1 U403 ( .A1(n759), .A2(KEYINPUT44), .ZN(n599) );
  XNOR2_X2 U404 ( .A(n397), .B(n424), .ZN(n719) );
  NAND2_X1 U405 ( .A1(n581), .A2(n373), .ZN(n565) );
  AND2_X1 U406 ( .A1(n548), .A2(n427), .ZN(n554) );
  NOR2_X1 U407 ( .A1(n368), .A2(n367), .ZN(n548) );
  INV_X1 U408 ( .A(n547), .ZN(n427) );
  XNOR2_X1 U409 ( .A(n490), .B(n489), .ZN(n546) );
  NOR2_X1 U410 ( .A1(n365), .A2(G902), .ZN(n490) );
  INV_X1 U411 ( .A(KEYINPUT88), .ZN(n502) );
  INV_X1 U412 ( .A(G110), .ZN(n386) );
  NAND2_X1 U413 ( .A1(n362), .A2(n422), .ZN(n620) );
  NAND2_X1 U414 ( .A1(n404), .A2(n571), .ZN(n475) );
  AND2_X1 U415 ( .A1(n662), .A2(n414), .ZN(n413) );
  XNOR2_X1 U416 ( .A(n360), .B(n562), .ZN(n415) );
  NAND2_X1 U417 ( .A1(n373), .A2(n374), .ZN(n372) );
  AND2_X1 U418 ( .A1(n437), .A2(KEYINPUT100), .ZN(n436) );
  INV_X1 U419 ( .A(n622), .ZN(n438) );
  NOR2_X1 U420 ( .A1(n647), .A2(n658), .ZN(n611) );
  NOR2_X1 U421 ( .A1(G953), .A2(G237), .ZN(n505) );
  INV_X1 U422 ( .A(G134), .ZN(n499) );
  XNOR2_X1 U423 ( .A(G137), .B(G140), .ZN(n516) );
  NAND2_X1 U424 ( .A1(n665), .A2(n417), .ZN(n575) );
  XNOR2_X1 U425 ( .A(n419), .B(n418), .ZN(n417) );
  INV_X1 U426 ( .A(KEYINPUT102), .ZN(n418) );
  XNOR2_X1 U427 ( .A(KEYINPUT71), .B(KEYINPUT34), .ZN(n596) );
  XNOR2_X1 U428 ( .A(n483), .B(n516), .ZN(n748) );
  XNOR2_X1 U429 ( .A(n480), .B(n482), .ZN(n435) );
  XOR2_X1 U430 ( .A(KEYINPUT24), .B(KEYINPUT90), .Z(n480) );
  XNOR2_X1 U431 ( .A(G128), .B(KEYINPUT80), .ZN(n479) );
  XNOR2_X1 U432 ( .A(n465), .B(n464), .ZN(n392) );
  XOR2_X1 U433 ( .A(KEYINPUT8), .B(KEYINPUT67), .Z(n464) );
  XNOR2_X1 U434 ( .A(n463), .B(n462), .ZN(n465) );
  INV_X1 U435 ( .A(KEYINPUT68), .ZN(n462) );
  XNOR2_X1 U436 ( .A(G140), .B(G131), .ZN(n407) );
  XNOR2_X1 U437 ( .A(n409), .B(n454), .ZN(n408) );
  XOR2_X1 U438 ( .A(KEYINPUT94), .B(KEYINPUT11), .Z(n454) );
  XNOR2_X1 U439 ( .A(n455), .B(n452), .ZN(n409) );
  INV_X1 U440 ( .A(KEYINPUT12), .ZN(n452) );
  XNOR2_X1 U441 ( .A(n516), .B(n517), .ZN(n448) );
  INV_X1 U442 ( .A(G104), .ZN(n517) );
  XNOR2_X1 U443 ( .A(n560), .B(n432), .ZN(n703) );
  INV_X1 U444 ( .A(KEYINPUT41), .ZN(n432) );
  NOR2_X1 U445 ( .A1(n682), .A2(n683), .ZN(n560) );
  XNOR2_X1 U446 ( .A(n556), .B(n555), .ZN(n572) );
  XNOR2_X1 U447 ( .A(n565), .B(n543), .ZN(n595) );
  AND2_X1 U448 ( .A1(n395), .A2(n521), .ZN(n561) );
  XNOR2_X1 U449 ( .A(n396), .B(KEYINPUT28), .ZN(n395) );
  NOR2_X1 U450 ( .A1(n564), .A2(n696), .ZN(n396) );
  XNOR2_X1 U451 ( .A(n604), .B(n603), .ZN(n610) );
  BUF_X1 U452 ( .A(n546), .Z(n366) );
  XNOR2_X1 U453 ( .A(n535), .B(n534), .ZN(n737) );
  INV_X1 U454 ( .A(KEYINPUT75), .ZN(n414) );
  AND2_X1 U455 ( .A1(n618), .A2(n476), .ZN(n477) );
  INV_X1 U456 ( .A(KEYINPUT83), .ZN(n391) );
  AND2_X1 U457 ( .A1(n449), .A2(n370), .ZN(n369) );
  OR2_X1 U458 ( .A1(n563), .A2(n372), .ZN(n371) );
  NAND2_X1 U459 ( .A1(KEYINPUT30), .A2(n559), .ZN(n370) );
  XNOR2_X1 U460 ( .A(G116), .B(G137), .ZN(n506) );
  NAND2_X1 U461 ( .A1(n436), .A2(n438), .ZN(n387) );
  AND2_X1 U462 ( .A1(n443), .A2(n353), .ZN(n440) );
  INV_X1 U463 ( .A(G237), .ZN(n538) );
  OR2_X1 U464 ( .A1(n546), .A2(n497), .ZN(n564) );
  XNOR2_X1 U465 ( .A(KEYINPUT74), .B(KEYINPUT16), .ZN(n530) );
  NAND2_X1 U466 ( .A1(G237), .A2(G234), .ZN(n495) );
  XOR2_X1 U467 ( .A(KEYINPUT98), .B(n652), .Z(n571) );
  AND2_X1 U468 ( .A1(n692), .A2(n366), .ZN(n621) );
  XNOR2_X1 U469 ( .A(n620), .B(KEYINPUT85), .ZN(n443) );
  XNOR2_X1 U470 ( .A(n634), .B(n633), .ZN(n635) );
  XNOR2_X1 U471 ( .A(n484), .B(n434), .ZN(n433) );
  XNOR2_X1 U472 ( .A(n435), .B(n481), .ZN(n434) );
  XNOR2_X1 U473 ( .A(n405), .B(n456), .ZN(n723) );
  XNOR2_X1 U474 ( .A(n408), .B(n406), .ZN(n405) );
  XNOR2_X1 U475 ( .A(n453), .B(n407), .ZN(n406) );
  XNOR2_X1 U476 ( .A(n426), .B(n425), .ZN(n424) );
  XNOR2_X1 U477 ( .A(n515), .B(n518), .ZN(n425) );
  XNOR2_X1 U478 ( .A(n737), .B(n536), .ZN(n642) );
  AND2_X1 U479 ( .A1(n637), .A2(G953), .ZN(n736) );
  NAND2_X1 U480 ( .A1(n703), .A2(n561), .ZN(n431) );
  INV_X1 U481 ( .A(KEYINPUT40), .ZN(n429) );
  INV_X1 U482 ( .A(KEYINPUT36), .ZN(n389) );
  NOR2_X1 U483 ( .A1(n620), .A2(n606), .ZN(n607) );
  INV_X1 U484 ( .A(n366), .ZN(n605) );
  XNOR2_X1 U485 ( .A(n364), .B(KEYINPUT105), .ZN(n760) );
  AND2_X1 U486 ( .A1(n551), .A2(n597), .ZN(n364) );
  NOR2_X1 U487 ( .A1(n428), .A2(n366), .ZN(n608) );
  OR2_X1 U488 ( .A1(n547), .A2(n428), .ZN(n350) );
  INV_X1 U489 ( .A(n692), .ZN(n388) );
  OR2_X1 U490 ( .A1(n662), .A2(n414), .ZN(n351) );
  BUF_X1 U491 ( .A(n563), .Z(n696) );
  AND2_X1 U492 ( .A1(n399), .A2(n398), .ZN(n352) );
  INV_X1 U493 ( .A(KEYINPUT30), .ZN(n374) );
  AND2_X1 U494 ( .A1(n621), .A2(n442), .ZN(n353) );
  AND2_X1 U495 ( .A1(n382), .A2(n597), .ZN(n354) );
  NOR2_X1 U496 ( .A1(n366), .A2(n695), .ZN(n355) );
  INV_X1 U497 ( .A(n588), .ZN(n422) );
  INV_X1 U498 ( .A(KEYINPUT101), .ZN(n587) );
  XNOR2_X1 U499 ( .A(KEYINPUT64), .B(KEYINPUT45), .ZN(n356) );
  NAND2_X1 U500 ( .A1(n357), .A2(n352), .ZN(n359) );
  XNOR2_X1 U501 ( .A(n400), .B(KEYINPUT70), .ZN(n357) );
  NAND2_X1 U502 ( .A1(n358), .A2(n390), .ZN(n570) );
  NOR2_X1 U503 ( .A1(n412), .A2(n415), .ZN(n358) );
  XNOR2_X2 U504 ( .A(n359), .B(n356), .ZN(n740) );
  NAND2_X1 U505 ( .A1(n764), .A2(n761), .ZN(n360) );
  XNOR2_X1 U506 ( .A(n649), .B(n391), .ZN(n390) );
  NAND2_X1 U507 ( .A1(n420), .A2(n588), .ZN(n419) );
  NAND2_X1 U508 ( .A1(n552), .A2(KEYINPUT47), .ZN(n361) );
  NAND2_X1 U509 ( .A1(n401), .A2(KEYINPUT44), .ZN(n398) );
  INV_X1 U510 ( .A(n610), .ZN(n362) );
  XNOR2_X1 U511 ( .A(n365), .B(KEYINPUT124), .ZN(n733) );
  AND2_X1 U512 ( .A1(n563), .A2(KEYINPUT30), .ZN(n367) );
  NAND2_X1 U513 ( .A1(n371), .A2(n369), .ZN(n368) );
  INV_X1 U514 ( .A(n559), .ZN(n373) );
  XNOR2_X2 U515 ( .A(n514), .B(n513), .ZN(n563) );
  NAND2_X1 U516 ( .A1(n376), .A2(n388), .ZN(n375) );
  XNOR2_X1 U517 ( .A(n377), .B(n389), .ZN(n376) );
  NAND2_X1 U518 ( .A1(n567), .A2(n566), .ZN(n377) );
  INV_X1 U519 ( .A(n596), .ZN(n379) );
  INV_X1 U520 ( .A(n688), .ZN(n380) );
  NAND2_X1 U521 ( .A1(n688), .A2(n384), .ZN(n383) );
  AND2_X1 U522 ( .A1(n616), .A2(n596), .ZN(n384) );
  XNOR2_X2 U523 ( .A(n589), .B(KEYINPUT33), .ZN(n688) );
  NAND2_X1 U524 ( .A1(n554), .A2(n581), .ZN(n550) );
  NAND2_X1 U525 ( .A1(n385), .A2(n611), .ZN(n400) );
  XNOR2_X1 U526 ( .A(n599), .B(KEYINPUT66), .ZN(n385) );
  NAND2_X1 U527 ( .A1(n443), .A2(n621), .ZN(n437) );
  NAND2_X1 U528 ( .A1(n439), .A2(n387), .ZN(n399) );
  NAND2_X1 U529 ( .A1(n392), .A2(G221), .ZN(n484) );
  NAND2_X1 U530 ( .A1(n392), .A2(G217), .ZN(n468) );
  NAND2_X1 U531 ( .A1(n393), .A2(n410), .ZN(n412) );
  XNOR2_X2 U532 ( .A(n749), .B(G146), .ZN(n397) );
  XNOR2_X1 U533 ( .A(n397), .B(n511), .ZN(n634) );
  NAND2_X1 U534 ( .A1(n611), .A2(n612), .ZN(n401) );
  NAND2_X1 U535 ( .A1(n616), .A2(n601), .ZN(n604) );
  XNOR2_X1 U536 ( .A(n557), .B(KEYINPUT95), .ZN(n403) );
  INV_X1 U537 ( .A(n665), .ZN(n404) );
  OR2_X1 U538 ( .A1(n545), .A2(n414), .ZN(n410) );
  NAND2_X1 U539 ( .A1(n545), .A2(n413), .ZN(n411) );
  XNOR2_X2 U540 ( .A(n526), .B(n500), .ZN(n749) );
  XNOR2_X2 U541 ( .A(n498), .B(KEYINPUT4), .ZN(n526) );
  XNOR2_X1 U542 ( .A(n673), .B(n416), .ZN(n623) );
  INV_X1 U543 ( .A(KEYINPUT79), .ZN(n416) );
  XNOR2_X2 U544 ( .A(n632), .B(KEYINPUT81), .ZN(n673) );
  NAND2_X2 U545 ( .A1(n584), .A2(n583), .ZN(n632) );
  INV_X1 U546 ( .A(n564), .ZN(n420) );
  NAND2_X1 U547 ( .A1(n421), .A2(n588), .ZN(n589) );
  XNOR2_X1 U548 ( .A(n613), .B(n587), .ZN(n421) );
  NOR2_X2 U549 ( .A1(n585), .A2(n691), .ZN(n423) );
  XNOR2_X1 U550 ( .A(n531), .B(n448), .ZN(n426) );
  INV_X1 U551 ( .A(n696), .ZN(n428) );
  INV_X1 U552 ( .A(n437), .ZN(n650) );
  NOR2_X1 U553 ( .A1(n441), .A2(n440), .ZN(n439) );
  AND2_X1 U554 ( .A1(n622), .A2(n442), .ZN(n441) );
  INV_X1 U555 ( .A(KEYINPUT100), .ZN(n442) );
  NAND2_X1 U556 ( .A1(n623), .A2(n740), .ZN(n444) );
  NOR2_X1 U557 ( .A1(n632), .A2(n674), .ZN(n446) );
  BUF_X1 U558 ( .A(n585), .Z(n692) );
  XNOR2_X1 U559 ( .A(n568), .B(KEYINPUT1), .ZN(n585) );
  OR2_X1 U560 ( .A1(n568), .A2(n691), .ZN(n547) );
  AND2_X1 U561 ( .A1(n496), .A2(n709), .ZN(n449) );
  INV_X1 U562 ( .A(KEYINPUT23), .ZN(n478) );
  XNOR2_X1 U563 ( .A(n479), .B(n478), .ZN(n481) );
  XNOR2_X1 U564 ( .A(KEYINPUT10), .B(KEYINPUT69), .ZN(n450) );
  INV_X1 U565 ( .A(KEYINPUT77), .ZN(n586) );
  BUF_X1 U566 ( .A(n673), .Z(n750) );
  INV_X1 U567 ( .A(G122), .ZN(n451) );
  XNOR2_X1 U568 ( .A(n451), .B(G104), .ZN(n529) );
  XNOR2_X1 U569 ( .A(n483), .B(n529), .ZN(n456) );
  NAND2_X1 U570 ( .A1(G214), .A2(n505), .ZN(n453) );
  NOR2_X1 U571 ( .A1(G902), .A2(n723), .ZN(n458) );
  XNOR2_X1 U572 ( .A(KEYINPUT13), .B(G475), .ZN(n457) );
  XNOR2_X1 U573 ( .A(n458), .B(n457), .ZN(n557) );
  INV_X1 U574 ( .A(G116), .ZN(n459) );
  XNOR2_X1 U575 ( .A(n459), .B(G107), .ZN(n528) );
  XOR2_X1 U576 ( .A(n528), .B(KEYINPUT9), .Z(n461) );
  XNOR2_X1 U577 ( .A(G134), .B(KEYINPUT7), .ZN(n460) );
  XNOR2_X1 U578 ( .A(n461), .B(n460), .ZN(n470) );
  INV_X4 U579 ( .A(G953), .ZN(n751) );
  NAND2_X1 U580 ( .A1(G234), .A2(n751), .ZN(n463) );
  XNOR2_X1 U581 ( .A(G122), .B(KEYINPUT96), .ZN(n466) );
  XNOR2_X2 U582 ( .A(G143), .B(G128), .ZN(n498) );
  XNOR2_X1 U583 ( .A(n498), .B(n466), .ZN(n467) );
  XNOR2_X1 U584 ( .A(n468), .B(n467), .ZN(n469) );
  XNOR2_X1 U585 ( .A(n470), .B(n469), .ZN(n728) );
  NOR2_X1 U586 ( .A1(G902), .A2(n728), .ZN(n472) );
  INV_X1 U587 ( .A(G478), .ZN(n471) );
  XNOR2_X1 U588 ( .A(n472), .B(n471), .ZN(n558) );
  XNOR2_X2 U589 ( .A(n473), .B(KEYINPUT97), .ZN(n665) );
  INV_X1 U590 ( .A(KEYINPUT99), .ZN(n474) );
  INV_X1 U591 ( .A(KEYINPUT47), .ZN(n476) );
  XNOR2_X1 U592 ( .A(KEYINPUT76), .B(n477), .ZN(n545) );
  XOR2_X1 U593 ( .A(KEYINPUT25), .B(KEYINPUT92), .Z(n488) );
  XOR2_X1 U594 ( .A(KEYINPUT91), .B(KEYINPUT20), .Z(n486) );
  XNOR2_X1 U595 ( .A(G902), .B(KEYINPUT15), .ZN(n537) );
  NAND2_X1 U596 ( .A1(G234), .A2(n537), .ZN(n485) );
  XNOR2_X1 U597 ( .A(n486), .B(n485), .ZN(n491) );
  AND2_X1 U598 ( .A1(n491), .A2(G217), .ZN(n487) );
  XNOR2_X1 U599 ( .A(n488), .B(n487), .ZN(n489) );
  AND2_X1 U600 ( .A1(n491), .A2(G221), .ZN(n492) );
  XNOR2_X1 U601 ( .A(n492), .B(KEYINPUT21), .ZN(n695) );
  NOR2_X1 U602 ( .A1(G900), .A2(n751), .ZN(n493) );
  NAND2_X1 U603 ( .A1(n493), .A2(G902), .ZN(n494) );
  NAND2_X1 U604 ( .A1(n751), .A2(G952), .ZN(n591) );
  NAND2_X1 U605 ( .A1(n494), .A2(n591), .ZN(n496) );
  XNOR2_X1 U606 ( .A(n495), .B(KEYINPUT14), .ZN(n709) );
  NAND2_X1 U607 ( .A1(n695), .A2(n449), .ZN(n497) );
  XNOR2_X1 U608 ( .A(n499), .B(G131), .ZN(n500) );
  XNOR2_X1 U609 ( .A(G119), .B(G113), .ZN(n501) );
  XNOR2_X1 U610 ( .A(n501), .B(KEYINPUT3), .ZN(n504) );
  XNOR2_X1 U611 ( .A(n502), .B(G101), .ZN(n503) );
  XNOR2_X1 U612 ( .A(n504), .B(n503), .ZN(n534) );
  NAND2_X1 U613 ( .A1(n505), .A2(G210), .ZN(n507) );
  XNOR2_X1 U614 ( .A(n507), .B(n506), .ZN(n509) );
  XNOR2_X1 U615 ( .A(KEYINPUT78), .B(KEYINPUT5), .ZN(n508) );
  XNOR2_X1 U616 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U617 ( .A(n534), .B(n510), .ZN(n511) );
  INV_X1 U618 ( .A(KEYINPUT72), .ZN(n512) );
  XNOR2_X1 U619 ( .A(n512), .B(G472), .ZN(n513) );
  XNOR2_X1 U620 ( .A(G101), .B(G107), .ZN(n515) );
  NAND2_X1 U621 ( .A1(G227), .A2(n751), .ZN(n518) );
  INV_X1 U622 ( .A(G902), .ZN(n539) );
  NAND2_X1 U623 ( .A1(n719), .A2(n539), .ZN(n520) );
  INV_X1 U624 ( .A(G469), .ZN(n519) );
  XNOR2_X2 U625 ( .A(n520), .B(n519), .ZN(n568) );
  XOR2_X1 U626 ( .A(n568), .B(KEYINPUT106), .Z(n521) );
  NAND2_X1 U627 ( .A1(G224), .A2(n751), .ZN(n522) );
  XNOR2_X1 U628 ( .A(n522), .B(KEYINPUT18), .ZN(n525) );
  XNOR2_X1 U629 ( .A(KEYINPUT17), .B(n523), .ZN(n524) );
  XNOR2_X1 U630 ( .A(n525), .B(n524), .ZN(n527) );
  XNOR2_X1 U631 ( .A(n526), .B(n527), .ZN(n536) );
  XNOR2_X1 U632 ( .A(n529), .B(n528), .ZN(n533) );
  XNOR2_X1 U633 ( .A(n531), .B(n530), .ZN(n532) );
  XNOR2_X1 U634 ( .A(n533), .B(n532), .ZN(n535) );
  INV_X1 U635 ( .A(n537), .ZN(n629) );
  NAND2_X1 U636 ( .A1(n539), .A2(n538), .ZN(n542) );
  AND2_X1 U637 ( .A1(n542), .A2(G210), .ZN(n540) );
  XNOR2_X2 U638 ( .A(n541), .B(n540), .ZN(n581) );
  AND2_X1 U639 ( .A1(n542), .A2(G214), .ZN(n559) );
  INV_X1 U640 ( .A(KEYINPUT19), .ZN(n543) );
  INV_X1 U641 ( .A(n595), .ZN(n544) );
  NAND2_X1 U642 ( .A1(n546), .A2(n695), .ZN(n691) );
  INV_X1 U643 ( .A(KEYINPUT104), .ZN(n549) );
  XNOR2_X1 U644 ( .A(n550), .B(n549), .ZN(n551) );
  AND2_X1 U645 ( .A1(n557), .A2(n558), .ZN(n597) );
  NAND2_X1 U646 ( .A1(n618), .A2(n662), .ZN(n552) );
  INV_X1 U647 ( .A(KEYINPUT38), .ZN(n553) );
  XNOR2_X1 U648 ( .A(n581), .B(n553), .ZN(n680) );
  NAND2_X1 U649 ( .A1(n554), .A2(n680), .ZN(n556) );
  XOR2_X1 U650 ( .A(KEYINPUT84), .B(KEYINPUT39), .Z(n555) );
  OR2_X1 U651 ( .A1(n558), .A2(n557), .ZN(n682) );
  NAND2_X1 U652 ( .A1(n680), .A2(n373), .ZN(n683) );
  XNOR2_X1 U653 ( .A(KEYINPUT82), .B(KEYINPUT46), .ZN(n562) );
  XNOR2_X1 U654 ( .A(n575), .B(KEYINPUT107), .ZN(n567) );
  INV_X1 U655 ( .A(n565), .ZN(n566) );
  INV_X1 U656 ( .A(KEYINPUT48), .ZN(n569) );
  XNOR2_X1 U657 ( .A(n570), .B(n569), .ZN(n584) );
  OR2_X1 U658 ( .A1(n572), .A2(n571), .ZN(n574) );
  INV_X1 U659 ( .A(KEYINPUT109), .ZN(n573) );
  XNOR2_X1 U660 ( .A(n574), .B(n573), .ZN(n762) );
  INV_X1 U661 ( .A(n575), .ZN(n576) );
  NAND2_X1 U662 ( .A1(n576), .A2(n373), .ZN(n577) );
  XNOR2_X1 U663 ( .A(n577), .B(KEYINPUT103), .ZN(n578) );
  NAND2_X1 U664 ( .A1(n578), .A2(n692), .ZN(n580) );
  INV_X1 U665 ( .A(KEYINPUT43), .ZN(n579) );
  XNOR2_X1 U666 ( .A(n580), .B(n579), .ZN(n582) );
  OR2_X1 U667 ( .A1(n582), .A2(n581), .ZN(n670) );
  AND2_X1 U668 ( .A1(n762), .A2(n670), .ZN(n583) );
  NOR2_X1 U669 ( .A1(G898), .A2(n751), .ZN(n590) );
  XOR2_X1 U670 ( .A(KEYINPUT89), .B(n590), .Z(n738) );
  NAND2_X1 U671 ( .A1(n738), .A2(G902), .ZN(n592) );
  NAND2_X1 U672 ( .A1(n592), .A2(n591), .ZN(n593) );
  NAND2_X1 U673 ( .A1(n593), .A2(n709), .ZN(n594) );
  XNOR2_X2 U674 ( .A(n598), .B(KEYINPUT35), .ZN(n759) );
  INV_X1 U675 ( .A(n695), .ZN(n600) );
  NOR2_X1 U676 ( .A1(n682), .A2(n600), .ZN(n601) );
  INV_X1 U677 ( .A(KEYINPUT73), .ZN(n602) );
  XNOR2_X1 U678 ( .A(n602), .B(KEYINPUT22), .ZN(n603) );
  NAND2_X1 U679 ( .A1(n388), .A2(n605), .ZN(n606) );
  XNOR2_X1 U680 ( .A(n607), .B(KEYINPUT32), .ZN(n647) );
  NAND2_X1 U681 ( .A1(n608), .A2(n692), .ZN(n609) );
  NOR2_X1 U682 ( .A1(n610), .A2(n609), .ZN(n658) );
  INV_X1 U683 ( .A(n759), .ZN(n612) );
  XNOR2_X1 U684 ( .A(KEYINPUT93), .B(KEYINPUT31), .ZN(n615) );
  AND2_X1 U685 ( .A1(n613), .A2(n428), .ZN(n701) );
  NAND2_X1 U686 ( .A1(n701), .A2(n616), .ZN(n614) );
  XOR2_X1 U687 ( .A(n615), .B(n614), .Z(n667) );
  INV_X1 U688 ( .A(n616), .ZN(n617) );
  NOR2_X1 U689 ( .A1(n617), .A2(n350), .ZN(n653) );
  NOR2_X1 U690 ( .A1(n667), .A2(n653), .ZN(n619) );
  INV_X1 U691 ( .A(n618), .ZN(n684) );
  NOR2_X1 U692 ( .A1(n619), .A2(n684), .ZN(n622) );
  INV_X1 U693 ( .A(KEYINPUT65), .ZN(n624) );
  NAND2_X1 U694 ( .A1(n624), .A2(KEYINPUT2), .ZN(n626) );
  NAND2_X1 U695 ( .A1(n629), .A2(KEYINPUT2), .ZN(n625) );
  NAND2_X1 U696 ( .A1(n625), .A2(KEYINPUT65), .ZN(n628) );
  AND2_X1 U697 ( .A1(n626), .A2(n628), .ZN(n627) );
  INV_X1 U698 ( .A(n628), .ZN(n630) );
  OR2_X1 U699 ( .A1(n630), .A2(n629), .ZN(n631) );
  NAND2_X1 U700 ( .A1(n732), .A2(G472), .ZN(n636) );
  XNOR2_X1 U701 ( .A(KEYINPUT86), .B(KEYINPUT62), .ZN(n633) );
  XNOR2_X1 U702 ( .A(n636), .B(n635), .ZN(n638) );
  INV_X1 U703 ( .A(G952), .ZN(n637) );
  NOR2_X2 U704 ( .A1(n638), .A2(n736), .ZN(n640) );
  INV_X1 U705 ( .A(KEYINPUT63), .ZN(n639) );
  XNOR2_X1 U706 ( .A(n640), .B(n639), .ZN(G57) );
  NAND2_X1 U707 ( .A1(n732), .A2(G210), .ZN(n644) );
  XOR2_X1 U708 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n641) );
  XNOR2_X1 U709 ( .A(n644), .B(n643), .ZN(n645) );
  NOR2_X2 U710 ( .A1(n645), .A2(n736), .ZN(n646) );
  XNOR2_X1 U711 ( .A(n646), .B(KEYINPUT56), .ZN(G51) );
  XOR2_X1 U712 ( .A(G119), .B(n647), .Z(G21) );
  XOR2_X1 U713 ( .A(G125), .B(KEYINPUT37), .Z(n648) );
  XNOR2_X1 U714 ( .A(n649), .B(n648), .ZN(G27) );
  XOR2_X1 U715 ( .A(G101), .B(n650), .Z(G3) );
  NAND2_X1 U716 ( .A1(n653), .A2(n665), .ZN(n651) );
  XNOR2_X1 U717 ( .A(n651), .B(G104), .ZN(G6) );
  XNOR2_X1 U718 ( .A(G107), .B(KEYINPUT27), .ZN(n657) );
  XOR2_X1 U719 ( .A(KEYINPUT110), .B(KEYINPUT26), .Z(n655) );
  NAND2_X1 U720 ( .A1(n653), .A2(n652), .ZN(n654) );
  XNOR2_X1 U721 ( .A(n655), .B(n654), .ZN(n656) );
  XNOR2_X1 U722 ( .A(n657), .B(n656), .ZN(G9) );
  XOR2_X1 U723 ( .A(G110), .B(n658), .Z(G12) );
  XOR2_X1 U724 ( .A(KEYINPUT29), .B(KEYINPUT111), .Z(n660) );
  NAND2_X1 U725 ( .A1(n662), .A2(n652), .ZN(n659) );
  XNOR2_X1 U726 ( .A(n660), .B(n659), .ZN(n661) );
  XOR2_X1 U727 ( .A(G128), .B(n661), .Z(G30) );
  NAND2_X1 U728 ( .A1(n662), .A2(n665), .ZN(n663) );
  XNOR2_X1 U729 ( .A(n663), .B(KEYINPUT112), .ZN(n664) );
  XNOR2_X1 U730 ( .A(G146), .B(n664), .ZN(G48) );
  NAND2_X1 U731 ( .A1(n667), .A2(n665), .ZN(n666) );
  XNOR2_X1 U732 ( .A(G113), .B(n666), .ZN(G15) );
  XOR2_X1 U733 ( .A(G116), .B(KEYINPUT113), .Z(n669) );
  NAND2_X1 U734 ( .A1(n667), .A2(n652), .ZN(n668) );
  XNOR2_X1 U735 ( .A(n669), .B(n668), .ZN(G18) );
  XOR2_X1 U736 ( .A(G140), .B(n670), .Z(n671) );
  XNOR2_X1 U737 ( .A(n671), .B(KEYINPUT115), .ZN(G42) );
  NAND2_X1 U738 ( .A1(n688), .A2(n703), .ZN(n672) );
  XNOR2_X1 U739 ( .A(n672), .B(KEYINPUT120), .ZN(n679) );
  NAND2_X1 U740 ( .A1(n740), .A2(n750), .ZN(n675) );
  INV_X1 U741 ( .A(KEYINPUT2), .ZN(n674) );
  NAND2_X1 U742 ( .A1(n675), .A2(n674), .ZN(n677) );
  NAND2_X1 U743 ( .A1(n677), .A2(n676), .ZN(n678) );
  AND2_X1 U744 ( .A1(n679), .A2(n678), .ZN(n714) );
  XNOR2_X1 U745 ( .A(KEYINPUT52), .B(KEYINPUT119), .ZN(n708) );
  NOR2_X1 U746 ( .A1(n680), .A2(n373), .ZN(n681) );
  NOR2_X1 U747 ( .A1(n682), .A2(n681), .ZN(n686) );
  NOR2_X1 U748 ( .A1(n684), .A2(n683), .ZN(n685) );
  NOR2_X1 U749 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U750 ( .A(KEYINPUT117), .B(n687), .ZN(n689) );
  NAND2_X1 U751 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U752 ( .A(n690), .B(KEYINPUT118), .ZN(n706) );
  XOR2_X1 U753 ( .A(KEYINPUT116), .B(KEYINPUT50), .Z(n694) );
  NAND2_X1 U754 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U755 ( .A(n694), .B(n693), .ZN(n699) );
  XNOR2_X1 U756 ( .A(KEYINPUT49), .B(n355), .ZN(n697) );
  NAND2_X1 U757 ( .A1(n697), .A2(n696), .ZN(n698) );
  NOR2_X1 U758 ( .A1(n699), .A2(n698), .ZN(n700) );
  OR2_X1 U759 ( .A1(n701), .A2(n700), .ZN(n702) );
  XOR2_X1 U760 ( .A(KEYINPUT51), .B(n702), .Z(n704) );
  NAND2_X1 U761 ( .A1(n704), .A2(n703), .ZN(n705) );
  NAND2_X1 U762 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U763 ( .A(n708), .B(n707), .ZN(n711) );
  NAND2_X1 U764 ( .A1(n709), .A2(G952), .ZN(n710) );
  NOR2_X1 U765 ( .A1(n711), .A2(n710), .ZN(n712) );
  NOR2_X1 U766 ( .A1(n712), .A2(G953), .ZN(n713) );
  NAND2_X1 U767 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U768 ( .A(n715), .B(KEYINPUT121), .ZN(n716) );
  XNOR2_X1 U769 ( .A(n716), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U770 ( .A1(n349), .A2(G469), .ZN(n721) );
  XOR2_X1 U771 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n717) );
  XOR2_X1 U772 ( .A(n717), .B(KEYINPUT122), .Z(n718) );
  XNOR2_X1 U773 ( .A(n719), .B(n718), .ZN(n720) );
  XNOR2_X1 U774 ( .A(n721), .B(n720), .ZN(n722) );
  NOR2_X1 U775 ( .A1(n736), .A2(n722), .ZN(G54) );
  NAND2_X1 U776 ( .A1(n732), .A2(G475), .ZN(n725) );
  XNOR2_X1 U777 ( .A(n725), .B(n724), .ZN(n726) );
  NOR2_X2 U778 ( .A1(n726), .A2(n736), .ZN(n727) );
  XNOR2_X1 U779 ( .A(n727), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U780 ( .A1(n349), .A2(G478), .ZN(n730) );
  XOR2_X1 U781 ( .A(n728), .B(KEYINPUT123), .Z(n729) );
  XNOR2_X1 U782 ( .A(n730), .B(n729), .ZN(n731) );
  NOR2_X1 U783 ( .A1(n736), .A2(n731), .ZN(G63) );
  NAND2_X1 U784 ( .A1(n349), .A2(G217), .ZN(n734) );
  XNOR2_X1 U785 ( .A(n734), .B(n733), .ZN(n735) );
  NOR2_X1 U786 ( .A1(n736), .A2(n735), .ZN(G66) );
  XOR2_X1 U787 ( .A(KEYINPUT126), .B(n737), .Z(n739) );
  NOR2_X1 U788 ( .A1(n739), .A2(n738), .ZN(n747) );
  NAND2_X1 U789 ( .A1(n740), .A2(n751), .ZN(n745) );
  XOR2_X1 U790 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n742) );
  NAND2_X1 U791 ( .A1(G224), .A2(G953), .ZN(n741) );
  XNOR2_X1 U792 ( .A(n742), .B(n741), .ZN(n743) );
  NAND2_X1 U793 ( .A1(n743), .A2(G898), .ZN(n744) );
  NAND2_X1 U794 ( .A1(n745), .A2(n744), .ZN(n746) );
  XNOR2_X1 U795 ( .A(n747), .B(n746), .ZN(G69) );
  XOR2_X1 U796 ( .A(n749), .B(n748), .Z(n753) );
  XNOR2_X1 U797 ( .A(n750), .B(n753), .ZN(n752) );
  NAND2_X1 U798 ( .A1(n752), .A2(n751), .ZN(n758) );
  XOR2_X1 U799 ( .A(n753), .B(G227), .Z(n754) );
  NAND2_X1 U800 ( .A1(n754), .A2(G900), .ZN(n755) );
  XOR2_X1 U801 ( .A(KEYINPUT127), .B(n755), .Z(n756) );
  NAND2_X1 U802 ( .A1(G953), .A2(n756), .ZN(n757) );
  NAND2_X1 U803 ( .A1(n758), .A2(n757), .ZN(G72) );
  XOR2_X1 U804 ( .A(n759), .B(G122), .Z(G24) );
  XNOR2_X1 U805 ( .A(G143), .B(n760), .ZN(G45) );
  XNOR2_X1 U806 ( .A(G131), .B(n761), .ZN(G33) );
  XNOR2_X1 U807 ( .A(G134), .B(KEYINPUT114), .ZN(n763) );
  XNOR2_X1 U808 ( .A(n763), .B(n762), .ZN(G36) );
  XNOR2_X1 U809 ( .A(G137), .B(n764), .ZN(G39) );
endmodule

