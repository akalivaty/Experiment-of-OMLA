

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U546 ( .A1(n517), .A2(G2105), .ZN(n560) );
  AND2_X1 U547 ( .A1(n782), .A2(n781), .ZN(n792) );
  AND2_X1 U548 ( .A1(n760), .A2(n759), .ZN(n761) );
  XNOR2_X1 U549 ( .A(n510), .B(KEYINPUT93), .ZN(n509) );
  OR2_X1 U550 ( .A1(n751), .A2(n747), .ZN(n510) );
  NOR2_X1 U551 ( .A1(n702), .A2(n701), .ZN(n704) );
  INV_X1 U552 ( .A(KEYINPUT31), .ZN(n703) );
  XOR2_X1 U553 ( .A(KEYINPUT64), .B(G2104), .Z(n517) );
  NOR2_X1 U554 ( .A1(G651), .A2(n627), .ZN(n638) );
  NOR2_X1 U555 ( .A1(G2104), .A2(G2105), .ZN(n511) );
  XOR2_X1 U556 ( .A(KEYINPUT17), .B(n511), .Z(n979) );
  NAND2_X1 U557 ( .A1(G137), .A2(n979), .ZN(n514) );
  NAND2_X1 U558 ( .A1(G2105), .A2(G2104), .ZN(n512) );
  XNOR2_X1 U559 ( .A(n512), .B(KEYINPUT67), .ZN(n977) );
  NAND2_X1 U560 ( .A1(G113), .A2(n977), .ZN(n513) );
  NAND2_X1 U561 ( .A1(n514), .A2(n513), .ZN(n522) );
  XOR2_X1 U562 ( .A(KEYINPUT23), .B(KEYINPUT66), .Z(n516) );
  NAND2_X1 U563 ( .A1(G101), .A2(n560), .ZN(n515) );
  XNOR2_X1 U564 ( .A(n516), .B(n515), .ZN(n520) );
  NAND2_X1 U565 ( .A1(G2105), .A2(n517), .ZN(n518) );
  XNOR2_X2 U566 ( .A(n518), .B(KEYINPUT65), .ZN(n984) );
  NAND2_X1 U567 ( .A1(n984), .A2(G125), .ZN(n519) );
  NAND2_X1 U568 ( .A1(n520), .A2(n519), .ZN(n521) );
  NOR2_X1 U569 ( .A1(n522), .A2(n521), .ZN(G160) );
  NOR2_X1 U570 ( .A1(G543), .A2(G651), .ZN(n630) );
  NAND2_X1 U571 ( .A1(G90), .A2(n630), .ZN(n524) );
  XOR2_X1 U572 ( .A(G543), .B(KEYINPUT0), .Z(n627) );
  INV_X1 U573 ( .A(G651), .ZN(n526) );
  NOR2_X1 U574 ( .A1(n627), .A2(n526), .ZN(n634) );
  NAND2_X1 U575 ( .A1(G77), .A2(n634), .ZN(n523) );
  NAND2_X1 U576 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U577 ( .A(n525), .B(KEYINPUT9), .ZN(n529) );
  NOR2_X1 U578 ( .A1(G543), .A2(n526), .ZN(n527) );
  XOR2_X1 U579 ( .A(KEYINPUT1), .B(n527), .Z(n631) );
  NAND2_X1 U580 ( .A1(G64), .A2(n631), .ZN(n528) );
  NAND2_X1 U581 ( .A1(n529), .A2(n528), .ZN(n532) );
  NAND2_X1 U582 ( .A1(G52), .A2(n638), .ZN(n530) );
  XOR2_X1 U583 ( .A(KEYINPUT70), .B(n530), .Z(n531) );
  NOR2_X1 U584 ( .A1(n532), .A2(n531), .ZN(G171) );
  AND2_X1 U585 ( .A1(G452), .A2(G94), .ZN(G173) );
  BUF_X1 U586 ( .A(n560), .Z(n978) );
  NAND2_X1 U587 ( .A1(G99), .A2(n978), .ZN(n534) );
  NAND2_X1 U588 ( .A1(G135), .A2(n979), .ZN(n533) );
  NAND2_X1 U589 ( .A1(n534), .A2(n533), .ZN(n540) );
  NAND2_X1 U590 ( .A1(G123), .A2(n984), .ZN(n535) );
  XNOR2_X1 U591 ( .A(n535), .B(KEYINPUT78), .ZN(n536) );
  XNOR2_X1 U592 ( .A(n536), .B(KEYINPUT18), .ZN(n538) );
  NAND2_X1 U593 ( .A1(G111), .A2(n977), .ZN(n537) );
  NAND2_X1 U594 ( .A1(n538), .A2(n537), .ZN(n539) );
  NOR2_X1 U595 ( .A1(n540), .A2(n539), .ZN(n970) );
  XNOR2_X1 U596 ( .A(n970), .B(G2096), .ZN(n541) );
  XNOR2_X1 U597 ( .A(n541), .B(KEYINPUT79), .ZN(n542) );
  OR2_X1 U598 ( .A1(G2100), .A2(n542), .ZN(G156) );
  INV_X1 U599 ( .A(G57), .ZN(G237) );
  INV_X1 U600 ( .A(G82), .ZN(G220) );
  NAND2_X1 U601 ( .A1(G88), .A2(n630), .ZN(n544) );
  NAND2_X1 U602 ( .A1(G75), .A2(n634), .ZN(n543) );
  NAND2_X1 U603 ( .A1(n544), .A2(n543), .ZN(n548) );
  NAND2_X1 U604 ( .A1(G50), .A2(n638), .ZN(n546) );
  NAND2_X1 U605 ( .A1(G62), .A2(n631), .ZN(n545) );
  NAND2_X1 U606 ( .A1(n546), .A2(n545), .ZN(n547) );
  NOR2_X1 U607 ( .A1(n548), .A2(n547), .ZN(G166) );
  NAND2_X1 U608 ( .A1(G51), .A2(n638), .ZN(n550) );
  NAND2_X1 U609 ( .A1(G63), .A2(n631), .ZN(n549) );
  NAND2_X1 U610 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U611 ( .A(KEYINPUT6), .B(n551), .ZN(n557) );
  NAND2_X1 U612 ( .A1(n630), .A2(G89), .ZN(n552) );
  XNOR2_X1 U613 ( .A(n552), .B(KEYINPUT4), .ZN(n554) );
  NAND2_X1 U614 ( .A1(G76), .A2(n634), .ZN(n553) );
  NAND2_X1 U615 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U616 ( .A(n555), .B(KEYINPUT5), .Z(n556) );
  NOR2_X1 U617 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U618 ( .A(KEYINPUT75), .B(n558), .Z(n559) );
  XOR2_X1 U619 ( .A(KEYINPUT7), .B(n559), .Z(G168) );
  XOR2_X1 U620 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U621 ( .A1(n560), .A2(G102), .ZN(n563) );
  NAND2_X1 U622 ( .A1(G114), .A2(n977), .ZN(n561) );
  XOR2_X1 U623 ( .A(KEYINPUT85), .B(n561), .Z(n562) );
  NAND2_X1 U624 ( .A1(n563), .A2(n562), .ZN(n567) );
  NAND2_X1 U625 ( .A1(G138), .A2(n979), .ZN(n565) );
  NAND2_X1 U626 ( .A1(G126), .A2(n984), .ZN(n564) );
  NAND2_X1 U627 ( .A1(n565), .A2(n564), .ZN(n566) );
  NOR2_X1 U628 ( .A1(n567), .A2(n566), .ZN(G164) );
  NAND2_X1 U629 ( .A1(G7), .A2(G661), .ZN(n568) );
  XNOR2_X1 U630 ( .A(n568), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U631 ( .A(G223), .ZN(n813) );
  NAND2_X1 U632 ( .A1(n813), .A2(G567), .ZN(n569) );
  XOR2_X1 U633 ( .A(KEYINPUT11), .B(n569), .Z(G234) );
  NAND2_X1 U634 ( .A1(G56), .A2(n631), .ZN(n570) );
  XOR2_X1 U635 ( .A(KEYINPUT14), .B(n570), .Z(n576) );
  NAND2_X1 U636 ( .A1(n630), .A2(G81), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n571), .B(KEYINPUT12), .ZN(n573) );
  NAND2_X1 U638 ( .A1(G68), .A2(n634), .ZN(n572) );
  NAND2_X1 U639 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U640 ( .A(KEYINPUT13), .B(n574), .Z(n575) );
  NOR2_X1 U641 ( .A1(n576), .A2(n575), .ZN(n578) );
  NAND2_X1 U642 ( .A1(n638), .A2(G43), .ZN(n577) );
  NAND2_X1 U643 ( .A1(n578), .A2(n577), .ZN(n879) );
  INV_X1 U644 ( .A(G860), .ZN(n599) );
  OR2_X1 U645 ( .A1(n879), .A2(n599), .ZN(G153) );
  INV_X1 U646 ( .A(G868), .ZN(n650) );
  NOR2_X1 U647 ( .A1(n650), .A2(G171), .ZN(n579) );
  XNOR2_X1 U648 ( .A(n579), .B(KEYINPUT73), .ZN(n588) );
  NAND2_X1 U649 ( .A1(G79), .A2(n634), .ZN(n581) );
  NAND2_X1 U650 ( .A1(G54), .A2(n638), .ZN(n580) );
  NAND2_X1 U651 ( .A1(n581), .A2(n580), .ZN(n585) );
  NAND2_X1 U652 ( .A1(G92), .A2(n630), .ZN(n583) );
  NAND2_X1 U653 ( .A1(G66), .A2(n631), .ZN(n582) );
  NAND2_X1 U654 ( .A1(n583), .A2(n582), .ZN(n584) );
  NOR2_X1 U655 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U656 ( .A(n586), .B(KEYINPUT15), .ZN(n963) );
  NAND2_X1 U657 ( .A1(n650), .A2(n963), .ZN(n587) );
  NAND2_X1 U658 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U659 ( .A(KEYINPUT74), .B(n589), .ZN(G284) );
  NAND2_X1 U660 ( .A1(G53), .A2(n638), .ZN(n591) );
  NAND2_X1 U661 ( .A1(G65), .A2(n631), .ZN(n590) );
  NAND2_X1 U662 ( .A1(n591), .A2(n590), .ZN(n595) );
  NAND2_X1 U663 ( .A1(G91), .A2(n630), .ZN(n593) );
  NAND2_X1 U664 ( .A1(G78), .A2(n634), .ZN(n592) );
  NAND2_X1 U665 ( .A1(n593), .A2(n592), .ZN(n594) );
  NOR2_X1 U666 ( .A1(n595), .A2(n594), .ZN(n885) );
  XNOR2_X1 U667 ( .A(n885), .B(KEYINPUT71), .ZN(G299) );
  NOR2_X1 U668 ( .A1(G286), .A2(n650), .ZN(n596) );
  XNOR2_X1 U669 ( .A(n596), .B(KEYINPUT76), .ZN(n598) );
  NOR2_X1 U670 ( .A1(G299), .A2(G868), .ZN(n597) );
  NOR2_X1 U671 ( .A1(n598), .A2(n597), .ZN(G297) );
  NAND2_X1 U672 ( .A1(n599), .A2(G559), .ZN(n600) );
  INV_X1 U673 ( .A(n963), .ZN(n606) );
  NAND2_X1 U674 ( .A1(n600), .A2(n606), .ZN(n601) );
  XNOR2_X1 U675 ( .A(n601), .B(KEYINPUT77), .ZN(n602) );
  XOR2_X1 U676 ( .A(KEYINPUT16), .B(n602), .Z(G148) );
  NOR2_X1 U677 ( .A1(G868), .A2(n879), .ZN(n605) );
  NAND2_X1 U678 ( .A1(G868), .A2(n606), .ZN(n603) );
  NOR2_X1 U679 ( .A1(G559), .A2(n603), .ZN(n604) );
  NOR2_X1 U680 ( .A1(n605), .A2(n604), .ZN(G282) );
  NAND2_X1 U681 ( .A1(n606), .A2(G559), .ZN(n647) );
  XNOR2_X1 U682 ( .A(n879), .B(n647), .ZN(n607) );
  NOR2_X1 U683 ( .A1(n607), .A2(G860), .ZN(n615) );
  NAND2_X1 U684 ( .A1(G55), .A2(n638), .ZN(n609) );
  NAND2_X1 U685 ( .A1(G67), .A2(n631), .ZN(n608) );
  NAND2_X1 U686 ( .A1(n609), .A2(n608), .ZN(n610) );
  XNOR2_X1 U687 ( .A(KEYINPUT80), .B(n610), .ZN(n614) );
  NAND2_X1 U688 ( .A1(G93), .A2(n630), .ZN(n612) );
  NAND2_X1 U689 ( .A1(G80), .A2(n634), .ZN(n611) );
  NAND2_X1 U690 ( .A1(n612), .A2(n611), .ZN(n613) );
  OR2_X1 U691 ( .A1(n614), .A2(n613), .ZN(n651) );
  XOR2_X1 U692 ( .A(n615), .B(n651), .Z(G145) );
  NAND2_X1 U693 ( .A1(G47), .A2(n638), .ZN(n617) );
  NAND2_X1 U694 ( .A1(G60), .A2(n631), .ZN(n616) );
  NAND2_X1 U695 ( .A1(n617), .A2(n616), .ZN(n618) );
  XNOR2_X1 U696 ( .A(KEYINPUT69), .B(n618), .ZN(n623) );
  NAND2_X1 U697 ( .A1(G85), .A2(n630), .ZN(n620) );
  NAND2_X1 U698 ( .A1(G72), .A2(n634), .ZN(n619) );
  NAND2_X1 U699 ( .A1(n620), .A2(n619), .ZN(n621) );
  XOR2_X1 U700 ( .A(KEYINPUT68), .B(n621), .Z(n622) );
  NAND2_X1 U701 ( .A1(n623), .A2(n622), .ZN(G290) );
  NAND2_X1 U702 ( .A1(G49), .A2(n638), .ZN(n625) );
  NAND2_X1 U703 ( .A1(G74), .A2(G651), .ZN(n624) );
  NAND2_X1 U704 ( .A1(n625), .A2(n624), .ZN(n626) );
  NOR2_X1 U705 ( .A1(n631), .A2(n626), .ZN(n629) );
  NAND2_X1 U706 ( .A1(n627), .A2(G87), .ZN(n628) );
  NAND2_X1 U707 ( .A1(n629), .A2(n628), .ZN(G288) );
  NAND2_X1 U708 ( .A1(G86), .A2(n630), .ZN(n633) );
  NAND2_X1 U709 ( .A1(G61), .A2(n631), .ZN(n632) );
  NAND2_X1 U710 ( .A1(n633), .A2(n632), .ZN(n637) );
  NAND2_X1 U711 ( .A1(n634), .A2(G73), .ZN(n635) );
  XOR2_X1 U712 ( .A(KEYINPUT2), .B(n635), .Z(n636) );
  NOR2_X1 U713 ( .A1(n637), .A2(n636), .ZN(n640) );
  NAND2_X1 U714 ( .A1(n638), .A2(G48), .ZN(n639) );
  NAND2_X1 U715 ( .A1(n640), .A2(n639), .ZN(G305) );
  XOR2_X1 U716 ( .A(n651), .B(G290), .Z(n643) );
  XOR2_X1 U717 ( .A(KEYINPUT19), .B(G288), .Z(n641) );
  XNOR2_X1 U718 ( .A(G299), .B(n641), .ZN(n642) );
  XNOR2_X1 U719 ( .A(n643), .B(n642), .ZN(n644) );
  XNOR2_X1 U720 ( .A(G166), .B(n644), .ZN(n645) );
  XNOR2_X1 U721 ( .A(n645), .B(G305), .ZN(n646) );
  XNOR2_X1 U722 ( .A(n879), .B(n646), .ZN(n964) );
  XNOR2_X1 U723 ( .A(n964), .B(n647), .ZN(n648) );
  NAND2_X1 U724 ( .A1(n648), .A2(G868), .ZN(n649) );
  XOR2_X1 U725 ( .A(KEYINPUT81), .B(n649), .Z(n653) );
  NAND2_X1 U726 ( .A1(n651), .A2(n650), .ZN(n652) );
  NAND2_X1 U727 ( .A1(n653), .A2(n652), .ZN(G295) );
  NAND2_X1 U728 ( .A1(G2078), .A2(G2084), .ZN(n654) );
  XOR2_X1 U729 ( .A(KEYINPUT20), .B(n654), .Z(n655) );
  NAND2_X1 U730 ( .A1(G2090), .A2(n655), .ZN(n656) );
  XNOR2_X1 U731 ( .A(KEYINPUT21), .B(n656), .ZN(n657) );
  NAND2_X1 U732 ( .A1(n657), .A2(G2072), .ZN(n658) );
  XNOR2_X1 U733 ( .A(KEYINPUT82), .B(n658), .ZN(G158) );
  XOR2_X1 U734 ( .A(KEYINPUT72), .B(G132), .Z(G219) );
  XNOR2_X1 U735 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U736 ( .A1(G661), .A2(G483), .ZN(n667) );
  NOR2_X1 U737 ( .A1(G219), .A2(G220), .ZN(n660) );
  XNOR2_X1 U738 ( .A(KEYINPUT22), .B(KEYINPUT83), .ZN(n659) );
  XNOR2_X1 U739 ( .A(n660), .B(n659), .ZN(n661) );
  NOR2_X1 U740 ( .A1(n661), .A2(G218), .ZN(n662) );
  NAND2_X1 U741 ( .A1(G96), .A2(n662), .ZN(n818) );
  NAND2_X1 U742 ( .A1(G2106), .A2(n818), .ZN(n666) );
  NAND2_X1 U743 ( .A1(G69), .A2(G120), .ZN(n663) );
  NOR2_X1 U744 ( .A1(G237), .A2(n663), .ZN(n664) );
  NAND2_X1 U745 ( .A1(G108), .A2(n664), .ZN(n819) );
  NAND2_X1 U746 ( .A1(G567), .A2(n819), .ZN(n665) );
  NAND2_X1 U747 ( .A1(n666), .A2(n665), .ZN(n941) );
  NOR2_X1 U748 ( .A1(n667), .A2(n941), .ZN(n668) );
  XNOR2_X1 U749 ( .A(n668), .B(KEYINPUT84), .ZN(n816) );
  NAND2_X1 U750 ( .A1(G36), .A2(n816), .ZN(G176) );
  INV_X1 U751 ( .A(G166), .ZN(G303) );
  NAND2_X1 U752 ( .A1(G107), .A2(n977), .ZN(n670) );
  NAND2_X1 U753 ( .A1(G119), .A2(n984), .ZN(n669) );
  NAND2_X1 U754 ( .A1(n670), .A2(n669), .ZN(n671) );
  XNOR2_X1 U755 ( .A(KEYINPUT88), .B(n671), .ZN(n675) );
  NAND2_X1 U756 ( .A1(G95), .A2(n978), .ZN(n673) );
  NAND2_X1 U757 ( .A1(G131), .A2(n979), .ZN(n672) );
  NAND2_X1 U758 ( .A1(n673), .A2(n672), .ZN(n674) );
  NOR2_X1 U759 ( .A1(n675), .A2(n674), .ZN(n974) );
  INV_X1 U760 ( .A(G1991), .ZN(n829) );
  NOR2_X1 U761 ( .A1(n974), .A2(n829), .ZN(n685) );
  NAND2_X1 U762 ( .A1(G105), .A2(n978), .ZN(n676) );
  XOR2_X1 U763 ( .A(KEYINPUT89), .B(n676), .Z(n677) );
  XNOR2_X1 U764 ( .A(n677), .B(KEYINPUT38), .ZN(n679) );
  NAND2_X1 U765 ( .A1(G141), .A2(n979), .ZN(n678) );
  NAND2_X1 U766 ( .A1(n679), .A2(n678), .ZN(n683) );
  NAND2_X1 U767 ( .A1(G117), .A2(n977), .ZN(n681) );
  NAND2_X1 U768 ( .A1(G129), .A2(n984), .ZN(n680) );
  NAND2_X1 U769 ( .A1(n681), .A2(n680), .ZN(n682) );
  NOR2_X1 U770 ( .A1(n683), .A2(n682), .ZN(n972) );
  INV_X1 U771 ( .A(G1996), .ZN(n797) );
  NOR2_X1 U772 ( .A1(n972), .A2(n797), .ZN(n684) );
  NOR2_X1 U773 ( .A1(n685), .A2(n684), .ZN(n912) );
  INV_X1 U774 ( .A(n912), .ZN(n689) );
  NOR2_X1 U775 ( .A1(G164), .A2(G1384), .ZN(n696) );
  NAND2_X1 U776 ( .A1(G40), .A2(G160), .ZN(n688) );
  INV_X1 U777 ( .A(KEYINPUT87), .ZN(n687) );
  XNOR2_X1 U778 ( .A(n688), .B(n687), .ZN(n692) );
  NOR2_X1 U779 ( .A1(n696), .A2(n692), .ZN(n807) );
  NAND2_X1 U780 ( .A1(n689), .A2(n807), .ZN(n793) );
  XNOR2_X1 U781 ( .A(KEYINPUT86), .B(G1986), .ZN(n690) );
  XNOR2_X1 U782 ( .A(n690), .B(G290), .ZN(n897) );
  NAND2_X1 U783 ( .A1(n807), .A2(n897), .ZN(n691) );
  AND2_X1 U784 ( .A1(n793), .A2(n691), .ZN(n782) );
  INV_X1 U785 ( .A(n692), .ZN(n697) );
  NAND2_X2 U786 ( .A1(n697), .A2(n696), .ZN(n735) );
  NAND2_X2 U787 ( .A1(G8), .A2(n735), .ZN(n776) );
  NOR2_X2 U788 ( .A1(G1966), .A2(n776), .ZN(n751) );
  NOR2_X1 U789 ( .A1(G2084), .A2(n735), .ZN(n747) );
  NAND2_X1 U790 ( .A1(G8), .A2(n509), .ZN(n693) );
  XNOR2_X1 U791 ( .A(n693), .B(KEYINPUT30), .ZN(n694) );
  NOR2_X1 U792 ( .A1(G168), .A2(n694), .ZN(n695) );
  XNOR2_X1 U793 ( .A(n695), .B(KEYINPUT94), .ZN(n702) );
  NAND2_X1 U794 ( .A1(G1961), .A2(n735), .ZN(n699) );
  AND2_X1 U795 ( .A1(n697), .A2(n696), .ZN(n713) );
  XOR2_X1 U796 ( .A(G2078), .B(KEYINPUT25), .Z(n836) );
  NAND2_X1 U797 ( .A1(n713), .A2(n836), .ZN(n698) );
  NAND2_X1 U798 ( .A1(n699), .A2(n698), .ZN(n700) );
  XOR2_X1 U799 ( .A(KEYINPUT90), .B(n700), .Z(n705) );
  NOR2_X1 U800 ( .A1(n705), .A2(G171), .ZN(n701) );
  XNOR2_X1 U801 ( .A(n704), .B(n703), .ZN(n748) );
  NAND2_X1 U802 ( .A1(n705), .A2(G171), .ZN(n734) );
  NAND2_X1 U803 ( .A1(n713), .A2(G2072), .ZN(n706) );
  XNOR2_X1 U804 ( .A(n706), .B(KEYINPUT27), .ZN(n708) );
  AND2_X1 U805 ( .A1(G1956), .A2(n735), .ZN(n707) );
  NOR2_X1 U806 ( .A1(n708), .A2(n707), .ZN(n711) );
  NOR2_X1 U807 ( .A1(n885), .A2(n711), .ZN(n710) );
  XNOR2_X1 U808 ( .A(KEYINPUT91), .B(KEYINPUT28), .ZN(n709) );
  XNOR2_X1 U809 ( .A(n710), .B(n709), .ZN(n731) );
  NAND2_X1 U810 ( .A1(n885), .A2(n711), .ZN(n729) );
  XNOR2_X1 U811 ( .A(KEYINPUT26), .B(KEYINPUT92), .ZN(n719) );
  NOR2_X1 U812 ( .A1(G1996), .A2(n719), .ZN(n712) );
  NOR2_X1 U813 ( .A1(n712), .A2(n879), .ZN(n717) );
  NAND2_X1 U814 ( .A1(G1348), .A2(n735), .ZN(n715) );
  NAND2_X1 U815 ( .A1(n713), .A2(G2067), .ZN(n714) );
  NAND2_X1 U816 ( .A1(n715), .A2(n714), .ZN(n725) );
  NAND2_X1 U817 ( .A1(n963), .A2(n725), .ZN(n716) );
  NAND2_X1 U818 ( .A1(n717), .A2(n716), .ZN(n724) );
  INV_X1 U819 ( .A(G1341), .ZN(n880) );
  NAND2_X1 U820 ( .A1(n880), .A2(n719), .ZN(n718) );
  NAND2_X1 U821 ( .A1(n718), .A2(n735), .ZN(n722) );
  NOR2_X1 U822 ( .A1(n735), .A2(n797), .ZN(n720) );
  NAND2_X1 U823 ( .A1(n720), .A2(n719), .ZN(n721) );
  NAND2_X1 U824 ( .A1(n722), .A2(n721), .ZN(n723) );
  NOR2_X1 U825 ( .A1(n724), .A2(n723), .ZN(n727) );
  NOR2_X1 U826 ( .A1(n725), .A2(n963), .ZN(n726) );
  NOR2_X1 U827 ( .A1(n727), .A2(n726), .ZN(n728) );
  NAND2_X1 U828 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U829 ( .A1(n731), .A2(n730), .ZN(n732) );
  XOR2_X1 U830 ( .A(KEYINPUT29), .B(n732), .Z(n733) );
  NAND2_X1 U831 ( .A1(n734), .A2(n733), .ZN(n749) );
  INV_X1 U832 ( .A(G8), .ZN(n740) );
  NOR2_X1 U833 ( .A1(G1971), .A2(n776), .ZN(n737) );
  NOR2_X1 U834 ( .A1(G2090), .A2(n735), .ZN(n736) );
  NOR2_X1 U835 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U836 ( .A1(n738), .A2(G303), .ZN(n739) );
  OR2_X1 U837 ( .A1(n740), .A2(n739), .ZN(n742) );
  AND2_X1 U838 ( .A1(n749), .A2(n742), .ZN(n741) );
  NAND2_X1 U839 ( .A1(n748), .A2(n741), .ZN(n745) );
  INV_X1 U840 ( .A(n742), .ZN(n743) );
  OR2_X1 U841 ( .A1(n743), .A2(G286), .ZN(n744) );
  NAND2_X1 U842 ( .A1(n745), .A2(n744), .ZN(n746) );
  XNOR2_X1 U843 ( .A(n746), .B(KEYINPUT32), .ZN(n755) );
  NAND2_X1 U844 ( .A1(G8), .A2(n747), .ZN(n753) );
  AND2_X1 U845 ( .A1(n749), .A2(n748), .ZN(n750) );
  NOR2_X1 U846 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U847 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U848 ( .A1(n755), .A2(n754), .ZN(n772) );
  NOR2_X1 U849 ( .A1(G1976), .A2(G288), .ZN(n763) );
  NOR2_X1 U850 ( .A1(G1971), .A2(G303), .ZN(n756) );
  NOR2_X1 U851 ( .A1(n763), .A2(n756), .ZN(n876) );
  NAND2_X1 U852 ( .A1(n772), .A2(n876), .ZN(n760) );
  INV_X1 U853 ( .A(KEYINPUT33), .ZN(n758) );
  NAND2_X1 U854 ( .A1(G288), .A2(G1976), .ZN(n757) );
  XOR2_X1 U855 ( .A(KEYINPUT95), .B(n757), .Z(n875) );
  AND2_X1 U856 ( .A1(n758), .A2(n875), .ZN(n759) );
  INV_X1 U857 ( .A(n776), .ZN(n762) );
  NAND2_X1 U858 ( .A1(n761), .A2(n762), .ZN(n766) );
  NAND2_X1 U859 ( .A1(n763), .A2(n762), .ZN(n764) );
  NAND2_X1 U860 ( .A1(n764), .A2(KEYINPUT33), .ZN(n765) );
  NAND2_X1 U861 ( .A1(n766), .A2(n765), .ZN(n767) );
  XNOR2_X1 U862 ( .A(n767), .B(KEYINPUT96), .ZN(n768) );
  XOR2_X1 U863 ( .A(G1981), .B(G305), .Z(n888) );
  NAND2_X1 U864 ( .A1(n768), .A2(n888), .ZN(n780) );
  NAND2_X1 U865 ( .A1(G8), .A2(G166), .ZN(n769) );
  NOR2_X1 U866 ( .A1(G2090), .A2(n769), .ZN(n770) );
  XNOR2_X1 U867 ( .A(KEYINPUT97), .B(n770), .ZN(n771) );
  NAND2_X1 U868 ( .A1(n772), .A2(n771), .ZN(n773) );
  AND2_X1 U869 ( .A1(n773), .A2(n776), .ZN(n778) );
  NOR2_X1 U870 ( .A1(G1981), .A2(G305), .ZN(n774) );
  XOR2_X1 U871 ( .A(n774), .B(KEYINPUT24), .Z(n775) );
  NOR2_X1 U872 ( .A1(n776), .A2(n775), .ZN(n777) );
  NOR2_X1 U873 ( .A1(n778), .A2(n777), .ZN(n779) );
  NAND2_X1 U874 ( .A1(n780), .A2(n779), .ZN(n781) );
  NAND2_X1 U875 ( .A1(G104), .A2(n978), .ZN(n784) );
  NAND2_X1 U876 ( .A1(G140), .A2(n979), .ZN(n783) );
  NAND2_X1 U877 ( .A1(n784), .A2(n783), .ZN(n785) );
  XNOR2_X1 U878 ( .A(KEYINPUT34), .B(n785), .ZN(n790) );
  NAND2_X1 U879 ( .A1(G116), .A2(n977), .ZN(n787) );
  NAND2_X1 U880 ( .A1(G128), .A2(n984), .ZN(n786) );
  NAND2_X1 U881 ( .A1(n787), .A2(n786), .ZN(n788) );
  XOR2_X1 U882 ( .A(KEYINPUT35), .B(n788), .Z(n789) );
  NOR2_X1 U883 ( .A1(n790), .A2(n789), .ZN(n791) );
  XNOR2_X1 U884 ( .A(KEYINPUT36), .B(n791), .ZN(n995) );
  XNOR2_X1 U885 ( .A(G2067), .B(KEYINPUT37), .ZN(n804) );
  NOR2_X1 U886 ( .A1(n995), .A2(n804), .ZN(n931) );
  NAND2_X1 U887 ( .A1(n931), .A2(n807), .ZN(n802) );
  NAND2_X1 U888 ( .A1(n792), .A2(n802), .ZN(n810) );
  INV_X1 U889 ( .A(n793), .ZN(n796) );
  NOR2_X1 U890 ( .A1(G1986), .A2(G290), .ZN(n794) );
  AND2_X1 U891 ( .A1(n829), .A2(n974), .ZN(n914) );
  NOR2_X1 U892 ( .A1(n794), .A2(n914), .ZN(n795) );
  NOR2_X1 U893 ( .A1(n796), .A2(n795), .ZN(n798) );
  AND2_X1 U894 ( .A1(n797), .A2(n972), .ZN(n908) );
  NOR2_X1 U895 ( .A1(n798), .A2(n908), .ZN(n800) );
  XNOR2_X1 U896 ( .A(KEYINPUT39), .B(KEYINPUT98), .ZN(n799) );
  XNOR2_X1 U897 ( .A(n800), .B(n799), .ZN(n801) );
  NAND2_X1 U898 ( .A1(n802), .A2(n801), .ZN(n803) );
  XOR2_X1 U899 ( .A(KEYINPUT99), .B(n803), .Z(n805) );
  NAND2_X1 U900 ( .A1(n995), .A2(n804), .ZN(n929) );
  NAND2_X1 U901 ( .A1(n805), .A2(n929), .ZN(n806) );
  NAND2_X1 U902 ( .A1(n807), .A2(n806), .ZN(n808) );
  XNOR2_X1 U903 ( .A(n808), .B(KEYINPUT100), .ZN(n809) );
  NAND2_X1 U904 ( .A1(n810), .A2(n809), .ZN(n812) );
  XOR2_X1 U905 ( .A(KEYINPUT40), .B(KEYINPUT101), .Z(n811) );
  XNOR2_X1 U906 ( .A(n812), .B(n811), .ZN(G329) );
  NAND2_X1 U907 ( .A1(G2106), .A2(n813), .ZN(G217) );
  AND2_X1 U908 ( .A1(G15), .A2(G2), .ZN(n814) );
  NAND2_X1 U909 ( .A1(G661), .A2(n814), .ZN(G259) );
  NAND2_X1 U910 ( .A1(G3), .A2(G1), .ZN(n815) );
  XNOR2_X1 U911 ( .A(n815), .B(KEYINPUT104), .ZN(n817) );
  NAND2_X1 U912 ( .A1(n817), .A2(n816), .ZN(G188) );
  NOR2_X1 U913 ( .A1(n819), .A2(n818), .ZN(G325) );
  XNOR2_X1 U914 ( .A(KEYINPUT105), .B(G325), .ZN(G261) );
  INV_X1 U916 ( .A(G171), .ZN(G301) );
  NAND2_X1 U917 ( .A1(G100), .A2(n978), .ZN(n821) );
  NAND2_X1 U918 ( .A1(G136), .A2(n979), .ZN(n820) );
  NAND2_X1 U919 ( .A1(n821), .A2(n820), .ZN(n827) );
  NAND2_X1 U920 ( .A1(G124), .A2(n984), .ZN(n822) );
  XNOR2_X1 U921 ( .A(n822), .B(KEYINPUT44), .ZN(n825) );
  NAND2_X1 U922 ( .A1(G112), .A2(n977), .ZN(n823) );
  XOR2_X1 U923 ( .A(KEYINPUT111), .B(n823), .Z(n824) );
  NAND2_X1 U924 ( .A1(n825), .A2(n824), .ZN(n826) );
  NOR2_X1 U925 ( .A1(n827), .A2(n826), .ZN(G162) );
  XNOR2_X1 U926 ( .A(G2084), .B(G34), .ZN(n828) );
  XNOR2_X1 U927 ( .A(n828), .B(KEYINPUT54), .ZN(n847) );
  XNOR2_X1 U928 ( .A(G2090), .B(G35), .ZN(n844) );
  XNOR2_X1 U929 ( .A(n829), .B(G25), .ZN(n830) );
  NAND2_X1 U930 ( .A1(n830), .A2(G28), .ZN(n831) );
  XNOR2_X1 U931 ( .A(n831), .B(KEYINPUT117), .ZN(n835) );
  XNOR2_X1 U932 ( .A(G1996), .B(G32), .ZN(n833) );
  XNOR2_X1 U933 ( .A(G26), .B(G2067), .ZN(n832) );
  NOR2_X1 U934 ( .A1(n833), .A2(n832), .ZN(n834) );
  NAND2_X1 U935 ( .A1(n835), .A2(n834), .ZN(n841) );
  XOR2_X1 U936 ( .A(n836), .B(G27), .Z(n839) );
  XOR2_X1 U937 ( .A(KEYINPUT118), .B(G33), .Z(n837) );
  XNOR2_X1 U938 ( .A(G2072), .B(n837), .ZN(n838) );
  NAND2_X1 U939 ( .A1(n839), .A2(n838), .ZN(n840) );
  NOR2_X1 U940 ( .A1(n841), .A2(n840), .ZN(n842) );
  XNOR2_X1 U941 ( .A(KEYINPUT53), .B(n842), .ZN(n843) );
  NOR2_X1 U942 ( .A1(n844), .A2(n843), .ZN(n845) );
  XNOR2_X1 U943 ( .A(n845), .B(KEYINPUT119), .ZN(n846) );
  NOR2_X1 U944 ( .A1(n847), .A2(n846), .ZN(n848) );
  XOR2_X1 U945 ( .A(KEYINPUT55), .B(n848), .Z(n849) );
  XNOR2_X1 U946 ( .A(KEYINPUT120), .B(n849), .ZN(n850) );
  NOR2_X1 U947 ( .A1(G29), .A2(n850), .ZN(n905) );
  XNOR2_X1 U948 ( .A(n880), .B(G19), .ZN(n858) );
  XOR2_X1 U949 ( .A(G1981), .B(G6), .Z(n853) );
  XOR2_X1 U950 ( .A(G20), .B(KEYINPUT124), .Z(n851) );
  XNOR2_X1 U951 ( .A(G1956), .B(n851), .ZN(n852) );
  NAND2_X1 U952 ( .A1(n853), .A2(n852), .ZN(n856) );
  XOR2_X1 U953 ( .A(KEYINPUT59), .B(G1348), .Z(n854) );
  XNOR2_X1 U954 ( .A(G4), .B(n854), .ZN(n855) );
  NOR2_X1 U955 ( .A1(n856), .A2(n855), .ZN(n857) );
  NAND2_X1 U956 ( .A1(n858), .A2(n857), .ZN(n859) );
  XNOR2_X1 U957 ( .A(n859), .B(KEYINPUT60), .ZN(n871) );
  XOR2_X1 U958 ( .A(G1976), .B(G23), .Z(n863) );
  XNOR2_X1 U959 ( .A(G1971), .B(G22), .ZN(n861) );
  XNOR2_X1 U960 ( .A(G24), .B(G1986), .ZN(n860) );
  NOR2_X1 U961 ( .A1(n861), .A2(n860), .ZN(n862) );
  NAND2_X1 U962 ( .A1(n863), .A2(n862), .ZN(n865) );
  XNOR2_X1 U963 ( .A(KEYINPUT125), .B(KEYINPUT58), .ZN(n864) );
  XNOR2_X1 U964 ( .A(n865), .B(n864), .ZN(n869) );
  XNOR2_X1 U965 ( .A(G1966), .B(G21), .ZN(n867) );
  XNOR2_X1 U966 ( .A(G5), .B(G1961), .ZN(n866) );
  NOR2_X1 U967 ( .A1(n867), .A2(n866), .ZN(n868) );
  NAND2_X1 U968 ( .A1(n869), .A2(n868), .ZN(n870) );
  NOR2_X1 U969 ( .A1(n871), .A2(n870), .ZN(n872) );
  XOR2_X1 U970 ( .A(KEYINPUT61), .B(n872), .Z(n873) );
  NOR2_X1 U971 ( .A1(G16), .A2(n873), .ZN(n902) );
  XNOR2_X1 U972 ( .A(G1961), .B(KEYINPUT122), .ZN(n874) );
  XNOR2_X1 U973 ( .A(n874), .B(G301), .ZN(n878) );
  NAND2_X1 U974 ( .A1(n876), .A2(n875), .ZN(n877) );
  NOR2_X1 U975 ( .A1(n878), .A2(n877), .ZN(n895) );
  XNOR2_X1 U976 ( .A(n880), .B(n879), .ZN(n882) );
  NAND2_X1 U977 ( .A1(G1971), .A2(G303), .ZN(n881) );
  NAND2_X1 U978 ( .A1(n882), .A2(n881), .ZN(n884) );
  XNOR2_X1 U979 ( .A(G1348), .B(n963), .ZN(n883) );
  NOR2_X1 U980 ( .A1(n884), .A2(n883), .ZN(n887) );
  XNOR2_X1 U981 ( .A(n885), .B(G1956), .ZN(n886) );
  NAND2_X1 U982 ( .A1(n887), .A2(n886), .ZN(n893) );
  XNOR2_X1 U983 ( .A(G1966), .B(G168), .ZN(n889) );
  NAND2_X1 U984 ( .A1(n889), .A2(n888), .ZN(n890) );
  XNOR2_X1 U985 ( .A(n890), .B(KEYINPUT57), .ZN(n891) );
  XNOR2_X1 U986 ( .A(n891), .B(KEYINPUT121), .ZN(n892) );
  NOR2_X1 U987 ( .A1(n893), .A2(n892), .ZN(n894) );
  NAND2_X1 U988 ( .A1(n895), .A2(n894), .ZN(n896) );
  NOR2_X1 U989 ( .A1(n897), .A2(n896), .ZN(n899) );
  XOR2_X1 U990 ( .A(G16), .B(KEYINPUT56), .Z(n898) );
  NOR2_X1 U991 ( .A1(n899), .A2(n898), .ZN(n900) );
  XOR2_X1 U992 ( .A(KEYINPUT123), .B(n900), .Z(n901) );
  NOR2_X1 U993 ( .A1(n902), .A2(n901), .ZN(n903) );
  NAND2_X1 U994 ( .A1(G11), .A2(n903), .ZN(n904) );
  NOR2_X1 U995 ( .A1(n905), .A2(n904), .ZN(n906) );
  XNOR2_X1 U996 ( .A(n906), .B(KEYINPUT126), .ZN(n939) );
  XOR2_X1 U997 ( .A(G2090), .B(G162), .Z(n907) );
  NOR2_X1 U998 ( .A1(n908), .A2(n907), .ZN(n909) );
  XOR2_X1 U999 ( .A(KEYINPUT51), .B(n909), .Z(n916) );
  XOR2_X1 U1000 ( .A(G2084), .B(G160), .Z(n910) );
  NOR2_X1 U1001 ( .A1(n970), .A2(n910), .ZN(n911) );
  NAND2_X1 U1002 ( .A1(n912), .A2(n911), .ZN(n913) );
  NOR2_X1 U1003 ( .A1(n914), .A2(n913), .ZN(n915) );
  NAND2_X1 U1004 ( .A1(n916), .A2(n915), .ZN(n928) );
  NAND2_X1 U1005 ( .A1(G103), .A2(n978), .ZN(n918) );
  NAND2_X1 U1006 ( .A1(G139), .A2(n979), .ZN(n917) );
  NAND2_X1 U1007 ( .A1(n918), .A2(n917), .ZN(n923) );
  NAND2_X1 U1008 ( .A1(G115), .A2(n977), .ZN(n920) );
  NAND2_X1 U1009 ( .A1(G127), .A2(n984), .ZN(n919) );
  NAND2_X1 U1010 ( .A1(n920), .A2(n919), .ZN(n921) );
  XOR2_X1 U1011 ( .A(KEYINPUT47), .B(n921), .Z(n922) );
  NOR2_X1 U1012 ( .A1(n923), .A2(n922), .ZN(n969) );
  XOR2_X1 U1013 ( .A(G2072), .B(n969), .Z(n925) );
  XOR2_X1 U1014 ( .A(G164), .B(G2078), .Z(n924) );
  NOR2_X1 U1015 ( .A1(n925), .A2(n924), .ZN(n926) );
  XOR2_X1 U1016 ( .A(KEYINPUT50), .B(n926), .Z(n927) );
  NOR2_X1 U1017 ( .A1(n928), .A2(n927), .ZN(n933) );
  INV_X1 U1018 ( .A(n929), .ZN(n930) );
  NOR2_X1 U1019 ( .A1(n931), .A2(n930), .ZN(n932) );
  NAND2_X1 U1020 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1021 ( .A(KEYINPUT52), .B(n934), .ZN(n935) );
  XNOR2_X1 U1022 ( .A(KEYINPUT116), .B(n935), .ZN(n936) );
  OR2_X1 U1023 ( .A1(KEYINPUT55), .A2(n936), .ZN(n937) );
  NAND2_X1 U1024 ( .A1(G29), .A2(n937), .ZN(n938) );
  NAND2_X1 U1025 ( .A1(n939), .A2(n938), .ZN(n940) );
  XOR2_X1 U1026 ( .A(KEYINPUT62), .B(n940), .Z(G311) );
  XNOR2_X1 U1027 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1028 ( .A(G120), .ZN(G236) );
  INV_X1 U1029 ( .A(G96), .ZN(G221) );
  INV_X1 U1030 ( .A(G69), .ZN(G235) );
  XOR2_X1 U1031 ( .A(KEYINPUT106), .B(n941), .Z(G319) );
  XOR2_X1 U1032 ( .A(KEYINPUT107), .B(G2084), .Z(n943) );
  XNOR2_X1 U1033 ( .A(G2078), .B(G2067), .ZN(n942) );
  XNOR2_X1 U1034 ( .A(n943), .B(n942), .ZN(n944) );
  XOR2_X1 U1035 ( .A(n944), .B(G2678), .Z(n946) );
  XNOR2_X1 U1036 ( .A(G2072), .B(KEYINPUT42), .ZN(n945) );
  XNOR2_X1 U1037 ( .A(n946), .B(n945), .ZN(n950) );
  XOR2_X1 U1038 ( .A(G2100), .B(G2096), .Z(n948) );
  XNOR2_X1 U1039 ( .A(G2090), .B(KEYINPUT43), .ZN(n947) );
  XNOR2_X1 U1040 ( .A(n948), .B(n947), .ZN(n949) );
  XOR2_X1 U1041 ( .A(n950), .B(n949), .Z(G227) );
  XOR2_X1 U1042 ( .A(KEYINPUT41), .B(KEYINPUT110), .Z(n952) );
  XNOR2_X1 U1043 ( .A(G1956), .B(G1976), .ZN(n951) );
  XNOR2_X1 U1044 ( .A(n952), .B(n951), .ZN(n962) );
  XOR2_X1 U1045 ( .A(G2474), .B(KEYINPUT108), .Z(n954) );
  XNOR2_X1 U1046 ( .A(G1996), .B(KEYINPUT109), .ZN(n953) );
  XNOR2_X1 U1047 ( .A(n954), .B(n953), .ZN(n958) );
  XOR2_X1 U1048 ( .A(G1991), .B(G1981), .Z(n956) );
  XNOR2_X1 U1049 ( .A(G1961), .B(G1971), .ZN(n955) );
  XNOR2_X1 U1050 ( .A(n956), .B(n955), .ZN(n957) );
  XOR2_X1 U1051 ( .A(n958), .B(n957), .Z(n960) );
  XNOR2_X1 U1052 ( .A(G1966), .B(G1986), .ZN(n959) );
  XNOR2_X1 U1053 ( .A(n960), .B(n959), .ZN(n961) );
  XNOR2_X1 U1054 ( .A(n962), .B(n961), .ZN(G229) );
  XNOR2_X1 U1055 ( .A(G286), .B(n963), .ZN(n965) );
  XNOR2_X1 U1056 ( .A(n965), .B(n964), .ZN(n966) );
  XOR2_X1 U1057 ( .A(G301), .B(n966), .Z(n967) );
  NOR2_X1 U1058 ( .A1(G37), .A2(n967), .ZN(n968) );
  XOR2_X1 U1059 ( .A(KEYINPUT115), .B(n968), .Z(G397) );
  XNOR2_X1 U1060 ( .A(n969), .B(G162), .ZN(n971) );
  XNOR2_X1 U1061 ( .A(n971), .B(n970), .ZN(n973) );
  XOR2_X1 U1062 ( .A(n973), .B(n972), .Z(n976) );
  XNOR2_X1 U1063 ( .A(G164), .B(n974), .ZN(n975) );
  XNOR2_X1 U1064 ( .A(n976), .B(n975), .ZN(n992) );
  NAND2_X1 U1065 ( .A1(G118), .A2(n977), .ZN(n989) );
  XNOR2_X1 U1066 ( .A(KEYINPUT45), .B(KEYINPUT113), .ZN(n983) );
  NAND2_X1 U1067 ( .A1(G106), .A2(n978), .ZN(n981) );
  NAND2_X1 U1068 ( .A1(G142), .A2(n979), .ZN(n980) );
  NAND2_X1 U1069 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1070 ( .A(n983), .B(n982), .ZN(n987) );
  NAND2_X1 U1071 ( .A1(n984), .A2(G130), .ZN(n985) );
  XOR2_X1 U1072 ( .A(KEYINPUT112), .B(n985), .Z(n986) );
  NOR2_X1 U1073 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1074 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1075 ( .A(n990), .B(KEYINPUT48), .ZN(n991) );
  XOR2_X1 U1076 ( .A(n992), .B(n991), .Z(n994) );
  XNOR2_X1 U1077 ( .A(G160), .B(KEYINPUT46), .ZN(n993) );
  XNOR2_X1 U1078 ( .A(n994), .B(n993), .ZN(n996) );
  XOR2_X1 U1079 ( .A(n996), .B(n995), .Z(n997) );
  NOR2_X1 U1080 ( .A1(G37), .A2(n997), .ZN(n998) );
  XNOR2_X1 U1081 ( .A(KEYINPUT114), .B(n998), .ZN(G395) );
  XNOR2_X1 U1082 ( .A(G1341), .B(G2443), .ZN(n1008) );
  XOR2_X1 U1083 ( .A(G2451), .B(G2446), .Z(n1000) );
  XNOR2_X1 U1084 ( .A(G1348), .B(KEYINPUT102), .ZN(n999) );
  XNOR2_X1 U1085 ( .A(n1000), .B(n999), .ZN(n1004) );
  XOR2_X1 U1086 ( .A(G2438), .B(KEYINPUT103), .Z(n1002) );
  XNOR2_X1 U1087 ( .A(G2454), .B(G2435), .ZN(n1001) );
  XNOR2_X1 U1088 ( .A(n1002), .B(n1001), .ZN(n1003) );
  XOR2_X1 U1089 ( .A(n1004), .B(n1003), .Z(n1006) );
  XNOR2_X1 U1090 ( .A(G2430), .B(G2427), .ZN(n1005) );
  XNOR2_X1 U1091 ( .A(n1006), .B(n1005), .ZN(n1007) );
  XNOR2_X1 U1092 ( .A(n1008), .B(n1007), .ZN(n1009) );
  NAND2_X1 U1093 ( .A1(n1009), .A2(G14), .ZN(n1015) );
  NAND2_X1 U1094 ( .A1(n1015), .A2(G319), .ZN(n1012) );
  NOR2_X1 U1095 ( .A1(G227), .A2(G229), .ZN(n1010) );
  XNOR2_X1 U1096 ( .A(KEYINPUT49), .B(n1010), .ZN(n1011) );
  NOR2_X1 U1097 ( .A1(n1012), .A2(n1011), .ZN(n1014) );
  NOR2_X1 U1098 ( .A1(G397), .A2(G395), .ZN(n1013) );
  NAND2_X1 U1099 ( .A1(n1014), .A2(n1013), .ZN(G225) );
  INV_X1 U1100 ( .A(G225), .ZN(G308) );
  INV_X1 U1101 ( .A(G108), .ZN(G238) );
  INV_X1 U1102 ( .A(n1015), .ZN(G401) );
endmodule

