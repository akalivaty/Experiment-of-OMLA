

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737;

  AND2_X1 U369 ( .A1(n385), .A2(n572), .ZN(n629) );
  INV_X2 U370 ( .A(G953), .ZN(n729) );
  AND2_X2 U371 ( .A1(n377), .A2(n386), .ZN(n357) );
  NOR2_X2 U372 ( .A1(n735), .A2(n736), .ZN(n354) );
  XNOR2_X2 U373 ( .A(G143), .B(KEYINPUT64), .ZN(n435) );
  NOR2_X2 U374 ( .A1(n558), .A2(n559), .ZN(n392) );
  XNOR2_X2 U375 ( .A(n715), .B(n374), .ZN(n609) );
  XNOR2_X2 U376 ( .A(n429), .B(G104), .ZN(n428) );
  XNOR2_X2 U377 ( .A(n511), .B(n455), .ZN(n379) );
  XNOR2_X2 U378 ( .A(n562), .B(KEYINPUT35), .ZN(n733) );
  INV_X1 U379 ( .A(KEYINPUT75), .ZN(n391) );
  INV_X1 U380 ( .A(G146), .ZN(n394) );
  INV_X1 U381 ( .A(G134), .ZN(n432) );
  AND2_X1 U382 ( .A1(n413), .A2(n381), .ZN(n598) );
  OR2_X1 U383 ( .A1(n542), .A2(n543), .ZN(n386) );
  XNOR2_X1 U384 ( .A(n409), .B(n408), .ZN(n735) );
  XNOR2_X1 U385 ( .A(n368), .B(n367), .ZN(n736) );
  XNOR2_X1 U386 ( .A(n571), .B(n570), .ZN(n734) );
  XNOR2_X1 U387 ( .A(n380), .B(KEYINPUT41), .ZN(n675) );
  XNOR2_X1 U388 ( .A(n576), .B(KEYINPUT86), .ZN(n543) );
  XNOR2_X1 U389 ( .A(n662), .B(n388), .ZN(n378) );
  XNOR2_X1 U390 ( .A(n618), .B(KEYINPUT85), .ZN(n619) );
  NAND2_X2 U391 ( .A1(n421), .A2(n417), .ZN(n584) );
  XNOR2_X1 U392 ( .A(n460), .B(n434), .ZN(n452) );
  XNOR2_X1 U393 ( .A(n471), .B(n431), .ZN(n430) );
  XNOR2_X1 U394 ( .A(n435), .B(G128), .ZN(n460) );
  XNOR2_X1 U395 ( .A(n432), .B(KEYINPUT66), .ZN(n431) );
  AND2_X1 U396 ( .A1(n687), .A2(n600), .ZN(n347) );
  AND2_X2 U397 ( .A1(n687), .A2(n600), .ZN(n705) );
  XNOR2_X1 U398 ( .A(n354), .B(KEYINPUT46), .ZN(n377) );
  XNOR2_X1 U399 ( .A(n364), .B(n350), .ZN(n535) );
  OR2_X1 U400 ( .A1(n601), .A2(G902), .ZN(n364) );
  XNOR2_X1 U401 ( .A(n499), .B(KEYINPUT25), .ZN(n398) );
  XNOR2_X1 U402 ( .A(n550), .B(n438), .ZN(n655) );
  XNOR2_X1 U403 ( .A(n551), .B(KEYINPUT71), .ZN(n438) );
  INV_X1 U404 ( .A(KEYINPUT33), .ZN(n551) );
  XNOR2_X1 U405 ( .A(n425), .B(KEYINPUT39), .ZN(n545) );
  AND2_X1 U406 ( .A1(n378), .A2(n387), .ZN(n512) );
  NOR2_X1 U407 ( .A1(n543), .A2(n378), .ZN(n569) );
  OR2_X1 U408 ( .A1(n617), .A2(G902), .ZN(n393) );
  INV_X1 U409 ( .A(n633), .ZN(n401) );
  XNOR2_X1 U410 ( .A(KEYINPUT11), .B(KEYINPUT96), .ZN(n365) );
  NOR2_X1 U411 ( .A1(G953), .A2(G237), .ZN(n502) );
  NAND2_X1 U412 ( .A1(n361), .A2(n358), .ZN(n588) );
  AND2_X1 U413 ( .A1(n363), .A2(n362), .ZN(n361) );
  NAND2_X1 U414 ( .A1(n360), .A2(KEYINPUT78), .ZN(n359) );
  XNOR2_X1 U415 ( .A(n433), .B(KEYINPUT65), .ZN(n471) );
  INV_X1 U416 ( .A(G131), .ZN(n433) );
  OR2_X1 U417 ( .A1(G237), .A2(G902), .ZN(n514) );
  XNOR2_X1 U418 ( .A(KEYINPUT79), .B(KEYINPUT8), .ZN(n461) );
  INV_X1 U419 ( .A(KEYINPUT48), .ZN(n376) );
  XNOR2_X1 U420 ( .A(n399), .B(KEYINPUT73), .ZN(n356) );
  INV_X1 U421 ( .A(G902), .ZN(n419) );
  XNOR2_X1 U422 ( .A(G134), .B(G122), .ZN(n457) );
  XNOR2_X1 U423 ( .A(n465), .B(n407), .ZN(n406) );
  INV_X1 U424 ( .A(KEYINPUT99), .ZN(n407) );
  XNOR2_X1 U425 ( .A(G116), .B(G107), .ZN(n465) );
  XNOR2_X1 U426 ( .A(n476), .B(n349), .ZN(n601) );
  XNOR2_X1 U427 ( .A(G113), .B(G143), .ZN(n467) );
  XNOR2_X1 U428 ( .A(n640), .B(n404), .ZN(n544) );
  INV_X1 U429 ( .A(KEYINPUT101), .ZN(n404) );
  NAND2_X1 U430 ( .A1(n655), .A2(n583), .ZN(n437) );
  AND2_X1 U431 ( .A1(n520), .A2(n369), .ZN(n538) );
  XNOR2_X1 U432 ( .A(n371), .B(n370), .ZN(n369) );
  AND2_X1 U433 ( .A1(n416), .A2(n584), .ZN(n519) );
  XNOR2_X1 U434 ( .A(G478), .B(n466), .ZN(n536) );
  NOR2_X1 U435 ( .A1(n703), .A2(G902), .ZN(n466) );
  INV_X1 U436 ( .A(n535), .ZN(n522) );
  INV_X1 U437 ( .A(KEYINPUT6), .ZN(n388) );
  NAND2_X1 U438 ( .A1(n544), .A2(n403), .ZN(n363) );
  NAND2_X1 U439 ( .A1(n636), .A2(n403), .ZN(n362) );
  XNOR2_X1 U440 ( .A(G146), .B(G125), .ZN(n469) );
  NAND2_X1 U441 ( .A1(n402), .A2(n400), .ZN(n399) );
  AND2_X1 U442 ( .A1(n531), .A2(n401), .ZN(n400) );
  NOR2_X1 U443 ( .A1(n588), .A2(KEYINPUT47), .ZN(n529) );
  XOR2_X1 U444 ( .A(KEYINPUT74), .B(KEYINPUT94), .Z(n504) );
  XNOR2_X1 U445 ( .A(n447), .B(n415), .ZN(n508) );
  INV_X1 U446 ( .A(KEYINPUT3), .ZN(n415) );
  XNOR2_X1 U447 ( .A(n469), .B(KEYINPUT10), .ZN(n488) );
  XNOR2_X1 U448 ( .A(n472), .B(n365), .ZN(n439) );
  XNOR2_X1 U449 ( .A(G140), .B(KEYINPUT12), .ZN(n472) );
  XOR2_X1 U450 ( .A(G122), .B(G104), .Z(n468) );
  INV_X1 U451 ( .A(KEYINPUT103), .ZN(n397) );
  XOR2_X1 U452 ( .A(G137), .B(G140), .Z(n489) );
  XOR2_X1 U453 ( .A(KEYINPUT17), .B(KEYINPUT89), .Z(n441) );
  XNOR2_X1 U454 ( .A(n444), .B(KEYINPUT18), .ZN(n414) );
  INV_X1 U455 ( .A(KEYINPUT4), .ZN(n434) );
  INV_X1 U456 ( .A(KEYINPUT104), .ZN(n548) );
  XNOR2_X1 U457 ( .A(n533), .B(n534), .ZN(n651) );
  XNOR2_X1 U458 ( .A(n540), .B(KEYINPUT38), .ZN(n410) );
  INV_X1 U459 ( .A(n524), .ZN(n387) );
  AND2_X1 U460 ( .A1(n568), .A2(n424), .ZN(n416) );
  INV_X1 U461 ( .A(n518), .ZN(n424) );
  INV_X1 U462 ( .A(KEYINPUT30), .ZN(n370) );
  XOR2_X1 U463 ( .A(KEYINPUT24), .B(G110), .Z(n491) );
  XNOR2_X1 U464 ( .A(G119), .B(G128), .ZN(n490) );
  XNOR2_X1 U465 ( .A(KEYINPUT70), .B(KEYINPUT23), .ZN(n494) );
  NOR2_X1 U466 ( .A1(n646), .A2(n412), .ZN(n411) );
  INV_X1 U467 ( .A(n645), .ZN(n412) );
  XNOR2_X1 U468 ( .A(G107), .B(G110), .ZN(n427) );
  INV_X1 U469 ( .A(n489), .ZN(n426) );
  INV_X1 U470 ( .A(KEYINPUT19), .ZN(n389) );
  OR2_X1 U471 ( .A1(n379), .A2(n418), .ZN(n417) );
  AND2_X1 U472 ( .A1(n423), .A2(n422), .ZN(n421) );
  NAND2_X1 U473 ( .A1(n420), .A2(n419), .ZN(n418) );
  NOR2_X1 U474 ( .A1(n657), .A2(n658), .ZN(n664) );
  XNOR2_X1 U475 ( .A(n405), .B(n464), .ZN(n703) );
  XNOR2_X1 U476 ( .A(n463), .B(n406), .ZN(n405) );
  XNOR2_X1 U477 ( .A(n601), .B(KEYINPUT59), .ZN(n602) );
  XNOR2_X1 U478 ( .A(n611), .B(n610), .ZN(n612) );
  INV_X1 U479 ( .A(KEYINPUT42), .ZN(n408) );
  INV_X1 U480 ( .A(KEYINPUT40), .ZN(n367) );
  XNOR2_X1 U481 ( .A(n437), .B(n436), .ZN(n561) );
  INV_X1 U482 ( .A(KEYINPUT34), .ZN(n436) );
  AND2_X1 U483 ( .A1(n569), .A2(n658), .ZN(n384) );
  XNOR2_X1 U484 ( .A(n523), .B(KEYINPUT100), .ZN(n640) );
  INV_X1 U485 ( .A(n378), .ZN(n372) );
  XNOR2_X1 U486 ( .A(n700), .B(n699), .ZN(n701) );
  XNOR2_X1 U487 ( .A(KEYINPUT15), .B(G902), .ZN(n348) );
  XOR2_X1 U488 ( .A(n468), .B(n467), .Z(n349) );
  XOR2_X1 U489 ( .A(n478), .B(n477), .Z(n350) );
  XNOR2_X1 U490 ( .A(n450), .B(n449), .ZN(n351) );
  XNOR2_X1 U491 ( .A(n500), .B(n398), .ZN(n568) );
  INV_X1 U492 ( .A(n381), .ZN(n646) );
  XOR2_X1 U493 ( .A(KEYINPUT22), .B(KEYINPUT72), .Z(n352) );
  INV_X1 U494 ( .A(KEYINPUT78), .ZN(n403) );
  XNOR2_X2 U495 ( .A(n353), .B(n391), .ZN(n687) );
  NAND2_X1 U496 ( .A1(n599), .A2(n598), .ZN(n353) );
  NAND2_X1 U497 ( .A1(n651), .A2(n649), .ZN(n380) );
  XNOR2_X2 U498 ( .A(n355), .B(n376), .ZN(n413) );
  NAND2_X1 U499 ( .A1(n357), .A2(n356), .ZN(n355) );
  OR2_X1 U500 ( .A1(n544), .A2(n636), .ZN(n652) );
  OR2_X1 U501 ( .A1(n544), .A2(n359), .ZN(n358) );
  INV_X1 U502 ( .A(n636), .ZN(n360) );
  AND2_X1 U503 ( .A1(n366), .A2(n658), .ZN(n385) );
  NAND2_X1 U504 ( .A1(n384), .A2(n366), .ZN(n571) );
  AND2_X1 U505 ( .A1(n366), .A2(n372), .ZN(n577) );
  XNOR2_X2 U506 ( .A(n567), .B(n352), .ZN(n366) );
  NAND2_X1 U507 ( .A1(n545), .A2(n636), .ZN(n368) );
  NAND2_X1 U508 ( .A1(n662), .A2(n647), .ZN(n371) );
  XNOR2_X2 U509 ( .A(n373), .B(n508), .ZN(n715) );
  XNOR2_X2 U510 ( .A(n383), .B(n448), .ZN(n373) );
  XNOR2_X1 U511 ( .A(n452), .B(n375), .ZN(n374) );
  XNOR2_X1 U512 ( .A(n414), .B(n443), .ZN(n375) );
  XNOR2_X2 U513 ( .A(n428), .B(n427), .ZN(n383) );
  NAND2_X1 U514 ( .A1(n379), .A2(n456), .ZN(n423) );
  XNOR2_X1 U515 ( .A(n379), .B(n440), .ZN(n699) );
  NAND2_X1 U516 ( .A1(n675), .A2(n537), .ZN(n409) );
  INV_X1 U517 ( .A(n382), .ZN(n540) );
  NAND2_X1 U518 ( .A1(n382), .A2(n647), .ZN(n390) );
  XNOR2_X2 U519 ( .A(n451), .B(n351), .ZN(n382) );
  OR2_X1 U520 ( .A1(n517), .A2(n382), .ZN(n381) );
  XNOR2_X1 U521 ( .A(n383), .B(n426), .ZN(n454) );
  XNOR2_X1 U522 ( .A(n390), .B(n389), .ZN(n558) );
  INV_X1 U523 ( .A(n386), .ZN(n643) );
  XNOR2_X1 U524 ( .A(n392), .B(KEYINPUT0), .ZN(n566) );
  NAND2_X1 U525 ( .A1(n705), .A2(G210), .ZN(n613) );
  XNOR2_X2 U526 ( .A(n393), .B(G472), .ZN(n662) );
  XNOR2_X2 U527 ( .A(n721), .B(n394), .ZN(n511) );
  XNOR2_X2 U528 ( .A(n452), .B(n430), .ZN(n721) );
  XNOR2_X1 U529 ( .A(n395), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U530 ( .A1(n621), .A2(n696), .ZN(n395) );
  XNOR2_X1 U531 ( .A(n497), .B(n496), .ZN(n707) );
  NAND2_X1 U532 ( .A1(n591), .A2(n396), .ZN(n593) );
  XNOR2_X1 U533 ( .A(n590), .B(n397), .ZN(n396) );
  NAND2_X1 U534 ( .A1(n529), .A2(n634), .ZN(n402) );
  NAND2_X1 U535 ( .A1(n410), .A2(n647), .ZN(n533) );
  NOR2_X1 U536 ( .A1(n410), .A2(n647), .ZN(n648) );
  NAND2_X1 U537 ( .A1(n538), .A2(n410), .ZN(n425) );
  NAND2_X2 U538 ( .A1(n413), .A2(n411), .ZN(n727) );
  NOR2_X2 U539 ( .A1(n689), .A2(n597), .ZN(n599) );
  INV_X1 U540 ( .A(n456), .ZN(n420) );
  NAND2_X1 U541 ( .A1(n456), .A2(G902), .ZN(n422) );
  INV_X1 U542 ( .A(n568), .ZN(n658) );
  XNOR2_X2 U543 ( .A(G101), .B(KEYINPUT88), .ZN(n429) );
  NAND2_X1 U544 ( .A1(n547), .A2(n664), .ZN(n579) );
  XNOR2_X2 U545 ( .A(n584), .B(KEYINPUT1), .ZN(n547) );
  XNOR2_X1 U546 ( .A(n613), .B(n612), .ZN(n614) );
  XNOR2_X1 U547 ( .A(n603), .B(n602), .ZN(n605) );
  XNOR2_X1 U548 ( .A(n579), .B(n548), .ZN(n549) );
  XOR2_X1 U549 ( .A(n698), .B(n697), .Z(n440) );
  INV_X1 U550 ( .A(n469), .ZN(n442) );
  XNOR2_X1 U551 ( .A(n442), .B(n441), .ZN(n443) );
  INV_X1 U552 ( .A(G475), .ZN(n477) );
  XNOR2_X1 U553 ( .A(n475), .B(n474), .ZN(n476) );
  INV_X1 U554 ( .A(KEYINPUT90), .ZN(n449) );
  XNOR2_X1 U555 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U556 ( .A(n620), .B(n619), .ZN(n621) );
  INV_X1 U557 ( .A(KEYINPUT122), .ZN(n606) );
  XNOR2_X1 U558 ( .A(n606), .B(KEYINPUT60), .ZN(n607) );
  AND2_X1 U559 ( .A1(G224), .A2(n729), .ZN(n444) );
  XOR2_X1 U560 ( .A(G122), .B(KEYINPUT16), .Z(n448) );
  XOR2_X1 U561 ( .A(KEYINPUT69), .B(G119), .Z(n446) );
  XNOR2_X1 U562 ( .A(G116), .B(G113), .ZN(n445) );
  XNOR2_X1 U563 ( .A(n446), .B(n445), .ZN(n447) );
  NAND2_X1 U564 ( .A1(n609), .A2(n348), .ZN(n451) );
  NAND2_X1 U565 ( .A1(G210), .A2(n514), .ZN(n450) );
  NAND2_X1 U566 ( .A1(G227), .A2(n729), .ZN(n453) );
  XNOR2_X1 U567 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U568 ( .A(KEYINPUT68), .B(G469), .ZN(n456) );
  INV_X1 U569 ( .A(n547), .ZN(n576) );
  INV_X1 U570 ( .A(n576), .ZN(n665) );
  XOR2_X1 U571 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n458) );
  XNOR2_X1 U572 ( .A(n458), .B(n457), .ZN(n459) );
  XOR2_X1 U573 ( .A(n460), .B(n459), .Z(n464) );
  NAND2_X1 U574 ( .A1(n729), .A2(G234), .ZN(n462) );
  XNOR2_X1 U575 ( .A(n462), .B(n461), .ZN(n493) );
  NAND2_X1 U576 ( .A1(G217), .A2(n493), .ZN(n463) );
  NAND2_X1 U577 ( .A1(G214), .A2(n502), .ZN(n470) );
  XNOR2_X1 U578 ( .A(n470), .B(n488), .ZN(n475) );
  XNOR2_X1 U579 ( .A(n471), .B(KEYINPUT97), .ZN(n473) );
  XNOR2_X1 U580 ( .A(n473), .B(n439), .ZN(n474) );
  XNOR2_X1 U581 ( .A(KEYINPUT98), .B(KEYINPUT13), .ZN(n478) );
  AND2_X1 U582 ( .A1(n536), .A2(n522), .ZN(n636) );
  NAND2_X1 U583 ( .A1(G234), .A2(G237), .ZN(n479) );
  XNOR2_X1 U584 ( .A(n479), .B(KEYINPUT14), .ZN(n481) );
  NAND2_X1 U585 ( .A1(G902), .A2(n481), .ZN(n553) );
  NOR2_X1 U586 ( .A1(G900), .A2(n553), .ZN(n480) );
  NAND2_X1 U587 ( .A1(G953), .A2(n480), .ZN(n483) );
  NAND2_X1 U588 ( .A1(G952), .A2(n481), .ZN(n482) );
  XNOR2_X1 U589 ( .A(KEYINPUT91), .B(n482), .ZN(n681) );
  NAND2_X1 U590 ( .A1(n681), .A2(n729), .ZN(n552) );
  NAND2_X1 U591 ( .A1(n483), .A2(n552), .ZN(n487) );
  NAND2_X1 U592 ( .A1(G234), .A2(n348), .ZN(n484) );
  XNOR2_X1 U593 ( .A(KEYINPUT20), .B(n484), .ZN(n498) );
  NAND2_X1 U594 ( .A1(G221), .A2(n498), .ZN(n485) );
  XNOR2_X1 U595 ( .A(n485), .B(KEYINPUT21), .ZN(n486) );
  XNOR2_X1 U596 ( .A(KEYINPUT93), .B(n486), .ZN(n546) );
  NAND2_X1 U597 ( .A1(n487), .A2(n546), .ZN(n518) );
  XNOR2_X1 U598 ( .A(KEYINPUT67), .B(n518), .ZN(n501) );
  XNOR2_X1 U599 ( .A(n489), .B(n488), .ZN(n723) );
  XNOR2_X1 U600 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U601 ( .A(n723), .B(n492), .ZN(n497) );
  NAND2_X1 U602 ( .A1(n493), .A2(G221), .ZN(n495) );
  NOR2_X1 U603 ( .A1(G902), .A2(n707), .ZN(n500) );
  NAND2_X1 U604 ( .A1(n498), .A2(G217), .ZN(n499) );
  NAND2_X1 U605 ( .A1(n501), .A2(n658), .ZN(n524) );
  NAND2_X1 U606 ( .A1(n502), .A2(G210), .ZN(n503) );
  XNOR2_X1 U607 ( .A(n504), .B(n503), .ZN(n505) );
  XOR2_X1 U608 ( .A(n505), .B(G137), .Z(n507) );
  XNOR2_X1 U609 ( .A(G101), .B(KEYINPUT5), .ZN(n506) );
  XNOR2_X1 U610 ( .A(n507), .B(n506), .ZN(n509) );
  XNOR2_X1 U611 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U612 ( .A(n511), .B(n510), .ZN(n617) );
  NAND2_X1 U613 ( .A1(n636), .A2(n512), .ZN(n513) );
  XNOR2_X1 U614 ( .A(n513), .B(KEYINPUT105), .ZN(n515) );
  NAND2_X1 U615 ( .A1(G214), .A2(n514), .ZN(n647) );
  NAND2_X1 U616 ( .A1(n515), .A2(n647), .ZN(n539) );
  NOR2_X1 U617 ( .A1(n665), .A2(n539), .ZN(n516) );
  XNOR2_X1 U618 ( .A(n516), .B(KEYINPUT43), .ZN(n517) );
  XNOR2_X1 U619 ( .A(KEYINPUT76), .B(n519), .ZN(n520) );
  NOR2_X1 U620 ( .A1(n535), .A2(n536), .ZN(n560) );
  NAND2_X1 U621 ( .A1(n538), .A2(n560), .ZN(n521) );
  NOR2_X1 U622 ( .A1(n540), .A2(n521), .ZN(n633) );
  NOR2_X1 U623 ( .A1(n522), .A2(n536), .ZN(n523) );
  INV_X1 U624 ( .A(n662), .ZN(n580) );
  OR2_X1 U625 ( .A1(n580), .A2(n524), .ZN(n526) );
  XNOR2_X1 U626 ( .A(KEYINPUT107), .B(KEYINPUT28), .ZN(n525) );
  XNOR2_X1 U627 ( .A(n526), .B(n525), .ZN(n528) );
  XNOR2_X1 U628 ( .A(n584), .B(KEYINPUT106), .ZN(n527) );
  NAND2_X1 U629 ( .A1(n528), .A2(n527), .ZN(n532) );
  NOR2_X1 U630 ( .A1(n532), .A2(n558), .ZN(n634) );
  NAND2_X1 U631 ( .A1(n652), .A2(n634), .ZN(n530) );
  NAND2_X1 U632 ( .A1(n530), .A2(KEYINPUT47), .ZN(n531) );
  INV_X1 U633 ( .A(n532), .ZN(n537) );
  INV_X1 U634 ( .A(KEYINPUT108), .ZN(n534) );
  NAND2_X1 U635 ( .A1(n536), .A2(n535), .ZN(n563) );
  INV_X1 U636 ( .A(n563), .ZN(n649) );
  NOR2_X1 U637 ( .A1(n540), .A2(n539), .ZN(n541) );
  XOR2_X1 U638 ( .A(KEYINPUT36), .B(n541), .Z(n542) );
  NAND2_X1 U639 ( .A1(n545), .A2(n544), .ZN(n645) );
  INV_X1 U640 ( .A(n546), .ZN(n657) );
  NAND2_X1 U641 ( .A1(n549), .A2(n378), .ZN(n550) );
  INV_X1 U642 ( .A(n552), .ZN(n557) );
  INV_X1 U643 ( .A(n553), .ZN(n554) );
  NOR2_X1 U644 ( .A1(G898), .A2(n729), .ZN(n717) );
  NAND2_X1 U645 ( .A1(n554), .A2(n717), .ZN(n555) );
  XOR2_X1 U646 ( .A(KEYINPUT92), .B(n555), .Z(n556) );
  NOR2_X1 U647 ( .A1(n557), .A2(n556), .ZN(n559) );
  BUF_X1 U648 ( .A(n566), .Z(n583) );
  NAND2_X1 U649 ( .A1(n561), .A2(n560), .ZN(n562) );
  NOR2_X1 U650 ( .A1(n657), .A2(n563), .ZN(n564) );
  XNOR2_X1 U651 ( .A(n564), .B(KEYINPUT102), .ZN(n565) );
  NAND2_X1 U652 ( .A1(n566), .A2(n565), .ZN(n567) );
  INV_X1 U653 ( .A(KEYINPUT32), .ZN(n570) );
  AND2_X1 U654 ( .A1(n576), .A2(n580), .ZN(n572) );
  NOR2_X1 U655 ( .A1(n734), .A2(n629), .ZN(n573) );
  XNOR2_X1 U656 ( .A(n573), .B(KEYINPUT83), .ZN(n574) );
  NOR2_X2 U657 ( .A1(n733), .A2(n574), .ZN(n575) );
  XNOR2_X1 U658 ( .A(n575), .B(KEYINPUT44), .ZN(n591) );
  NAND2_X1 U659 ( .A1(n577), .A2(n576), .ZN(n578) );
  NOR2_X1 U660 ( .A1(n658), .A2(n578), .ZN(n622) );
  NOR2_X1 U661 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U662 ( .A(KEYINPUT95), .B(n581), .Z(n672) );
  NAND2_X1 U663 ( .A1(n583), .A2(n672), .ZN(n582) );
  XNOR2_X1 U664 ( .A(n582), .B(KEYINPUT31), .ZN(n639) );
  AND2_X1 U665 ( .A1(n584), .A2(n583), .ZN(n585) );
  NAND2_X1 U666 ( .A1(n664), .A2(n585), .ZN(n586) );
  NOR2_X1 U667 ( .A1(n662), .A2(n586), .ZN(n625) );
  NOR2_X1 U668 ( .A1(n639), .A2(n625), .ZN(n587) );
  NOR2_X1 U669 ( .A1(n588), .A2(n587), .ZN(n589) );
  NOR2_X1 U670 ( .A1(n622), .A2(n589), .ZN(n590) );
  XNOR2_X1 U671 ( .A(KEYINPUT45), .B(KEYINPUT81), .ZN(n592) );
  XNOR2_X2 U672 ( .A(n593), .B(n592), .ZN(n689) );
  NOR2_X1 U673 ( .A1(n727), .A2(n689), .ZN(n594) );
  NOR2_X1 U674 ( .A1(KEYINPUT2), .A2(n594), .ZN(n595) );
  NOR2_X2 U675 ( .A1(n595), .A2(n348), .ZN(n600) );
  NAND2_X1 U676 ( .A1(KEYINPUT2), .A2(n645), .ZN(n596) );
  XOR2_X1 U677 ( .A(KEYINPUT77), .B(n596), .Z(n597) );
  NAND2_X1 U678 ( .A1(n705), .A2(G475), .ZN(n603) );
  NOR2_X1 U679 ( .A1(G952), .A2(n729), .ZN(n604) );
  XNOR2_X1 U680 ( .A(KEYINPUT87), .B(n604), .ZN(n696) );
  NAND2_X1 U681 ( .A1(n605), .A2(n696), .ZN(n608) );
  XNOR2_X1 U682 ( .A(n608), .B(n607), .ZN(G60) );
  XNOR2_X1 U683 ( .A(n609), .B(KEYINPUT54), .ZN(n611) );
  XOR2_X1 U684 ( .A(KEYINPUT55), .B(KEYINPUT84), .Z(n610) );
  NAND2_X1 U685 ( .A1(n614), .A2(n696), .ZN(n616) );
  XOR2_X1 U686 ( .A(KEYINPUT82), .B(KEYINPUT56), .Z(n615) );
  XNOR2_X1 U687 ( .A(n616), .B(n615), .ZN(G51) );
  NAND2_X1 U688 ( .A1(n705), .A2(G472), .ZN(n620) );
  XNOR2_X1 U689 ( .A(KEYINPUT62), .B(n617), .ZN(n618) );
  XNOR2_X1 U690 ( .A(G101), .B(n622), .ZN(n623) );
  XNOR2_X1 U691 ( .A(n623), .B(KEYINPUT109), .ZN(G3) );
  NAND2_X1 U692 ( .A1(n625), .A2(n636), .ZN(n624) );
  XNOR2_X1 U693 ( .A(n624), .B(G104), .ZN(G6) );
  XOR2_X1 U694 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n627) );
  NAND2_X1 U695 ( .A1(n625), .A2(n640), .ZN(n626) );
  XNOR2_X1 U696 ( .A(n627), .B(n626), .ZN(n628) );
  XNOR2_X1 U697 ( .A(G107), .B(n628), .ZN(G9) );
  XOR2_X1 U698 ( .A(G110), .B(n629), .Z(G12) );
  XOR2_X1 U699 ( .A(KEYINPUT110), .B(KEYINPUT29), .Z(n631) );
  NAND2_X1 U700 ( .A1(n634), .A2(n640), .ZN(n630) );
  XNOR2_X1 U701 ( .A(n631), .B(n630), .ZN(n632) );
  XNOR2_X1 U702 ( .A(G128), .B(n632), .ZN(G30) );
  XOR2_X1 U703 ( .A(G143), .B(n633), .Z(G45) );
  NAND2_X1 U704 ( .A1(n634), .A2(n636), .ZN(n635) );
  XNOR2_X1 U705 ( .A(n635), .B(G146), .ZN(G48) );
  XOR2_X1 U706 ( .A(G113), .B(KEYINPUT111), .Z(n638) );
  NAND2_X1 U707 ( .A1(n639), .A2(n636), .ZN(n637) );
  XNOR2_X1 U708 ( .A(n638), .B(n637), .ZN(G15) );
  NAND2_X1 U709 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U710 ( .A(n641), .B(KEYINPUT112), .ZN(n642) );
  XNOR2_X1 U711 ( .A(G116), .B(n642), .ZN(G18) );
  XNOR2_X1 U712 ( .A(G125), .B(n643), .ZN(n644) );
  XNOR2_X1 U713 ( .A(n644), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U714 ( .A(G134), .B(n645), .ZN(G36) );
  XOR2_X1 U715 ( .A(G140), .B(n646), .Z(G42) );
  NAND2_X1 U716 ( .A1(n655), .A2(n675), .ZN(n684) );
  XOR2_X1 U717 ( .A(KEYINPUT118), .B(n648), .Z(n650) );
  NAND2_X1 U718 ( .A1(n650), .A2(n649), .ZN(n654) );
  NAND2_X1 U719 ( .A1(n652), .A2(n651), .ZN(n653) );
  NAND2_X1 U720 ( .A1(n654), .A2(n653), .ZN(n656) );
  NAND2_X1 U721 ( .A1(n656), .A2(n655), .ZN(n678) );
  XOR2_X1 U722 ( .A(KEYINPUT49), .B(KEYINPUT113), .Z(n660) );
  NAND2_X1 U723 ( .A1(n658), .A2(n657), .ZN(n659) );
  XNOR2_X1 U724 ( .A(n660), .B(n659), .ZN(n661) );
  NOR2_X1 U725 ( .A1(n662), .A2(n661), .ZN(n663) );
  XOR2_X1 U726 ( .A(KEYINPUT114), .B(n663), .Z(n670) );
  XNOR2_X1 U727 ( .A(KEYINPUT50), .B(KEYINPUT116), .ZN(n667) );
  NOR2_X1 U728 ( .A1(n665), .A2(n664), .ZN(n666) );
  XNOR2_X1 U729 ( .A(n667), .B(n666), .ZN(n668) );
  XOR2_X1 U730 ( .A(KEYINPUT115), .B(n668), .Z(n669) );
  NOR2_X1 U731 ( .A1(n670), .A2(n669), .ZN(n671) );
  NOR2_X1 U732 ( .A1(n672), .A2(n671), .ZN(n673) );
  XOR2_X1 U733 ( .A(KEYINPUT51), .B(n673), .Z(n674) );
  XNOR2_X1 U734 ( .A(KEYINPUT117), .B(n674), .ZN(n676) );
  NAND2_X1 U735 ( .A1(n676), .A2(n675), .ZN(n677) );
  NAND2_X1 U736 ( .A1(n678), .A2(n677), .ZN(n679) );
  XNOR2_X1 U737 ( .A(n679), .B(KEYINPUT52), .ZN(n680) );
  XOR2_X1 U738 ( .A(KEYINPUT119), .B(n680), .Z(n682) );
  NAND2_X1 U739 ( .A1(n682), .A2(n681), .ZN(n683) );
  NAND2_X1 U740 ( .A1(n684), .A2(n683), .ZN(n693) );
  INV_X1 U741 ( .A(KEYINPUT2), .ZN(n685) );
  NAND2_X1 U742 ( .A1(n685), .A2(n727), .ZN(n686) );
  XNOR2_X1 U743 ( .A(n686), .B(KEYINPUT80), .ZN(n688) );
  NAND2_X1 U744 ( .A1(n688), .A2(n687), .ZN(n691) );
  INV_X1 U745 ( .A(n689), .ZN(n712) );
  NOR2_X1 U746 ( .A1(n712), .A2(KEYINPUT2), .ZN(n690) );
  NOR2_X1 U747 ( .A1(n691), .A2(n690), .ZN(n692) );
  NOR2_X1 U748 ( .A1(n693), .A2(n692), .ZN(n694) );
  NAND2_X1 U749 ( .A1(n729), .A2(n694), .ZN(n695) );
  XOR2_X1 U750 ( .A(KEYINPUT53), .B(n695), .Z(G75) );
  INV_X1 U751 ( .A(n696), .ZN(n709) );
  NAND2_X1 U752 ( .A1(n347), .A2(G469), .ZN(n700) );
  XOR2_X1 U753 ( .A(KEYINPUT121), .B(KEYINPUT120), .Z(n698) );
  XNOR2_X1 U754 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n697) );
  NOR2_X1 U755 ( .A1(n709), .A2(n701), .ZN(G54) );
  NAND2_X1 U756 ( .A1(G478), .A2(n347), .ZN(n702) );
  XNOR2_X1 U757 ( .A(n703), .B(n702), .ZN(n704) );
  NOR2_X1 U758 ( .A1(n709), .A2(n704), .ZN(G63) );
  NAND2_X1 U759 ( .A1(G217), .A2(n347), .ZN(n706) );
  XNOR2_X1 U760 ( .A(n707), .B(n706), .ZN(n708) );
  NOR2_X1 U761 ( .A1(n709), .A2(n708), .ZN(G66) );
  NAND2_X1 U762 ( .A1(G953), .A2(G224), .ZN(n710) );
  XNOR2_X1 U763 ( .A(KEYINPUT61), .B(n710), .ZN(n711) );
  NAND2_X1 U764 ( .A1(n711), .A2(G898), .ZN(n714) );
  NAND2_X1 U765 ( .A1(n712), .A2(n729), .ZN(n713) );
  NAND2_X1 U766 ( .A1(n714), .A2(n713), .ZN(n720) );
  XOR2_X1 U767 ( .A(n715), .B(KEYINPUT123), .Z(n716) );
  NOR2_X1 U768 ( .A1(n717), .A2(n716), .ZN(n718) );
  XOR2_X1 U769 ( .A(KEYINPUT124), .B(n718), .Z(n719) );
  XOR2_X1 U770 ( .A(n720), .B(n719), .Z(G69) );
  XOR2_X1 U771 ( .A(n721), .B(KEYINPUT125), .Z(n722) );
  XNOR2_X1 U772 ( .A(n723), .B(n722), .ZN(n728) );
  XNOR2_X1 U773 ( .A(G227), .B(n728), .ZN(n724) );
  NAND2_X1 U774 ( .A1(n724), .A2(G900), .ZN(n725) );
  NAND2_X1 U775 ( .A1(n725), .A2(G953), .ZN(n726) );
  XNOR2_X1 U776 ( .A(n726), .B(KEYINPUT126), .ZN(n732) );
  XNOR2_X1 U777 ( .A(n728), .B(n727), .ZN(n730) );
  NAND2_X1 U778 ( .A1(n730), .A2(n729), .ZN(n731) );
  NAND2_X1 U779 ( .A1(n732), .A2(n731), .ZN(G72) );
  XOR2_X1 U780 ( .A(n733), .B(G122), .Z(G24) );
  XOR2_X1 U781 ( .A(G119), .B(n734), .Z(G21) );
  XOR2_X1 U782 ( .A(G137), .B(n735), .Z(G39) );
  XNOR2_X1 U783 ( .A(G131), .B(KEYINPUT127), .ZN(n737) );
  XNOR2_X1 U784 ( .A(n737), .B(n736), .ZN(G33) );
endmodule

