//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 0 1 1 0 1 0 1 1 1 1 0 1 0 1 1 0 1 1 1 0 1 1 1 1 0 0 1 1 0 0 1 1 0 1 0 0 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n706, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n751, new_n752, new_n753, new_n754, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n763, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n779, new_n780, new_n781,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n861, new_n862, new_n863,
    new_n864, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n923, new_n924,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n971, new_n972,
    new_n973, new_n974, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988;
  INV_X1    g000(.A(KEYINPUT86), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT77), .ZN(new_n203));
  NAND2_X1  g002(.A1(G226gat), .A2(G233gat), .ZN(new_n204));
  INV_X1    g003(.A(G183gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(KEYINPUT27), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT27), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(G183gat), .ZN(new_n208));
  INV_X1    g007(.A(G190gat), .ZN(new_n209));
  AND4_X1   g008(.A1(KEYINPUT28), .A2(new_n206), .A3(new_n208), .A4(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT65), .ZN(new_n211));
  AOI21_X1  g010(.A(G190gat), .B1(new_n206), .B2(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(KEYINPUT27), .B(G183gat), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n212), .B1(new_n211), .B2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT28), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n210), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(G183gat), .A2(G190gat), .ZN(new_n217));
  OAI21_X1  g016(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n218));
  XNOR2_X1  g017(.A(new_n218), .B(KEYINPUT66), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT26), .ZN(new_n220));
  INV_X1    g019(.A(G169gat), .ZN(new_n221));
  INV_X1    g020(.A(G176gat), .ZN(new_n222));
  NAND4_X1  g021(.A1(new_n220), .A2(new_n221), .A3(new_n222), .A4(KEYINPUT67), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT67), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n224), .B1(G169gat), .B2(G176gat), .ZN(new_n225));
  NOR3_X1   g024(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n223), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n217), .B1(new_n219), .B2(new_n227), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n216), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT64), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n205), .A2(G190gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n209), .A2(G183gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(KEYINPUT24), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT23), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n235), .A2(new_n221), .A3(new_n222), .ZN(new_n236));
  OAI21_X1  g035(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  AND2_X1   g037(.A1(G183gat), .A2(G190gat), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT24), .ZN(new_n240));
  AOI22_X1  g039(.A1(new_n239), .A2(new_n240), .B1(G169gat), .B2(G176gat), .ZN(new_n241));
  AND4_X1   g040(.A1(KEYINPUT25), .A2(new_n234), .A3(new_n238), .A4(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(G169gat), .A2(G176gat), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n243), .B1(new_n217), .B2(KEYINPUT24), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n244), .B1(new_n233), .B2(KEYINPUT24), .ZN(new_n245));
  AOI21_X1  g044(.A(KEYINPUT25), .B1(new_n245), .B2(new_n238), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n230), .B1(new_n242), .B2(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(G183gat), .B(G190gat), .ZN(new_n248));
  OAI211_X1 g047(.A(new_n241), .B(new_n238), .C1(new_n240), .C2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT25), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n245), .A2(KEYINPUT25), .A3(new_n238), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n251), .A2(KEYINPUT64), .A3(new_n252), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n229), .B1(new_n247), .B2(new_n253), .ZN(new_n254));
  OAI211_X1 g053(.A(KEYINPUT75), .B(new_n204), .C1(new_n254), .C2(KEYINPUT29), .ZN(new_n255));
  INV_X1    g054(.A(new_n204), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT66), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n218), .B(new_n257), .ZN(new_n258));
  OR2_X1    g057(.A1(new_n225), .A2(new_n226), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n258), .A2(new_n259), .A3(new_n223), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n206), .A2(new_n208), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(KEYINPUT65), .ZN(new_n262));
  AOI21_X1  g061(.A(KEYINPUT28), .B1(new_n262), .B2(new_n212), .ZN(new_n263));
  OAI211_X1 g062(.A(new_n260), .B(new_n217), .C1(new_n263), .C2(new_n210), .ZN(new_n264));
  AND3_X1   g063(.A1(new_n251), .A2(KEYINPUT64), .A3(new_n252), .ZN(new_n265));
  AOI21_X1  g064(.A(KEYINPUT64), .B1(new_n251), .B2(new_n252), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n264), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT29), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n256), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT75), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n251), .A2(new_n252), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n264), .A2(new_n271), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n270), .B1(new_n272), .B2(new_n256), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n255), .B1(new_n269), .B2(new_n273), .ZN(new_n274));
  AOI21_X1  g073(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n275));
  OR2_X1    g074(.A1(new_n275), .A2(KEYINPUT73), .ZN(new_n276));
  XNOR2_X1  g075(.A(G197gat), .B(G204gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n275), .A2(KEYINPUT73), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n276), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT74), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  XOR2_X1   g080(.A(G211gat), .B(G218gat), .Z(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(new_n282), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n279), .A2(new_n280), .A3(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n274), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n204), .A2(new_n268), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n288), .B1(new_n264), .B2(new_n271), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n289), .B1(new_n254), .B2(new_n256), .ZN(new_n290));
  OAI21_X1  g089(.A(KEYINPUT76), .B1(new_n290), .B2(new_n286), .ZN(new_n291));
  INV_X1    g090(.A(new_n289), .ZN(new_n292));
  OAI211_X1 g091(.A(new_n256), .B(new_n264), .C1(new_n265), .C2(new_n266), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT76), .ZN(new_n295));
  AND3_X1   g094(.A1(new_n279), .A2(new_n280), .A3(new_n284), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n284), .B1(new_n279), .B2(new_n280), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n294), .A2(new_n295), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n291), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n287), .A2(new_n300), .ZN(new_n301));
  XNOR2_X1  g100(.A(G8gat), .B(G36gat), .ZN(new_n302));
  XNOR2_X1  g101(.A(G64gat), .B(G92gat), .ZN(new_n303));
  XOR2_X1   g102(.A(new_n302), .B(new_n303), .Z(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n203), .B1(new_n301), .B2(new_n305), .ZN(new_n306));
  AOI211_X1 g105(.A(KEYINPUT77), .B(new_n304), .C1(new_n287), .C2(new_n300), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT30), .ZN(new_n308));
  AOI22_X1  g107(.A1(new_n286), .A2(new_n274), .B1(new_n291), .B2(new_n299), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n308), .B1(new_n309), .B2(new_n304), .ZN(new_n310));
  AND4_X1   g109(.A1(new_n308), .A2(new_n287), .A3(new_n300), .A4(new_n304), .ZN(new_n311));
  OAI22_X1  g110(.A1(new_n306), .A2(new_n307), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(G127gat), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n313), .A2(KEYINPUT68), .A3(G134gat), .ZN(new_n314));
  XNOR2_X1  g113(.A(G113gat), .B(G120gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n313), .A2(G134gat), .ZN(new_n316));
  INV_X1    g115(.A(G134gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(G127gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  OAI221_X1 g118(.A(new_n314), .B1(new_n315), .B2(KEYINPUT1), .C1(KEYINPUT68), .C2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT69), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n316), .A2(new_n318), .A3(KEYINPUT69), .ZN(new_n323));
  INV_X1    g122(.A(new_n315), .ZN(new_n324));
  XOR2_X1   g123(.A(KEYINPUT70), .B(KEYINPUT1), .Z(new_n325));
  NAND4_X1  g124(.A1(new_n322), .A2(new_n323), .A3(new_n324), .A4(new_n325), .ZN(new_n326));
  AND2_X1   g125(.A1(new_n320), .A2(new_n326), .ZN(new_n327));
  XOR2_X1   g126(.A(G141gat), .B(G148gat), .Z(new_n328));
  INV_X1    g127(.A(G155gat), .ZN(new_n329));
  INV_X1    g128(.A(G162gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(G155gat), .A2(G162gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(KEYINPUT2), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n328), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  XNOR2_X1  g134(.A(G141gat), .B(G148gat), .ZN(new_n336));
  OAI211_X1 g135(.A(new_n332), .B(new_n331), .C1(new_n336), .C2(KEYINPUT2), .ZN(new_n337));
  AND2_X1   g136(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n327), .A2(KEYINPUT4), .A3(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT4), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n320), .A2(new_n326), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n335), .A2(new_n337), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n340), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(KEYINPUT3), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT3), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n335), .A2(new_n337), .A3(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n344), .A2(new_n341), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(G225gat), .A2(G233gat), .ZN(new_n348));
  NAND4_X1  g147(.A1(new_n339), .A2(new_n343), .A3(new_n347), .A4(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n341), .A2(new_n342), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n338), .A2(new_n320), .A3(new_n326), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n348), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  XOR2_X1   g151(.A(KEYINPUT78), .B(KEYINPUT5), .Z(new_n353));
  OAI21_X1  g152(.A(new_n349), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  XOR2_X1   g153(.A(G1gat), .B(G29gat), .Z(new_n355));
  XNOR2_X1  g154(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n356));
  XNOR2_X1  g155(.A(new_n355), .B(new_n356), .ZN(new_n357));
  XNOR2_X1  g156(.A(G57gat), .B(G85gat), .ZN(new_n358));
  XNOR2_X1  g157(.A(new_n357), .B(new_n358), .ZN(new_n359));
  OAI211_X1 g158(.A(new_n354), .B(new_n359), .C1(new_n349), .C2(new_n353), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n339), .A2(new_n347), .A3(new_n343), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT39), .ZN(new_n362));
  INV_X1    g161(.A(new_n348), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n361), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(new_n359), .ZN(new_n365));
  AND2_X1   g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n350), .A2(new_n351), .A3(new_n348), .ZN(new_n367));
  XNOR2_X1  g166(.A(new_n367), .B(KEYINPUT82), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n362), .B1(new_n361), .B2(new_n363), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  AND2_X1   g169(.A1(new_n366), .A2(new_n370), .ZN(new_n371));
  XNOR2_X1  g170(.A(KEYINPUT83), .B(KEYINPUT40), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n360), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n366), .A2(new_n370), .A3(KEYINPUT40), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT84), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n371), .A2(KEYINPUT84), .A3(KEYINPUT40), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n373), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n312), .A2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n354), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n349), .A2(new_n353), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n365), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT6), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n382), .A2(new_n383), .A3(new_n360), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n287), .A2(new_n300), .A3(new_n304), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n380), .A2(new_n381), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n386), .A2(KEYINPUT6), .A3(new_n359), .ZN(new_n387));
  AND3_X1   g186(.A1(new_n384), .A2(new_n385), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n274), .A2(new_n298), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT37), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n390), .B1(new_n294), .B2(new_n286), .ZN(new_n391));
  AOI21_X1  g190(.A(KEYINPUT38), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  OAI211_X1 g191(.A(new_n392), .B(new_n305), .C1(KEYINPUT37), .C2(new_n301), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n295), .B1(new_n294), .B2(new_n298), .ZN(new_n394));
  AOI211_X1 g193(.A(KEYINPUT76), .B(new_n286), .C1(new_n292), .C2(new_n293), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n204), .B1(new_n254), .B2(KEYINPUT29), .ZN(new_n397));
  INV_X1    g196(.A(new_n273), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n298), .B1(new_n399), .B2(new_n255), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n305), .B1(new_n396), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n305), .A2(KEYINPUT37), .ZN(new_n402));
  AOI22_X1  g201(.A1(new_n401), .A2(new_n402), .B1(KEYINPUT37), .B2(new_n301), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT38), .ZN(new_n404));
  OAI211_X1 g203(.A(new_n388), .B(new_n393), .C1(new_n403), .C2(new_n404), .ZN(new_n405));
  XNOR2_X1  g204(.A(G78gat), .B(G106gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(KEYINPUT31), .B(G50gat), .ZN(new_n407));
  XNOR2_X1  g206(.A(new_n406), .B(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(G228gat), .A2(G233gat), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n279), .A2(new_n284), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n276), .A2(new_n282), .A3(new_n277), .A4(new_n278), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n411), .A2(new_n268), .A3(new_n412), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n338), .B1(new_n413), .B2(new_n345), .ZN(new_n414));
  AOI22_X1  g213(.A1(new_n283), .A2(new_n285), .B1(new_n268), .B2(new_n346), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n410), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(G22gat), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n283), .A2(new_n268), .A3(new_n285), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n338), .B1(new_n418), .B2(new_n345), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n346), .A2(new_n268), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n286), .A2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(new_n410), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  OAI211_X1 g222(.A(new_n416), .B(new_n417), .C1(new_n419), .C2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(KEYINPUT3), .B1(new_n298), .B2(new_n268), .ZN(new_n426));
  OAI211_X1 g225(.A(new_n422), .B(new_n421), .C1(new_n426), .C2(new_n338), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n417), .B1(new_n427), .B2(new_n416), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n409), .B1(new_n425), .B2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT80), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n423), .A2(new_n419), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n413), .A2(new_n345), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(new_n342), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n422), .B1(new_n433), .B2(new_n421), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n430), .B1(new_n431), .B2(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n427), .A2(KEYINPUT80), .A3(new_n416), .ZN(new_n436));
  AND3_X1   g235(.A1(new_n435), .A2(G22gat), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n424), .A2(KEYINPUT81), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT81), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n427), .A2(new_n439), .A3(new_n417), .A4(new_n416), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n438), .A2(new_n440), .A3(new_n408), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n429), .B1(new_n437), .B2(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n379), .A2(new_n405), .A3(new_n442), .ZN(new_n443));
  OAI21_X1  g242(.A(KEYINPUT77), .B1(new_n309), .B2(new_n304), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n301), .A2(new_n203), .A3(new_n305), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n385), .A2(KEYINPUT30), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n309), .A2(new_n308), .A3(new_n304), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n384), .A2(new_n387), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n446), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n442), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT34), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n267), .A2(new_n327), .ZN(new_n455));
  OAI211_X1 g254(.A(new_n341), .B(new_n264), .C1(new_n265), .C2(new_n266), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(G227gat), .A2(G233gat), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n454), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT71), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n457), .A2(new_n454), .A3(new_n458), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n459), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(new_n458), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n455), .A2(new_n463), .A3(new_n456), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(KEYINPUT32), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT33), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  XOR2_X1   g266(.A(G15gat), .B(G43gat), .Z(new_n468));
  XNOR2_X1  g267(.A(G71gat), .B(G99gat), .ZN(new_n469));
  XNOR2_X1  g268(.A(new_n468), .B(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n465), .A2(new_n467), .A3(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(new_n470), .ZN(new_n472));
  OAI211_X1 g271(.A(new_n464), .B(KEYINPUT32), .C1(new_n466), .C2(new_n472), .ZN(new_n473));
  NAND4_X1  g272(.A1(new_n457), .A2(KEYINPUT71), .A3(new_n454), .A4(new_n458), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n462), .A2(new_n471), .A3(new_n473), .A4(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n471), .A2(new_n473), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n461), .A2(new_n460), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n457), .A2(new_n458), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(KEYINPUT34), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n477), .A2(new_n474), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n476), .A2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT72), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n475), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT36), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n476), .A2(new_n480), .A3(KEYINPUT72), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n475), .A2(new_n481), .A3(KEYINPUT36), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  AND3_X1   g287(.A1(new_n443), .A2(new_n453), .A3(new_n488), .ZN(new_n489));
  AND3_X1   g288(.A1(new_n446), .A2(new_n449), .A3(new_n450), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n475), .A2(new_n481), .A3(new_n442), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(KEYINPUT85), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT85), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n475), .A2(new_n481), .A3(new_n442), .A4(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n490), .A2(new_n492), .A3(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT35), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n442), .A2(new_n496), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n451), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n483), .A2(new_n485), .ZN(new_n499));
  AOI22_X1  g298(.A1(new_n495), .A2(KEYINPUT35), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n202), .B1(new_n489), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n495), .A2(KEYINPUT35), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n498), .A2(new_n499), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n443), .A2(new_n453), .A3(new_n488), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n504), .A2(KEYINPUT86), .A3(new_n505), .ZN(new_n506));
  XOR2_X1   g305(.A(G57gat), .B(G64gat), .Z(new_n507));
  INV_X1    g306(.A(KEYINPUT9), .ZN(new_n508));
  INV_X1    g307(.A(G71gat), .ZN(new_n509));
  INV_X1    g308(.A(G78gat), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n507), .A2(new_n511), .ZN(new_n512));
  XOR2_X1   g311(.A(G71gat), .B(G78gat), .Z(new_n513));
  OR2_X1    g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n512), .A2(new_n513), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT21), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(G231gat), .A2(G233gat), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n518), .B(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n520), .B(G127gat), .ZN(new_n521));
  XNOR2_X1  g320(.A(G15gat), .B(G22gat), .ZN(new_n522));
  INV_X1    g321(.A(G1gat), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n522), .A2(KEYINPUT16), .A3(new_n523), .ZN(new_n524));
  OR2_X1    g323(.A1(KEYINPUT89), .A2(G8gat), .ZN(new_n525));
  OAI211_X1 g324(.A(new_n524), .B(new_n525), .C1(new_n523), .C2(new_n522), .ZN(new_n526));
  NAND2_X1  g325(.A1(KEYINPUT89), .A2(G8gat), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n526), .B(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(new_n528), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n529), .B1(new_n517), .B2(new_n516), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n521), .B(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n532), .B(new_n329), .ZN(new_n533));
  XOR2_X1   g332(.A(G183gat), .B(G211gat), .Z(new_n534));
  XNOR2_X1  g333(.A(new_n533), .B(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  OR2_X1    g335(.A1(new_n531), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n531), .A2(new_n536), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(KEYINPUT14), .B(G29gat), .ZN(new_n540));
  INV_X1    g339(.A(G36gat), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(G29gat), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n543), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  AOI21_X1  g344(.A(KEYINPUT15), .B1(G43gat), .B2(G50gat), .ZN(new_n546));
  XNOR2_X1  g345(.A(KEYINPUT87), .B(G43gat), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n546), .B1(new_n547), .B2(G50gat), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(G43gat), .B(G50gat), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(KEYINPUT15), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n545), .A2(KEYINPUT15), .A3(new_n550), .ZN(new_n553));
  AND2_X1   g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT88), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n554), .A2(new_n555), .A3(KEYINPUT17), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n552), .A2(new_n555), .A3(new_n553), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT17), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(G85gat), .A2(G92gat), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n561), .B(KEYINPUT7), .ZN(new_n562));
  XNOR2_X1  g361(.A(G99gat), .B(G106gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(G99gat), .A2(G106gat), .ZN(new_n564));
  INV_X1    g363(.A(G85gat), .ZN(new_n565));
  INV_X1    g364(.A(G92gat), .ZN(new_n566));
  AOI22_X1  g365(.A1(KEYINPUT8), .A2(new_n564), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  AND3_X1   g366(.A1(new_n562), .A2(new_n563), .A3(new_n567), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n563), .B1(new_n562), .B2(new_n567), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n570), .A2(KEYINPUT92), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT92), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n572), .B1(new_n568), .B2(new_n569), .ZN(new_n573));
  AND2_X1   g372(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n560), .A2(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(G190gat), .B(G218gat), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(KEYINPUT93), .ZN(new_n577));
  AND2_X1   g376(.A1(G232gat), .A2(G233gat), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n578), .A2(KEYINPUT41), .ZN(new_n579));
  AND2_X1   g378(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n552), .A2(new_n553), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n580), .B1(new_n574), .B2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n576), .A2(KEYINPUT93), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n575), .A2(new_n583), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n571), .A2(new_n573), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n587), .B1(new_n556), .B2(new_n559), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n584), .B1(new_n588), .B2(new_n582), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n578), .A2(KEYINPUT41), .ZN(new_n590));
  XNOR2_X1  g389(.A(G134gat), .B(G162gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n590), .B(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n586), .A2(new_n589), .A3(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n592), .B1(new_n586), .B2(new_n589), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(G230gat), .A2(G233gat), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n516), .A2(new_n570), .ZN(new_n599));
  OAI211_X1 g398(.A(new_n514), .B(new_n515), .C1(new_n568), .C2(new_n569), .ZN(new_n600));
  AOI21_X1  g399(.A(KEYINPUT10), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n514), .A2(KEYINPUT10), .A3(new_n515), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n602), .B1(new_n571), .B2(new_n573), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n598), .B1(new_n601), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n599), .A2(new_n600), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n604), .B1(new_n598), .B2(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(G120gat), .B(G148gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(G176gat), .B(G204gat), .ZN(new_n608));
  XOR2_X1   g407(.A(new_n607), .B(new_n608), .Z(new_n609));
  XNOR2_X1  g408(.A(new_n606), .B(new_n609), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n539), .A2(new_n597), .A3(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(G113gat), .B(G141gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(G197gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(KEYINPUT11), .B(G169gat), .ZN(new_n614));
  XOR2_X1   g413(.A(new_n613), .B(new_n614), .Z(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(KEYINPUT12), .ZN(new_n616));
  AND2_X1   g415(.A1(new_n557), .A2(new_n558), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n557), .A2(new_n558), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n529), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(G229gat), .A2(G233gat), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n554), .A2(new_n528), .ZN(new_n621));
  NAND4_X1  g420(.A1(new_n619), .A2(KEYINPUT18), .A3(new_n620), .A4(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n622), .A2(KEYINPUT90), .ZN(new_n623));
  INV_X1    g422(.A(new_n621), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n624), .B1(new_n560), .B2(new_n529), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT90), .ZN(new_n626));
  NAND4_X1  g425(.A1(new_n625), .A2(new_n626), .A3(KEYINPUT18), .A4(new_n620), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n623), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n619), .A2(new_n620), .A3(new_n621), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT18), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n529), .A2(new_n581), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n631), .A2(new_n621), .ZN(new_n632));
  XOR2_X1   g431(.A(new_n620), .B(KEYINPUT13), .Z(new_n633));
  AOI22_X1  g432(.A1(new_n629), .A2(new_n630), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n616), .B1(new_n628), .B2(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n628), .A2(new_n616), .A3(new_n634), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n636), .A2(KEYINPUT91), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT91), .ZN(new_n638));
  NAND4_X1  g437(.A1(new_n628), .A2(new_n638), .A3(new_n616), .A4(new_n634), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n635), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n611), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n501), .A2(new_n506), .A3(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n642), .A2(new_n450), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(new_n523), .ZN(G1324gat));
  INV_X1    g443(.A(KEYINPUT42), .ZN(new_n645));
  INV_X1    g444(.A(new_n312), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n642), .A2(new_n646), .ZN(new_n647));
  XOR2_X1   g446(.A(KEYINPUT16), .B(G8gat), .Z(new_n648));
  AOI21_X1  g447(.A(new_n645), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  OAI21_X1  g448(.A(G8gat), .B1(new_n642), .B2(new_n646), .ZN(new_n650));
  NOR2_X1   g449(.A1(KEYINPUT94), .A2(KEYINPUT42), .ZN(new_n651));
  MUX2_X1   g450(.A(KEYINPUT94), .B(new_n651), .S(new_n648), .Z(new_n652));
  AOI22_X1  g451(.A1(new_n649), .A2(new_n650), .B1(new_n647), .B2(new_n652), .ZN(G1325gat));
  NOR2_X1   g452(.A1(new_n488), .A2(KEYINPUT95), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT95), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n655), .B1(new_n486), .B2(new_n487), .ZN(new_n656));
  OR2_X1    g455(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  OAI21_X1  g456(.A(G15gat), .B1(new_n642), .B2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n499), .ZN(new_n659));
  OR2_X1    g458(.A1(new_n659), .A2(G15gat), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n658), .B1(new_n642), .B2(new_n660), .ZN(G1326gat));
  NOR2_X1   g460(.A1(new_n642), .A2(new_n442), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT96), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n662), .A2(new_n663), .ZN(new_n666));
  OR3_X1    g465(.A1(new_n665), .A2(KEYINPUT97), .A3(new_n666), .ZN(new_n667));
  OAI21_X1  g466(.A(KEYINPUT97), .B1(new_n665), .B2(new_n666), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g468(.A(KEYINPUT43), .B(G22gat), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n669), .B(new_n671), .ZN(G1327gat));
  NAND3_X1  g471(.A1(new_n501), .A2(new_n506), .A3(new_n596), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n673), .A2(KEYINPUT44), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT99), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n675), .B1(new_n594), .B2(new_n595), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n586), .A2(new_n589), .ZN(new_n677));
  INV_X1    g476(.A(new_n592), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n679), .A2(KEYINPUT99), .A3(new_n593), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n676), .A2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n682), .A2(KEYINPUT44), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  OAI211_X1 g483(.A(new_n443), .B(new_n453), .C1(new_n654), .C2(new_n656), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n684), .B1(new_n685), .B2(new_n504), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n674), .A2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT100), .ZN(new_n689));
  INV_X1    g488(.A(new_n610), .ZN(new_n690));
  NOR3_X1   g489(.A1(new_n539), .A2(new_n640), .A3(new_n690), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(KEYINPUT98), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n688), .A2(new_n689), .A3(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n450), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n686), .B1(new_n673), .B2(KEYINPUT44), .ZN(new_n696));
  OAI21_X1  g495(.A(KEYINPUT100), .B1(new_n696), .B2(new_n692), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n694), .A2(new_n695), .A3(new_n697), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n543), .B1(new_n698), .B2(KEYINPUT101), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n699), .B1(KEYINPUT101), .B2(new_n698), .ZN(new_n700));
  NAND4_X1  g499(.A1(new_n501), .A2(new_n506), .A3(new_n596), .A4(new_n691), .ZN(new_n701));
  INV_X1    g500(.A(new_n701), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n702), .A2(new_n543), .A3(new_n695), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(KEYINPUT45), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n700), .A2(new_n704), .ZN(G1328gat));
  NOR3_X1   g504(.A1(new_n701), .A2(G36gat), .A3(new_n646), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n706), .B(KEYINPUT46), .ZN(new_n707));
  AND3_X1   g506(.A1(new_n694), .A2(new_n312), .A3(new_n697), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n707), .B1(new_n708), .B2(new_n541), .ZN(G1329gat));
  INV_X1    g508(.A(new_n657), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n694), .A2(new_n710), .A3(new_n697), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(new_n547), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT47), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n659), .A2(new_n547), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n701), .A2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT102), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NOR3_X1   g517(.A1(new_n701), .A2(KEYINPUT102), .A3(new_n715), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n713), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n712), .A2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT103), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n688), .A2(new_n710), .A3(new_n693), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(new_n547), .ZN(new_n725));
  INV_X1    g524(.A(new_n716), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(KEYINPUT47), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n722), .A2(new_n723), .A3(new_n728), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n720), .B1(new_n711), .B2(new_n547), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n713), .B1(new_n725), .B2(new_n726), .ZN(new_n731));
  OAI21_X1  g530(.A(KEYINPUT103), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n729), .A2(new_n732), .ZN(G1330gat));
  INV_X1    g532(.A(G50gat), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n452), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n735), .B1(new_n702), .B2(KEYINPUT104), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n736), .B1(KEYINPUT104), .B2(new_n702), .ZN(new_n737));
  NOR3_X1   g536(.A1(new_n696), .A2(new_n442), .A3(new_n692), .ZN(new_n738));
  OAI211_X1 g537(.A(new_n737), .B(KEYINPUT48), .C1(new_n734), .C2(new_n738), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n694), .A2(new_n452), .A3(new_n697), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(G50gat), .ZN(new_n741));
  AND2_X1   g540(.A1(new_n741), .A2(new_n737), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n739), .B1(new_n742), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g542(.A1(new_n685), .A2(new_n504), .ZN(new_n744));
  INV_X1    g543(.A(new_n539), .ZN(new_n745));
  INV_X1    g544(.A(new_n640), .ZN(new_n746));
  NOR4_X1   g545(.A1(new_n745), .A2(new_n746), .A3(new_n596), .A4(new_n610), .ZN(new_n747));
  AND2_X1   g546(.A1(new_n744), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(new_n695), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g549(.A(new_n646), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n748), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(KEYINPUT105), .ZN(new_n753));
  NOR2_X1   g552(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n753), .B(new_n754), .ZN(G1333gat));
  INV_X1    g554(.A(new_n748), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n509), .B1(new_n756), .B2(new_n659), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n657), .A2(new_n509), .ZN(new_n758));
  AND3_X1   g557(.A1(new_n748), .A2(KEYINPUT106), .A3(new_n758), .ZN(new_n759));
  AOI21_X1  g558(.A(KEYINPUT106), .B1(new_n748), .B2(new_n758), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n757), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g561(.A1(new_n748), .A2(new_n452), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g563(.A1(new_n746), .A2(new_n539), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n688), .A2(new_n690), .A3(new_n765), .ZN(new_n766));
  OAI21_X1  g565(.A(G85gat), .B1(new_n766), .B2(new_n450), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n744), .A2(new_n596), .A3(new_n765), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT51), .ZN(new_n769));
  OR2_X1    g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n768), .A2(new_n769), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT107), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n770), .A2(KEYINPUT107), .A3(new_n771), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n774), .A2(new_n690), .A3(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n695), .A2(new_n565), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n767), .B1(new_n776), .B2(new_n777), .ZN(G1336gat));
  NAND4_X1  g577(.A1(new_n772), .A2(new_n566), .A3(new_n312), .A4(new_n690), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n766), .A2(new_n646), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n779), .B1(new_n780), .B2(new_n566), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n781), .B(KEYINPUT52), .ZN(G1337gat));
  OAI21_X1  g581(.A(G99gat), .B1(new_n766), .B2(new_n657), .ZN(new_n783));
  OR2_X1    g582(.A1(new_n659), .A2(G99gat), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n783), .B1(new_n776), .B2(new_n784), .ZN(G1338gat));
  OAI21_X1  g584(.A(G106gat), .B1(new_n766), .B2(new_n442), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT109), .ZN(new_n787));
  OR3_X1    g586(.A1(new_n442), .A2(G106gat), .A3(new_n610), .ZN(new_n788));
  INV_X1    g587(.A(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n772), .A2(KEYINPUT108), .A3(new_n789), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n786), .A2(new_n787), .A3(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT53), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n787), .A2(KEYINPUT53), .ZN(new_n793));
  AOI22_X1  g592(.A1(new_n772), .A2(new_n789), .B1(KEYINPUT108), .B2(new_n793), .ZN(new_n794));
  AOI22_X1  g593(.A1(new_n791), .A2(new_n792), .B1(new_n786), .B2(new_n794), .ZN(G1339gat));
  INV_X1    g594(.A(KEYINPUT114), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT10), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n605), .A2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(new_n603), .ZN(new_n799));
  INV_X1    g598(.A(new_n598), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n798), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT110), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n798), .A2(new_n799), .A3(KEYINPUT110), .A4(new_n800), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n803), .A2(new_n804), .A3(KEYINPUT54), .A4(new_n604), .ZN(new_n805));
  INV_X1    g604(.A(new_n604), .ZN(new_n806));
  XNOR2_X1  g605(.A(KEYINPUT111), .B(KEYINPUT54), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n609), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n805), .A2(KEYINPUT55), .A3(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(KEYINPUT112), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT112), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n805), .A2(new_n811), .A3(KEYINPUT55), .A4(new_n808), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(KEYINPUT55), .B1(new_n805), .B2(new_n808), .ZN(new_n814));
  INV_X1    g613(.A(new_n606), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n814), .B1(new_n815), .B2(new_n609), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n813), .A2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  OAI22_X1  g617(.A1(new_n625), .A2(new_n620), .B1(new_n632), .B2(new_n633), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(new_n615), .ZN(new_n820));
  INV_X1    g619(.A(new_n820), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n821), .B1(new_n637), .B2(new_n639), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT113), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n818), .A2(new_n822), .A3(new_n823), .A4(new_n681), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n637), .A2(new_n639), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(new_n820), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n681), .A2(new_n813), .A3(new_n816), .ZN(new_n827));
  OAI21_X1  g626(.A(KEYINPUT113), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n824), .A2(new_n828), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n640), .A2(new_n817), .ZN(new_n830));
  AOI211_X1 g629(.A(new_n610), .B(new_n821), .C1(new_n637), .C2(new_n639), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n682), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n539), .B1(new_n829), .B2(new_n832), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n611), .A2(new_n746), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n796), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(new_n834), .ZN(new_n836));
  OAI22_X1  g635(.A1(new_n826), .A2(new_n610), .B1(new_n640), .B2(new_n817), .ZN(new_n837));
  AOI22_X1  g636(.A1(new_n828), .A2(new_n824), .B1(new_n837), .B2(new_n682), .ZN(new_n838));
  OAI211_X1 g637(.A(KEYINPUT114), .B(new_n836), .C1(new_n838), .C2(new_n539), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n835), .A2(new_n839), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n840), .A2(new_n450), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n492), .A2(new_n494), .ZN(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n843), .A2(new_n312), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(G113gat), .B1(new_n846), .B2(new_n746), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n312), .A2(new_n450), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n659), .A2(new_n452), .ZN(new_n849));
  NAND4_X1  g648(.A1(new_n835), .A2(new_n839), .A3(new_n848), .A4(new_n849), .ZN(new_n850));
  XNOR2_X1  g649(.A(new_n850), .B(KEYINPUT115), .ZN(new_n851));
  AND2_X1   g650(.A1(new_n746), .A2(G113gat), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n847), .B1(new_n851), .B2(new_n852), .ZN(G1340gat));
  INV_X1    g652(.A(G120gat), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n846), .A2(new_n854), .A3(new_n690), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT116), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n851), .A2(new_n690), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n856), .B1(new_n857), .B2(G120gat), .ZN(new_n858));
  AOI211_X1 g657(.A(KEYINPUT116), .B(new_n854), .C1(new_n851), .C2(new_n690), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n855), .B1(new_n858), .B2(new_n859), .ZN(G1341gat));
  NOR3_X1   g659(.A1(new_n845), .A2(KEYINPUT117), .A3(new_n745), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n861), .A2(G127gat), .ZN(new_n862));
  OAI21_X1  g661(.A(KEYINPUT117), .B1(new_n845), .B2(new_n745), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n745), .A2(new_n313), .ZN(new_n864));
  AOI22_X1  g663(.A1(new_n862), .A2(new_n863), .B1(new_n851), .B2(new_n864), .ZN(G1342gat));
  AND4_X1   g664(.A1(new_n317), .A2(new_n841), .A3(new_n596), .A4(new_n844), .ZN(new_n866));
  XNOR2_X1  g665(.A(new_n866), .B(KEYINPUT56), .ZN(new_n867));
  AOI211_X1 g666(.A(KEYINPUT118), .B(new_n317), .C1(new_n851), .C2(new_n596), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT118), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n851), .A2(new_n596), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n869), .B1(new_n870), .B2(G134gat), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n867), .B1(new_n868), .B2(new_n871), .ZN(G1343gat));
  INV_X1    g671(.A(G141gat), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n657), .A2(new_n848), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n835), .A2(new_n839), .A3(new_n452), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT57), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  AOI22_X1  g676(.A1(new_n828), .A2(new_n824), .B1(new_n837), .B2(new_n597), .ZN(new_n878));
  OAI21_X1  g677(.A(KEYINPUT119), .B1(new_n878), .B2(new_n539), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n837), .A2(new_n597), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n829), .A2(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT119), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n881), .A2(new_n882), .A3(new_n745), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n879), .A2(new_n883), .A3(new_n836), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n452), .A2(KEYINPUT57), .ZN(new_n885));
  INV_X1    g684(.A(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n874), .B1(new_n877), .B2(new_n887), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n873), .B1(new_n888), .B2(new_n746), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n710), .A2(new_n442), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(new_n646), .ZN(new_n891));
  NOR3_X1   g690(.A1(new_n840), .A2(new_n891), .A3(new_n450), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n746), .A2(new_n873), .ZN(new_n893));
  XOR2_X1   g692(.A(new_n893), .B(KEYINPUT120), .Z(new_n894));
  AND2_X1   g693(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  OAI21_X1  g694(.A(KEYINPUT58), .B1(new_n889), .B2(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(KEYINPUT121), .B1(new_n888), .B2(new_n746), .ZN(new_n897));
  AOI22_X1  g696(.A1(new_n875), .A2(new_n876), .B1(new_n884), .B2(new_n886), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT121), .ZN(new_n899));
  NOR4_X1   g698(.A1(new_n898), .A2(new_n899), .A3(new_n640), .A4(new_n874), .ZN(new_n900));
  NOR3_X1   g699(.A1(new_n897), .A2(new_n900), .A3(new_n873), .ZN(new_n901));
  OR2_X1    g700(.A1(new_n895), .A2(KEYINPUT58), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n896), .B1(new_n901), .B2(new_n902), .ZN(G1344gat));
  INV_X1    g702(.A(G148gat), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n892), .A2(new_n904), .A3(new_n690), .ZN(new_n905));
  AOI211_X1 g704(.A(KEYINPUT59), .B(new_n904), .C1(new_n888), .C2(new_n690), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT59), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n818), .A2(new_n596), .A3(new_n822), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n880), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n834), .B1(new_n909), .B2(new_n745), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n876), .B1(new_n910), .B2(new_n442), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n911), .B1(new_n840), .B2(new_n885), .ZN(new_n912));
  NAND4_X1  g711(.A1(new_n912), .A2(new_n690), .A3(new_n657), .A4(new_n848), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n907), .B1(new_n913), .B2(G148gat), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n905), .B1(new_n906), .B2(new_n914), .ZN(G1345gat));
  NAND3_X1  g714(.A1(new_n892), .A2(new_n329), .A3(new_n539), .ZN(new_n916));
  NOR3_X1   g715(.A1(new_n898), .A2(new_n745), .A3(new_n874), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n916), .B1(new_n917), .B2(new_n329), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT122), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  OAI211_X1 g719(.A(KEYINPUT122), .B(new_n916), .C1(new_n917), .C2(new_n329), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(G1346gat));
  NAND3_X1  g721(.A1(new_n892), .A2(new_n330), .A3(new_n596), .ZN(new_n923));
  NOR3_X1   g722(.A1(new_n898), .A2(new_n682), .A3(new_n874), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n923), .B1(new_n924), .B2(new_n330), .ZN(G1347gat));
  NOR2_X1   g724(.A1(new_n646), .A2(new_n695), .ZN(new_n926));
  NAND4_X1  g725(.A1(new_n835), .A2(new_n839), .A3(new_n849), .A4(new_n926), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT123), .ZN(new_n928));
  OR2_X1    g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n927), .A2(new_n928), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n929), .A2(new_n746), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(G169gat), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT124), .ZN(new_n933));
  NOR4_X1   g732(.A1(new_n840), .A2(new_n695), .A3(new_n646), .A4(new_n843), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n934), .A2(new_n221), .A3(new_n746), .ZN(new_n935));
  AND3_X1   g734(.A1(new_n932), .A2(new_n933), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n933), .B1(new_n932), .B2(new_n935), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n936), .A2(new_n937), .ZN(G1348gat));
  NAND3_X1  g737(.A1(new_n934), .A2(new_n222), .A3(new_n690), .ZN(new_n939));
  XNOR2_X1  g738(.A(new_n927), .B(KEYINPUT123), .ZN(new_n940));
  AND2_X1   g739(.A1(new_n940), .A2(new_n690), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n939), .B1(new_n941), .B2(new_n222), .ZN(G1349gat));
  INV_X1    g741(.A(KEYINPUT60), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n745), .A2(new_n261), .ZN(new_n944));
  AOI21_X1  g743(.A(KEYINPUT125), .B1(new_n934), .B2(new_n944), .ZN(new_n945));
  AND2_X1   g744(.A1(new_n940), .A2(new_n539), .ZN(new_n946));
  OAI211_X1 g745(.A(new_n943), .B(new_n945), .C1(new_n946), .C2(new_n205), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n205), .B1(new_n940), .B2(new_n539), .ZN(new_n948));
  INV_X1    g747(.A(new_n945), .ZN(new_n949));
  OAI21_X1  g748(.A(KEYINPUT60), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n947), .A2(new_n950), .ZN(G1350gat));
  NAND3_X1  g750(.A1(new_n934), .A2(new_n209), .A3(new_n681), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT61), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n940), .A2(new_n596), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n953), .B1(new_n954), .B2(G190gat), .ZN(new_n955));
  AOI211_X1 g754(.A(KEYINPUT61), .B(new_n209), .C1(new_n940), .C2(new_n596), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n952), .B1(new_n955), .B2(new_n956), .ZN(G1351gat));
  INV_X1    g756(.A(new_n840), .ZN(new_n958));
  NAND4_X1  g757(.A1(new_n958), .A2(new_n450), .A3(new_n312), .A4(new_n890), .ZN(new_n959));
  INV_X1    g758(.A(new_n959), .ZN(new_n960));
  AOI21_X1  g759(.A(G197gat), .B1(new_n960), .B2(new_n746), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n912), .A2(KEYINPUT126), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT126), .ZN(new_n963));
  OAI211_X1 g762(.A(new_n911), .B(new_n963), .C1(new_n840), .C2(new_n885), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n657), .A2(new_n926), .ZN(new_n965));
  INV_X1    g764(.A(new_n965), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n962), .A2(new_n964), .A3(new_n966), .ZN(new_n967));
  INV_X1    g766(.A(new_n967), .ZN(new_n968));
  AND2_X1   g767(.A1(new_n746), .A2(G197gat), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n961), .B1(new_n968), .B2(new_n969), .ZN(G1352gat));
  OAI21_X1  g769(.A(G204gat), .B1(new_n967), .B2(new_n610), .ZN(new_n971));
  OR2_X1    g770(.A1(new_n610), .A2(G204gat), .ZN(new_n972));
  OAI21_X1  g771(.A(KEYINPUT62), .B1(new_n959), .B2(new_n972), .ZN(new_n973));
  OR3_X1    g772(.A1(new_n959), .A2(KEYINPUT62), .A3(new_n972), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n971), .A2(new_n973), .A3(new_n974), .ZN(G1353gat));
  INV_X1    g774(.A(G211gat), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n966), .A2(new_n539), .ZN(new_n977));
  INV_X1    g776(.A(new_n977), .ZN(new_n978));
  AOI21_X1  g777(.A(new_n976), .B1(new_n912), .B2(new_n978), .ZN(new_n979));
  XNOR2_X1  g778(.A(new_n979), .B(KEYINPUT63), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n960), .A2(new_n976), .A3(new_n539), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n980), .A2(new_n981), .ZN(G1354gat));
  INV_X1    g781(.A(G218gat), .ZN(new_n983));
  NOR2_X1   g782(.A1(new_n597), .A2(new_n983), .ZN(new_n984));
  NAND4_X1  g783(.A1(new_n962), .A2(new_n964), .A3(new_n966), .A4(new_n984), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n983), .B1(new_n959), .B2(new_n682), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g786(.A(KEYINPUT127), .ZN(new_n988));
  XNOR2_X1  g787(.A(new_n987), .B(new_n988), .ZN(G1355gat));
endmodule


