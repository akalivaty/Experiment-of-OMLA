//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 1 1 1 1 1 0 1 0 1 1 1 0 0 0 0 0 0 0 1 1 0 0 0 0 1 1 1 0 1 0 0 1 0 1 1 1 1 0 1 0 0 0 1 1 1 0 1 1 1 1 0 1 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:43 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n752, new_n753, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n763, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011;
  INV_X1    g000(.A(G134), .ZN(new_n187));
  OAI21_X1  g001(.A(KEYINPUT11), .B1(new_n187), .B2(G137), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT11), .ZN(new_n189));
  INV_X1    g003(.A(G137), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n189), .A2(new_n190), .A3(G134), .ZN(new_n191));
  AOI22_X1  g005(.A1(new_n188), .A2(new_n191), .B1(new_n187), .B2(G137), .ZN(new_n192));
  INV_X1    g006(.A(G131), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n192), .B(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT65), .ZN(new_n195));
  INV_X1    g009(.A(G146), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n195), .B1(G143), .B2(new_n196), .ZN(new_n197));
  XNOR2_X1  g011(.A(KEYINPUT64), .B(G143), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n197), .B1(new_n198), .B2(new_n196), .ZN(new_n199));
  INV_X1    g013(.A(G143), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(KEYINPUT64), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT64), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G143), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n201), .A2(new_n203), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n204), .A2(new_n195), .A3(G146), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n199), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(KEYINPUT0), .A2(G128), .ZN(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n198), .A2(new_n196), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n200), .A2(G146), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n208), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  OR2_X1    g026(.A1(KEYINPUT0), .A2(G128), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n194), .A2(new_n209), .A3(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G119), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G116), .ZN(new_n217));
  INV_X1    g031(.A(G116), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G119), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  XNOR2_X1  g034(.A(KEYINPUT2), .B(G113), .ZN(new_n221));
  OR2_X1    g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n220), .A2(new_n221), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT68), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n222), .A2(KEYINPUT68), .A3(new_n223), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n192), .A2(new_n193), .ZN(new_n229));
  OR3_X1    g043(.A1(new_n190), .A2(KEYINPUT66), .A3(G134), .ZN(new_n230));
  OAI21_X1  g044(.A(KEYINPUT66), .B1(new_n190), .B2(G134), .ZN(new_n231));
  OAI211_X1 g045(.A(new_n230), .B(new_n231), .C1(new_n187), .C2(G137), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(G131), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT1), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(G128), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n235), .B1(new_n199), .B2(new_n205), .ZN(new_n236));
  OAI21_X1  g050(.A(KEYINPUT1), .B1(new_n200), .B2(G146), .ZN(new_n237));
  AOI22_X1  g051(.A1(new_n210), .A2(new_n211), .B1(G128), .B2(new_n237), .ZN(new_n238));
  OAI211_X1 g052(.A(new_n229), .B(new_n233), .C1(new_n236), .C2(new_n238), .ZN(new_n239));
  AND3_X1   g053(.A1(new_n215), .A2(new_n228), .A3(new_n239), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n240), .A2(KEYINPUT28), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  XNOR2_X1  g056(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n243));
  XNOR2_X1  g057(.A(new_n243), .B(G101), .ZN(new_n244));
  INV_X1    g058(.A(G237), .ZN(new_n245));
  INV_X1    g059(.A(G953), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n245), .A2(new_n246), .A3(G210), .ZN(new_n247));
  XNOR2_X1  g061(.A(new_n244), .B(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(new_n235), .ZN(new_n249));
  NOR3_X1   g063(.A1(new_n198), .A2(KEYINPUT65), .A3(new_n196), .ZN(new_n250));
  OAI21_X1  g064(.A(KEYINPUT65), .B1(new_n200), .B2(G146), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n251), .B1(new_n204), .B2(G146), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n249), .B1(new_n250), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n210), .A2(new_n211), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n237), .A2(G128), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n253), .A2(new_n256), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n257), .A2(KEYINPUT67), .A3(new_n229), .A4(new_n233), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT67), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n239), .A2(new_n259), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n258), .A2(new_n260), .A3(new_n215), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n240), .B1(new_n261), .B2(new_n224), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT28), .ZN(new_n263));
  OAI211_X1 g077(.A(new_n242), .B(new_n248), .C1(new_n262), .C2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT29), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n215), .A2(KEYINPUT30), .A3(new_n239), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT30), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n267), .B1(new_n261), .B2(new_n268), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n240), .B1(new_n269), .B2(new_n224), .ZN(new_n270));
  OAI211_X1 g084(.A(new_n264), .B(new_n265), .C1(new_n270), .C2(new_n248), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n215), .A2(new_n239), .ZN(new_n272));
  XOR2_X1   g086(.A(new_n272), .B(new_n228), .Z(new_n273));
  AOI21_X1  g087(.A(new_n241), .B1(new_n273), .B2(KEYINPUT28), .ZN(new_n274));
  INV_X1    g088(.A(new_n248), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n275), .A2(new_n265), .ZN(new_n276));
  AOI21_X1  g090(.A(G902), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n271), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(G472), .ZN(new_n279));
  NOR2_X1   g093(.A1(G472), .A2(G902), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n261), .A2(new_n268), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n282), .A2(new_n224), .A3(new_n266), .ZN(new_n283));
  INV_X1    g097(.A(new_n240), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n283), .A2(new_n284), .A3(new_n248), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n242), .B1(new_n262), .B2(new_n263), .ZN(new_n286));
  AOI22_X1  g100(.A1(new_n285), .A2(KEYINPUT31), .B1(new_n286), .B2(new_n275), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT31), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n270), .A2(new_n288), .A3(new_n248), .ZN(new_n289));
  AOI211_X1 g103(.A(KEYINPUT32), .B(new_n281), .C1(new_n287), .C2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT32), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n285), .A2(KEYINPUT31), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n286), .A2(new_n275), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n292), .A2(new_n289), .A3(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n291), .B1(new_n294), .B2(new_n280), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n279), .B1(new_n290), .B2(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(G214), .B1(G237), .B2(G902), .ZN(new_n297));
  INV_X1    g111(.A(G104), .ZN(new_n298));
  INV_X1    g112(.A(G107), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(KEYINPUT75), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT75), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(G107), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n300), .B1(new_n304), .B2(new_n298), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(G101), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT3), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(G104), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n308), .B1(new_n301), .B2(new_n303), .ZN(new_n309));
  OAI21_X1  g123(.A(G107), .B1(new_n298), .B2(KEYINPUT3), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n298), .A2(KEYINPUT3), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n309), .A2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(G101), .ZN(new_n314));
  AOI21_X1  g128(.A(KEYINPUT76), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT76), .ZN(new_n316));
  NOR4_X1   g130(.A1(new_n309), .A2(new_n312), .A3(new_n316), .A4(G101), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n306), .B1(new_n315), .B2(new_n317), .ZN(new_n318));
  OR2_X1    g132(.A1(new_n217), .A2(KEYINPUT5), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n217), .A2(new_n219), .A3(KEYINPUT5), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n319), .A2(G113), .A3(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT78), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n319), .A2(KEYINPUT78), .A3(new_n320), .A4(G113), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n323), .A2(new_n222), .A3(new_n324), .ZN(new_n325));
  OAI21_X1  g139(.A(KEYINPUT79), .B1(new_n318), .B2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(new_n325), .ZN(new_n327));
  AND2_X1   g141(.A1(new_n305), .A2(G101), .ZN(new_n328));
  XNOR2_X1  g142(.A(KEYINPUT75), .B(G107), .ZN(new_n329));
  OAI211_X1 g143(.A(new_n311), .B(new_n310), .C1(new_n329), .C2(new_n308), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n316), .B1(new_n330), .B2(G101), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n313), .A2(KEYINPUT76), .A3(new_n314), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n328), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT79), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n327), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n326), .A2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT77), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT4), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n330), .A2(new_n338), .A3(G101), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n331), .A2(new_n332), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n338), .B1(new_n330), .B2(G101), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n340), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n337), .B1(new_n343), .B2(new_n224), .ZN(new_n344));
  OAI21_X1  g158(.A(G101), .B1(new_n309), .B2(new_n312), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(KEYINPUT4), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n346), .B1(new_n331), .B2(new_n332), .ZN(new_n347));
  INV_X1    g161(.A(new_n224), .ZN(new_n348));
  NOR4_X1   g162(.A1(new_n347), .A2(KEYINPUT77), .A3(new_n348), .A4(new_n340), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n336), .B1(new_n344), .B2(new_n349), .ZN(new_n350));
  XOR2_X1   g164(.A(G110), .B(G122), .Z(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(new_n351), .ZN(new_n353));
  OAI211_X1 g167(.A(new_n336), .B(new_n353), .C1(new_n344), .C2(new_n349), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n352), .A2(KEYINPUT6), .A3(new_n354), .ZN(new_n355));
  AOI22_X1  g169(.A1(new_n208), .A2(new_n206), .B1(new_n212), .B2(new_n213), .ZN(new_n356));
  INV_X1    g170(.A(G125), .ZN(new_n357));
  OAI21_X1  g171(.A(KEYINPUT80), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n209), .A2(new_n214), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT80), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n359), .A2(new_n360), .A3(G125), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n253), .A2(new_n357), .A3(new_n256), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n358), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(G224), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n364), .A2(G953), .ZN(new_n365));
  XNOR2_X1  g179(.A(new_n363), .B(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT6), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n350), .A2(new_n367), .A3(new_n351), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n355), .A2(new_n366), .A3(new_n368), .ZN(new_n369));
  OAI21_X1  g183(.A(G210), .B1(G237), .B2(G902), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n342), .B1(new_n315), .B2(new_n317), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n371), .A2(new_n224), .A3(new_n339), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(KEYINPUT77), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n343), .A2(new_n337), .A3(new_n224), .ZN(new_n374));
  AOI22_X1  g188(.A1(new_n373), .A2(new_n374), .B1(new_n326), .B2(new_n335), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n363), .A2(new_n365), .ZN(new_n376));
  AOI22_X1  g190(.A1(new_n375), .A2(new_n353), .B1(new_n376), .B2(KEYINPUT7), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n333), .A2(new_n325), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n321), .A2(new_n222), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n378), .B1(new_n333), .B2(new_n379), .ZN(new_n380));
  XOR2_X1   g194(.A(new_n351), .B(KEYINPUT8), .Z(new_n381));
  OAI21_X1  g195(.A(KEYINPUT7), .B1(new_n364), .B2(G953), .ZN(new_n382));
  AOI22_X1  g196(.A1(new_n380), .A2(new_n381), .B1(new_n363), .B2(new_n382), .ZN(new_n383));
  AOI21_X1  g197(.A(G902), .B1(new_n377), .B2(new_n383), .ZN(new_n384));
  AND3_X1   g198(.A1(new_n369), .A2(new_n370), .A3(new_n384), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n370), .B1(new_n369), .B2(new_n384), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n297), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(G469), .ZN(new_n388));
  INV_X1    g202(.A(G902), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT10), .ZN(new_n390));
  INV_X1    g204(.A(new_n206), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n210), .A2(KEYINPUT1), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(G128), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n236), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n390), .B1(new_n318), .B2(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n371), .A2(new_n356), .A3(new_n339), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n333), .A2(KEYINPUT10), .A3(new_n257), .ZN(new_n397));
  INV_X1    g211(.A(new_n194), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n395), .A2(new_n396), .A3(new_n397), .A4(new_n398), .ZN(new_n399));
  XOR2_X1   g213(.A(G110), .B(G140), .Z(new_n400));
  XNOR2_X1  g214(.A(new_n400), .B(KEYINPUT73), .ZN(new_n401));
  AND2_X1   g215(.A1(new_n246), .A2(G227), .ZN(new_n402));
  XNOR2_X1  g216(.A(new_n401), .B(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n399), .A2(new_n403), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n318), .A2(new_n394), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n333), .A2(new_n257), .ZN(new_n406));
  OAI211_X1 g220(.A(KEYINPUT12), .B(new_n194), .C1(new_n405), .C2(new_n406), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n194), .B1(new_n405), .B2(new_n406), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT12), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n404), .B1(new_n407), .B2(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n395), .A2(new_n396), .A3(new_n397), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(new_n194), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n403), .B1(new_n413), .B2(new_n399), .ZN(new_n414));
  OAI211_X1 g228(.A(new_n388), .B(new_n389), .C1(new_n411), .C2(new_n414), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n388), .A2(new_n389), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  AND2_X1   g231(.A1(new_n399), .A2(new_n403), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(new_n413), .ZN(new_n419));
  AND3_X1   g233(.A1(new_n395), .A2(new_n396), .A3(new_n397), .ZN(new_n420));
  AOI22_X1  g234(.A1(new_n410), .A2(new_n407), .B1(new_n420), .B2(new_n398), .ZN(new_n421));
  XOR2_X1   g235(.A(new_n403), .B(KEYINPUT74), .Z(new_n422));
  OAI211_X1 g236(.A(new_n419), .B(G469), .C1(new_n421), .C2(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n415), .A2(new_n417), .A3(new_n423), .ZN(new_n424));
  XOR2_X1   g238(.A(KEYINPUT9), .B(G234), .Z(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  OAI21_X1  g240(.A(G221), .B1(new_n426), .B2(G902), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n424), .A2(new_n427), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n387), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT25), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT16), .ZN(new_n431));
  INV_X1    g245(.A(G140), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(G125), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n357), .A2(G140), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n433), .A2(new_n434), .A3(KEYINPUT70), .ZN(new_n435));
  OR3_X1    g249(.A1(new_n357), .A2(KEYINPUT70), .A3(G140), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n431), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n433), .A2(KEYINPUT16), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n196), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(new_n438), .ZN(new_n440));
  NOR3_X1   g254(.A1(new_n357), .A2(KEYINPUT70), .A3(G140), .ZN(new_n441));
  XNOR2_X1  g255(.A(G125), .B(G140), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n441), .B1(new_n442), .B2(KEYINPUT70), .ZN(new_n443));
  OAI211_X1 g257(.A(G146), .B(new_n440), .C1(new_n443), .C2(new_n431), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n439), .A2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(G128), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(G119), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n216), .A2(G128), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n449), .A2(KEYINPUT69), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT69), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n451), .B1(new_n447), .B2(new_n448), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  XOR2_X1   g267(.A(KEYINPUT24), .B(G110), .Z(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT23), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n447), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n446), .A2(KEYINPUT23), .A3(G119), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n457), .A2(new_n448), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(G110), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n445), .A2(new_n455), .A3(new_n460), .ZN(new_n461));
  OAI22_X1  g275(.A1(new_n453), .A2(new_n454), .B1(G110), .B2(new_n459), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n442), .A2(new_n196), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n462), .A2(new_n444), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(KEYINPUT72), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT72), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n461), .A2(new_n464), .A3(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n246), .A2(G221), .A3(G234), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n469), .B(KEYINPUT71), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT22), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n470), .B(new_n471), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n472), .B(G137), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n466), .A2(new_n468), .A3(new_n473), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n472), .B(new_n190), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n475), .A2(KEYINPUT72), .A3(new_n465), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n430), .B1(new_n477), .B2(new_n389), .ZN(new_n478));
  AOI211_X1 g292(.A(KEYINPUT25), .B(G902), .C1(new_n474), .C2(new_n476), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(G217), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n481), .B1(G234), .B2(new_n389), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n482), .A2(G902), .ZN(new_n483));
  AOI22_X1  g297(.A1(new_n480), .A2(new_n482), .B1(new_n477), .B2(new_n483), .ZN(new_n484));
  XNOR2_X1  g298(.A(G113), .B(G122), .ZN(new_n485));
  XNOR2_X1  g299(.A(new_n485), .B(new_n298), .ZN(new_n486));
  INV_X1    g300(.A(G214), .ZN(new_n487));
  NOR3_X1   g301(.A1(new_n487), .A2(G237), .A3(G953), .ZN(new_n488));
  OAI21_X1  g302(.A(KEYINPUT81), .B1(new_n198), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(G143), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT81), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n245), .A2(new_n246), .A3(G214), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n202), .A2(G143), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n200), .A2(KEYINPUT64), .ZN(new_n494));
  OAI211_X1 g308(.A(new_n491), .B(new_n492), .C1(new_n493), .C2(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n489), .A2(new_n490), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(G131), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT17), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n489), .A2(new_n193), .A3(new_n495), .A4(new_n490), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n497), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  AND2_X1   g314(.A1(new_n439), .A2(new_n444), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n496), .A2(KEYINPUT17), .A3(G131), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n500), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  AND3_X1   g317(.A1(new_n496), .A2(KEYINPUT18), .A3(G131), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT82), .ZN(new_n505));
  NAND2_X1  g319(.A1(KEYINPUT18), .A2(G131), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n489), .A2(new_n506), .A3(new_n495), .A4(new_n490), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n435), .A2(new_n436), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n463), .B1(new_n508), .B2(new_n196), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  NOR3_X1   g324(.A1(new_n504), .A2(new_n505), .A3(new_n510), .ZN(new_n511));
  AND2_X1   g325(.A1(new_n507), .A2(new_n509), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n496), .A2(KEYINPUT18), .A3(G131), .ZN(new_n513));
  AOI21_X1  g327(.A(KEYINPUT82), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  OAI211_X1 g328(.A(new_n486), .B(new_n503), .C1(new_n511), .C2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT85), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n505), .B1(new_n504), .B2(new_n510), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n512), .A2(KEYINPUT82), .A3(new_n513), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n486), .B1(new_n520), .B2(new_n503), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n517), .A2(new_n521), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n503), .B1(new_n511), .B2(new_n514), .ZN(new_n523));
  INV_X1    g337(.A(new_n486), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n523), .A2(KEYINPUT85), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(new_n389), .ZN(new_n526));
  OAI21_X1  g340(.A(KEYINPUT86), .B1(new_n522), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n523), .A2(new_n524), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n528), .A2(new_n516), .A3(new_n515), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT86), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n529), .A2(new_n530), .A3(new_n389), .A4(new_n525), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n527), .A2(G475), .A3(new_n531), .ZN(new_n532));
  NOR3_X1   g346(.A1(new_n426), .A2(new_n481), .A3(G953), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n204), .A2(G128), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n446), .A2(G143), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n187), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n446), .B1(new_n201), .B2(new_n203), .ZN(new_n538));
  INV_X1    g352(.A(new_n536), .ZN(new_n539));
  NOR3_X1   g353(.A1(new_n538), .A2(G134), .A3(new_n539), .ZN(new_n540));
  OAI21_X1  g354(.A(KEYINPUT90), .B1(new_n537), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n535), .A2(new_n187), .A3(new_n536), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT90), .ZN(new_n543));
  OAI21_X1  g357(.A(G134), .B1(new_n538), .B2(new_n539), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n541), .A2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(G122), .ZN(new_n547));
  OAI21_X1  g361(.A(KEYINPUT88), .B1(new_n547), .B2(G116), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT88), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n549), .A2(new_n218), .A3(G122), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  XNOR2_X1  g365(.A(KEYINPUT87), .B(G122), .ZN(new_n552));
  OAI211_X1 g366(.A(new_n551), .B(new_n304), .C1(new_n218), .C2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(KEYINPUT91), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n547), .A2(KEYINPUT87), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT87), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(G122), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n218), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT91), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n559), .A2(new_n560), .A3(new_n304), .A4(new_n551), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT14), .ZN(new_n562));
  AND3_X1   g376(.A1(new_n548), .A2(new_n550), .A3(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n562), .B1(new_n548), .B2(new_n550), .ZN(new_n564));
  NOR3_X1   g378(.A1(new_n563), .A2(new_n564), .A3(new_n558), .ZN(new_n565));
  OAI211_X1 g379(.A(new_n554), .B(new_n561), .C1(new_n565), .C2(new_n299), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n546), .A2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT13), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n568), .B1(new_n446), .B2(G143), .ZN(new_n569));
  OAI21_X1  g383(.A(KEYINPUT89), .B1(new_n538), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n538), .A2(KEYINPUT13), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT89), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n536), .A2(KEYINPUT13), .ZN(new_n573));
  OAI211_X1 g387(.A(new_n572), .B(new_n573), .C1(new_n198), .C2(new_n446), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n570), .A2(new_n571), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(G134), .ZN(new_n576));
  INV_X1    g390(.A(new_n551), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n329), .B1(new_n577), .B2(new_n558), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(new_n553), .ZN(new_n579));
  AND3_X1   g393(.A1(new_n576), .A2(new_n579), .A3(new_n542), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n534), .B1(new_n567), .B2(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n576), .A2(new_n579), .A3(new_n542), .ZN(new_n582));
  OAI211_X1 g396(.A(new_n582), .B(new_n533), .C1(new_n566), .C2(new_n546), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(new_n389), .ZN(new_n585));
  INV_X1    g399(.A(G478), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n586), .A2(KEYINPUT15), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n585), .B(new_n588), .ZN(new_n589));
  NOR2_X1   g403(.A1(G475), .A2(G902), .ZN(new_n590));
  INV_X1    g404(.A(new_n515), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n497), .A2(new_n499), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(KEYINPUT83), .ZN(new_n593));
  INV_X1    g407(.A(new_n442), .ZN(new_n594));
  MUX2_X1   g408(.A(new_n594), .B(new_n508), .S(KEYINPUT19), .Z(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(new_n196), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT83), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n497), .A2(new_n597), .A3(new_n499), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n593), .A2(new_n444), .A3(new_n596), .A4(new_n598), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n486), .B1(new_n599), .B2(new_n520), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n590), .B1(new_n591), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(KEYINPUT20), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT84), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT20), .ZN(new_n604));
  OAI211_X1 g418(.A(new_n604), .B(new_n590), .C1(new_n591), .C2(new_n600), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n602), .A2(new_n603), .A3(new_n605), .ZN(new_n606));
  OR2_X1    g420(.A1(new_n605), .A2(new_n603), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n532), .A2(new_n589), .A3(new_n606), .A4(new_n607), .ZN(new_n608));
  AND2_X1   g422(.A1(new_n246), .A2(G952), .ZN(new_n609));
  INV_X1    g423(.A(G234), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n609), .B1(new_n610), .B2(new_n245), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  OAI211_X1 g426(.A(G902), .B(G953), .C1(new_n610), .C2(new_n245), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n613), .B(KEYINPUT92), .ZN(new_n614));
  XNOR2_X1  g428(.A(KEYINPUT21), .B(G898), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n612), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n608), .A2(new_n616), .ZN(new_n617));
  AND4_X1   g431(.A1(new_n296), .A2(new_n429), .A3(new_n484), .A4(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(new_n314), .ZN(G3));
  NAND2_X1  g433(.A1(new_n294), .A2(new_n280), .ZN(new_n620));
  AOI21_X1  g434(.A(G902), .B1(new_n287), .B2(new_n289), .ZN(new_n621));
  INV_X1    g435(.A(G472), .ZN(new_n622));
  OAI211_X1 g436(.A(new_n484), .B(new_n620), .C1(new_n621), .C2(new_n622), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n623), .A2(new_n428), .ZN(new_n624));
  INV_X1    g438(.A(new_n616), .ZN(new_n625));
  OAI211_X1 g439(.A(new_n297), .B(new_n625), .C1(new_n385), .C2(new_n386), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT33), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT93), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n627), .B1(new_n583), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n584), .A2(new_n629), .ZN(new_n630));
  OAI211_X1 g444(.A(new_n581), .B(new_n583), .C1(new_n628), .C2(new_n627), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n632), .A2(G478), .A3(new_n389), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT94), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n585), .A2(new_n586), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n632), .A2(KEYINPUT94), .A3(G478), .A4(new_n389), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n635), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n532), .A2(new_n607), .A3(new_n606), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n626), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n624), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT34), .B(G104), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(KEYINPUT95), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n642), .B(new_n644), .ZN(G6));
  INV_X1    g459(.A(new_n589), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n602), .A2(new_n605), .ZN(new_n647));
  AND3_X1   g461(.A1(new_n646), .A2(new_n647), .A3(new_n532), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  OAI21_X1  g463(.A(KEYINPUT96), .B1(new_n626), .B2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n297), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n369), .A2(new_n384), .ZN(new_n652));
  INV_X1    g466(.A(new_n370), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n369), .A2(new_n370), .A3(new_n384), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n651), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT96), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n656), .A2(new_n657), .A3(new_n625), .A4(new_n648), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n650), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(new_n624), .ZN(new_n660));
  XOR2_X1   g474(.A(KEYINPUT35), .B(G107), .Z(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G9));
  AOI21_X1  g476(.A(new_n281), .B1(new_n287), .B2(new_n289), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n294), .A2(new_n389), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n663), .B1(new_n664), .B2(G472), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n480), .A2(new_n482), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT36), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n475), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(KEYINPUT97), .ZN(new_n669));
  OR2_X1    g483(.A1(new_n669), .A2(new_n465), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n669), .A2(new_n465), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n670), .A2(new_n671), .A3(new_n483), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n666), .A2(new_n672), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n429), .A2(new_n617), .A3(new_n665), .A4(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(KEYINPUT98), .B(KEYINPUT37), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G110), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n674), .B(new_n676), .ZN(G12));
  INV_X1    g491(.A(new_n428), .ZN(new_n678));
  AND4_X1   g492(.A1(new_n296), .A2(new_n656), .A3(new_n678), .A4(new_n673), .ZN(new_n679));
  INV_X1    g493(.A(G900), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n612), .B1(new_n614), .B2(new_n680), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n649), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G128), .ZN(G30));
  AND2_X1   g498(.A1(new_n666), .A2(new_n672), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n685), .A2(new_n297), .A3(new_n646), .A4(new_n639), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT99), .ZN(new_n687));
  OR2_X1    g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n270), .A2(new_n275), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n389), .B1(new_n273), .B2(new_n248), .ZN(new_n690));
  OAI21_X1  g504(.A(G472), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  OAI21_X1  g505(.A(new_n691), .B1(new_n290), .B2(new_n295), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n385), .A2(new_n386), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(KEYINPUT38), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT38), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n695), .B1(new_n385), .B2(new_n386), .ZN(new_n696));
  AND2_X1   g510(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n686), .A2(new_n687), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n688), .A2(new_n692), .A3(new_n697), .A4(new_n698), .ZN(new_n699));
  XOR2_X1   g513(.A(new_n681), .B(KEYINPUT39), .Z(new_n700));
  NAND2_X1  g514(.A1(new_n678), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(KEYINPUT40), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(new_n204), .ZN(G45));
  NAND2_X1  g518(.A1(new_n620), .A2(KEYINPUT32), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n663), .A2(new_n291), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n685), .B1(new_n707), .B2(new_n279), .ZN(new_n708));
  INV_X1    g522(.A(new_n681), .ZN(new_n709));
  AND3_X1   g523(.A1(new_n638), .A2(new_n639), .A3(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT100), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n710), .A2(new_n711), .A3(new_n656), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n638), .A2(new_n639), .A3(new_n709), .ZN(new_n713));
  OAI21_X1  g527(.A(KEYINPUT100), .B1(new_n713), .B2(new_n387), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n708), .A2(new_n712), .A3(new_n714), .A4(new_n678), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G146), .ZN(G48));
  INV_X1    g530(.A(new_n414), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n410), .A2(new_n407), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(new_n418), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n388), .B1(new_n720), .B2(new_n389), .ZN(new_n721));
  INV_X1    g535(.A(new_n415), .ZN(new_n722));
  INV_X1    g536(.A(new_n427), .ZN(new_n723));
  NOR3_X1   g537(.A1(new_n721), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  AND3_X1   g538(.A1(new_n296), .A2(new_n484), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(new_n641), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(KEYINPUT101), .ZN(new_n727));
  XOR2_X1   g541(.A(KEYINPUT41), .B(G113), .Z(new_n728));
  XNOR2_X1  g542(.A(new_n727), .B(new_n728), .ZN(G15));
  NAND2_X1  g543(.A1(new_n659), .A2(new_n725), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G116), .ZN(G18));
  AND3_X1   g545(.A1(new_n656), .A2(KEYINPUT102), .A3(new_n724), .ZN(new_n732));
  AOI21_X1  g546(.A(KEYINPUT102), .B1(new_n656), .B2(new_n724), .ZN(new_n733));
  OAI211_X1 g547(.A(new_n617), .B(new_n708), .C1(new_n732), .C2(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(KEYINPUT103), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G119), .ZN(G21));
  NOR2_X1   g550(.A1(new_n274), .A2(new_n248), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n288), .B1(new_n270), .B2(new_n248), .ZN(new_n738));
  OAI21_X1  g552(.A(KEYINPUT105), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT105), .ZN(new_n740));
  OAI211_X1 g554(.A(new_n292), .B(new_n740), .C1(new_n248), .C2(new_n274), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n739), .A2(new_n741), .A3(new_n289), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n280), .B(KEYINPUT104), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n664), .A2(G472), .ZN(new_n745));
  AND4_X1   g559(.A1(new_n484), .A2(new_n744), .A3(new_n724), .A4(new_n745), .ZN(new_n746));
  AND3_X1   g560(.A1(new_n639), .A2(KEYINPUT106), .A3(new_n646), .ZN(new_n747));
  AOI21_X1  g561(.A(KEYINPUT106), .B1(new_n639), .B2(new_n646), .ZN(new_n748));
  NOR3_X1   g562(.A1(new_n747), .A2(new_n626), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n746), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G122), .ZN(G24));
  AND3_X1   g565(.A1(new_n744), .A2(new_n745), .A3(new_n673), .ZN(new_n752));
  OAI211_X1 g566(.A(new_n710), .B(new_n752), .C1(new_n732), .C2(new_n733), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G125), .ZN(G27));
  NOR3_X1   g568(.A1(new_n385), .A2(new_n386), .A3(new_n651), .ZN(new_n755));
  AND3_X1   g569(.A1(new_n296), .A2(new_n484), .A3(new_n755), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n756), .A2(KEYINPUT42), .A3(new_n678), .A4(new_n710), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT42), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n296), .A2(new_n755), .A3(new_n484), .A4(new_n678), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n758), .B1(new_n759), .B2(new_n713), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n757), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G131), .ZN(G33));
  NOR3_X1   g576(.A1(new_n759), .A2(new_n649), .A3(new_n681), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(new_n187), .ZN(G36));
  OAI21_X1  g578(.A(new_n419), .B1(new_n421), .B2(new_n422), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT45), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  OAI211_X1 g581(.A(new_n419), .B(KEYINPUT45), .C1(new_n421), .C2(new_n422), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n767), .A2(G469), .A3(new_n768), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n769), .A2(KEYINPUT46), .A3(new_n417), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT107), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n769), .A2(KEYINPUT107), .A3(KEYINPUT46), .A4(new_n417), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n772), .A2(new_n415), .A3(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT108), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n772), .A2(KEYINPUT108), .A3(new_n415), .A4(new_n773), .ZN(new_n777));
  INV_X1    g591(.A(new_n769), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n778), .A2(new_n416), .ZN(new_n779));
  OAI211_X1 g593(.A(new_n776), .B(new_n777), .C1(KEYINPUT46), .C2(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(new_n427), .ZN(new_n781));
  INV_X1    g595(.A(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(new_n755), .ZN(new_n783));
  AND3_X1   g597(.A1(new_n532), .A2(new_n607), .A3(new_n606), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(new_n638), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT43), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n784), .A2(KEYINPUT43), .A3(new_n638), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n665), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(new_n673), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT44), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n783), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n789), .A2(KEYINPUT44), .A3(new_n673), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n782), .A2(new_n700), .A3(new_n792), .A4(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(G137), .ZN(G39));
  INV_X1    g609(.A(KEYINPUT47), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n781), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n780), .A2(KEYINPUT47), .A3(new_n427), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NOR3_X1   g613(.A1(new_n783), .A2(new_n296), .A3(new_n484), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n799), .A2(new_n710), .A3(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(G140), .ZN(G42));
  AOI21_X1  g616(.A(new_n611), .B1(new_n787), .B2(new_n788), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n755), .A2(new_n724), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n744), .A2(new_n745), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n805), .A2(new_n685), .A3(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n484), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n803), .A2(new_n809), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n810), .A2(new_n783), .ZN(new_n811));
  XOR2_X1   g625(.A(new_n811), .B(KEYINPUT114), .Z(new_n812));
  OR2_X1    g626(.A1(new_n721), .A2(new_n722), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n813), .A2(new_n427), .ZN(new_n814));
  INV_X1    g628(.A(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n797), .A2(new_n798), .A3(new_n815), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n807), .B1(new_n812), .B2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(new_n692), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n804), .A2(new_n484), .A3(new_n612), .A4(new_n818), .ZN(new_n819));
  OR3_X1    g633(.A1(new_n819), .A2(new_n639), .A3(new_n638), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n724), .A2(new_n651), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n697), .B1(KEYINPUT115), .B2(new_n821), .ZN(new_n822));
  OR2_X1    g636(.A1(new_n821), .A2(KEYINPUT115), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n822), .A2(new_n809), .A3(new_n803), .A4(new_n823), .ZN(new_n824));
  XOR2_X1   g638(.A(new_n824), .B(KEYINPUT50), .Z(new_n825));
  NAND4_X1  g639(.A1(new_n817), .A2(KEYINPUT51), .A3(new_n820), .A4(new_n825), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n826), .B(KEYINPUT116), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n817), .A2(new_n820), .A3(new_n825), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT51), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT53), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n747), .A2(new_n748), .A3(new_n387), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT110), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n673), .B1(new_n707), .B2(new_n691), .ZN(new_n834));
  AND3_X1   g648(.A1(new_n424), .A2(new_n427), .A3(new_n709), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n832), .A2(new_n833), .A3(new_n834), .A4(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n639), .A2(new_n646), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT106), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n639), .A2(KEYINPUT106), .A3(new_n646), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n839), .A2(new_n656), .A3(new_n840), .A4(new_n835), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n692), .A2(new_n685), .ZN(new_n842));
  OAI21_X1  g656(.A(KEYINPUT110), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  AND2_X1   g657(.A1(new_n836), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n296), .A2(new_n673), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n713), .A2(new_n387), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n845), .B1(new_n711), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n710), .A2(new_n656), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n428), .B1(new_n848), .B2(KEYINPUT100), .ZN(new_n849));
  AOI22_X1  g663(.A1(new_n847), .A2(new_n849), .B1(new_n682), .B2(new_n679), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n844), .A2(KEYINPUT52), .A3(new_n753), .A4(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT52), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n753), .A2(new_n683), .A3(new_n715), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n836), .A2(new_n843), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n852), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  AND2_X1   g669(.A1(new_n851), .A2(new_n855), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n656), .A2(new_n617), .A3(new_n678), .A4(new_n665), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n639), .A2(new_n589), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n656), .A2(new_n625), .A3(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n665), .A2(new_n678), .A3(new_n484), .ZN(new_n860));
  OAI22_X1  g674(.A1(new_n857), .A2(new_n685), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT109), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n642), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n784), .A2(new_n646), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n626), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n865), .A2(new_n624), .ZN(new_n866));
  AOI21_X1  g680(.A(KEYINPUT109), .B1(new_n674), .B2(new_n866), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n863), .A2(new_n618), .A3(new_n867), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n532), .A2(new_n647), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n296), .A2(new_n589), .A3(new_n869), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n870), .B1(new_n640), .B2(new_n806), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n871), .A2(new_n673), .A3(new_n755), .A4(new_n835), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n763), .B1(new_n757), .B2(new_n760), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n730), .A2(new_n734), .A3(new_n726), .A4(new_n750), .ZN(new_n874));
  INV_X1    g688(.A(new_n874), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n868), .A2(new_n872), .A3(new_n873), .A4(new_n875), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n831), .B1(new_n856), .B2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(new_n763), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n761), .A2(new_n872), .A3(KEYINPUT53), .A4(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT113), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n874), .A2(new_n880), .ZN(new_n881));
  AOI22_X1  g695(.A1(new_n659), .A2(new_n725), .B1(new_n746), .B2(new_n749), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n882), .A2(KEYINPUT113), .A3(new_n726), .A4(new_n734), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n879), .B1(new_n881), .B2(new_n883), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n851), .A2(KEYINPUT111), .A3(new_n855), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT111), .ZN(new_n886));
  OAI211_X1 g700(.A(new_n886), .B(new_n852), .C1(new_n853), .C2(new_n854), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n884), .A2(new_n885), .A3(new_n868), .A4(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT54), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n877), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n890), .A2(KEYINPUT112), .ZN(new_n891));
  INV_X1    g705(.A(new_n876), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n892), .A2(new_n831), .A3(new_n887), .A4(new_n885), .ZN(new_n893));
  OAI21_X1  g707(.A(KEYINPUT53), .B1(new_n856), .B2(new_n876), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n893), .A2(KEYINPUT54), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n891), .A2(new_n895), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n893), .A2(KEYINPUT112), .A3(KEYINPUT54), .A4(new_n894), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n827), .A2(new_n830), .A3(new_n896), .A4(new_n897), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n732), .A2(new_n733), .ZN(new_n899));
  OAI221_X1 g713(.A(new_n609), .B1(new_n819), .B2(new_n640), .C1(new_n810), .C2(new_n899), .ZN(new_n900));
  XOR2_X1   g714(.A(new_n900), .B(KEYINPUT117), .Z(new_n901));
  NAND2_X1  g715(.A1(new_n296), .A2(new_n484), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n805), .A2(new_n902), .ZN(new_n903));
  OR2_X1    g717(.A1(new_n903), .A2(KEYINPUT48), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n903), .A2(KEYINPUT48), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n901), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(KEYINPUT118), .ZN(new_n907));
  OAI22_X1  g721(.A1(new_n898), .A2(new_n907), .B1(G952), .B2(G953), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n813), .B(KEYINPUT49), .ZN(new_n909));
  NOR4_X1   g723(.A1(new_n909), .A2(new_n808), .A3(new_n651), .A4(new_n785), .ZN(new_n910));
  INV_X1    g724(.A(new_n697), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n910), .A2(new_n427), .A3(new_n818), .A4(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n908), .A2(new_n912), .ZN(G75));
  AOI21_X1  g727(.A(new_n389), .B1(new_n877), .B2(new_n888), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(G210), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT56), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(KEYINPUT55), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n355), .A2(new_n368), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n919), .B(new_n366), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n920), .B(KEYINPUT119), .ZN(new_n921));
  INV_X1    g735(.A(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT55), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n915), .A2(new_n923), .A3(new_n916), .ZN(new_n924));
  AND3_X1   g738(.A1(new_n918), .A2(new_n922), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n922), .B1(new_n918), .B2(new_n924), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n246), .A2(G952), .ZN(new_n927));
  NOR3_X1   g741(.A1(new_n925), .A2(new_n926), .A3(new_n927), .ZN(G51));
  NAND2_X1  g742(.A1(new_n877), .A2(new_n888), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n929), .A2(KEYINPUT54), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(new_n890), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT57), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n931), .B1(new_n932), .B2(new_n416), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n417), .A2(KEYINPUT57), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n720), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n914), .A2(new_n778), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n927), .B1(new_n935), .B2(new_n936), .ZN(G54));
  NAND3_X1  g751(.A1(new_n914), .A2(KEYINPUT58), .A3(G475), .ZN(new_n938));
  OR2_X1    g752(.A1(new_n591), .A2(new_n600), .ZN(new_n939));
  INV_X1    g753(.A(new_n939), .ZN(new_n940));
  AND2_X1   g754(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n938), .A2(new_n940), .ZN(new_n942));
  NOR3_X1   g756(.A1(new_n941), .A2(new_n942), .A3(new_n927), .ZN(G60));
  NAND2_X1  g757(.A1(G478), .A2(G902), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n944), .B(KEYINPUT59), .Z(new_n945));
  AOI21_X1  g759(.A(new_n945), .B1(new_n630), .B2(new_n631), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n927), .B1(new_n931), .B2(new_n946), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n945), .B1(new_n896), .B2(new_n897), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n947), .B1(new_n948), .B2(new_n632), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT120), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  OAI211_X1 g765(.A(new_n947), .B(KEYINPUT120), .C1(new_n948), .C2(new_n632), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n951), .A2(new_n952), .ZN(G63));
  NAND2_X1  g767(.A1(G217), .A2(G902), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(KEYINPUT121), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n955), .B(KEYINPUT60), .ZN(new_n956));
  AND2_X1   g770(.A1(new_n929), .A2(new_n956), .ZN(new_n957));
  AND3_X1   g771(.A1(new_n957), .A2(new_n670), .A3(new_n671), .ZN(new_n958));
  INV_X1    g772(.A(new_n927), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n477), .B(KEYINPUT123), .ZN(new_n960));
  INV_X1    g774(.A(new_n960), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n959), .B1(new_n957), .B2(new_n961), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n958), .A2(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT122), .ZN(new_n964));
  OAI211_X1 g778(.A(new_n964), .B(new_n959), .C1(new_n957), .C2(new_n961), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT61), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n963), .B(new_n967), .ZN(G66));
  NAND2_X1  g782(.A1(new_n868), .A2(new_n875), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n969), .A2(new_n246), .ZN(new_n970));
  OAI21_X1  g784(.A(G953), .B1(new_n615), .B2(new_n364), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n919), .B1(G898), .B2(new_n246), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n972), .B(new_n973), .ZN(G69));
  XNOR2_X1  g788(.A(new_n269), .B(new_n595), .ZN(new_n975));
  NAND2_X1  g789(.A1(G900), .A2(G953), .ZN(new_n976));
  OR2_X1    g790(.A1(new_n873), .A2(KEYINPUT124), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n873), .A2(KEYINPUT124), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n853), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NOR4_X1   g793(.A1(new_n902), .A2(new_n387), .A3(new_n748), .A4(new_n747), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n782), .A2(new_n700), .A3(new_n980), .ZN(new_n981));
  NAND4_X1  g795(.A1(new_n801), .A2(new_n794), .A3(new_n979), .A4(new_n981), .ZN(new_n982));
  OAI211_X1 g796(.A(new_n975), .B(new_n976), .C1(new_n982), .C2(G953), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT62), .ZN(new_n984));
  OR3_X1    g798(.A1(new_n703), .A2(new_n984), .A3(new_n853), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n984), .B1(new_n703), .B2(new_n853), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n701), .B1(new_n640), .B2(new_n864), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n988), .A2(new_n756), .ZN(new_n989));
  NAND4_X1  g803(.A1(new_n801), .A2(new_n987), .A3(new_n794), .A4(new_n989), .ZN(new_n990));
  INV_X1    g804(.A(new_n990), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n991), .A2(G953), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n983), .B1(new_n992), .B2(new_n975), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n246), .B1(G227), .B2(G900), .ZN(new_n994));
  XNOR2_X1  g808(.A(new_n993), .B(new_n994), .ZN(G72));
  NAND2_X1  g809(.A1(G472), .A2(G902), .ZN(new_n996));
  XOR2_X1   g810(.A(new_n996), .B(KEYINPUT63), .Z(new_n997));
  OAI21_X1  g811(.A(new_n997), .B1(new_n990), .B2(new_n969), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n998), .A2(KEYINPUT125), .ZN(new_n999));
  INV_X1    g813(.A(KEYINPUT125), .ZN(new_n1000));
  OAI211_X1 g814(.A(new_n1000), .B(new_n997), .C1(new_n990), .C2(new_n969), .ZN(new_n1001));
  AND3_X1   g815(.A1(new_n999), .A2(new_n689), .A3(new_n1001), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n997), .B1(new_n982), .B2(new_n969), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n1003), .A2(new_n270), .A3(new_n275), .ZN(new_n1004));
  XNOR2_X1  g818(.A(new_n270), .B(new_n248), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1005), .A2(new_n997), .ZN(new_n1006));
  XNOR2_X1  g820(.A(new_n1006), .B(KEYINPUT126), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n893), .A2(new_n894), .A3(new_n1007), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n1004), .A2(new_n959), .A3(new_n1008), .ZN(new_n1009));
  OR3_X1    g823(.A1(new_n1002), .A2(new_n1009), .A3(KEYINPUT127), .ZN(new_n1010));
  OAI21_X1  g824(.A(KEYINPUT127), .B1(new_n1002), .B2(new_n1009), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1010), .A2(new_n1011), .ZN(G57));
endmodule


