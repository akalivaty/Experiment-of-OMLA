//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 1 0 0 1 1 0 0 0 0 1 0 0 1 1 0 0 0 0 0 0 1 1 1 0 1 0 0 0 1 1 1 0 1 0 1 1 0 0 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:44 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n712, new_n713, new_n714, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n730, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n795, new_n796, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062;
  INV_X1    g000(.A(G953), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G227), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT76), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n188), .B(new_n189), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n190), .B(G110), .ZN(new_n191));
  OR2_X1    g005(.A1(new_n191), .A2(G140), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(G140), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G104), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G107), .ZN(new_n196));
  OR2_X1    g010(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n197));
  INV_X1    g011(.A(G107), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G104), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n196), .B1(new_n197), .B2(new_n199), .ZN(new_n200));
  NOR2_X1   g014(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n195), .A2(G107), .ZN(new_n202));
  NAND2_X1  g016(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n201), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  OAI21_X1  g018(.A(G101), .B1(new_n200), .B2(new_n204), .ZN(new_n205));
  AND2_X1   g019(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n197), .B1(new_n199), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G101), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n202), .A2(new_n201), .ZN(new_n209));
  NAND4_X1  g023(.A1(new_n207), .A2(new_n208), .A3(new_n196), .A4(new_n209), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n205), .A2(KEYINPUT4), .A3(new_n210), .ZN(new_n211));
  XNOR2_X1  g025(.A(G143), .B(G146), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n212), .A2(KEYINPUT0), .A3(G128), .ZN(new_n213));
  XNOR2_X1  g027(.A(KEYINPUT0), .B(G128), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n213), .B1(new_n212), .B2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT4), .ZN(new_n217));
  OAI211_X1 g031(.A(new_n217), .B(G101), .C1(new_n200), .C2(new_n204), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n211), .A2(new_n216), .A3(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT79), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n211), .A2(KEYINPUT79), .A3(new_n216), .A4(new_n218), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G137), .ZN(new_n224));
  OAI21_X1  g038(.A(KEYINPUT65), .B1(new_n224), .B2(G134), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT65), .ZN(new_n226));
  INV_X1    g040(.A(G134), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n226), .A2(new_n227), .A3(G137), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n225), .A2(new_n228), .ZN(new_n229));
  OAI211_X1 g043(.A(KEYINPUT64), .B(KEYINPUT11), .C1(new_n227), .C2(G137), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n224), .A2(G134), .ZN(new_n232));
  AOI21_X1  g046(.A(KEYINPUT11), .B1(new_n232), .B2(KEYINPUT64), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n229), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(G131), .ZN(new_n235));
  INV_X1    g049(.A(G131), .ZN(new_n236));
  OAI211_X1 g050(.A(new_n236), .B(new_n229), .C1(new_n231), .C2(new_n233), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  XNOR2_X1  g052(.A(new_n238), .B(KEYINPUT80), .ZN(new_n239));
  INV_X1    g053(.A(G128), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n240), .A2(KEYINPUT1), .ZN(new_n241));
  INV_X1    g055(.A(G146), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G143), .ZN(new_n243));
  INV_X1    g057(.A(G143), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G146), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n241), .A2(new_n243), .A3(new_n245), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n244), .A2(KEYINPUT1), .A3(G146), .ZN(new_n247));
  OAI211_X1 g061(.A(new_n246), .B(new_n247), .C1(G128), .C2(new_n212), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n199), .A2(new_n196), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G101), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n248), .A2(new_n210), .A3(new_n250), .ZN(new_n251));
  OR2_X1    g065(.A1(new_n251), .A2(KEYINPUT10), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(KEYINPUT10), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n223), .A2(new_n239), .A3(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT81), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n223), .A2(new_n256), .A3(new_n254), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(new_n238), .ZN(new_n258));
  AOI22_X1  g072(.A1(new_n221), .A2(new_n222), .B1(new_n253), .B2(new_n252), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n259), .A2(new_n256), .ZN(new_n260));
  OAI211_X1 g074(.A(new_n194), .B(new_n255), .C1(new_n258), .C2(new_n260), .ZN(new_n261));
  AND3_X1   g075(.A1(new_n248), .A2(new_n210), .A3(new_n250), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n248), .B1(new_n210), .B2(new_n250), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n238), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(KEYINPUT12), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT12), .ZN(new_n266));
  OAI211_X1 g080(.A(new_n238), .B(new_n266), .C1(new_n262), .C2(new_n263), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT77), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n270), .B1(new_n192), .B2(new_n193), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(G140), .ZN(new_n273));
  XNOR2_X1  g087(.A(new_n191), .B(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(new_n270), .ZN(new_n275));
  AOI22_X1  g089(.A1(new_n269), .A2(new_n255), .B1(new_n272), .B2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  AOI21_X1  g091(.A(G902), .B1(new_n261), .B2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(G469), .ZN(new_n279));
  OAI21_X1  g093(.A(KEYINPUT82), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT82), .ZN(new_n281));
  AND3_X1   g095(.A1(new_n223), .A2(new_n254), .A3(new_n239), .ZN(new_n282));
  INV_X1    g096(.A(new_n238), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n283), .B1(new_n259), .B2(new_n256), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n223), .A2(new_n254), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(KEYINPUT81), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n282), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n276), .B1(new_n287), .B2(new_n194), .ZN(new_n288));
  OAI211_X1 g102(.A(new_n281), .B(G469), .C1(new_n288), .C2(G902), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n268), .B1(new_n259), .B2(new_n239), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(new_n194), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n291), .B1(new_n287), .B2(new_n194), .ZN(new_n292));
  INV_X1    g106(.A(G902), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n292), .A2(new_n279), .A3(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n280), .A2(new_n289), .A3(new_n294), .ZN(new_n295));
  OAI21_X1  g109(.A(G214), .B1(G237), .B2(G902), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT5), .ZN(new_n298));
  INV_X1    g112(.A(G119), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n298), .A2(new_n299), .A3(G116), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT67), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n301), .B1(new_n299), .B2(G116), .ZN(new_n302));
  INV_X1    g116(.A(G116), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n303), .A2(KEYINPUT67), .A3(G119), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n299), .A2(G116), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  OAI211_X1 g121(.A(G113), .B(new_n300), .C1(new_n307), .C2(new_n298), .ZN(new_n308));
  AOI22_X1  g122(.A1(new_n302), .A2(new_n304), .B1(G116), .B2(new_n299), .ZN(new_n309));
  XOR2_X1   g123(.A(KEYINPUT2), .B(G113), .Z(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n308), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n210), .A2(new_n250), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND4_X1  g128(.A1(new_n308), .A2(new_n210), .A3(new_n250), .A4(new_n311), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  XNOR2_X1  g130(.A(G110), .B(G122), .ZN(new_n317));
  XOR2_X1   g131(.A(new_n317), .B(KEYINPUT8), .Z(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n316), .A2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(G125), .ZN(new_n321));
  OR2_X1    g135(.A1(new_n212), .A2(new_n214), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n321), .B1(new_n322), .B2(new_n213), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n248), .A2(G125), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(G224), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n327), .A2(G953), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT7), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n324), .A2(new_n326), .A3(new_n330), .ZN(new_n331));
  OAI22_X1  g145(.A1(new_n323), .A2(new_n325), .B1(new_n329), .B2(new_n328), .ZN(new_n332));
  AND2_X1   g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT83), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n320), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n318), .B1(new_n314), .B2(new_n315), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n331), .A2(new_n332), .ZN(new_n337));
  OAI21_X1  g151(.A(KEYINPUT83), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(new_n310), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT66), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n307), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n310), .B1(new_n309), .B2(KEYINPUT66), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n343), .A2(new_n211), .A3(new_n218), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n344), .A2(new_n315), .A3(new_n317), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n335), .A2(new_n338), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n344), .A2(new_n315), .ZN(new_n347));
  INV_X1    g161(.A(new_n317), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n349), .A2(KEYINPUT6), .A3(new_n345), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n324), .A2(new_n326), .ZN(new_n351));
  XNOR2_X1  g165(.A(new_n351), .B(new_n328), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT6), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n347), .A2(new_n353), .A3(new_n348), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n350), .A2(new_n352), .A3(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n346), .A2(new_n355), .A3(new_n293), .ZN(new_n356));
  OAI21_X1  g170(.A(G210), .B1(G237), .B2(G902), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n346), .A2(new_n355), .A3(new_n293), .A4(new_n357), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n297), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  XOR2_X1   g175(.A(KEYINPUT9), .B(G234), .Z(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  OAI21_X1  g177(.A(G221), .B1(new_n363), .B2(G902), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n295), .A2(new_n361), .A3(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT30), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n215), .B1(new_n235), .B2(new_n237), .ZN(new_n367));
  INV_X1    g181(.A(new_n232), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n224), .A2(G134), .ZN(new_n369));
  OAI21_X1  g183(.A(G131), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  AND3_X1   g184(.A1(new_n237), .A2(new_n248), .A3(new_n370), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n366), .B1(new_n367), .B2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(new_n237), .ZN(new_n373));
  OAI21_X1  g187(.A(KEYINPUT64), .B1(new_n227), .B2(G137), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT11), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(new_n230), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n236), .B1(new_n377), .B2(new_n229), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n216), .B1(new_n373), .B2(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n237), .A2(new_n248), .A3(new_n370), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n379), .A2(KEYINPUT30), .A3(new_n380), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n372), .A2(new_n381), .A3(new_n343), .ZN(new_n382));
  INV_X1    g196(.A(G237), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n383), .A2(new_n187), .A3(G210), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT27), .ZN(new_n385));
  XNOR2_X1  g199(.A(new_n384), .B(new_n385), .ZN(new_n386));
  XNOR2_X1  g200(.A(new_n386), .B(KEYINPUT26), .ZN(new_n387));
  XNOR2_X1  g201(.A(new_n387), .B(new_n208), .ZN(new_n388));
  INV_X1    g202(.A(new_n343), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n379), .A2(new_n389), .A3(new_n380), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n382), .A2(new_n388), .A3(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT68), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND4_X1  g207(.A1(new_n382), .A2(KEYINPUT68), .A3(new_n388), .A4(new_n390), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n393), .A2(KEYINPUT31), .A3(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT31), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n391), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT28), .ZN(new_n399));
  OR2_X1    g213(.A1(new_n390), .A2(new_n399), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n343), .B1(new_n367), .B2(new_n371), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n390), .A2(new_n399), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n400), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n388), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n398), .A2(new_n405), .ZN(new_n406));
  NOR2_X1   g220(.A1(G472), .A2(G902), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n406), .A2(KEYINPUT32), .A3(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT32), .ZN(new_n409));
  AOI22_X1  g223(.A1(new_n395), .A2(new_n397), .B1(new_n404), .B2(new_n403), .ZN(new_n410));
  INV_X1    g224(.A(new_n407), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n409), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT29), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n413), .B1(new_n403), .B2(new_n404), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n382), .A2(new_n390), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n416), .A2(new_n388), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n293), .B1(new_n414), .B2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT70), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n401), .A2(new_n419), .ZN(new_n420));
  OAI211_X1 g234(.A(KEYINPUT70), .B(new_n343), .C1(new_n367), .C2(new_n371), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT69), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n390), .A2(new_n423), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n379), .A2(new_n389), .A3(KEYINPUT69), .A4(new_n380), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n399), .B1(new_n422), .B2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n402), .ZN(new_n428));
  NOR4_X1   g242(.A1(new_n427), .A2(new_n413), .A3(new_n404), .A4(new_n428), .ZN(new_n429));
  OAI21_X1  g243(.A(G472), .B1(new_n418), .B2(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n408), .A2(new_n412), .A3(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(G217), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n432), .B1(G234), .B2(new_n293), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  OR3_X1    g248(.A1(new_n299), .A2(KEYINPUT71), .A3(G128), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n299), .A2(G128), .ZN(new_n436));
  AOI21_X1  g250(.A(KEYINPUT71), .B1(new_n299), .B2(G128), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n435), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  OR2_X1    g252(.A1(KEYINPUT24), .A2(G110), .ZN(new_n439));
  NAND2_X1  g253(.A1(KEYINPUT24), .A2(G110), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n439), .A2(KEYINPUT72), .A3(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(KEYINPUT72), .B1(new_n439), .B2(new_n440), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n438), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(KEYINPUT74), .ZN(new_n445));
  INV_X1    g259(.A(new_n443), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(new_n441), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT74), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n447), .A2(new_n448), .A3(new_n438), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n436), .A2(KEYINPUT23), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT23), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n451), .B1(new_n299), .B2(G128), .ZN(new_n452));
  OAI211_X1 g266(.A(new_n450), .B(new_n452), .C1(G119), .C2(new_n240), .ZN(new_n453));
  OR2_X1    g267(.A1(new_n453), .A2(G110), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n445), .A2(new_n449), .A3(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(KEYINPUT73), .A2(G125), .A3(G140), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  AOI21_X1  g271(.A(G140), .B1(KEYINPUT73), .B2(G125), .ZN(new_n458));
  OAI21_X1  g272(.A(KEYINPUT16), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NOR3_X1   g273(.A1(new_n321), .A2(KEYINPUT16), .A3(G140), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n459), .A2(G146), .A3(new_n461), .ZN(new_n462));
  XNOR2_X1  g276(.A(G125), .B(G140), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(new_n242), .ZN(new_n464));
  AND2_X1   g278(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n455), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n453), .A2(G110), .ZN(new_n467));
  AOI21_X1  g281(.A(G146), .B1(new_n459), .B2(new_n461), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT16), .ZN(new_n469));
  NAND2_X1  g283(.A1(KEYINPUT73), .A2(G125), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(new_n273), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n469), .B1(new_n471), .B2(new_n456), .ZN(new_n472));
  NOR3_X1   g286(.A1(new_n472), .A2(new_n242), .A3(new_n460), .ZN(new_n473));
  OAI221_X1 g287(.A(new_n467), .B1(new_n447), .B2(new_n438), .C1(new_n468), .C2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n466), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n187), .A2(G221), .A3(G234), .ZN(new_n476));
  XNOR2_X1  g290(.A(new_n476), .B(KEYINPUT22), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n477), .B(G137), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n475), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n466), .A2(new_n474), .A3(new_n478), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n480), .A2(new_n293), .A3(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT25), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n480), .A2(KEYINPUT25), .A3(new_n293), .A4(new_n481), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n434), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT75), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n480), .A2(new_n481), .ZN(new_n489));
  NOR3_X1   g303(.A1(new_n489), .A2(G902), .A3(new_n433), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n487), .A2(new_n488), .A3(new_n491), .ZN(new_n492));
  OAI21_X1  g306(.A(KEYINPUT75), .B1(new_n486), .B2(new_n490), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n431), .A2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(G475), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT88), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n497), .B1(new_n473), .B2(new_n468), .ZN(new_n498));
  NOR2_X1   g312(.A1(G237), .A2(G953), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT84), .ZN(new_n500));
  NAND4_X1  g314(.A1(new_n499), .A2(new_n500), .A3(new_n244), .A4(G214), .ZN(new_n501));
  XNOR2_X1  g315(.A(KEYINPUT84), .B(G143), .ZN(new_n502));
  INV_X1    g316(.A(G214), .ZN(new_n503));
  NOR3_X1   g317(.A1(new_n503), .A2(G237), .A3(G953), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n501), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(new_n236), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT17), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n499), .A2(G214), .ZN(new_n508));
  NAND2_X1  g322(.A1(KEYINPUT84), .A2(G143), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n500), .A2(new_n244), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n511), .A2(G131), .A3(new_n501), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n506), .A2(new_n507), .A3(new_n512), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n242), .B1(new_n472), .B2(new_n460), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n514), .A2(new_n462), .A3(KEYINPUT88), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n505), .A2(new_n236), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(KEYINPUT17), .ZN(new_n517));
  NAND4_X1  g331(.A1(new_n498), .A2(new_n513), .A3(new_n515), .A4(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT18), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n519), .A2(KEYINPUT85), .ZN(new_n520));
  AOI21_X1  g334(.A(G131), .B1(new_n511), .B2(new_n501), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n520), .B1(new_n516), .B2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(new_n520), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n505), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n471), .A2(G146), .A3(new_n456), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n464), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n522), .A2(new_n524), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n518), .A2(new_n527), .ZN(new_n528));
  XNOR2_X1  g342(.A(G113), .B(G122), .ZN(new_n529));
  XNOR2_X1  g343(.A(new_n529), .B(new_n195), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n518), .A2(new_n527), .A3(new_n530), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n496), .B1(new_n534), .B2(new_n293), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT20), .ZN(new_n537));
  XOR2_X1   g351(.A(KEYINPUT86), .B(KEYINPUT19), .Z(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(new_n463), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n471), .A2(KEYINPUT19), .A3(new_n456), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n539), .A2(new_n242), .A3(new_n540), .ZN(new_n541));
  OAI211_X1 g355(.A(new_n462), .B(new_n541), .C1(new_n516), .C2(new_n521), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n527), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(new_n531), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT87), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n523), .B1(new_n506), .B2(new_n512), .ZN(new_n547));
  INV_X1    g361(.A(new_n524), .ZN(new_n548));
  INV_X1    g362(.A(new_n526), .ZN(new_n549));
  NOR3_X1   g363(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n542), .ZN(new_n551));
  OAI211_X1 g365(.A(KEYINPUT87), .B(new_n531), .C1(new_n550), .C2(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n546), .A2(new_n533), .A3(new_n552), .ZN(new_n553));
  NOR2_X1   g367(.A1(G475), .A2(G902), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n537), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n552), .A2(new_n533), .ZN(new_n556));
  AOI21_X1  g370(.A(KEYINPUT87), .B1(new_n543), .B2(new_n531), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n537), .B(new_n554), .C1(new_n556), .C2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n536), .B1(new_n555), .B2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT91), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n240), .A2(G143), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(KEYINPUT13), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT13), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n564), .B1(new_n240), .B2(G143), .ZN(new_n565));
  OAI211_X1 g379(.A(new_n563), .B(new_n565), .C1(G128), .C2(new_n244), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(G134), .ZN(new_n567));
  XNOR2_X1  g381(.A(G116), .B(G122), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n568), .B(new_n198), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n244), .A2(G128), .ZN(new_n570));
  OR3_X1    g384(.A1(new_n562), .A2(new_n570), .A3(G134), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n567), .A2(new_n569), .A3(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT89), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n567), .A2(new_n569), .A3(KEYINPUT89), .A4(new_n571), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(G122), .ZN(new_n577));
  OR3_X1    g391(.A1(new_n577), .A2(KEYINPUT14), .A3(G116), .ZN(new_n578));
  OR2_X1    g392(.A1(new_n578), .A2(KEYINPUT90), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n577), .A2(G116), .ZN(new_n580));
  OAI21_X1  g394(.A(KEYINPUT14), .B1(new_n577), .B2(G116), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n578), .A2(KEYINPUT90), .ZN(new_n582));
  NAND4_X1  g396(.A1(new_n579), .A2(new_n580), .A3(new_n581), .A4(new_n582), .ZN(new_n583));
  OAI21_X1  g397(.A(G134), .B1(new_n562), .B2(new_n570), .ZN(new_n584));
  AOI22_X1  g398(.A1(new_n583), .A2(G107), .B1(new_n571), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n568), .A2(new_n198), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NOR3_X1   g401(.A1(new_n363), .A2(new_n432), .A3(G953), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n576), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n588), .B1(new_n576), .B2(new_n587), .ZN(new_n591));
  OAI211_X1 g405(.A(new_n561), .B(new_n293), .C1(new_n590), .C2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(G478), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n593), .A2(KEYINPUT15), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n592), .B(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(G234), .A2(G237), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n596), .A2(G952), .A3(new_n187), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n597), .B(KEYINPUT92), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  XOR2_X1   g413(.A(KEYINPUT21), .B(G898), .Z(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n596), .A2(G902), .A3(G953), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n599), .B1(new_n601), .B2(new_n603), .ZN(new_n604));
  NOR3_X1   g418(.A1(new_n560), .A2(new_n595), .A3(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  NOR3_X1   g420(.A1(new_n365), .A2(new_n495), .A3(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(new_n208), .ZN(G3));
  INV_X1    g422(.A(new_n365), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n576), .A2(new_n587), .ZN(new_n610));
  INV_X1    g424(.A(new_n588), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(new_n589), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT33), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n612), .A2(KEYINPUT33), .A3(new_n589), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n593), .A2(G902), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n615), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n613), .A2(new_n293), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(new_n593), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n560), .A2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n406), .A2(new_n407), .ZN(new_n624));
  OAI21_X1  g438(.A(G472), .B1(new_n410), .B2(G902), .ZN(new_n625));
  INV_X1    g439(.A(new_n604), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n494), .A2(new_n624), .A3(new_n625), .A4(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n609), .A2(new_n623), .A3(new_n628), .ZN(new_n629));
  XOR2_X1   g443(.A(KEYINPUT34), .B(G104), .Z(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G6));
  OAI21_X1  g445(.A(new_n554), .B1(new_n556), .B2(new_n557), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(KEYINPUT20), .ZN(new_n633));
  AND3_X1   g447(.A1(new_n633), .A2(KEYINPUT93), .A3(new_n558), .ZN(new_n634));
  AOI21_X1  g448(.A(KEYINPUT93), .B1(new_n633), .B2(new_n558), .ZN(new_n635));
  OAI211_X1 g449(.A(new_n595), .B(new_n536), .C1(new_n634), .C2(new_n635), .ZN(new_n636));
  NOR3_X1   g450(.A1(new_n365), .A2(new_n627), .A3(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(KEYINPUT35), .B(G107), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G9));
  AND2_X1   g453(.A1(new_n625), .A2(new_n624), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n433), .A2(G902), .ZN(new_n642));
  OR2_X1    g456(.A1(new_n475), .A2(KEYINPUT94), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n479), .A2(KEYINPUT36), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n475), .A2(KEYINPUT94), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n643), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n644), .B1(new_n643), .B2(new_n645), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n642), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT95), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  OAI211_X1 g465(.A(KEYINPUT95), .B(new_n642), .C1(new_n647), .C2(new_n648), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n651), .A2(new_n487), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n653), .A2(new_n605), .ZN(new_n654));
  NOR3_X1   g468(.A1(new_n365), .A2(new_n641), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(KEYINPUT37), .B(G110), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(KEYINPUT96), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n655), .B(new_n657), .ZN(G12));
  INV_X1    g472(.A(KEYINPUT98), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n598), .B(KEYINPUT97), .ZN(new_n660));
  INV_X1    g474(.A(G900), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n660), .B1(new_n661), .B2(new_n603), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n659), .B1(new_n636), .B2(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT93), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n664), .B1(new_n555), .B2(new_n559), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n633), .A2(KEYINPUT93), .A3(new_n558), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n535), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(new_n662), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n667), .A2(KEYINPUT98), .A3(new_n595), .A4(new_n668), .ZN(new_n669));
  AND3_X1   g483(.A1(new_n663), .A2(new_n653), .A3(new_n669), .ZN(new_n670));
  AND4_X1   g484(.A1(new_n431), .A2(new_n295), .A3(new_n361), .A4(new_n364), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G128), .ZN(G30));
  NAND2_X1  g487(.A1(new_n393), .A2(new_n394), .ZN(new_n674));
  AOI22_X1  g488(.A1(new_n420), .A2(new_n421), .B1(new_n424), .B2(new_n425), .ZN(new_n675));
  OAI21_X1  g489(.A(KEYINPUT100), .B1(new_n675), .B2(new_n388), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n422), .A2(new_n426), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT100), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n677), .A2(new_n678), .A3(new_n404), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n674), .A2(new_n676), .A3(new_n679), .A4(G472), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT101), .ZN(new_n681));
  NAND2_X1  g495(.A1(G472), .A2(G902), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n680), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n681), .B1(new_n680), .B2(new_n682), .ZN(new_n685));
  OAI211_X1 g499(.A(new_n408), .B(new_n412), .C1(new_n684), .C2(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT102), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n680), .A2(new_n682), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(KEYINPUT101), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(new_n683), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n691), .A2(KEYINPUT102), .A3(new_n412), .A4(new_n408), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n653), .B1(new_n688), .B2(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT40), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n662), .B(KEYINPUT39), .ZN(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n295), .A2(new_n694), .A3(new_n364), .A4(new_n696), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n295), .A2(new_n364), .A3(new_n696), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(KEYINPUT40), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n560), .A2(new_n595), .A3(new_n296), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT38), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT99), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n359), .A2(new_n702), .A3(new_n360), .ZN(new_n703));
  INV_X1    g517(.A(new_n703), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n702), .B1(new_n359), .B2(new_n360), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n701), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(new_n705), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n707), .A2(KEYINPUT38), .A3(new_n703), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n700), .B1(new_n706), .B2(new_n708), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n693), .A2(new_n697), .A3(new_n699), .A4(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G143), .ZN(G45));
  NAND3_X1  g525(.A1(new_n560), .A2(new_n621), .A3(new_n668), .ZN(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(new_n653), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n671), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G146), .ZN(G48));
  NAND2_X1  g531(.A1(KEYINPUT103), .A2(G469), .ZN(new_n718));
  INV_X1    g532(.A(new_n718), .ZN(new_n719));
  NOR3_X1   g533(.A1(new_n282), .A2(new_n274), .A3(new_n268), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n255), .B1(new_n258), .B2(new_n260), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n720), .B1(new_n721), .B2(new_n274), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n719), .B1(new_n722), .B2(G902), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n292), .A2(new_n293), .A3(new_n718), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n723), .A2(new_n361), .A3(new_n724), .A4(new_n364), .ZN(new_n725));
  NOR3_X1   g539(.A1(new_n495), .A2(new_n604), .A3(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(new_n623), .ZN(new_n727));
  XNOR2_X1  g541(.A(KEYINPUT41), .B(G113), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n727), .B(new_n728), .ZN(G15));
  INV_X1    g543(.A(new_n636), .ZN(new_n730));
  AND2_X1   g544(.A1(new_n726), .A2(new_n730), .ZN(new_n731));
  XOR2_X1   g545(.A(KEYINPUT104), .B(G116), .Z(new_n732));
  XNOR2_X1  g546(.A(new_n731), .B(new_n732), .ZN(G18));
  NOR3_X1   g547(.A1(new_n722), .A2(G902), .A3(new_n719), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n718), .B1(new_n292), .B2(new_n293), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n736), .A2(KEYINPUT105), .A3(new_n361), .A4(new_n364), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT105), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n725), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(new_n654), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n740), .A2(new_n431), .A3(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G119), .ZN(G21));
  NOR2_X1   g557(.A1(new_n486), .A2(new_n490), .ZN(new_n744));
  OAI21_X1  g558(.A(KEYINPUT106), .B1(new_n427), .B2(new_n428), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT106), .ZN(new_n746));
  OAI211_X1 g560(.A(new_n746), .B(new_n402), .C1(new_n675), .C2(new_n399), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n745), .A2(new_n404), .A3(new_n747), .ZN(new_n748));
  AND2_X1   g562(.A1(new_n748), .A2(new_n398), .ZN(new_n749));
  OAI211_X1 g563(.A(new_n625), .B(new_n744), .C1(new_n749), .C2(new_n411), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n723), .A2(new_n364), .A3(new_n724), .ZN(new_n751));
  NOR3_X1   g565(.A1(new_n750), .A2(new_n604), .A3(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(new_n594), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n592), .B(new_n753), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n535), .B1(new_n633), .B2(new_n558), .ZN(new_n755));
  OAI21_X1  g569(.A(KEYINPUT107), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT107), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n560), .A2(new_n595), .A3(new_n757), .ZN(new_n758));
  AND3_X1   g572(.A1(new_n756), .A2(new_n758), .A3(new_n361), .ZN(new_n759));
  AND3_X1   g573(.A1(new_n752), .A2(KEYINPUT108), .A3(new_n759), .ZN(new_n760));
  AOI21_X1  g574(.A(KEYINPUT108), .B1(new_n752), .B2(new_n759), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(new_n577), .ZN(G24));
  OAI21_X1  g577(.A(new_n625), .B1(new_n749), .B2(new_n411), .ZN(new_n764));
  INV_X1    g578(.A(new_n764), .ZN(new_n765));
  AND2_X1   g579(.A1(new_n725), .A2(new_n738), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n725), .A2(new_n738), .ZN(new_n767));
  OAI211_X1 g581(.A(new_n715), .B(new_n765), .C1(new_n766), .C2(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G125), .ZN(G27));
  NOR3_X1   g583(.A1(new_n722), .A2(G469), .A3(G902), .ZN(new_n770));
  AND3_X1   g584(.A1(new_n192), .A2(new_n270), .A3(new_n193), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n771), .A2(new_n271), .ZN(new_n772));
  OAI21_X1  g586(.A(KEYINPUT109), .B1(new_n290), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n272), .A2(new_n275), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT109), .ZN(new_n775));
  OAI211_X1 g589(.A(new_n774), .B(new_n775), .C1(new_n282), .C2(new_n268), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n261), .A2(new_n773), .A3(new_n776), .A4(G469), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n279), .A2(new_n293), .ZN(new_n778));
  INV_X1    g592(.A(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  OAI21_X1  g594(.A(KEYINPUT110), .B1(new_n770), .B2(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n359), .A2(new_n296), .A3(new_n360), .ZN(new_n782));
  INV_X1    g596(.A(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT110), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n294), .A2(new_n784), .A3(new_n779), .A4(new_n777), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n781), .A2(new_n364), .A3(new_n783), .A4(new_n785), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n786), .A2(new_n495), .ZN(new_n787));
  AOI21_X1  g601(.A(KEYINPUT42), .B1(new_n787), .B2(new_n713), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n431), .A2(new_n744), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT42), .ZN(new_n790));
  NOR4_X1   g604(.A1(new_n786), .A2(new_n789), .A3(new_n790), .A4(new_n712), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n788), .A2(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(KEYINPUT111), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(new_n236), .ZN(G33));
  AND2_X1   g608(.A1(new_n663), .A2(new_n669), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n787), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(G134), .ZN(G36));
  INV_X1    g611(.A(new_n364), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n261), .A2(new_n773), .A3(new_n776), .A4(KEYINPUT45), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(G469), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n288), .A2(KEYINPUT45), .ZN(new_n801));
  OAI21_X1  g615(.A(KEYINPUT112), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT45), .ZN(new_n803));
  INV_X1    g617(.A(new_n261), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n803), .B1(new_n804), .B2(new_n276), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT112), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n805), .A2(new_n806), .A3(G469), .A4(new_n799), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n802), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n808), .A2(new_n779), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT46), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n770), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  AOI211_X1 g625(.A(new_n810), .B(new_n778), .C1(new_n802), .C2(new_n807), .ZN(new_n812));
  INV_X1    g626(.A(new_n812), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n798), .B1(new_n811), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n755), .A2(new_n621), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT43), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n815), .B(new_n816), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n641), .A2(KEYINPUT44), .A3(new_n817), .A4(new_n653), .ZN(new_n818));
  AND2_X1   g632(.A1(new_n818), .A2(new_n783), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n641), .A2(new_n653), .A3(new_n817), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT44), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n814), .A2(new_n696), .A3(new_n819), .A4(new_n822), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n823), .B(G137), .ZN(G39));
  AOI21_X1  g638(.A(new_n778), .B1(new_n802), .B2(new_n807), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n294), .B1(new_n825), .B2(KEYINPUT46), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n364), .B1(new_n826), .B2(new_n812), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n827), .A2(KEYINPUT47), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT47), .ZN(new_n829));
  OAI211_X1 g643(.A(new_n829), .B(new_n364), .C1(new_n826), .C2(new_n812), .ZN(new_n830));
  NOR4_X1   g644(.A1(new_n431), .A2(new_n494), .A3(new_n712), .A4(new_n782), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n828), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n832), .B(G140), .ZN(G42));
  NAND2_X1  g647(.A1(new_n187), .A2(G952), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n817), .A2(new_n660), .ZN(new_n835));
  INV_X1    g649(.A(new_n751), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(new_n783), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(new_n789), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  XOR2_X1   g654(.A(new_n840), .B(KEYINPUT48), .Z(new_n841));
  NAND2_X1  g655(.A1(new_n688), .A2(new_n692), .ZN(new_n842));
  INV_X1    g656(.A(new_n842), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n837), .B1(new_n493), .B2(new_n492), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n843), .A2(new_n599), .A3(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n845), .A2(KEYINPUT118), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT118), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n843), .A2(new_n844), .A3(new_n847), .A4(new_n599), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  AOI211_X1 g663(.A(new_n834), .B(new_n841), .C1(new_n623), .C2(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(new_n750), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n851), .A2(new_n836), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n852), .A2(new_n835), .ZN(new_n853));
  AND2_X1   g667(.A1(new_n706), .A2(new_n708), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n853), .A2(new_n297), .A3(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT50), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(KEYINPUT117), .ZN(new_n857));
  INV_X1    g671(.A(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n853), .A2(new_n297), .A3(new_n854), .A4(new_n857), .ZN(new_n860));
  INV_X1    g674(.A(new_n653), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n764), .A2(new_n861), .ZN(new_n862));
  AOI22_X1  g676(.A1(new_n859), .A2(new_n860), .B1(new_n862), .B2(new_n838), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n560), .A2(new_n621), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n846), .A2(new_n848), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n835), .A2(new_n750), .A3(new_n782), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n828), .A2(new_n830), .ZN(new_n868));
  INV_X1    g682(.A(new_n736), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n868), .B1(new_n364), .B2(new_n869), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n866), .B1(new_n867), .B2(new_n870), .ZN(new_n871));
  XOR2_X1   g685(.A(KEYINPUT116), .B(KEYINPUT51), .Z(new_n872));
  OAI21_X1  g686(.A(new_n850), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(new_n866), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT51), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT119), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n870), .B(new_n876), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n875), .B1(new_n877), .B2(new_n867), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n873), .B1(new_n874), .B2(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT53), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n295), .A2(new_n364), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n861), .A2(new_n595), .A3(new_n662), .ZN(new_n882));
  AND2_X1   g696(.A1(new_n667), .A2(new_n783), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n881), .A2(new_n431), .A3(new_n882), .A4(new_n883), .ZN(new_n884));
  AND3_X1   g698(.A1(new_n781), .A2(new_n364), .A3(new_n785), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n885), .A2(new_n713), .A3(new_n783), .A4(new_n862), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(new_n887), .ZN(new_n888));
  AND2_X1   g702(.A1(new_n759), .A2(new_n668), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n842), .A2(new_n889), .A3(new_n861), .A4(new_n885), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n671), .B1(new_n670), .B2(new_n715), .ZN(new_n891));
  AND4_X1   g705(.A1(KEYINPUT52), .A2(new_n890), .A3(new_n891), .A4(new_n768), .ZN(new_n892));
  AOI211_X1 g706(.A(new_n714), .B(new_n764), .C1(new_n737), .C2(new_n739), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n431), .A2(new_n295), .A3(new_n361), .A4(new_n364), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n663), .A2(new_n653), .A3(new_n669), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n894), .B1(new_n895), .B2(new_n714), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n893), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g711(.A(KEYINPUT52), .B1(new_n897), .B2(new_n890), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n888), .B1(new_n892), .B2(new_n898), .ZN(new_n899));
  AND3_X1   g713(.A1(new_n431), .A2(new_n494), .A3(new_n626), .ZN(new_n900));
  INV_X1    g714(.A(new_n725), .ZN(new_n901));
  OAI211_X1 g715(.A(new_n900), .B(new_n901), .C1(new_n623), .C2(new_n730), .ZN(new_n902));
  OAI211_X1 g716(.A(new_n742), .B(new_n902), .C1(new_n760), .C2(new_n761), .ZN(new_n903));
  INV_X1    g717(.A(new_n903), .ZN(new_n904));
  AND2_X1   g718(.A1(new_n787), .A2(new_n795), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n787), .A2(new_n713), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(new_n790), .ZN(new_n907));
  INV_X1    g721(.A(new_n791), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n905), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n595), .A2(new_n755), .ZN(new_n910));
  NOR3_X1   g724(.A1(new_n365), .A2(new_n627), .A3(new_n910), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n655), .A2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT113), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n607), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(new_n629), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n609), .A2(new_n640), .A3(new_n741), .ZN(new_n916));
  INV_X1    g730(.A(new_n910), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n609), .A2(new_n628), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n915), .B1(new_n919), .B2(KEYINPUT113), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n904), .A2(new_n909), .A3(new_n914), .A4(new_n920), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n880), .B1(new_n899), .B2(new_n921), .ZN(new_n922));
  OAI21_X1  g736(.A(KEYINPUT113), .B1(new_n655), .B2(new_n911), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n916), .A2(new_n918), .A3(new_n913), .ZN(new_n924));
  INV_X1    g738(.A(new_n607), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n923), .A2(new_n924), .A3(new_n925), .A4(new_n629), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n796), .B1(new_n788), .B2(new_n791), .ZN(new_n927));
  NOR3_X1   g741(.A1(new_n926), .A2(new_n927), .A3(new_n903), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n890), .A2(new_n891), .A3(new_n768), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT52), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n897), .A2(KEYINPUT52), .A3(new_n890), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n887), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n928), .A2(new_n933), .A3(KEYINPUT53), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n922), .A2(KEYINPUT115), .A3(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT115), .ZN(new_n936));
  OAI211_X1 g750(.A(new_n936), .B(new_n880), .C1(new_n899), .C2(new_n921), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT54), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n740), .A2(new_n660), .A3(new_n851), .A4(new_n817), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT114), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n922), .A2(new_n942), .A3(new_n934), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n928), .A2(new_n933), .A3(KEYINPUT114), .A4(KEYINPUT53), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n943), .A2(KEYINPUT54), .A3(new_n944), .ZN(new_n945));
  NAND4_X1  g759(.A1(new_n879), .A2(new_n940), .A3(new_n941), .A4(new_n945), .ZN(new_n946));
  OR2_X1    g760(.A1(G952), .A2(G953), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  AND2_X1   g762(.A1(new_n869), .A2(KEYINPUT49), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n869), .A2(KEYINPUT49), .ZN(new_n950));
  NOR3_X1   g764(.A1(new_n949), .A2(new_n950), .A3(new_n815), .ZN(new_n951));
  NOR4_X1   g765(.A1(new_n486), .A2(new_n490), .A3(new_n297), .A4(new_n798), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n951), .A2(new_n843), .A3(new_n854), .A4(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n948), .A2(new_n953), .ZN(G75));
  NAND4_X1  g768(.A1(new_n935), .A2(G210), .A3(G902), .A4(new_n937), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n350), .A2(new_n354), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n956), .B(new_n352), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n957), .B(KEYINPUT120), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n958), .B(KEYINPUT55), .Z(new_n959));
  XNOR2_X1  g773(.A(KEYINPUT121), .B(KEYINPUT56), .ZN(new_n960));
  AND3_X1   g774(.A1(new_n955), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT56), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n959), .B1(new_n955), .B2(new_n962), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n187), .A2(G952), .ZN(new_n964));
  NOR3_X1   g778(.A1(new_n961), .A2(new_n963), .A3(new_n964), .ZN(G51));
  XNOR2_X1  g779(.A(new_n778), .B(KEYINPUT57), .ZN(new_n966));
  AND3_X1   g780(.A1(new_n935), .A2(KEYINPUT54), .A3(new_n937), .ZN(new_n967));
  AOI21_X1  g781(.A(KEYINPUT54), .B1(new_n935), .B2(new_n937), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n966), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n969), .A2(new_n292), .ZN(new_n970));
  OR3_X1    g784(.A1(new_n938), .A2(new_n293), .A3(new_n808), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n964), .B1(new_n970), .B2(new_n971), .ZN(G54));
  NAND4_X1  g786(.A1(new_n935), .A2(KEYINPUT58), .A3(G902), .A4(new_n937), .ZN(new_n973));
  INV_X1    g787(.A(new_n553), .ZN(new_n974));
  OR3_X1    g788(.A1(new_n973), .A2(new_n496), .A3(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(new_n964), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n974), .B1(new_n973), .B2(new_n496), .ZN(new_n977));
  AND3_X1   g791(.A1(new_n975), .A2(new_n976), .A3(new_n977), .ZN(G60));
  AND2_X1   g792(.A1(new_n615), .A2(new_n616), .ZN(new_n979));
  NAND2_X1  g793(.A1(G478), .A2(G902), .ZN(new_n980));
  XOR2_X1   g794(.A(new_n980), .B(KEYINPUT59), .Z(new_n981));
  INV_X1    g795(.A(new_n981), .ZN(new_n982));
  OAI211_X1 g796(.A(new_n979), .B(new_n982), .C1(new_n967), .C2(new_n968), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n981), .B1(new_n940), .B2(new_n945), .ZN(new_n984));
  OAI211_X1 g798(.A(new_n983), .B(new_n976), .C1(new_n984), .C2(new_n979), .ZN(new_n985));
  INV_X1    g799(.A(new_n985), .ZN(G63));
  XNOR2_X1  g800(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n432), .A2(new_n293), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n987), .B(new_n988), .ZN(new_n989));
  INV_X1    g803(.A(new_n989), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n489), .B1(new_n938), .B2(new_n990), .ZN(new_n991));
  OR2_X1    g805(.A1(new_n647), .A2(new_n648), .ZN(new_n992));
  NAND4_X1  g806(.A1(new_n935), .A2(new_n992), .A3(new_n937), .A4(new_n989), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n991), .A2(new_n976), .A3(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT61), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND4_X1  g810(.A1(new_n991), .A2(KEYINPUT61), .A3(new_n976), .A4(new_n993), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n996), .A2(new_n997), .ZN(G66));
  OAI21_X1  g812(.A(G953), .B1(new_n601), .B2(new_n327), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n926), .A2(new_n903), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n999), .B1(new_n1000), .B2(G953), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n956), .B1(G898), .B2(new_n187), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n1001), .B(new_n1002), .ZN(G69));
  INV_X1    g817(.A(KEYINPUT124), .ZN(new_n1004));
  INV_X1    g818(.A(KEYINPUT123), .ZN(new_n1005));
  INV_X1    g819(.A(new_n698), .ZN(new_n1006));
  INV_X1    g820(.A(new_n495), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n622), .A2(new_n910), .ZN(new_n1008));
  NAND4_X1  g822(.A1(new_n1006), .A2(new_n1007), .A3(new_n783), .A4(new_n1008), .ZN(new_n1009));
  AND3_X1   g823(.A1(new_n897), .A2(KEYINPUT62), .A3(new_n710), .ZN(new_n1010));
  AOI21_X1  g824(.A(KEYINPUT62), .B1(new_n897), .B2(new_n710), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n1009), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n832), .A2(new_n823), .ZN(new_n1013));
  OAI21_X1  g827(.A(new_n1005), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  AND2_X1   g828(.A1(new_n832), .A2(new_n823), .ZN(new_n1015));
  INV_X1    g829(.A(new_n1009), .ZN(new_n1016));
  INV_X1    g830(.A(KEYINPUT62), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n842), .A2(new_n861), .ZN(new_n1018));
  NAND3_X1  g832(.A1(new_n699), .A2(new_n697), .A3(new_n709), .ZN(new_n1019));
  NOR2_X1   g833(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g834(.A1(new_n672), .A2(new_n716), .A3(new_n768), .ZN(new_n1021));
  OAI21_X1  g835(.A(new_n1017), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g836(.A1(new_n897), .A2(KEYINPUT62), .A3(new_n710), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n1016), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g838(.A1(new_n1015), .A2(new_n1024), .A3(KEYINPUT123), .ZN(new_n1025));
  AOI21_X1  g839(.A(G953), .B1(new_n1014), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n372), .A2(new_n381), .ZN(new_n1027));
  AND2_X1   g841(.A1(new_n539), .A2(new_n540), .ZN(new_n1028));
  XNOR2_X1  g842(.A(new_n1027), .B(new_n1028), .ZN(new_n1029));
  INV_X1    g843(.A(new_n1029), .ZN(new_n1030));
  OAI21_X1  g844(.A(new_n1004), .B1(new_n1026), .B2(new_n1030), .ZN(new_n1031));
  NOR3_X1   g845(.A1(new_n1012), .A2(new_n1005), .A3(new_n1013), .ZN(new_n1032));
  AOI21_X1  g846(.A(KEYINPUT123), .B1(new_n1015), .B2(new_n1024), .ZN(new_n1033));
  OAI21_X1  g847(.A(new_n187), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g848(.A1(new_n1034), .A2(KEYINPUT124), .A3(new_n1029), .ZN(new_n1035));
  AND2_X1   g849(.A1(new_n1031), .A2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g850(.A(new_n1029), .B1(G900), .B2(G953), .ZN(new_n1037));
  NAND4_X1  g851(.A1(new_n814), .A2(new_n696), .A3(new_n759), .A4(new_n839), .ZN(new_n1038));
  INV_X1    g852(.A(KEYINPUT125), .ZN(new_n1039));
  OAI21_X1  g853(.A(new_n909), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  NOR2_X1   g854(.A1(new_n1040), .A2(new_n1021), .ZN(new_n1041));
  NAND2_X1  g855(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1042));
  NAND3_X1  g856(.A1(new_n1041), .A2(new_n1015), .A3(new_n1042), .ZN(new_n1043));
  OAI21_X1  g857(.A(new_n1037), .B1(new_n1043), .B2(G953), .ZN(new_n1044));
  AOI21_X1  g858(.A(new_n187), .B1(G227), .B2(G900), .ZN(new_n1045));
  INV_X1    g859(.A(new_n1045), .ZN(new_n1046));
  OAI211_X1 g860(.A(new_n1036), .B(new_n1044), .C1(KEYINPUT126), .C2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g861(.A1(new_n1031), .A2(new_n1035), .A3(new_n1044), .ZN(new_n1048));
  NAND3_X1  g862(.A1(new_n1031), .A2(new_n1035), .A3(KEYINPUT126), .ZN(new_n1049));
  NAND3_X1  g863(.A1(new_n1048), .A2(new_n1049), .A3(new_n1045), .ZN(new_n1050));
  NAND2_X1  g864(.A1(new_n1047), .A2(new_n1050), .ZN(G72));
  NAND4_X1  g865(.A1(new_n1041), .A2(new_n1000), .A3(new_n1015), .A4(new_n1042), .ZN(new_n1052));
  XOR2_X1   g866(.A(new_n682), .B(KEYINPUT63), .Z(new_n1053));
  NAND2_X1  g867(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g868(.A(KEYINPUT127), .ZN(new_n1055));
  NOR2_X1   g869(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g870(.A(KEYINPUT127), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1057));
  NOR4_X1   g871(.A1(new_n1056), .A2(new_n1057), .A3(new_n388), .A4(new_n415), .ZN(new_n1058));
  OAI21_X1  g872(.A(new_n674), .B1(new_n388), .B2(new_n416), .ZN(new_n1059));
  AND4_X1   g873(.A1(new_n944), .A2(new_n943), .A3(new_n1053), .A4(new_n1059), .ZN(new_n1060));
  NAND3_X1  g874(.A1(new_n1014), .A2(new_n1000), .A3(new_n1025), .ZN(new_n1061));
  AOI211_X1 g875(.A(new_n404), .B(new_n416), .C1(new_n1061), .C2(new_n1053), .ZN(new_n1062));
  NOR4_X1   g876(.A1(new_n1058), .A2(new_n964), .A3(new_n1060), .A4(new_n1062), .ZN(G57));
endmodule


