

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724;

  NOR2_X1 U369 ( .A1(n618), .A2(n698), .ZN(n619) );
  NOR2_X1 U370 ( .A1(n625), .A2(n698), .ZN(n626) );
  XNOR2_X1 U371 ( .A(n463), .B(KEYINPUT32), .ZN(n721) );
  XNOR2_X1 U372 ( .A(n510), .B(n509), .ZN(n701) );
  INV_X1 U373 ( .A(G953), .ZN(n713) );
  NOR2_X1 U374 ( .A1(n602), .A2(n698), .ZN(n604) );
  NOR2_X1 U375 ( .A1(n608), .A2(n698), .ZN(n610) );
  XNOR2_X2 U376 ( .A(n408), .B(G134), .ZN(n434) );
  XNOR2_X2 U377 ( .A(n710), .B(G146), .ZN(n457) );
  XNOR2_X2 U378 ( .A(n434), .B(n433), .ZN(n710) );
  XNOR2_X2 U379 ( .A(n376), .B(n375), .ZN(n582) );
  NOR2_X1 U380 ( .A1(n586), .A2(n585), .ZN(n712) );
  AND2_X1 U381 ( .A1(n506), .A2(n505), .ZN(n507) );
  AND2_X1 U382 ( .A1(n480), .A2(n462), .ZN(n463) );
  AND2_X1 U383 ( .A1(n461), .A2(n349), .ZN(n462) );
  XNOR2_X1 U384 ( .A(n469), .B(n468), .ZN(n484) );
  XNOR2_X2 U385 ( .A(n386), .B(n352), .ZN(n490) );
  XNOR2_X2 U386 ( .A(n477), .B(n476), .ZN(n613) );
  NOR2_X1 U387 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U388 ( .A(n348), .B(n374), .ZN(n375) );
  INV_X1 U389 ( .A(G119), .ZN(n353) );
  XNOR2_X1 U390 ( .A(n437), .B(G472), .ZN(n539) );
  XNOR2_X1 U391 ( .A(n447), .B(n351), .ZN(n605) );
  AND2_X1 U392 ( .A1(n588), .A2(n712), .ZN(n587) );
  INV_X1 U393 ( .A(KEYINPUT18), .ZN(n366) );
  XNOR2_X1 U394 ( .A(n561), .B(n560), .ZN(n680) );
  AND2_X1 U395 ( .A1(n601), .A2(G953), .ZN(n698) );
  XNOR2_X1 U396 ( .A(n526), .B(n525), .ZN(n527) );
  XNOR2_X1 U397 ( .A(KEYINPUT36), .B(KEYINPUT85), .ZN(n525) );
  NOR2_X1 U398 ( .A1(n493), .A2(n494), .ZN(n640) );
  XOR2_X1 U399 ( .A(KEYINPUT78), .B(KEYINPUT88), .Z(n348) );
  XOR2_X1 U400 ( .A(n460), .B(KEYINPUT104), .Z(n349) );
  XNOR2_X1 U401 ( .A(KEYINPUT48), .B(KEYINPUT81), .ZN(n350) );
  XOR2_X1 U402 ( .A(n446), .B(n445), .Z(n351) );
  XOR2_X1 U403 ( .A(n385), .B(KEYINPUT0), .Z(n352) );
  INV_X1 U404 ( .A(n634), .ZN(n500) );
  INV_X1 U405 ( .A(KEYINPUT71), .ZN(n354) );
  OR2_X1 U406 ( .A1(n721), .A2(n466), .ZN(n467) );
  XOR2_X1 U407 ( .A(KEYINPUT69), .B(KEYINPUT10), .Z(n387) );
  XNOR2_X1 U408 ( .A(n570), .B(KEYINPUT46), .ZN(n571) );
  XNOR2_X1 U409 ( .A(KEYINPUT3), .B(G101), .ZN(n357) );
  XNOR2_X1 U410 ( .A(n387), .B(G140), .ZN(n389) );
  XNOR2_X1 U411 ( .A(n367), .B(n366), .ZN(n368) );
  XNOR2_X1 U412 ( .A(n449), .B(KEYINPUT25), .ZN(n450) );
  XNOR2_X1 U413 ( .A(n389), .B(n388), .ZN(n708) );
  XNOR2_X1 U414 ( .A(n369), .B(n368), .ZN(n371) );
  XNOR2_X1 U415 ( .A(n451), .B(n450), .ZN(n489) );
  INV_X1 U416 ( .A(KEYINPUT38), .ZN(n559) );
  XNOR2_X1 U417 ( .A(n575), .B(n350), .ZN(n586) );
  XNOR2_X1 U418 ( .A(n582), .B(n559), .ZN(n650) );
  NOR2_X1 U419 ( .A1(n565), .A2(n650), .ZN(n567) );
  BUF_X1 U420 ( .A(n539), .Z(n528) );
  XNOR2_X1 U421 ( .A(n426), .B(n425), .ZN(n480) );
  NAND2_X1 U422 ( .A1(KEYINPUT71), .A2(n353), .ZN(n356) );
  NAND2_X1 U423 ( .A1(n354), .A2(G119), .ZN(n355) );
  NAND2_X1 U424 ( .A1(n356), .A2(n355), .ZN(n358) );
  XNOR2_X1 U425 ( .A(n358), .B(n357), .ZN(n360) );
  XNOR2_X1 U426 ( .A(G113), .B(G116), .ZN(n359) );
  XNOR2_X1 U427 ( .A(n360), .B(n359), .ZN(n430) );
  XNOR2_X1 U428 ( .A(n430), .B(G122), .ZN(n363) );
  XNOR2_X1 U429 ( .A(G110), .B(G107), .ZN(n361) );
  XNOR2_X1 U430 ( .A(n361), .B(G104), .ZN(n455) );
  XOR2_X1 U431 ( .A(n455), .B(KEYINPUT16), .Z(n362) );
  XNOR2_X1 U432 ( .A(n363), .B(n362), .ZN(n699) );
  XOR2_X1 U433 ( .A(KEYINPUT75), .B(KEYINPUT17), .Z(n365) );
  XNOR2_X1 U434 ( .A(KEYINPUT4), .B(KEYINPUT87), .ZN(n364) );
  XNOR2_X1 U435 ( .A(n365), .B(n364), .ZN(n369) );
  NAND2_X1 U436 ( .A1(G224), .A2(n713), .ZN(n367) );
  XNOR2_X2 U437 ( .A(G143), .B(G128), .ZN(n408) );
  XOR2_X1 U438 ( .A(G146), .B(G125), .Z(n388) );
  XNOR2_X1 U439 ( .A(n408), .B(n388), .ZN(n370) );
  XNOR2_X1 U440 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X1 U441 ( .A(n699), .B(n372), .ZN(n614) );
  INV_X1 U442 ( .A(KEYINPUT15), .ZN(n373) );
  XNOR2_X1 U443 ( .A(n373), .B(G902), .ZN(n513) );
  NOR2_X1 U444 ( .A1(n614), .A2(n513), .ZN(n376) );
  OR2_X1 U445 ( .A1(G237), .A2(G902), .ZN(n377) );
  NAND2_X1 U446 ( .A1(G210), .A2(n377), .ZN(n374) );
  INV_X1 U447 ( .A(n582), .ZN(n524) );
  NAND2_X1 U448 ( .A1(n377), .A2(G214), .ZN(n378) );
  XNOR2_X1 U449 ( .A(KEYINPUT89), .B(n378), .ZN(n651) );
  INV_X1 U450 ( .A(n651), .ZN(n540) );
  NAND2_X1 U451 ( .A1(n524), .A2(n540), .ZN(n379) );
  XNOR2_X1 U452 ( .A(n379), .B(KEYINPUT19), .ZN(n535) );
  OR2_X1 U453 ( .A1(G898), .A2(n713), .ZN(n700) );
  NAND2_X1 U454 ( .A1(G234), .A2(G237), .ZN(n380) );
  XNOR2_X1 U455 ( .A(KEYINPUT14), .B(n380), .ZN(n381) );
  NAND2_X1 U456 ( .A1(G902), .A2(n381), .ZN(n516) );
  OR2_X1 U457 ( .A1(n700), .A2(n516), .ZN(n383) );
  NAND2_X1 U458 ( .A1(G952), .A2(n381), .ZN(n678) );
  NOR2_X1 U459 ( .A1(G953), .A2(n678), .ZN(n382) );
  XOR2_X1 U460 ( .A(KEYINPUT90), .B(n382), .Z(n519) );
  NAND2_X1 U461 ( .A1(n383), .A2(n519), .ZN(n384) );
  NAND2_X1 U462 ( .A1(n535), .A2(n384), .ZN(n386) );
  INV_X1 U463 ( .A(KEYINPUT67), .ZN(n385) );
  XNOR2_X1 U464 ( .A(KEYINPUT13), .B(G475), .ZN(n404) );
  XOR2_X1 U465 ( .A(KEYINPUT11), .B(G122), .Z(n391) );
  XNOR2_X1 U466 ( .A(G131), .B(G143), .ZN(n390) );
  XNOR2_X1 U467 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U468 ( .A(n708), .B(n392), .ZN(n402) );
  XOR2_X1 U469 ( .A(KEYINPUT96), .B(G104), .Z(n394) );
  XNOR2_X1 U470 ( .A(G113), .B(KEYINPUT94), .ZN(n393) );
  XNOR2_X1 U471 ( .A(n394), .B(n393), .ZN(n398) );
  XOR2_X1 U472 ( .A(KEYINPUT97), .B(KEYINPUT98), .Z(n396) );
  XNOR2_X1 U473 ( .A(KEYINPUT95), .B(KEYINPUT12), .ZN(n395) );
  XNOR2_X1 U474 ( .A(n396), .B(n395), .ZN(n397) );
  XOR2_X1 U475 ( .A(n398), .B(n397), .Z(n400) );
  NOR2_X1 U476 ( .A1(G953), .A2(G237), .ZN(n427) );
  NAND2_X1 U477 ( .A1(G214), .A2(n427), .ZN(n399) );
  XNOR2_X1 U478 ( .A(n400), .B(n399), .ZN(n401) );
  XNOR2_X1 U479 ( .A(n402), .B(n401), .ZN(n622) );
  NOR2_X1 U480 ( .A1(G902), .A2(n622), .ZN(n403) );
  XNOR2_X1 U481 ( .A(n404), .B(n403), .ZN(n492) );
  XOR2_X1 U482 ( .A(KEYINPUT8), .B(KEYINPUT68), .Z(n406) );
  NAND2_X1 U483 ( .A1(G234), .A2(n713), .ZN(n405) );
  XNOR2_X1 U484 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U485 ( .A(KEYINPUT80), .B(n407), .ZN(n441) );
  NAND2_X1 U486 ( .A1(G217), .A2(n441), .ZN(n409) );
  XNOR2_X1 U487 ( .A(n409), .B(n434), .ZN(n416) );
  XOR2_X1 U488 ( .A(G107), .B(KEYINPUT101), .Z(n411) );
  XNOR2_X1 U489 ( .A(KEYINPUT7), .B(KEYINPUT9), .ZN(n410) );
  XNOR2_X1 U490 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U491 ( .A(n412), .B(KEYINPUT100), .Z(n414) );
  XNOR2_X1 U492 ( .A(G116), .B(G122), .ZN(n413) );
  XNOR2_X1 U493 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U494 ( .A(n416), .B(n415), .ZN(n694) );
  INV_X1 U495 ( .A(G902), .ZN(n436) );
  NAND2_X1 U496 ( .A1(n694), .A2(n436), .ZN(n417) );
  XNOR2_X1 U497 ( .A(n417), .B(G478), .ZN(n494) );
  NOR2_X1 U498 ( .A1(n492), .A2(n494), .ZN(n418) );
  XNOR2_X1 U499 ( .A(KEYINPUT102), .B(n418), .ZN(n653) );
  INV_X1 U500 ( .A(n513), .ZN(n419) );
  NAND2_X1 U501 ( .A1(n419), .A2(G234), .ZN(n420) );
  XNOR2_X1 U502 ( .A(n420), .B(KEYINPUT20), .ZN(n448) );
  NAND2_X1 U503 ( .A1(n448), .A2(G221), .ZN(n421) );
  XOR2_X1 U504 ( .A(KEYINPUT21), .B(n421), .Z(n662) );
  INV_X1 U505 ( .A(KEYINPUT93), .ZN(n422) );
  XNOR2_X1 U506 ( .A(n662), .B(n422), .ZN(n487) );
  NAND2_X1 U507 ( .A1(n653), .A2(n487), .ZN(n423) );
  XNOR2_X1 U508 ( .A(n423), .B(KEYINPUT103), .ZN(n424) );
  NAND2_X1 U509 ( .A1(n490), .A2(n424), .ZN(n426) );
  XNOR2_X1 U510 ( .A(KEYINPUT65), .B(KEYINPUT22), .ZN(n425) );
  NAND2_X1 U511 ( .A1(n427), .A2(G210), .ZN(n428) );
  XNOR2_X1 U512 ( .A(n428), .B(KEYINPUT5), .ZN(n429) );
  XNOR2_X1 U513 ( .A(n430), .B(n429), .ZN(n435) );
  XNOR2_X1 U514 ( .A(G137), .B(G131), .ZN(n432) );
  INV_X1 U515 ( .A(KEYINPUT4), .ZN(n431) );
  XNOR2_X1 U516 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U517 ( .A(n435), .B(n457), .ZN(n598) );
  NAND2_X1 U518 ( .A1(n598), .A2(n436), .ZN(n437) );
  XNOR2_X1 U519 ( .A(n528), .B(KEYINPUT6), .ZN(n521) );
  XOR2_X1 U520 ( .A(KEYINPUT77), .B(n521), .Z(n461) );
  XOR2_X1 U521 ( .A(KEYINPUT74), .B(KEYINPUT23), .Z(n439) );
  XNOR2_X1 U522 ( .A(G119), .B(G110), .ZN(n438) );
  XNOR2_X1 U523 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U524 ( .A(n708), .B(n440), .ZN(n447) );
  NAND2_X1 U525 ( .A1(n441), .A2(G221), .ZN(n446) );
  XOR2_X1 U526 ( .A(KEYINPUT91), .B(KEYINPUT24), .Z(n443) );
  XNOR2_X1 U527 ( .A(G137), .B(G128), .ZN(n442) );
  XNOR2_X1 U528 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U529 ( .A(n444), .B(KEYINPUT92), .Z(n445) );
  NOR2_X1 U530 ( .A1(n605), .A2(G902), .ZN(n451) );
  NAND2_X1 U531 ( .A1(G217), .A2(n448), .ZN(n449) );
  INV_X1 U532 ( .A(n489), .ZN(n515) );
  XNOR2_X1 U533 ( .A(G140), .B(G101), .ZN(n453) );
  NAND2_X1 U534 ( .A1(n713), .A2(G227), .ZN(n452) );
  XNOR2_X1 U535 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U536 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U537 ( .A(n457), .B(n456), .ZN(n690) );
  OR2_X1 U538 ( .A1(n690), .A2(G902), .ZN(n459) );
  XNOR2_X1 U539 ( .A(KEYINPUT70), .B(G469), .ZN(n458) );
  XNOR2_X2 U540 ( .A(n459), .B(n458), .ZN(n532) );
  XNOR2_X2 U541 ( .A(n532), .B(KEYINPUT1), .ZN(n659) );
  NAND2_X1 U542 ( .A1(n515), .A2(n659), .ZN(n460) );
  INV_X1 U543 ( .A(n515), .ZN(n663) );
  NOR2_X1 U544 ( .A1(n663), .A2(n528), .ZN(n464) );
  INV_X1 U545 ( .A(n659), .ZN(n579) );
  AND2_X1 U546 ( .A1(n464), .A2(n579), .ZN(n465) );
  AND2_X1 U547 ( .A1(n480), .A2(n465), .ZN(n634) );
  INV_X1 U548 ( .A(KEYINPUT44), .ZN(n504) );
  NAND2_X1 U549 ( .A1(n500), .A2(n504), .ZN(n466) );
  NAND2_X1 U550 ( .A1(n467), .A2(KEYINPUT84), .ZN(n479) );
  AND2_X1 U551 ( .A1(n489), .A2(n487), .ZN(n660) );
  NAND2_X1 U552 ( .A1(n660), .A2(n659), .ZN(n469) );
  INV_X1 U553 ( .A(KEYINPUT73), .ZN(n468) );
  XNOR2_X1 U554 ( .A(n484), .B(KEYINPUT105), .ZN(n471) );
  INV_X1 U555 ( .A(n521), .ZN(n470) );
  NAND2_X1 U556 ( .A1(n471), .A2(n470), .ZN(n472) );
  XNOR2_X2 U557 ( .A(n472), .B(KEYINPUT33), .ZN(n679) );
  NAND2_X1 U558 ( .A1(n679), .A2(n490), .ZN(n474) );
  INV_X1 U559 ( .A(KEYINPUT34), .ZN(n473) );
  XNOR2_X1 U560 ( .A(n474), .B(n473), .ZN(n475) );
  AND2_X1 U561 ( .A1(n494), .A2(n492), .ZN(n548) );
  NAND2_X1 U562 ( .A1(n475), .A2(n548), .ZN(n477) );
  XNOR2_X1 U563 ( .A(KEYINPUT76), .B(KEYINPUT35), .ZN(n476) );
  INV_X1 U564 ( .A(n613), .ZN(n478) );
  NAND2_X1 U565 ( .A1(n479), .A2(n478), .ZN(n499) );
  NAND2_X1 U566 ( .A1(n521), .A2(n480), .ZN(n481) );
  XNOR2_X1 U567 ( .A(n481), .B(KEYINPUT83), .ZN(n483) );
  AND2_X1 U568 ( .A1(n579), .A2(n663), .ZN(n482) );
  AND2_X1 U569 ( .A1(n483), .A2(n482), .ZN(n627) );
  INV_X1 U570 ( .A(n528), .ZN(n666) );
  OR2_X1 U571 ( .A1(n484), .A2(n666), .ZN(n670) );
  INV_X1 U572 ( .A(n670), .ZN(n485) );
  NAND2_X1 U573 ( .A1(n490), .A2(n485), .ZN(n486) );
  XNOR2_X1 U574 ( .A(n486), .B(KEYINPUT31), .ZN(n643) );
  AND2_X1 U575 ( .A1(n487), .A2(n532), .ZN(n488) );
  AND2_X1 U576 ( .A1(n489), .A2(n488), .ZN(n538) );
  NAND2_X1 U577 ( .A1(n490), .A2(n538), .ZN(n491) );
  NOR2_X1 U578 ( .A1(n528), .A2(n491), .ZN(n630) );
  NOR2_X1 U579 ( .A1(n643), .A2(n630), .ZN(n496) );
  XNOR2_X1 U580 ( .A(n492), .B(KEYINPUT99), .ZN(n493) );
  NAND2_X1 U581 ( .A1(n494), .A2(n493), .ZN(n576) );
  INV_X1 U582 ( .A(n576), .ZN(n642) );
  NOR2_X1 U583 ( .A1(n640), .A2(n642), .ZN(n550) );
  XOR2_X1 U584 ( .A(n550), .B(KEYINPUT79), .Z(n495) );
  NOR2_X1 U585 ( .A1(n496), .A2(n495), .ZN(n497) );
  NOR2_X1 U586 ( .A1(n627), .A2(n497), .ZN(n498) );
  NAND2_X1 U587 ( .A1(n499), .A2(n498), .ZN(n508) );
  NAND2_X1 U588 ( .A1(n500), .A2(KEYINPUT44), .ZN(n501) );
  NOR2_X1 U589 ( .A1(n721), .A2(n501), .ZN(n503) );
  NAND2_X1 U590 ( .A1(n613), .A2(KEYINPUT84), .ZN(n502) );
  NAND2_X1 U591 ( .A1(n503), .A2(n502), .ZN(n506) );
  NAND2_X1 U592 ( .A1(n504), .A2(KEYINPUT84), .ZN(n505) );
  NOR2_X2 U593 ( .A1(n508), .A2(n507), .ZN(n510) );
  XOR2_X1 U594 ( .A(KEYINPUT64), .B(KEYINPUT45), .Z(n509) );
  NAND2_X1 U595 ( .A1(n513), .A2(KEYINPUT2), .ZN(n512) );
  INV_X1 U596 ( .A(KEYINPUT66), .ZN(n511) );
  NAND2_X1 U597 ( .A1(n512), .A2(n511), .ZN(n589) );
  INV_X1 U598 ( .A(n589), .ZN(n514) );
  OR2_X1 U599 ( .A1(n514), .A2(n513), .ZN(n588) );
  NAND2_X1 U600 ( .A1(n515), .A2(n662), .ZN(n530) );
  NOR2_X1 U601 ( .A1(G900), .A2(n516), .ZN(n517) );
  NAND2_X1 U602 ( .A1(G953), .A2(n517), .ZN(n518) );
  NAND2_X1 U603 ( .A1(n519), .A2(n518), .ZN(n545) );
  NAND2_X1 U604 ( .A1(n540), .A2(n545), .ZN(n520) );
  NOR2_X1 U605 ( .A1(n521), .A2(n520), .ZN(n522) );
  NAND2_X1 U606 ( .A1(n640), .A2(n522), .ZN(n523) );
  NOR2_X1 U607 ( .A1(n530), .A2(n523), .ZN(n578) );
  NAND2_X1 U608 ( .A1(n578), .A2(n524), .ZN(n526) );
  NAND2_X1 U609 ( .A1(n527), .A2(n659), .ZN(n612) );
  INV_X1 U610 ( .A(n550), .ZN(n648) );
  NAND2_X1 U611 ( .A1(n528), .A2(n545), .ZN(n529) );
  NOR2_X1 U612 ( .A1(n530), .A2(n529), .ZN(n531) );
  XOR2_X1 U613 ( .A(KEYINPUT28), .B(n531), .Z(n534) );
  XOR2_X1 U614 ( .A(KEYINPUT110), .B(n532), .Z(n533) );
  NOR2_X1 U615 ( .A1(n534), .A2(n533), .ZN(n562) );
  NAND2_X1 U616 ( .A1(n562), .A2(n535), .ZN(n555) );
  INV_X1 U617 ( .A(n555), .ZN(n638) );
  NAND2_X1 U618 ( .A1(n648), .A2(n638), .ZN(n536) );
  NAND2_X1 U619 ( .A1(n536), .A2(KEYINPUT47), .ZN(n537) );
  AND2_X1 U620 ( .A1(n612), .A2(n537), .ZN(n558) );
  XNOR2_X1 U621 ( .A(n538), .B(KEYINPUT107), .ZN(n544) );
  NAND2_X1 U622 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U623 ( .A(n541), .B(KEYINPUT108), .ZN(n542) );
  XNOR2_X1 U624 ( .A(n542), .B(KEYINPUT30), .ZN(n543) );
  NOR2_X1 U625 ( .A1(n544), .A2(n543), .ZN(n546) );
  NAND2_X1 U626 ( .A1(n546), .A2(n545), .ZN(n565) );
  NOR2_X1 U627 ( .A1(n582), .A2(n565), .ZN(n547) );
  NAND2_X1 U628 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U629 ( .A(KEYINPUT109), .B(n549), .ZN(n720) );
  AND2_X1 U630 ( .A1(n550), .A2(KEYINPUT79), .ZN(n553) );
  OR2_X1 U631 ( .A1(n550), .A2(KEYINPUT79), .ZN(n551) );
  NOR2_X1 U632 ( .A1(KEYINPUT47), .A2(n551), .ZN(n552) );
  NOR2_X1 U633 ( .A1(n553), .A2(n552), .ZN(n554) );
  NOR2_X1 U634 ( .A1(n555), .A2(n554), .ZN(n556) );
  NOR2_X1 U635 ( .A1(n720), .A2(n556), .ZN(n557) );
  NAND2_X1 U636 ( .A1(n558), .A2(n557), .ZN(n574) );
  XOR2_X1 U637 ( .A(KEYINPUT112), .B(KEYINPUT42), .Z(n564) );
  XOR2_X1 U638 ( .A(KEYINPUT41), .B(KEYINPUT111), .Z(n561) );
  NOR2_X1 U639 ( .A1(n651), .A2(n650), .ZN(n649) );
  NAND2_X1 U640 ( .A1(n649), .A2(n653), .ZN(n560) );
  NAND2_X1 U641 ( .A1(n562), .A2(n680), .ZN(n563) );
  XNOR2_X1 U642 ( .A(n564), .B(n563), .ZN(n723) );
  INV_X1 U643 ( .A(n640), .ZN(n568) );
  XNOR2_X1 U644 ( .A(KEYINPUT72), .B(KEYINPUT39), .ZN(n566) );
  XNOR2_X1 U645 ( .A(n567), .B(n566), .ZN(n577) );
  NOR2_X1 U646 ( .A1(n568), .A2(n577), .ZN(n569) );
  XNOR2_X1 U647 ( .A(n569), .B(KEYINPUT40), .ZN(n722) );
  NOR2_X1 U648 ( .A1(n723), .A2(n722), .ZN(n572) );
  INV_X1 U649 ( .A(KEYINPUT82), .ZN(n570) );
  XNOR2_X1 U650 ( .A(n572), .B(n571), .ZN(n573) );
  NOR2_X1 U651 ( .A1(n577), .A2(n576), .ZN(n645) );
  INV_X1 U652 ( .A(n645), .ZN(n584) );
  XNOR2_X1 U653 ( .A(KEYINPUT106), .B(n578), .ZN(n580) );
  NAND2_X1 U654 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U655 ( .A(n581), .B(KEYINPUT43), .ZN(n583) );
  NAND2_X1 U656 ( .A1(n583), .A2(n582), .ZN(n646) );
  NAND2_X1 U657 ( .A1(n584), .A2(n646), .ZN(n585) );
  NAND2_X1 U658 ( .A1(n701), .A2(n587), .ZN(n594) );
  INV_X1 U659 ( .A(n588), .ZN(n592) );
  NAND2_X1 U660 ( .A1(KEYINPUT66), .A2(KEYINPUT2), .ZN(n590) );
  AND2_X1 U661 ( .A1(n590), .A2(n589), .ZN(n591) );
  OR2_X1 U662 ( .A1(n592), .A2(n591), .ZN(n593) );
  NAND2_X1 U663 ( .A1(n594), .A2(n593), .ZN(n596) );
  AND2_X2 U664 ( .A1(n712), .A2(n701), .ZN(n647) );
  NAND2_X1 U665 ( .A1(n647), .A2(KEYINPUT2), .ZN(n595) );
  AND2_X2 U666 ( .A1(n596), .A2(n595), .ZN(n687) );
  NAND2_X1 U667 ( .A1(n687), .A2(G472), .ZN(n600) );
  XOR2_X1 U668 ( .A(KEYINPUT86), .B(KEYINPUT62), .Z(n597) );
  XNOR2_X1 U669 ( .A(n598), .B(n597), .ZN(n599) );
  XNOR2_X1 U670 ( .A(n600), .B(n599), .ZN(n602) );
  INV_X1 U671 ( .A(G952), .ZN(n601) );
  INV_X1 U672 ( .A(KEYINPUT63), .ZN(n603) );
  XNOR2_X1 U673 ( .A(n604), .B(n603), .ZN(G57) );
  NAND2_X1 U674 ( .A1(n687), .A2(G217), .ZN(n607) );
  XNOR2_X1 U675 ( .A(n605), .B(KEYINPUT122), .ZN(n606) );
  XNOR2_X1 U676 ( .A(n607), .B(n606), .ZN(n608) );
  INV_X1 U677 ( .A(KEYINPUT123), .ZN(n609) );
  XNOR2_X1 U678 ( .A(n610), .B(n609), .ZN(G66) );
  XOR2_X1 U679 ( .A(G125), .B(KEYINPUT37), .Z(n611) );
  XNOR2_X1 U680 ( .A(n612), .B(n611), .ZN(G27) );
  XOR2_X1 U681 ( .A(n613), .B(G122), .Z(G24) );
  NAND2_X1 U682 ( .A1(n687), .A2(G210), .ZN(n617) );
  XOR2_X1 U683 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n615) );
  XNOR2_X1 U684 ( .A(n614), .B(n615), .ZN(n616) );
  XNOR2_X1 U685 ( .A(n617), .B(n616), .ZN(n618) );
  XNOR2_X1 U686 ( .A(n619), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U687 ( .A1(n687), .A2(G475), .ZN(n624) );
  XNOR2_X1 U688 ( .A(KEYINPUT119), .B(KEYINPUT120), .ZN(n620) );
  XNOR2_X1 U689 ( .A(n620), .B(KEYINPUT59), .ZN(n621) );
  XNOR2_X1 U690 ( .A(n622), .B(n621), .ZN(n623) );
  XNOR2_X1 U691 ( .A(n624), .B(n623), .ZN(n625) );
  XNOR2_X1 U692 ( .A(n626), .B(KEYINPUT60), .ZN(G60) );
  XNOR2_X1 U693 ( .A(G101), .B(n627), .ZN(n628) );
  XNOR2_X1 U694 ( .A(n628), .B(KEYINPUT113), .ZN(G3) );
  NAND2_X1 U695 ( .A1(n630), .A2(n640), .ZN(n629) );
  XNOR2_X1 U696 ( .A(n629), .B(G104), .ZN(G6) );
  XOR2_X1 U697 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n632) );
  NAND2_X1 U698 ( .A1(n630), .A2(n642), .ZN(n631) );
  XNOR2_X1 U699 ( .A(n632), .B(n631), .ZN(n633) );
  XNOR2_X1 U700 ( .A(G107), .B(n633), .ZN(G9) );
  XOR2_X1 U701 ( .A(G110), .B(n634), .Z(G12) );
  XOR2_X1 U702 ( .A(KEYINPUT29), .B(KEYINPUT114), .Z(n636) );
  NAND2_X1 U703 ( .A1(n638), .A2(n642), .ZN(n635) );
  XNOR2_X1 U704 ( .A(n636), .B(n635), .ZN(n637) );
  XNOR2_X1 U705 ( .A(G128), .B(n637), .ZN(G30) );
  NAND2_X1 U706 ( .A1(n638), .A2(n640), .ZN(n639) );
  XNOR2_X1 U707 ( .A(n639), .B(G146), .ZN(G48) );
  NAND2_X1 U708 ( .A1(n643), .A2(n640), .ZN(n641) );
  XNOR2_X1 U709 ( .A(n641), .B(G113), .ZN(G15) );
  NAND2_X1 U710 ( .A1(n643), .A2(n642), .ZN(n644) );
  XNOR2_X1 U711 ( .A(n644), .B(G116), .ZN(G18) );
  XOR2_X1 U712 ( .A(G134), .B(n645), .Z(G36) );
  XNOR2_X1 U713 ( .A(G140), .B(n646), .ZN(G42) );
  XNOR2_X1 U714 ( .A(n647), .B(KEYINPUT2), .ZN(n684) );
  XOR2_X1 U715 ( .A(KEYINPUT117), .B(KEYINPUT52), .Z(n676) );
  NAND2_X1 U716 ( .A1(n649), .A2(n648), .ZN(n656) );
  NAND2_X1 U717 ( .A1(n651), .A2(n650), .ZN(n652) );
  XOR2_X1 U718 ( .A(KEYINPUT115), .B(n652), .Z(n654) );
  NAND2_X1 U719 ( .A1(n654), .A2(n653), .ZN(n655) );
  NAND2_X1 U720 ( .A1(n656), .A2(n655), .ZN(n657) );
  NAND2_X1 U721 ( .A1(n679), .A2(n657), .ZN(n658) );
  XNOR2_X1 U722 ( .A(n658), .B(KEYINPUT116), .ZN(n674) );
  NOR2_X1 U723 ( .A1(n660), .A2(n659), .ZN(n661) );
  XNOR2_X1 U724 ( .A(n661), .B(KEYINPUT50), .ZN(n668) );
  NOR2_X1 U725 ( .A1(n663), .A2(n662), .ZN(n664) );
  XNOR2_X1 U726 ( .A(n664), .B(KEYINPUT49), .ZN(n665) );
  NAND2_X1 U727 ( .A1(n666), .A2(n665), .ZN(n667) );
  OR2_X1 U728 ( .A1(n668), .A2(n667), .ZN(n669) );
  AND2_X1 U729 ( .A1(n670), .A2(n669), .ZN(n671) );
  XNOR2_X1 U730 ( .A(KEYINPUT51), .B(n671), .ZN(n672) );
  NAND2_X1 U731 ( .A1(n672), .A2(n680), .ZN(n673) );
  NAND2_X1 U732 ( .A1(n674), .A2(n673), .ZN(n675) );
  XOR2_X1 U733 ( .A(n676), .B(n675), .Z(n677) );
  NOR2_X1 U734 ( .A1(n678), .A2(n677), .ZN(n682) );
  AND2_X1 U735 ( .A1(n680), .A2(n679), .ZN(n681) );
  NOR2_X1 U736 ( .A1(n682), .A2(n681), .ZN(n683) );
  NAND2_X1 U737 ( .A1(n684), .A2(n683), .ZN(n685) );
  NOR2_X1 U738 ( .A1(n685), .A2(G953), .ZN(n686) );
  XNOR2_X1 U739 ( .A(n686), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U740 ( .A1(n687), .A2(G469), .ZN(n692) );
  XOR2_X1 U741 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n688) );
  XNOR2_X1 U742 ( .A(n688), .B(KEYINPUT118), .ZN(n689) );
  XNOR2_X1 U743 ( .A(n690), .B(n689), .ZN(n691) );
  XNOR2_X1 U744 ( .A(n692), .B(n691), .ZN(n693) );
  NOR2_X1 U745 ( .A1(n698), .A2(n693), .ZN(G54) );
  NAND2_X1 U746 ( .A1(n687), .A2(G478), .ZN(n696) );
  XNOR2_X1 U747 ( .A(n694), .B(KEYINPUT121), .ZN(n695) );
  XNOR2_X1 U748 ( .A(n696), .B(n695), .ZN(n697) );
  NOR2_X1 U749 ( .A1(n698), .A2(n697), .ZN(G63) );
  NAND2_X1 U750 ( .A1(n700), .A2(n699), .ZN(n707) );
  AND2_X1 U751 ( .A1(n701), .A2(n713), .ZN(n705) );
  NAND2_X1 U752 ( .A1(G953), .A2(G224), .ZN(n702) );
  XNOR2_X1 U753 ( .A(KEYINPUT61), .B(n702), .ZN(n703) );
  AND2_X1 U754 ( .A1(n703), .A2(G898), .ZN(n704) );
  NOR2_X1 U755 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U756 ( .A(n707), .B(n706), .ZN(G69) );
  XNOR2_X1 U757 ( .A(n708), .B(KEYINPUT124), .ZN(n709) );
  XNOR2_X1 U758 ( .A(n710), .B(n709), .ZN(n715) );
  XOR2_X1 U759 ( .A(KEYINPUT125), .B(n715), .Z(n711) );
  XNOR2_X1 U760 ( .A(n712), .B(n711), .ZN(n714) );
  NAND2_X1 U761 ( .A1(n714), .A2(n713), .ZN(n719) );
  XOR2_X1 U762 ( .A(G227), .B(n715), .Z(n716) );
  NAND2_X1 U763 ( .A1(n716), .A2(G900), .ZN(n717) );
  NAND2_X1 U764 ( .A1(n717), .A2(G953), .ZN(n718) );
  NAND2_X1 U765 ( .A1(n719), .A2(n718), .ZN(G72) );
  XOR2_X1 U766 ( .A(G143), .B(n720), .Z(G45) );
  XOR2_X1 U767 ( .A(G119), .B(n721), .Z(G21) );
  XOR2_X1 U768 ( .A(n722), .B(G131), .Z(G33) );
  XOR2_X1 U769 ( .A(n723), .B(G137), .Z(n724) );
  XNOR2_X1 U770 ( .A(KEYINPUT126), .B(n724), .ZN(G39) );
endmodule

