//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 0 1 1 0 0 0 1 0 1 1 0 1 1 0 0 1 1 1 0 1 0 0 1 0 1 0 0 1 1 1 0 0 0 0 0 0 1 0 0 1 1 1 0 0 0 1 1 1 0 1 1 1 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:07 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n615, new_n616, new_n617,
    new_n618, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n641, new_n642, new_n643, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n713, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965;
  INV_X1    g000(.A(KEYINPUT69), .ZN(new_n187));
  INV_X1    g001(.A(G119), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G116), .ZN(new_n189));
  INV_X1    g003(.A(G116), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G119), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n189), .A2(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT2), .B(G113), .ZN(new_n193));
  XOR2_X1   g007(.A(new_n192), .B(new_n193), .Z(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n196));
  INV_X1    g010(.A(G137), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G134), .ZN(new_n198));
  NOR2_X1   g012(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n196), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G131), .ZN(new_n201));
  INV_X1    g015(.A(G134), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G137), .ZN(new_n203));
  NAND4_X1  g017(.A1(new_n197), .A2(KEYINPUT65), .A3(KEYINPUT11), .A4(G134), .ZN(new_n204));
  NAND4_X1  g018(.A1(new_n200), .A2(new_n201), .A3(new_n203), .A4(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(KEYINPUT66), .ZN(new_n206));
  AND2_X1   g020(.A1(new_n204), .A2(new_n203), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT66), .ZN(new_n208));
  NAND4_X1  g022(.A1(new_n207), .A2(new_n208), .A3(new_n201), .A4(new_n200), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n206), .A2(new_n209), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n201), .B1(new_n198), .B2(new_n203), .ZN(new_n211));
  XOR2_X1   g025(.A(new_n211), .B(KEYINPUT67), .Z(new_n212));
  INV_X1    g026(.A(KEYINPUT64), .ZN(new_n213));
  INV_X1    g027(.A(G143), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n213), .B1(new_n214), .B2(G146), .ZN(new_n215));
  INV_X1    g029(.A(G146), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n216), .A2(KEYINPUT64), .A3(G143), .ZN(new_n217));
  INV_X1    g031(.A(G128), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n218), .A2(KEYINPUT1), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n214), .A2(G146), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n215), .A2(new_n217), .A3(new_n219), .A4(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n216), .A2(G143), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n218), .B1(new_n222), .B2(KEYINPUT1), .ZN(new_n223));
  XNOR2_X1  g037(.A(G143), .B(G146), .ZN(new_n224));
  NOR3_X1   g038(.A1(new_n223), .A2(new_n224), .A3(KEYINPUT68), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT68), .ZN(new_n226));
  OAI21_X1  g040(.A(KEYINPUT1), .B1(new_n214), .B2(G146), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(G128), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n222), .A2(new_n220), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n226), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n221), .B1(new_n225), .B2(new_n230), .ZN(new_n231));
  AND3_X1   g045(.A1(new_n210), .A2(new_n212), .A3(new_n231), .ZN(new_n232));
  AND3_X1   g046(.A1(new_n215), .A2(new_n217), .A3(new_n220), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n233), .A2(KEYINPUT0), .A3(G128), .ZN(new_n234));
  NAND2_X1  g048(.A1(KEYINPUT0), .A2(G128), .ZN(new_n235));
  OR2_X1    g049(.A1(KEYINPUT0), .A2(G128), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n229), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n234), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n207), .A2(new_n200), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G131), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n238), .B1(new_n210), .B2(new_n240), .ZN(new_n241));
  NOR3_X1   g055(.A1(new_n232), .A2(new_n241), .A3(KEYINPUT30), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT30), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n210), .A2(new_n240), .ZN(new_n244));
  AND2_X1   g058(.A1(new_n234), .A2(new_n237), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n210), .A2(new_n212), .A3(new_n231), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n243), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  OAI211_X1 g062(.A(new_n187), .B(new_n195), .C1(new_n242), .C2(new_n248), .ZN(new_n249));
  NOR2_X1   g063(.A1(G237), .A2(G953), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(G210), .ZN(new_n251));
  XOR2_X1   g065(.A(new_n251), .B(KEYINPUT27), .Z(new_n252));
  XNOR2_X1  g066(.A(KEYINPUT26), .B(G101), .ZN(new_n253));
  XNOR2_X1  g067(.A(new_n252), .B(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  OAI21_X1  g069(.A(KEYINPUT30), .B1(new_n232), .B2(new_n241), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n246), .A2(new_n243), .A3(new_n247), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n194), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  AOI22_X1  g072(.A1(new_n206), .A2(new_n209), .B1(G131), .B2(new_n239), .ZN(new_n259));
  OAI211_X1 g073(.A(new_n247), .B(new_n194), .C1(new_n259), .C2(new_n238), .ZN(new_n260));
  AND2_X1   g074(.A1(new_n260), .A2(new_n187), .ZN(new_n261));
  OAI211_X1 g075(.A(new_n249), .B(new_n255), .C1(new_n258), .C2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(KEYINPUT31), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT70), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT28), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n195), .B1(new_n232), .B2(new_n241), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n266), .B1(new_n267), .B2(new_n260), .ZN(new_n268));
  AND2_X1   g082(.A1(new_n260), .A2(new_n266), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n254), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT71), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  OAI211_X1 g086(.A(KEYINPUT71), .B(new_n254), .C1(new_n268), .C2(new_n269), .ZN(new_n273));
  AND2_X1   g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n262), .A2(KEYINPUT70), .A3(KEYINPUT31), .ZN(new_n275));
  OR2_X1    g089(.A1(new_n258), .A2(new_n261), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT31), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n276), .A2(new_n277), .A3(new_n255), .A4(new_n249), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n265), .A2(new_n274), .A3(new_n275), .A4(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(G472), .ZN(new_n280));
  INV_X1    g094(.A(G902), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n279), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT32), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n279), .A2(KEYINPUT32), .A3(new_n280), .A4(new_n281), .ZN(new_n285));
  NOR3_X1   g099(.A1(new_n268), .A2(new_n269), .A3(new_n254), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n276), .A2(new_n249), .ZN(new_n287));
  AOI211_X1 g101(.A(KEYINPUT29), .B(new_n286), .C1(new_n287), .C2(new_n254), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n286), .A2(KEYINPUT29), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(new_n281), .ZN(new_n290));
  OAI21_X1  g104(.A(G472), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n284), .A2(new_n285), .A3(new_n291), .ZN(new_n292));
  XNOR2_X1  g106(.A(KEYINPUT9), .B(G234), .ZN(new_n293));
  OAI21_X1  g107(.A(G221), .B1(new_n293), .B2(G902), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(G469), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT77), .ZN(new_n297));
  INV_X1    g111(.A(G104), .ZN(new_n298));
  OAI21_X1  g112(.A(KEYINPUT3), .B1(new_n298), .B2(G107), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT3), .ZN(new_n300));
  INV_X1    g114(.A(G107), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n300), .A2(new_n301), .A3(G104), .ZN(new_n302));
  INV_X1    g116(.A(G101), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n298), .A2(G107), .ZN(new_n304));
  NAND4_X1  g118(.A1(new_n299), .A2(new_n302), .A3(new_n303), .A4(new_n304), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n298), .A2(G107), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n301), .A2(G104), .ZN(new_n307));
  OAI21_X1  g121(.A(G101), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  AND2_X1   g122(.A1(new_n305), .A2(new_n308), .ZN(new_n309));
  NAND4_X1  g123(.A1(new_n231), .A2(new_n297), .A3(KEYINPUT10), .A4(new_n309), .ZN(new_n310));
  OAI21_X1  g124(.A(KEYINPUT68), .B1(new_n223), .B2(new_n224), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n228), .A2(new_n226), .A3(new_n229), .ZN(new_n312));
  AOI22_X1  g126(.A1(new_n311), .A2(new_n312), .B1(new_n233), .B2(new_n219), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n305), .A2(new_n308), .A3(KEYINPUT10), .ZN(new_n314));
  OAI21_X1  g128(.A(KEYINPUT77), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n310), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n299), .A2(new_n302), .A3(new_n304), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT76), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND4_X1  g133(.A1(new_n299), .A2(new_n302), .A3(KEYINPUT76), .A4(new_n304), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT4), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n321), .A2(new_n322), .A3(G101), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n303), .B1(new_n319), .B2(new_n320), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n305), .A2(KEYINPUT4), .ZN(new_n325));
  OAI211_X1 g139(.A(new_n245), .B(new_n323), .C1(new_n324), .C2(new_n325), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n221), .B1(new_n233), .B2(new_n223), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(new_n309), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT10), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n316), .A2(new_n259), .A3(new_n326), .A4(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT80), .ZN(new_n332));
  XNOR2_X1  g146(.A(G110), .B(G140), .ZN(new_n333));
  INV_X1    g147(.A(G227), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n334), .A2(G953), .ZN(new_n335));
  XOR2_X1   g149(.A(new_n333), .B(new_n335), .Z(new_n336));
  AND3_X1   g150(.A1(new_n331), .A2(new_n332), .A3(new_n336), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n332), .B1(new_n331), .B2(new_n336), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT78), .ZN(new_n339));
  AOI21_X1  g153(.A(KEYINPUT12), .B1(new_n244), .B2(new_n339), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n328), .B1(new_n231), .B2(new_n309), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(new_n244), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  OAI211_X1 g157(.A(new_n341), .B(new_n244), .C1(new_n339), .C2(KEYINPUT12), .ZN(new_n344));
  AND2_X1   g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NOR3_X1   g159(.A1(new_n337), .A2(new_n338), .A3(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n316), .A2(new_n326), .A3(new_n330), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(new_n244), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n336), .B1(new_n348), .B2(new_n331), .ZN(new_n349));
  OAI211_X1 g163(.A(new_n296), .B(new_n281), .C1(new_n346), .C2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(KEYINPUT81), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n331), .A2(new_n336), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(KEYINPUT80), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n331), .A2(new_n332), .A3(new_n336), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n343), .A2(new_n344), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(new_n349), .ZN(new_n357));
  AOI21_X1  g171(.A(G902), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT81), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n358), .A2(new_n359), .A3(new_n296), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n351), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n355), .A2(new_n331), .ZN(new_n362));
  INV_X1    g176(.A(new_n336), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n348), .A2(new_n336), .A3(new_n331), .ZN(new_n365));
  AOI21_X1  g179(.A(G902), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NOR3_X1   g180(.A1(new_n366), .A2(KEYINPUT79), .A3(new_n296), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT79), .ZN(new_n368));
  AND3_X1   g182(.A1(new_n348), .A2(new_n336), .A3(new_n331), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n336), .B1(new_n355), .B2(new_n331), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n281), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n368), .B1(new_n371), .B2(G469), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n367), .A2(new_n372), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n295), .B1(new_n361), .B2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(G475), .ZN(new_n375));
  INV_X1    g189(.A(G237), .ZN(new_n376));
  INV_X1    g190(.A(G953), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n376), .A2(new_n377), .A3(G214), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(new_n214), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n250), .A2(G143), .A3(G214), .ZN(new_n380));
  NAND2_X1  g194(.A1(KEYINPUT18), .A2(G131), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n379), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(KEYINPUT86), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT86), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n379), .A2(new_n384), .A3(new_n380), .A4(new_n381), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT18), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n379), .A2(new_n380), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(G131), .ZN(new_n389));
  INV_X1    g203(.A(G140), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(G125), .ZN(new_n391));
  INV_X1    g205(.A(G125), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(G140), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT73), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n391), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n390), .A2(KEYINPUT73), .A3(G125), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n395), .A2(G146), .A3(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT85), .ZN(new_n398));
  XNOR2_X1  g212(.A(G125), .B(G140), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(new_n216), .ZN(new_n400));
  AND3_X1   g214(.A1(new_n397), .A2(new_n398), .A3(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n398), .B1(new_n397), .B2(new_n400), .ZN(new_n402));
  OAI221_X1 g216(.A(new_n386), .B1(new_n387), .B2(new_n389), .C1(new_n401), .C2(new_n402), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n395), .A2(KEYINPUT16), .A3(new_n396), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT16), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n391), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(G146), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT17), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n379), .A2(new_n201), .A3(new_n380), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n389), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n404), .A2(new_n216), .A3(new_n406), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n388), .A2(KEYINPUT17), .A3(G131), .ZN(new_n413));
  NAND4_X1  g227(.A1(new_n408), .A2(new_n411), .A3(new_n412), .A4(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n403), .A2(new_n414), .ZN(new_n415));
  XNOR2_X1  g229(.A(G113), .B(G122), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n416), .B(new_n298), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n415), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n403), .A2(new_n417), .A3(new_n414), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n375), .B1(new_n421), .B2(new_n281), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  AND3_X1   g237(.A1(new_n403), .A2(new_n417), .A3(new_n414), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT87), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT19), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n399), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  AOI22_X1  g241(.A1(new_n395), .A2(new_n396), .B1(new_n399), .B2(KEYINPUT87), .ZN(new_n428));
  OAI211_X1 g242(.A(new_n216), .B(new_n427), .C1(new_n428), .C2(new_n426), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT88), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n429), .A2(new_n408), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n389), .A2(new_n410), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n430), .B1(new_n429), .B2(new_n408), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n403), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n424), .B1(new_n435), .B2(new_n418), .ZN(new_n436));
  NOR2_X1   g250(.A1(G475), .A2(G902), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  NOR3_X1   g252(.A1(new_n436), .A2(KEYINPUT20), .A3(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT20), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n435), .A2(new_n418), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(new_n420), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n440), .B1(new_n442), .B2(new_n437), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n423), .B1(new_n439), .B2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT89), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(KEYINPUT20), .B1(new_n436), .B2(new_n438), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n442), .A2(new_n440), .A3(new_n437), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n449), .A2(KEYINPUT89), .A3(new_n423), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n446), .A2(new_n450), .ZN(new_n451));
  AOI21_X1  g265(.A(KEYINPUT13), .B1(new_n218), .B2(G143), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n452), .A2(new_n202), .ZN(new_n453));
  XNOR2_X1  g267(.A(G128), .B(G143), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n453), .B(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n190), .A2(G122), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n190), .A2(G122), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT90), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  OAI21_X1  g275(.A(KEYINPUT90), .B1(new_n457), .B2(new_n458), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(new_n301), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n463), .A2(new_n301), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n455), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n454), .B(new_n202), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n456), .B1(new_n458), .B2(KEYINPUT14), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT91), .ZN(new_n470));
  OAI22_X1  g284(.A1(new_n469), .A2(new_n470), .B1(KEYINPUT14), .B2(new_n456), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n471), .B1(new_n470), .B2(new_n469), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n464), .B(new_n468), .C1(new_n472), .C2(new_n301), .ZN(new_n473));
  INV_X1    g287(.A(G217), .ZN(new_n474));
  NOR3_X1   g288(.A1(new_n293), .A2(new_n474), .A3(G953), .ZN(new_n475));
  AND3_X1   g289(.A1(new_n467), .A2(new_n473), .A3(new_n475), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n475), .B1(new_n467), .B2(new_n473), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n281), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(G478), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n479), .A2(KEYINPUT15), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n478), .B(new_n481), .ZN(new_n482));
  AND2_X1   g296(.A1(new_n377), .A2(G952), .ZN(new_n483));
  INV_X1    g297(.A(G234), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n483), .B1(new_n484), .B2(new_n376), .ZN(new_n485));
  XOR2_X1   g299(.A(new_n485), .B(KEYINPUT92), .Z(new_n486));
  OAI211_X1 g300(.A(G902), .B(G953), .C1(new_n484), .C2(new_n376), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n487), .B(KEYINPUT93), .ZN(new_n488));
  XOR2_X1   g302(.A(KEYINPUT21), .B(G898), .Z(new_n489));
  OAI21_X1  g303(.A(new_n486), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n482), .A2(new_n490), .ZN(new_n491));
  OAI21_X1  g305(.A(G214), .B1(G237), .B2(G902), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n234), .A2(G125), .A3(new_n237), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n493), .B1(new_n313), .B2(G125), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n377), .A2(G224), .ZN(new_n495));
  XOR2_X1   g309(.A(new_n495), .B(KEYINPUT83), .Z(new_n496));
  NAND3_X1  g310(.A1(new_n494), .A2(KEYINPUT7), .A3(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT84), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT7), .ZN(new_n499));
  INV_X1    g313(.A(new_n495), .ZN(new_n500));
  OAI221_X1 g314(.A(new_n493), .B1(new_n499), .B2(new_n500), .C1(new_n313), .C2(G125), .ZN(new_n501));
  OR2_X1    g315(.A1(new_n192), .A2(new_n193), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT5), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n503), .A2(new_n188), .A3(G116), .ZN(new_n504));
  OAI211_X1 g318(.A(G113), .B(new_n504), .C1(new_n192), .C2(new_n503), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n305), .A2(new_n308), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n309), .A2(new_n502), .A3(new_n505), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  XOR2_X1   g324(.A(KEYINPUT82), .B(KEYINPUT8), .Z(new_n511));
  XNOR2_X1  g325(.A(G110), .B(G122), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n511), .B(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n497), .A2(new_n498), .A3(new_n501), .A4(new_n514), .ZN(new_n515));
  OAI211_X1 g329(.A(new_n195), .B(new_n323), .C1(new_n324), .C2(new_n325), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n516), .A2(new_n509), .A3(new_n512), .ZN(new_n517));
  AND2_X1   g331(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n497), .A2(new_n501), .A3(new_n514), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(KEYINPUT84), .ZN(new_n520));
  AOI21_X1  g334(.A(G902), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  OAI21_X1  g335(.A(G210), .B1(G237), .B2(G902), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n512), .B1(new_n516), .B2(new_n509), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n524), .A2(KEYINPUT6), .A3(new_n517), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n494), .B(new_n495), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n517), .A2(KEYINPUT6), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(new_n523), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n525), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  AND3_X1   g343(.A1(new_n521), .A2(new_n522), .A3(new_n529), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n522), .B1(new_n521), .B2(new_n529), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n492), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NOR3_X1   g346(.A1(new_n451), .A2(new_n491), .A3(new_n532), .ZN(new_n533));
  AND2_X1   g347(.A1(new_n374), .A2(new_n533), .ZN(new_n534));
  XNOR2_X1  g348(.A(KEYINPUT22), .B(G137), .ZN(new_n535));
  AND3_X1   g349(.A1(new_n377), .A2(G221), .A3(G234), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n535), .B(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n408), .A2(new_n412), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT23), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n539), .B1(new_n188), .B2(G128), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n188), .A2(G128), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n218), .A2(KEYINPUT23), .A3(G119), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(G110), .ZN(new_n544));
  OR3_X1    g358(.A1(new_n188), .A2(KEYINPUT72), .A3(G128), .ZN(new_n545));
  OAI21_X1  g359(.A(KEYINPUT72), .B1(new_n188), .B2(G128), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n545), .A2(new_n541), .A3(new_n546), .ZN(new_n547));
  XNOR2_X1  g361(.A(KEYINPUT24), .B(G110), .ZN(new_n548));
  OAI211_X1 g362(.A(new_n538), .B(new_n544), .C1(new_n547), .C2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n547), .A2(new_n548), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n550), .B1(G110), .B2(new_n543), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n551), .A2(new_n408), .A3(new_n400), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n537), .B1(new_n549), .B2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n549), .A2(new_n552), .A3(new_n537), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n474), .B1(G234), .B2(new_n281), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n557), .A2(G902), .ZN(new_n558));
  XOR2_X1   g372(.A(new_n558), .B(KEYINPUT74), .Z(new_n559));
  NAND2_X1  g373(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  XOR2_X1   g374(.A(new_n560), .B(KEYINPUT75), .Z(new_n561));
  INV_X1    g375(.A(KEYINPUT25), .ZN(new_n562));
  INV_X1    g376(.A(new_n555), .ZN(new_n563));
  OAI211_X1 g377(.A(new_n562), .B(new_n281), .C1(new_n563), .C2(new_n553), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(new_n557), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n562), .B1(new_n556), .B2(new_n281), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n561), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n292), .A2(new_n534), .A3(new_n568), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n569), .B(G101), .ZN(G3));
  INV_X1    g384(.A(new_n282), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n280), .B1(new_n279), .B2(new_n281), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  OR2_X1    g387(.A1(new_n476), .A2(new_n477), .ZN(new_n574));
  XOR2_X1   g388(.A(new_n574), .B(KEYINPUT33), .Z(new_n575));
  NAND2_X1  g389(.A1(new_n281), .A2(G478), .ZN(new_n576));
  INV_X1    g390(.A(new_n478), .ZN(new_n577));
  XOR2_X1   g391(.A(KEYINPUT94), .B(G478), .Z(new_n578));
  OAI22_X1  g392(.A1(new_n575), .A2(new_n576), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n451), .A2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n492), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n521), .A2(new_n529), .ZN(new_n582));
  INV_X1    g396(.A(new_n522), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n521), .A2(new_n529), .A3(new_n522), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n581), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(new_n490), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n580), .A2(new_n587), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n573), .A2(new_n568), .A3(new_n374), .A4(new_n588), .ZN(new_n589));
  XOR2_X1   g403(.A(KEYINPUT34), .B(G104), .Z(new_n590));
  XNOR2_X1  g404(.A(new_n589), .B(new_n590), .ZN(G6));
  NAND2_X1  g405(.A1(new_n279), .A2(new_n281), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(G472), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n593), .A2(new_n374), .A3(new_n282), .A4(new_n568), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT96), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n439), .A2(KEYINPUT95), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n596), .B(new_n443), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n482), .A2(new_n422), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n595), .B1(new_n599), .B2(new_n587), .ZN(new_n600));
  INV_X1    g414(.A(new_n587), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n601), .A2(KEYINPUT96), .A3(new_n597), .A4(new_n598), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n594), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(KEYINPUT35), .B(G107), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n603), .B(new_n604), .ZN(G9));
  NAND2_X1  g419(.A1(new_n549), .A2(new_n552), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n537), .A2(KEYINPUT36), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n606), .B(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(new_n559), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n609), .B1(new_n565), .B2(new_n566), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n610), .B(KEYINPUT97), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n534), .A2(new_n573), .A3(new_n611), .ZN(new_n612));
  XOR2_X1   g426(.A(KEYINPUT37), .B(G110), .Z(new_n613));
  XNOR2_X1  g427(.A(new_n612), .B(new_n613), .ZN(G12));
  AND2_X1   g428(.A1(new_n611), .A2(new_n586), .ZN(new_n615));
  OR2_X1    g429(.A1(new_n488), .A2(G900), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n599), .B1(new_n486), .B2(new_n616), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n292), .A2(new_n374), .A3(new_n615), .A4(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(G128), .ZN(G30));
  NAND2_X1  g433(.A1(new_n616), .A2(new_n486), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n620), .B(KEYINPUT39), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n374), .A2(new_n621), .ZN(new_n622));
  XOR2_X1   g436(.A(new_n622), .B(KEYINPUT40), .Z(new_n623));
  AOI21_X1  g437(.A(new_n255), .B1(new_n267), .B2(new_n260), .ZN(new_n624));
  XOR2_X1   g438(.A(new_n624), .B(KEYINPUT99), .Z(new_n625));
  INV_X1    g439(.A(new_n262), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n281), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(G472), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n284), .A2(new_n628), .A3(new_n285), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n584), .A2(new_n585), .ZN(new_n630));
  XNOR2_X1  g444(.A(KEYINPUT98), .B(KEYINPUT38), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n610), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n632), .A2(new_n492), .A3(new_n633), .ZN(new_n634));
  AOI21_X1  g448(.A(KEYINPUT89), .B1(new_n449), .B2(new_n423), .ZN(new_n635));
  AOI211_X1 g449(.A(new_n445), .B(new_n422), .C1(new_n447), .C2(new_n448), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NOR3_X1   g451(.A1(new_n634), .A2(new_n637), .A3(new_n482), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n623), .A2(new_n629), .A3(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(G143), .ZN(G45));
  NAND3_X1  g454(.A1(new_n451), .A2(new_n579), .A3(new_n620), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n292), .A2(new_n374), .A3(new_n615), .A4(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(G146), .ZN(G48));
  NAND2_X1  g458(.A1(new_n356), .A2(new_n357), .ZN(new_n645));
  AND3_X1   g459(.A1(new_n645), .A2(KEYINPUT100), .A3(new_n281), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n358), .A2(KEYINPUT100), .ZN(new_n647));
  OAI21_X1  g461(.A(G469), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(new_n361), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n649), .A2(new_n295), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n292), .A2(new_n568), .A3(new_n588), .A4(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(KEYINPUT41), .B(G113), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G15));
  NAND2_X1  g467(.A1(new_n602), .A2(new_n600), .ZN(new_n654));
  AND4_X1   g468(.A1(new_n292), .A2(new_n654), .A3(new_n568), .A4(new_n650), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(new_n190), .ZN(G18));
  NOR3_X1   g470(.A1(new_n635), .A2(new_n636), .A3(new_n491), .ZN(new_n657));
  AND4_X1   g471(.A1(new_n294), .A2(new_n657), .A3(new_n648), .A4(new_n361), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n292), .A2(new_n615), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G119), .ZN(G21));
  OAI21_X1  g474(.A(KEYINPUT101), .B1(new_n637), .B2(new_n482), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT101), .ZN(new_n662));
  INV_X1    g476(.A(new_n482), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n451), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n532), .B1(new_n661), .B2(new_n664), .ZN(new_n665));
  AND4_X1   g479(.A1(new_n294), .A2(new_n648), .A3(new_n361), .A4(new_n490), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n280), .A2(new_n281), .ZN(new_n667));
  AND2_X1   g481(.A1(new_n263), .A2(new_n270), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n667), .B1(new_n668), .B2(new_n278), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n572), .A2(new_n669), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n665), .A2(new_n666), .A3(new_n568), .A4(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G122), .ZN(G24));
  NOR3_X1   g486(.A1(new_n649), .A2(new_n295), .A3(new_n532), .ZN(new_n673));
  NOR3_X1   g487(.A1(new_n572), .A2(new_n633), .A3(new_n669), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n673), .A2(new_n642), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G125), .ZN(G27));
  OAI211_X1 g490(.A(new_n272), .B(new_n273), .C1(new_n262), .C2(KEYINPUT31), .ZN(new_n677));
  AOI21_X1  g491(.A(KEYINPUT70), .B1(new_n262), .B2(KEYINPUT31), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  AOI21_X1  g493(.A(G902), .B1(new_n679), .B2(new_n275), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n680), .A2(KEYINPUT105), .A3(KEYINPUT32), .A4(new_n280), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT105), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n285), .A2(new_n682), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n681), .A2(new_n683), .A3(new_n284), .A4(new_n291), .ZN(new_n684));
  AND3_X1   g498(.A1(new_n684), .A2(KEYINPUT42), .A3(new_n568), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n630), .A2(new_n581), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(new_n294), .ZN(new_n687));
  AND4_X1   g501(.A1(new_n359), .A2(new_n645), .A3(new_n296), .A4(new_n281), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n359), .B1(new_n358), .B2(new_n296), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT103), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n365), .B(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT102), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n692), .B1(new_n362), .B2(new_n363), .ZN(new_n693));
  AOI211_X1 g507(.A(KEYINPUT102), .B(new_n336), .C1(new_n355), .C2(new_n331), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  AOI21_X1  g509(.A(G902), .B1(new_n691), .B2(new_n695), .ZN(new_n696));
  OAI22_X1  g510(.A1(new_n688), .A2(new_n689), .B1(new_n696), .B2(new_n296), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT104), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  OAI211_X1 g513(.A(new_n361), .B(KEYINPUT104), .C1(new_n296), .C2(new_n696), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n687), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(new_n642), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n685), .A2(KEYINPUT106), .A3(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT106), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n684), .A2(KEYINPUT42), .A3(new_n568), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n705), .B1(new_n706), .B2(new_n702), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT42), .ZN(new_n708));
  AND2_X1   g522(.A1(new_n292), .A2(new_n568), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n709), .A2(new_n642), .A3(new_n701), .ZN(new_n710));
  AOI22_X1  g524(.A1(new_n704), .A2(new_n707), .B1(new_n708), .B2(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(new_n201), .ZN(G33));
  NAND4_X1  g526(.A1(new_n701), .A2(new_n292), .A3(new_n568), .A4(new_n617), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G134), .ZN(G36));
  XNOR2_X1  g528(.A(new_n451), .B(KEYINPUT107), .ZN(new_n715));
  AND2_X1   g529(.A1(new_n715), .A2(new_n579), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(KEYINPUT43), .ZN(new_n717));
  AND2_X1   g531(.A1(new_n637), .A2(new_n579), .ZN(new_n718));
  OR2_X1    g532(.A1(new_n718), .A2(KEYINPUT43), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n573), .A2(new_n633), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n720), .A2(KEYINPUT44), .A3(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(KEYINPUT108), .ZN(new_n723));
  AOI21_X1  g537(.A(KEYINPUT44), .B1(new_n720), .B2(new_n721), .ZN(new_n724));
  INV_X1    g538(.A(new_n686), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n691), .A2(new_n695), .A3(KEYINPUT45), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n369), .A2(new_n370), .ZN(new_n727));
  OAI211_X1 g541(.A(new_n726), .B(G469), .C1(KEYINPUT45), .C2(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(G469), .A2(G902), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n728), .A2(KEYINPUT46), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(new_n361), .ZN(new_n731));
  AOI21_X1  g545(.A(KEYINPUT46), .B1(new_n728), .B2(new_n729), .ZN(new_n732));
  OR2_X1    g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n733), .A2(new_n294), .A3(new_n621), .ZN(new_n734));
  NOR3_X1   g548(.A1(new_n724), .A2(new_n725), .A3(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n723), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(KEYINPUT109), .B(G137), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n736), .B(new_n737), .ZN(G39));
  NOR4_X1   g552(.A1(new_n292), .A2(new_n568), .A3(new_n641), .A4(new_n725), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n733), .A2(KEYINPUT47), .A3(new_n294), .ZN(new_n740));
  INV_X1    g554(.A(new_n740), .ZN(new_n741));
  AOI21_X1  g555(.A(KEYINPUT47), .B1(new_n733), .B2(new_n294), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n739), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G140), .ZN(G42));
  NOR3_X1   g558(.A1(new_n629), .A2(new_n567), .A3(new_n561), .ZN(new_n745));
  XOR2_X1   g559(.A(new_n649), .B(KEYINPUT49), .Z(new_n746));
  NOR3_X1   g560(.A1(new_n632), .A2(new_n295), .A3(new_n581), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n745), .A2(new_n746), .A3(new_n716), .A4(new_n747), .ZN(new_n748));
  AND3_X1   g562(.A1(new_n569), .A2(new_n659), .A3(new_n671), .ZN(new_n749));
  INV_X1    g563(.A(new_n588), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n593), .A2(new_n282), .A3(new_n611), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n374), .A2(new_n533), .ZN(new_n752));
  OAI22_X1  g566(.A1(new_n594), .A2(new_n750), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n446), .A2(new_n450), .A3(new_n663), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT110), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n446), .A2(KEYINPUT110), .A3(new_n450), .A4(new_n663), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(new_n601), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n594), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n753), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n709), .A2(new_n654), .A3(new_n650), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n749), .A2(new_n651), .A3(new_n761), .A4(new_n762), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n701), .A2(new_n642), .A3(new_n674), .ZN(new_n764));
  AND3_X1   g578(.A1(new_n482), .A2(new_n423), .A3(new_n620), .ZN(new_n765));
  AND4_X1   g579(.A1(new_n597), .A2(new_n611), .A3(new_n686), .A4(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n292), .A2(new_n374), .A3(new_n766), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n713), .A2(new_n764), .A3(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT111), .ZN(new_n769));
  AND2_X1   g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n763), .A2(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT112), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n710), .A2(new_n708), .ZN(new_n773));
  AOI21_X1  g587(.A(KEYINPUT106), .B1(new_n685), .B2(new_n703), .ZN(new_n774));
  NOR3_X1   g588(.A1(new_n706), .A2(new_n705), .A3(new_n702), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n773), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n713), .A2(new_n764), .A3(KEYINPUT111), .A4(new_n767), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n771), .A2(new_n772), .A3(new_n776), .A4(new_n777), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n587), .B1(new_n756), .B2(new_n757), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n573), .A2(new_n779), .A3(new_n568), .A4(new_n374), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n651), .A2(new_n589), .A3(new_n612), .A4(new_n780), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n781), .A2(new_n655), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n768), .A2(new_n769), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n782), .A2(new_n783), .A3(new_n777), .A4(new_n749), .ZN(new_n784));
  OAI21_X1  g598(.A(KEYINPUT112), .B1(new_n784), .B2(new_n711), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n778), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n699), .A2(new_n700), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n620), .B(KEYINPUT113), .ZN(new_n788));
  NOR3_X1   g602(.A1(new_n610), .A2(new_n295), .A3(new_n788), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n629), .A2(new_n665), .A3(new_n787), .A4(new_n789), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n618), .A2(new_n643), .A3(new_n790), .A4(new_n675), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(KEYINPUT114), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT52), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT114), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n791), .B(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n796), .A2(KEYINPUT52), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n794), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n786), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(KEYINPUT53), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT53), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n791), .A2(new_n793), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n802), .B1(new_n792), .B2(new_n793), .ZN(new_n803));
  INV_X1    g617(.A(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n786), .A2(new_n801), .A3(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n800), .A2(KEYINPUT54), .A3(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT115), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n771), .A2(new_n776), .A3(new_n777), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n808), .A2(new_n801), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n809), .A2(new_n804), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT54), .ZN(new_n811));
  AOI22_X1  g625(.A1(new_n778), .A2(new_n785), .B1(new_n794), .B2(new_n797), .ZN(new_n812));
  OAI211_X1 g626(.A(new_n810), .B(new_n811), .C1(new_n812), .C2(KEYINPUT53), .ZN(new_n813));
  AND3_X1   g627(.A1(new_n806), .A2(new_n807), .A3(new_n813), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n807), .B1(new_n806), .B2(new_n813), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n486), .B1(new_n717), .B2(new_n719), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n649), .A2(new_n687), .ZN(new_n817));
  AND2_X1   g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(new_n674), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n649), .A2(new_n687), .A3(new_n486), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n745), .A2(new_n820), .ZN(new_n821));
  OR3_X1    g635(.A1(new_n821), .A2(new_n451), .A3(new_n579), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n819), .A2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(new_n486), .ZN(new_n824));
  AND2_X1   g638(.A1(new_n670), .A2(new_n568), .ZN(new_n825));
  NOR4_X1   g639(.A1(new_n632), .A2(new_n649), .A3(new_n295), .A4(new_n492), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n720), .A2(new_n824), .A3(new_n825), .A4(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT50), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT118), .ZN(new_n830));
  XNOR2_X1  g644(.A(new_n829), .B(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n827), .A2(new_n828), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT117), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n832), .B(new_n833), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n823), .B1(new_n831), .B2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT116), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT51), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n831), .A2(new_n834), .ZN(new_n839));
  INV_X1    g653(.A(new_n823), .ZN(new_n840));
  INV_X1    g654(.A(new_n742), .ZN(new_n841));
  OAI211_X1 g655(.A(new_n841), .B(new_n740), .C1(new_n294), .C2(new_n649), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n842), .A2(new_n825), .A3(new_n686), .A4(new_n816), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n839), .A2(new_n840), .A3(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n837), .A2(new_n838), .A3(new_n844), .ZN(new_n845));
  OAI211_X1 g659(.A(new_n835), .B(new_n843), .C1(new_n836), .C2(KEYINPUT51), .ZN(new_n846));
  AND2_X1   g660(.A1(new_n684), .A2(new_n568), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n818), .A2(new_n847), .ZN(new_n848));
  OR2_X1    g662(.A1(new_n848), .A2(KEYINPUT119), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n848), .A2(KEYINPUT119), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n849), .A2(KEYINPUT48), .A3(new_n850), .ZN(new_n851));
  AOI21_X1  g665(.A(KEYINPUT48), .B1(new_n849), .B2(new_n850), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n816), .A2(new_n825), .A3(new_n673), .ZN(new_n853));
  OAI211_X1 g667(.A(new_n853), .B(new_n483), .C1(new_n580), .C2(new_n821), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n851), .A2(new_n852), .A3(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n845), .A2(new_n846), .A3(new_n855), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n814), .A2(new_n815), .A3(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(G952), .A2(G953), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n748), .B1(new_n857), .B2(new_n858), .ZN(G75));
  NAND2_X1  g673(.A1(new_n525), .A2(new_n528), .ZN(new_n860));
  XNOR2_X1  g674(.A(new_n860), .B(new_n526), .ZN(new_n861));
  INV_X1    g675(.A(new_n861), .ZN(new_n862));
  AOI21_X1  g676(.A(KEYINPUT53), .B1(new_n786), .B2(new_n798), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n803), .A2(new_n808), .A3(new_n801), .ZN(new_n864));
  OAI211_X1 g678(.A(G210), .B(G902), .C1(new_n863), .C2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT55), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT120), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n867), .A2(KEYINPUT56), .ZN(new_n868));
  AND3_X1   g682(.A1(new_n865), .A2(new_n866), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n866), .B1(new_n865), .B2(new_n868), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n862), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n865), .A2(new_n868), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n872), .A2(KEYINPUT55), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n865), .A2(new_n866), .A3(new_n868), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n873), .A2(new_n861), .A3(new_n874), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n377), .A2(G952), .ZN(new_n876));
  INV_X1    g690(.A(new_n876), .ZN(new_n877));
  AND3_X1   g691(.A1(new_n871), .A2(new_n875), .A3(new_n877), .ZN(G51));
  XOR2_X1   g692(.A(new_n729), .B(KEYINPUT57), .Z(new_n879));
  NAND2_X1  g693(.A1(new_n799), .A2(new_n801), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n811), .B1(new_n880), .B2(new_n810), .ZN(new_n881));
  INV_X1    g695(.A(new_n813), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n879), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n883), .A2(new_n645), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n880), .A2(new_n810), .ZN(new_n885));
  XOR2_X1   g699(.A(new_n728), .B(KEYINPUT121), .Z(new_n886));
  NAND3_X1  g700(.A1(new_n885), .A2(G902), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n876), .B1(new_n884), .B2(new_n887), .ZN(G54));
  AND2_X1   g702(.A1(KEYINPUT58), .A2(G475), .ZN(new_n889));
  OAI211_X1 g703(.A(G902), .B(new_n889), .C1(new_n863), .C2(new_n864), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n876), .B1(new_n890), .B2(new_n436), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n885), .A2(G902), .A3(new_n442), .A4(new_n889), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT122), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n893), .B(new_n894), .ZN(G60));
  INV_X1    g709(.A(new_n575), .ZN(new_n896));
  XNOR2_X1  g710(.A(KEYINPUT123), .B(KEYINPUT59), .ZN(new_n897));
  NAND2_X1  g711(.A1(G478), .A2(G902), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n897), .B(new_n898), .ZN(new_n899));
  OAI211_X1 g713(.A(new_n896), .B(new_n899), .C1(new_n881), .C2(new_n882), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(new_n877), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n899), .B1(new_n814), .B2(new_n815), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n901), .B1(new_n902), .B2(new_n575), .ZN(G63));
  NAND2_X1  g717(.A1(G217), .A2(G902), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT60), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n904), .B(new_n905), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n885), .A2(new_n608), .A3(new_n906), .ZN(new_n907));
  AND2_X1   g721(.A1(new_n885), .A2(new_n906), .ZN(new_n908));
  OAI211_X1 g722(.A(new_n877), .B(new_n907), .C1(new_n908), .C2(new_n556), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT61), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n885), .A2(new_n906), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n912), .A2(new_n555), .A3(new_n554), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n913), .A2(KEYINPUT61), .A3(new_n877), .A4(new_n907), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n911), .A2(new_n914), .ZN(G66));
  NAND3_X1  g729(.A1(new_n489), .A2(G224), .A3(G953), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n916), .B1(new_n763), .B2(G953), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n860), .B1(G898), .B2(new_n377), .ZN(new_n918));
  XOR2_X1   g732(.A(new_n917), .B(new_n918), .Z(G69));
  NAND3_X1  g733(.A1(new_n756), .A2(new_n580), .A3(new_n757), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n622), .A2(new_n725), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n709), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n743), .A2(new_n922), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n923), .B1(new_n723), .B2(new_n735), .ZN(new_n924));
  AND3_X1   g738(.A1(new_n618), .A2(new_n643), .A3(new_n675), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n639), .A2(new_n925), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n926), .B(KEYINPUT62), .ZN(new_n927));
  INV_X1    g741(.A(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n924), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n929), .A2(new_n377), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n256), .A2(new_n257), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n427), .B1(new_n428), .B2(new_n426), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n931), .B(new_n932), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n930), .A2(KEYINPUT124), .A3(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT124), .ZN(new_n935));
  AOI21_X1  g749(.A(G953), .B1(new_n924), .B2(new_n928), .ZN(new_n936));
  INV_X1    g750(.A(new_n933), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n935), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(new_n734), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n939), .A2(new_n665), .A3(new_n847), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n925), .A2(new_n713), .A3(new_n743), .A4(new_n940), .ZN(new_n941));
  AOI211_X1 g755(.A(new_n711), .B(new_n941), .C1(new_n723), .C2(new_n735), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n942), .A2(new_n377), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n933), .B1(G900), .B2(G953), .ZN(new_n944));
  AOI22_X1  g758(.A1(new_n934), .A2(new_n938), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT125), .ZN(new_n946));
  INV_X1    g760(.A(G900), .ZN(new_n947));
  OAI21_X1  g761(.A(G953), .B1(new_n334), .B2(new_n947), .ZN(new_n948));
  AND3_X1   g762(.A1(new_n945), .A2(new_n946), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n946), .B1(new_n945), .B2(new_n948), .ZN(new_n950));
  OAI22_X1  g764(.A1(new_n949), .A2(new_n950), .B1(new_n948), .B2(new_n945), .ZN(G72));
  INV_X1    g765(.A(new_n287), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n942), .A2(new_n254), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n287), .A2(new_n255), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n953), .B1(new_n929), .B2(new_n954), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n955), .A2(new_n749), .A3(new_n782), .ZN(new_n956));
  XOR2_X1   g770(.A(KEYINPUT126), .B(KEYINPUT63), .Z(new_n957));
  NOR2_X1   g771(.A1(new_n280), .A2(new_n281), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n957), .B(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n287), .B(new_n254), .ZN(new_n961));
  OAI211_X1 g775(.A(new_n956), .B(new_n877), .C1(new_n960), .C2(new_n961), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n800), .A2(new_n805), .A3(new_n960), .A4(new_n961), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n963), .A2(KEYINPUT127), .ZN(new_n964));
  OR2_X1    g778(.A1(new_n963), .A2(KEYINPUT127), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n962), .B1(new_n964), .B2(new_n965), .ZN(G57));
endmodule


