//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 0 0 0 1 0 1 0 1 0 0 0 0 1 1 0 1 1 0 0 0 1 1 0 1 1 0 0 1 1 0 0 0 1 0 0 1 1 0 0 1 0 1 1 1 0 1 1 1 1 0 0 1 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:18 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n566, new_n567, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n582, new_n583, new_n584, new_n585, new_n586, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n612, new_n613,
    new_n614, new_n615, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n635, new_n636, new_n639,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n851, new_n852, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1228;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT65), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  NOR2_X1   g027(.A1(new_n451), .A2(new_n452), .ZN(G325));
  INV_X1    g028(.A(G325), .ZN(G261));
  NAND2_X1  g029(.A1(new_n451), .A2(G2106), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n452), .A2(G567), .ZN(new_n456));
  XOR2_X1   g031(.A(new_n456), .B(KEYINPUT66), .Z(new_n457));
  NAND2_X1  g032(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  NAND2_X1  g034(.A1(G101), .A2(G2104), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT67), .ZN(new_n461));
  AND3_X1   g036(.A1(new_n461), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n462));
  AOI21_X1  g037(.A(KEYINPUT3), .B1(new_n461), .B2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G137), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n460), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  XNOR2_X1  g043(.A(KEYINPUT3), .B(G2104), .ZN(new_n469));
  AOI22_X1  g044(.A1(new_n469), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n470));
  OR2_X1    g045(.A1(new_n470), .A2(new_n467), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(G160));
  INV_X1    g048(.A(KEYINPUT3), .ZN(new_n474));
  INV_X1    g049(.A(G2104), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n474), .B1(new_n475), .B2(KEYINPUT67), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n461), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(new_n467), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n478), .A2(G2105), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  OR2_X1    g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G112), .C2(new_n467), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n481), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  INV_X1    g063(.A(G138), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n489), .A2(G2105), .ZN(new_n490));
  AOI21_X1  g065(.A(KEYINPUT4), .B1(new_n469), .B2(new_n490), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n467), .A2(KEYINPUT4), .A3(G138), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n492), .B1(new_n476), .B2(new_n477), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(G126), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n495), .B1(new_n476), .B2(new_n477), .ZN(new_n496));
  AND2_X1   g071(.A1(G114), .A2(G2104), .ZN(new_n497));
  OAI21_X1  g072(.A(G2105), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n475), .A2(G2105), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(G102), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n494), .A2(new_n498), .A3(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(G164));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  XOR2_X1   g078(.A(KEYINPUT68), .B(G651), .Z(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(KEYINPUT6), .ZN(new_n505));
  OR2_X1    g080(.A1(KEYINPUT6), .A2(G651), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n503), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G50), .ZN(new_n508));
  INV_X1    g083(.A(G88), .ZN(new_n509));
  AND2_X1   g084(.A1(KEYINPUT69), .A2(G543), .ZN(new_n510));
  NOR2_X1   g085(.A1(KEYINPUT69), .A2(G543), .ZN(new_n511));
  OAI21_X1  g086(.A(KEYINPUT5), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT5), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n512), .A2(KEYINPUT70), .B1(new_n513), .B2(G543), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT70), .ZN(new_n515));
  OAI211_X1 g090(.A(new_n515), .B(KEYINPUT5), .C1(new_n510), .C2(new_n511), .ZN(new_n516));
  XNOR2_X1  g091(.A(KEYINPUT68), .B(G651), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT6), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n506), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n514), .A2(new_n516), .A3(new_n519), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n508), .B1(new_n509), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n514), .A2(G62), .A3(new_n516), .ZN(new_n522));
  NAND2_X1  g097(.A1(G75), .A2(G543), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n517), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n521), .A2(new_n524), .ZN(G166));
  NAND2_X1  g100(.A1(new_n512), .A2(KEYINPUT70), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n513), .A2(G543), .ZN(new_n527));
  AND2_X1   g102(.A1(G63), .A2(G651), .ZN(new_n528));
  NAND4_X1  g103(.A1(new_n526), .A2(new_n516), .A3(new_n527), .A4(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT71), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND4_X1  g106(.A1(new_n514), .A2(KEYINPUT71), .A3(new_n516), .A4(new_n528), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n535));
  XOR2_X1   g110(.A(new_n535), .B(KEYINPUT7), .Z(new_n536));
  INV_X1    g111(.A(new_n536), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n519), .A2(G51), .A3(G543), .ZN(new_n538));
  INV_X1    g113(.A(G89), .ZN(new_n539));
  OAI211_X1 g114(.A(new_n537), .B(new_n538), .C1(new_n520), .C2(new_n539), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n534), .A2(new_n540), .ZN(G168));
  NAND3_X1  g116(.A1(new_n514), .A2(G64), .A3(new_n516), .ZN(new_n542));
  NAND2_X1  g117(.A1(G77), .A2(G543), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n517), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND4_X1  g119(.A1(new_n514), .A2(G90), .A3(new_n516), .A4(new_n519), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n519), .A2(G52), .A3(G543), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n544), .A2(new_n547), .ZN(G171));
  NAND4_X1  g123(.A1(new_n514), .A2(G81), .A3(new_n516), .A4(new_n519), .ZN(new_n549));
  XNOR2_X1  g124(.A(KEYINPUT72), .B(G43), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n519), .A2(G543), .A3(new_n550), .ZN(new_n551));
  AND2_X1   g126(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  NAND4_X1  g127(.A1(new_n526), .A2(G56), .A3(new_n516), .A4(new_n527), .ZN(new_n553));
  NAND2_X1  g128(.A1(G68), .A2(G543), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(new_n504), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n552), .A2(new_n556), .A3(KEYINPUT73), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT73), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n549), .A2(new_n551), .ZN(new_n559));
  AOI21_X1  g134(.A(new_n517), .B1(new_n553), .B2(new_n554), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n557), .A2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G860), .ZN(G153));
  NAND4_X1  g139(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g140(.A1(G1), .A2(G3), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT8), .ZN(new_n567));
  NAND4_X1  g142(.A1(G319), .A2(G483), .A3(G661), .A4(new_n567), .ZN(G188));
  NAND3_X1  g143(.A1(new_n514), .A2(G65), .A3(new_n516), .ZN(new_n569));
  NAND2_X1  g144(.A1(G78), .A2(G543), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n519), .A2(G53), .A3(G543), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n572), .A2(KEYINPUT74), .A3(KEYINPUT9), .ZN(new_n573));
  NAND2_X1  g148(.A1(KEYINPUT74), .A2(KEYINPUT9), .ZN(new_n574));
  NAND4_X1  g149(.A1(new_n519), .A2(G53), .A3(G543), .A4(new_n574), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n571), .A2(G651), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT75), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n520), .A2(new_n577), .ZN(new_n578));
  NAND4_X1  g153(.A1(new_n514), .A2(KEYINPUT75), .A3(new_n516), .A4(new_n519), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n578), .A2(G91), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n576), .A2(new_n580), .ZN(G299));
  INV_X1    g156(.A(new_n544), .ZN(new_n582));
  INV_X1    g157(.A(new_n547), .ZN(new_n583));
  AOI21_X1  g158(.A(KEYINPUT76), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT76), .ZN(new_n585));
  NOR3_X1   g160(.A1(new_n544), .A2(new_n547), .A3(new_n585), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n584), .A2(new_n586), .ZN(G301));
  OAI21_X1  g162(.A(KEYINPUT77), .B1(new_n534), .B2(new_n540), .ZN(new_n588));
  INV_X1    g163(.A(new_n520), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n589), .A2(G89), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT77), .ZN(new_n591));
  AND2_X1   g166(.A1(new_n538), .A2(new_n537), .ZN(new_n592));
  NAND4_X1  g167(.A1(new_n590), .A2(new_n533), .A3(new_n591), .A4(new_n592), .ZN(new_n593));
  AND2_X1   g168(.A1(new_n588), .A2(new_n593), .ZN(G286));
  INV_X1    g169(.A(G166), .ZN(G303));
  NAND2_X1  g170(.A1(new_n514), .A2(new_n516), .ZN(new_n596));
  INV_X1    g171(.A(G74), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n519), .A2(G49), .A3(G543), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT78), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND4_X1  g176(.A1(new_n519), .A2(KEYINPUT78), .A3(G49), .A4(G543), .ZN(new_n602));
  AOI22_X1  g177(.A1(G651), .A2(new_n598), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n578), .A2(G87), .A3(new_n579), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(G288));
  NAND2_X1  g180(.A1(G73), .A2(G543), .ZN(new_n606));
  INV_X1    g181(.A(G61), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n596), .B2(new_n607), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n608), .A2(new_n504), .B1(G48), .B2(new_n507), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n578), .A2(G86), .A3(new_n579), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n609), .A2(new_n610), .ZN(G305));
  XOR2_X1   g186(.A(KEYINPUT79), .B(G47), .Z(new_n612));
  AOI22_X1  g187(.A1(new_n589), .A2(G85), .B1(new_n507), .B2(new_n612), .ZN(new_n613));
  AND2_X1   g188(.A1(new_n514), .A2(new_n516), .ZN(new_n614));
  AOI22_X1  g189(.A1(new_n614), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n613), .B1(new_n517), .B2(new_n615), .ZN(G290));
  INV_X1    g191(.A(G868), .ZN(new_n617));
  NOR2_X1   g192(.A1(G301), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g193(.A(KEYINPUT81), .B(G66), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n514), .A2(new_n516), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(G79), .A2(G543), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(KEYINPUT80), .Z(new_n622));
  NAND2_X1  g197(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n623), .A2(G651), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n507), .A2(G54), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n578), .A2(G92), .A3(new_n579), .ZN(new_n627));
  INV_X1    g202(.A(KEYINPUT10), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND4_X1  g204(.A1(new_n578), .A2(KEYINPUT10), .A3(G92), .A4(new_n579), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n626), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT82), .ZN(new_n632));
  AOI21_X1  g207(.A(new_n618), .B1(new_n632), .B2(new_n617), .ZN(G284));
  AOI21_X1  g208(.A(new_n618), .B1(new_n632), .B2(new_n617), .ZN(G321));
  NOR2_X1   g209(.A1(G286), .A2(new_n617), .ZN(new_n635));
  XNOR2_X1  g210(.A(G299), .B(KEYINPUT83), .ZN(new_n636));
  AOI21_X1  g211(.A(new_n635), .B1(new_n617), .B2(new_n636), .ZN(G297));
  AOI21_X1  g212(.A(new_n635), .B1(new_n617), .B2(new_n636), .ZN(G280));
  INV_X1    g213(.A(G559), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n632), .B1(new_n639), .B2(G860), .ZN(G148));
  INV_X1    g215(.A(KEYINPUT82), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n631), .B(new_n641), .ZN(new_n642));
  OR3_X1    g217(.A1(new_n642), .A2(KEYINPUT84), .A3(G559), .ZN(new_n643));
  OAI21_X1  g218(.A(KEYINPUT84), .B1(new_n642), .B2(G559), .ZN(new_n644));
  AOI21_X1  g219(.A(new_n617), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n645), .A2(KEYINPUT85), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n645), .A2(KEYINPUT85), .ZN(new_n647));
  OAI211_X1 g222(.A(new_n646), .B(new_n647), .C1(G868), .C2(new_n563), .ZN(G323));
  XNOR2_X1  g223(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g224(.A1(new_n469), .A2(new_n499), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT12), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT13), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(G2100), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n480), .A2(G135), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n483), .A2(G123), .ZN(new_n655));
  NOR2_X1   g230(.A1(G99), .A2(G2105), .ZN(new_n656));
  OAI21_X1  g231(.A(G2104), .B1(new_n467), .B2(G111), .ZN(new_n657));
  OAI211_X1 g232(.A(new_n654), .B(new_n655), .C1(new_n656), .C2(new_n657), .ZN(new_n658));
  INV_X1    g233(.A(G2096), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n653), .A2(new_n660), .ZN(G156));
  XNOR2_X1  g236(.A(G2451), .B(G2454), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT16), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n663), .B(KEYINPUT86), .Z(new_n664));
  INV_X1    g239(.A(KEYINPUT14), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2427), .B(G2438), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(G2430), .ZN(new_n667));
  XNOR2_X1  g242(.A(KEYINPUT15), .B(G2435), .ZN(new_n668));
  AOI21_X1  g243(.A(new_n665), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  OAI21_X1  g244(.A(new_n669), .B1(new_n668), .B2(new_n667), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n664), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1341), .B(G1348), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT87), .ZN(new_n673));
  XNOR2_X1  g248(.A(G2443), .B(G2446), .ZN(new_n674));
  XOR2_X1   g249(.A(new_n673), .B(new_n674), .Z(new_n675));
  OR2_X1    g250(.A1(new_n671), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n671), .A2(new_n675), .ZN(new_n677));
  AND3_X1   g252(.A1(new_n676), .A2(G14), .A3(new_n677), .ZN(G401));
  XOR2_X1   g253(.A(G2072), .B(G2078), .Z(new_n679));
  XOR2_X1   g254(.A(new_n679), .B(KEYINPUT17), .Z(new_n680));
  XOR2_X1   g255(.A(G2084), .B(G2090), .Z(new_n681));
  XNOR2_X1  g256(.A(G2067), .B(G2678), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n680), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n681), .A2(new_n682), .ZN(new_n684));
  INV_X1    g259(.A(new_n681), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n685), .A2(new_n679), .ZN(new_n686));
  OAI211_X1 g261(.A(new_n683), .B(new_n684), .C1(new_n682), .C2(new_n686), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n684), .A2(new_n679), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT18), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(new_n659), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(G2100), .ZN(G227));
  XNOR2_X1  g267(.A(G1971), .B(G1976), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT19), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1956), .B(G2474), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1961), .B(G1966), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n694), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n695), .A2(new_n696), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n694), .A2(KEYINPUT89), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n700), .B(new_n701), .Z(new_n702));
  NOR3_X1   g277(.A1(new_n694), .A2(new_n695), .A3(new_n696), .ZN(new_n703));
  XNOR2_X1  g278(.A(KEYINPUT88), .B(KEYINPUT20), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n702), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(G1986), .ZN(new_n707));
  XOR2_X1   g282(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(G1991), .B(G1996), .ZN(new_n710));
  INV_X1    g285(.A(G1981), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n709), .B(new_n712), .ZN(G229));
  NOR2_X1   g288(.A1(G4), .A2(G16), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n714), .B1(new_n632), .B2(G16), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(G1348), .ZN(new_n716));
  XNOR2_X1  g291(.A(KEYINPUT31), .B(G11), .ZN(new_n717));
  XOR2_X1   g292(.A(KEYINPUT96), .B(G28), .Z(new_n718));
  NOR2_X1   g293(.A1(new_n718), .A2(KEYINPUT30), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n718), .A2(KEYINPUT30), .ZN(new_n720));
  INV_X1    g295(.A(G29), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  OAI221_X1 g297(.A(new_n717), .B1(new_n719), .B2(new_n722), .C1(new_n658), .C2(new_n721), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT97), .ZN(new_n724));
  INV_X1    g299(.A(G16), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n725), .A2(G21), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G168), .B2(new_n725), .ZN(new_n727));
  XNOR2_X1  g302(.A(KEYINPUT95), .B(G1966), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n727), .B(new_n728), .Z(new_n729));
  NAND2_X1  g304(.A1(new_n725), .A2(G5), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(G171), .B2(new_n725), .ZN(new_n731));
  AOI211_X1 g306(.A(new_n724), .B(new_n729), .C1(G1961), .C2(new_n731), .ZN(new_n732));
  OR2_X1    g307(.A1(new_n732), .A2(KEYINPUT98), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n721), .A2(G32), .ZN(new_n734));
  NAND3_X1  g309(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n735));
  INV_X1    g310(.A(KEYINPUT26), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND4_X1  g312(.A1(KEYINPUT26), .A2(G117), .A3(G2104), .A4(G2105), .ZN(new_n738));
  AOI22_X1  g313(.A1(new_n737), .A2(new_n738), .B1(new_n499), .B2(G105), .ZN(new_n739));
  INV_X1    g314(.A(G141), .ZN(new_n740));
  INV_X1    g315(.A(G129), .ZN(new_n741));
  OAI221_X1 g316(.A(new_n739), .B1(new_n479), .B2(new_n740), .C1(new_n741), .C2(new_n482), .ZN(new_n742));
  INV_X1    g317(.A(KEYINPUT94), .ZN(new_n743));
  OR2_X1    g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n742), .A2(new_n743), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(new_n746), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n734), .B1(new_n747), .B2(new_n721), .ZN(new_n748));
  XNOR2_X1  g323(.A(KEYINPUT27), .B(G1996), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  NOR2_X1   g325(.A1(G164), .A2(new_n721), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(G27), .B2(new_n721), .ZN(new_n752));
  INV_X1    g327(.A(G2078), .ZN(new_n753));
  AND2_X1   g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n752), .A2(new_n753), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n721), .A2(G26), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(KEYINPUT28), .Z(new_n757));
  NAND2_X1  g332(.A1(new_n480), .A2(G140), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n483), .A2(G128), .ZN(new_n759));
  OR2_X1    g334(.A1(G104), .A2(G2105), .ZN(new_n760));
  OAI211_X1 g335(.A(new_n760), .B(G2104), .C1(G116), .C2(new_n467), .ZN(new_n761));
  NAND3_X1  g336(.A1(new_n758), .A2(new_n759), .A3(new_n761), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n757), .B1(new_n762), .B2(G29), .ZN(new_n763));
  INV_X1    g338(.A(G2067), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  NOR3_X1   g340(.A1(new_n754), .A2(new_n755), .A3(new_n765), .ZN(new_n766));
  OAI211_X1 g341(.A(new_n750), .B(new_n766), .C1(G1961), .C2(new_n731), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n563), .A2(new_n725), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(new_n725), .B2(G19), .ZN(new_n769));
  INV_X1    g344(.A(new_n769), .ZN(new_n770));
  AND2_X1   g345(.A1(new_n770), .A2(G1341), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n770), .A2(G1341), .ZN(new_n772));
  NOR3_X1   g347(.A1(new_n767), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n732), .A2(KEYINPUT98), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n721), .A2(G33), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n467), .A2(G103), .A3(G2104), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT25), .Z(new_n777));
  INV_X1    g352(.A(G139), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n777), .B1(new_n479), .B2(new_n778), .ZN(new_n779));
  INV_X1    g354(.A(KEYINPUT93), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  AOI22_X1  g356(.A1(new_n469), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n782));
  OR2_X1    g357(.A1(new_n782), .A2(new_n467), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  INV_X1    g359(.A(new_n784), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n775), .B1(new_n785), .B2(new_n721), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n786), .A2(G2072), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n721), .A2(G35), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G162), .B2(new_n721), .ZN(new_n789));
  XNOR2_X1  g364(.A(KEYINPUT99), .B(KEYINPUT29), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(G2090), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n789), .B(new_n791), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n721), .B1(KEYINPUT24), .B2(G34), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(KEYINPUT24), .B2(G34), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(new_n472), .B2(G29), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(G2084), .ZN(new_n796));
  NAND3_X1  g371(.A1(new_n787), .A2(new_n792), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n725), .A2(G20), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT23), .ZN(new_n799));
  INV_X1    g374(.A(G299), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n799), .B1(new_n800), .B2(new_n725), .ZN(new_n801));
  XNOR2_X1  g376(.A(KEYINPUT100), .B(G1956), .ZN(new_n802));
  INV_X1    g377(.A(new_n802), .ZN(new_n803));
  AND2_X1   g378(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n801), .A2(new_n803), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n786), .A2(G2072), .ZN(new_n806));
  NOR4_X1   g381(.A1(new_n797), .A2(new_n804), .A3(new_n805), .A4(new_n806), .ZN(new_n807));
  NAND4_X1  g382(.A1(new_n733), .A2(new_n773), .A3(new_n774), .A4(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n725), .A2(G22), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(G166), .B2(new_n725), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n810), .A2(G1971), .ZN(new_n811));
  AND2_X1   g386(.A1(new_n810), .A2(G1971), .ZN(new_n812));
  XOR2_X1   g387(.A(KEYINPUT33), .B(G1976), .Z(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT91), .ZN(new_n814));
  INV_X1    g389(.A(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n725), .A2(G23), .ZN(new_n816));
  INV_X1    g391(.A(G288), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n816), .B1(new_n817), .B2(new_n725), .ZN(new_n818));
  AOI211_X1 g393(.A(new_n811), .B(new_n812), .C1(new_n815), .C2(new_n818), .ZN(new_n819));
  MUX2_X1   g394(.A(G6), .B(G305), .S(G16), .Z(new_n820));
  XOR2_X1   g395(.A(KEYINPUT32), .B(G1981), .Z(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  OR2_X1    g397(.A1(new_n818), .A2(new_n815), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n819), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT92), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND4_X1  g401(.A1(new_n819), .A2(KEYINPUT92), .A3(new_n822), .A4(new_n823), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT34), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n826), .A2(KEYINPUT34), .A3(new_n827), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n721), .A2(G25), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n480), .A2(G131), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n483), .A2(G119), .ZN(new_n834));
  OR2_X1    g409(.A1(G95), .A2(G2105), .ZN(new_n835));
  OAI211_X1 g410(.A(new_n835), .B(G2104), .C1(G107), .C2(new_n467), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n833), .A2(new_n834), .A3(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(new_n837), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n832), .B1(new_n838), .B2(new_n721), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT90), .ZN(new_n840));
  XOR2_X1   g415(.A(KEYINPUT35), .B(G1991), .Z(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  MUX2_X1   g417(.A(G24), .B(G290), .S(G16), .Z(new_n843));
  OAI21_X1  g418(.A(new_n842), .B1(G1986), .B2(new_n843), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n844), .B1(G1986), .B2(new_n843), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n830), .A2(new_n831), .A3(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n846), .A2(KEYINPUT36), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT36), .ZN(new_n848));
  NAND4_X1  g423(.A1(new_n830), .A2(new_n848), .A3(new_n831), .A4(new_n845), .ZN(new_n849));
  AOI211_X1 g424(.A(new_n716), .B(new_n808), .C1(new_n847), .C2(new_n849), .ZN(G311));
  NAND2_X1  g425(.A1(new_n847), .A2(new_n849), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n808), .A2(new_n716), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(G150));
  XOR2_X1   g428(.A(KEYINPUT103), .B(G55), .Z(new_n854));
  NAND2_X1  g429(.A1(new_n507), .A2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(G93), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n855), .B1(new_n856), .B2(new_n520), .ZN(new_n857));
  NAND4_X1  g432(.A1(new_n526), .A2(G67), .A3(new_n516), .A4(new_n527), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT102), .ZN(new_n859));
  NAND2_X1  g434(.A1(G80), .A2(G543), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n858), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n858), .A2(new_n860), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n517), .B1(new_n862), .B2(KEYINPUT102), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n857), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(G860), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(KEYINPUT37), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n632), .A2(G559), .ZN(new_n868));
  XOR2_X1   g443(.A(KEYINPUT101), .B(KEYINPUT38), .Z(new_n869));
  XNOR2_X1  g444(.A(new_n868), .B(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n862), .A2(KEYINPUT102), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n871), .A2(new_n861), .A3(new_n504), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n552), .A2(new_n556), .ZN(new_n873));
  AOI22_X1  g448(.A1(new_n589), .A2(G93), .B1(new_n507), .B2(new_n854), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n875), .B1(new_n562), .B2(new_n864), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n876), .A2(KEYINPUT104), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT104), .ZN(new_n878));
  OAI211_X1 g453(.A(new_n875), .B(new_n878), .C1(new_n562), .C2(new_n864), .ZN(new_n879));
  AND2_X1   g454(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n870), .B(new_n880), .ZN(new_n881));
  AND2_X1   g456(.A1(new_n881), .A2(KEYINPUT39), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n865), .B1(new_n881), .B2(KEYINPUT39), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n867), .B1(new_n882), .B2(new_n883), .ZN(G145));
  OR3_X1    g459(.A1(new_n467), .A2(KEYINPUT107), .A3(G118), .ZN(new_n885));
  OAI21_X1  g460(.A(KEYINPUT107), .B1(new_n467), .B2(G118), .ZN(new_n886));
  OR2_X1    g461(.A1(G106), .A2(G2105), .ZN(new_n887));
  NAND4_X1  g462(.A1(new_n885), .A2(G2104), .A3(new_n886), .A4(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(G142), .ZN(new_n889));
  INV_X1    g464(.A(G130), .ZN(new_n890));
  OAI221_X1 g465(.A(new_n888), .B1(new_n479), .B2(new_n889), .C1(new_n890), .C2(new_n482), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(new_n651), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(new_n838), .ZN(new_n893));
  OAI21_X1  g468(.A(KEYINPUT105), .B1(new_n491), .B2(new_n493), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n475), .A2(KEYINPUT3), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n474), .A2(G2104), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n490), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT4), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  AND3_X1   g474(.A1(new_n467), .A2(KEYINPUT4), .A3(G138), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n900), .B1(new_n462), .B2(new_n463), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT105), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n899), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  NAND4_X1  g478(.A1(new_n894), .A2(new_n903), .A3(new_n498), .A4(new_n500), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n762), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n744), .A2(new_n745), .A3(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n906), .B1(new_n744), .B2(new_n745), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n905), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n909), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n911), .A2(new_n904), .A3(new_n907), .ZN(new_n912));
  OR2_X1    g487(.A1(new_n784), .A2(KEYINPUT106), .ZN(new_n913));
  AND3_X1   g488(.A1(new_n910), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n784), .A2(KEYINPUT106), .ZN(new_n915));
  AOI22_X1  g490(.A1(new_n910), .A2(new_n912), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  OAI211_X1 g491(.A(KEYINPUT108), .B(new_n893), .C1(new_n914), .C2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n910), .A2(new_n912), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n913), .A2(new_n915), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  OR2_X1    g495(.A1(new_n893), .A2(KEYINPUT108), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n893), .A2(KEYINPUT108), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n910), .A2(new_n912), .A3(new_n913), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n920), .A2(new_n921), .A3(new_n922), .A4(new_n923), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n658), .B(new_n472), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n925), .B(new_n487), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n917), .A2(new_n924), .A3(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(G37), .ZN(new_n928));
  AND2_X1   g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n926), .B1(new_n917), .B2(new_n924), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n930), .A2(KEYINPUT109), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT109), .ZN(new_n932));
  AOI211_X1 g507(.A(new_n932), .B(new_n926), .C1(new_n917), .C2(new_n924), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n929), .B1(new_n931), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(KEYINPUT110), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT110), .ZN(new_n936));
  OAI211_X1 g511(.A(new_n929), .B(new_n936), .C1(new_n931), .C2(new_n933), .ZN(new_n937));
  AND3_X1   g512(.A1(new_n935), .A2(KEYINPUT40), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(KEYINPUT40), .B1(new_n935), .B2(new_n937), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n938), .A2(new_n939), .ZN(G395));
  NAND2_X1  g515(.A1(new_n643), .A2(new_n644), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(new_n880), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n877), .A2(new_n879), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n643), .A2(new_n644), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n629), .A2(new_n630), .ZN(new_n946));
  INV_X1    g521(.A(new_n626), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(new_n800), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n631), .A2(G299), .ZN(new_n950));
  AND2_X1   g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n945), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n948), .A2(KEYINPUT111), .A3(new_n800), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT111), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n955), .B1(new_n631), .B2(G299), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n954), .A2(new_n950), .A3(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT41), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n958), .B1(new_n631), .B2(G299), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n949), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n942), .A2(new_n944), .A3(new_n962), .ZN(new_n963));
  XNOR2_X1  g538(.A(new_n817), .B(G305), .ZN(new_n964));
  XNOR2_X1  g539(.A(G290), .B(G166), .ZN(new_n965));
  XNOR2_X1  g540(.A(new_n964), .B(new_n965), .ZN(new_n966));
  XNOR2_X1  g541(.A(new_n966), .B(KEYINPUT42), .ZN(new_n967));
  AND3_X1   g542(.A1(new_n953), .A2(new_n963), .A3(new_n967), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n967), .B1(new_n953), .B2(new_n963), .ZN(new_n969));
  OAI21_X1  g544(.A(G868), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n970), .B1(G868), .B2(new_n864), .ZN(G295));
  OAI21_X1  g546(.A(new_n970), .B1(G868), .B2(new_n864), .ZN(G331));
  NAND3_X1  g547(.A1(new_n588), .A2(G171), .A3(new_n593), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT112), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(G301), .A2(G168), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n588), .A2(KEYINPUT112), .A3(G171), .A4(new_n593), .ZN(new_n977));
  AND3_X1   g552(.A1(new_n975), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n951), .B1(new_n880), .B2(new_n978), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n975), .A2(new_n976), .A3(new_n977), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n943), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(KEYINPUT113), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT113), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n943), .A2(new_n980), .A3(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n979), .A2(new_n982), .A3(new_n984), .ZN(new_n985));
  AOI22_X1  g560(.A1(new_n974), .A2(new_n973), .B1(G301), .B2(G168), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n986), .A2(new_n877), .A3(new_n879), .A4(new_n977), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n981), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n962), .A2(new_n988), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n985), .A2(new_n989), .A3(new_n966), .ZN(new_n990));
  AND2_X1   g565(.A1(new_n990), .A2(new_n928), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n979), .A2(new_n981), .ZN(new_n992));
  AND3_X1   g567(.A1(new_n943), .A2(new_n983), .A3(new_n980), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n983), .B1(new_n943), .B2(new_n980), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n943), .A2(new_n980), .ZN(new_n995));
  NOR3_X1   g570(.A1(new_n993), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  AND2_X1   g571(.A1(new_n954), .A2(new_n956), .ZN(new_n997));
  AOI22_X1  g572(.A1(new_n952), .A2(new_n958), .B1(new_n997), .B2(new_n960), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n992), .B1(new_n996), .B2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(new_n966), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n991), .A2(new_n1001), .A3(KEYINPUT114), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT114), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n982), .A2(new_n987), .A3(new_n984), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n997), .A2(new_n960), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1005), .B1(KEYINPUT41), .B2(new_n951), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n966), .B1(new_n1007), .B2(new_n992), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n990), .A2(new_n928), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1003), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1002), .A2(new_n1010), .A3(KEYINPUT43), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n985), .A2(new_n989), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(new_n1000), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT43), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n1013), .A2(new_n1014), .A3(new_n928), .A4(new_n990), .ZN(new_n1015));
  AND2_X1   g590(.A1(new_n1015), .A2(KEYINPUT44), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1011), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT44), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1014), .B1(new_n991), .B2(new_n1013), .ZN(new_n1019));
  NOR3_X1   g594(.A1(new_n1008), .A2(new_n1009), .A3(KEYINPUT43), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1018), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1017), .A2(new_n1021), .ZN(G397));
  XOR2_X1   g597(.A(KEYINPUT115), .B(G1384), .Z(new_n1023));
  AOI21_X1  g598(.A(KEYINPUT116), .B1(new_n904), .B2(new_n1023), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1024), .A2(KEYINPUT45), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n904), .A2(KEYINPUT116), .A3(new_n1023), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n468), .A2(new_n471), .A3(G40), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1029), .ZN(new_n1030));
  XNOR2_X1  g605(.A(new_n762), .B(G2067), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1031), .B1(new_n746), .B2(G1996), .ZN(new_n1032));
  INV_X1    g607(.A(G1996), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n747), .A2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1030), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1035));
  XNOR2_X1  g610(.A(new_n1035), .B(KEYINPUT117), .ZN(new_n1036));
  XOR2_X1   g611(.A(new_n837), .B(new_n841), .Z(new_n1037));
  AOI21_X1  g612(.A(new_n1036), .B1(new_n1029), .B2(new_n1037), .ZN(new_n1038));
  NOR3_X1   g613(.A1(new_n1030), .A2(G1986), .A3(G290), .ZN(new_n1039));
  XOR2_X1   g614(.A(new_n1039), .B(KEYINPUT48), .Z(new_n1040));
  NAND2_X1  g615(.A1(new_n906), .A2(new_n764), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n838), .A2(new_n841), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1041), .B1(new_n1036), .B2(new_n1042), .ZN(new_n1043));
  AOI22_X1  g618(.A1(new_n1038), .A2(new_n1040), .B1(new_n1043), .B2(new_n1029), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1029), .B1(new_n746), .B2(new_n1031), .ZN(new_n1045));
  XOR2_X1   g620(.A(new_n1045), .B(KEYINPUT126), .Z(new_n1046));
  NAND2_X1  g621(.A1(new_n1029), .A2(new_n1033), .ZN(new_n1047));
  XOR2_X1   g622(.A(new_n1047), .B(KEYINPUT46), .Z(new_n1048));
  OR3_X1    g623(.A1(new_n1046), .A2(new_n1048), .A3(KEYINPUT127), .ZN(new_n1049));
  OAI21_X1  g624(.A(KEYINPUT127), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1049), .A2(KEYINPUT47), .A3(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1044), .A2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g627(.A(KEYINPUT47), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(G8), .ZN(new_n1055));
  INV_X1    g630(.A(G1384), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n501), .A2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1028), .B1(new_n1057), .B2(KEYINPUT50), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT50), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n904), .A2(new_n1059), .A3(new_n1056), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1061), .A2(G2090), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT45), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1057), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1028), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n904), .A2(KEYINPUT45), .A3(new_n1023), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1065), .A2(new_n1066), .A3(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(G1971), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1055), .B1(new_n1063), .B2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g646(.A(G8), .B1(new_n521), .B2(new_n524), .ZN(new_n1072));
  XNOR2_X1  g647(.A(new_n1072), .B(KEYINPUT55), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1071), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(G1976), .ZN(new_n1076));
  AOI21_X1  g651(.A(KEYINPUT52), .B1(G288), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n904), .A2(new_n1056), .ZN(new_n1078));
  OAI21_X1  g653(.A(G8), .B1(new_n1078), .B2(new_n1028), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1079), .ZN(new_n1080));
  OAI211_X1 g655(.A(new_n1077), .B(new_n1080), .C1(new_n1076), .C2(G288), .ZN(new_n1081));
  NOR2_X1   g656(.A1(G288), .A2(new_n1076), .ZN(new_n1082));
  OAI21_X1  g657(.A(KEYINPUT52), .B1(new_n1082), .B2(new_n1079), .ZN(new_n1083));
  AND2_X1   g658(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n589), .A2(G86), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n711), .B1(new_n609), .B2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n609), .A2(new_n711), .A3(new_n610), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT118), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n609), .A2(KEYINPUT118), .A3(new_n711), .A4(new_n610), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1086), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  AND2_X1   g666(.A1(new_n1091), .A2(KEYINPUT49), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1080), .B1(new_n1091), .B2(KEYINPUT49), .ZN(new_n1093));
  OAI211_X1 g668(.A(new_n1075), .B(new_n1084), .C1(new_n1092), .C2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1028), .B1(new_n1078), .B2(KEYINPUT50), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n501), .A2(new_n1059), .A3(new_n1056), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1070), .B1(new_n1097), .B2(G2090), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1074), .B1(G8), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(G2084), .ZN(new_n1100));
  AND3_X1   g675(.A1(new_n1058), .A2(new_n1100), .A3(new_n1060), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT120), .ZN(new_n1102));
  NOR3_X1   g677(.A1(new_n491), .A2(KEYINPUT105), .A3(new_n493), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n902), .B1(new_n899), .B2(new_n901), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  AND2_X1   g680(.A1(new_n498), .A2(new_n500), .ZN(new_n1106));
  AOI21_X1  g681(.A(G1384), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  OAI211_X1 g682(.A(new_n1102), .B(new_n1066), .C1(new_n1107), .C2(KEYINPUT45), .ZN(new_n1108));
  AOI21_X1  g683(.A(KEYINPUT45), .B1(new_n904), .B2(new_n1056), .ZN(new_n1109));
  OAI21_X1  g684(.A(KEYINPUT120), .B1(new_n1109), .B2(new_n1028), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n501), .A2(KEYINPUT45), .A3(new_n1056), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1108), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1101), .B1(new_n1112), .B2(new_n728), .ZN(new_n1113));
  OR3_X1    g688(.A1(new_n1113), .A2(new_n1055), .A3(G286), .ZN(new_n1114));
  NOR3_X1   g689(.A1(new_n1094), .A2(new_n1099), .A3(new_n1114), .ZN(new_n1115));
  OAI21_X1  g690(.A(KEYINPUT63), .B1(new_n1071), .B2(new_n1074), .ZN(new_n1116));
  OR2_X1    g691(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1117));
  OAI22_X1  g692(.A1(new_n1115), .A2(KEYINPUT63), .B1(new_n1094), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT119), .ZN(new_n1119));
  OAI211_X1 g694(.A(new_n1076), .B(new_n817), .C1(new_n1092), .C2(new_n1093), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(new_n1080), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1070), .ZN(new_n1124));
  OAI21_X1  g699(.A(G8), .B1(new_n1124), .B2(new_n1062), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1125), .A2(new_n1073), .ZN(new_n1126));
  OAI211_X1 g701(.A(new_n1126), .B(new_n1084), .C1(new_n1092), .C2(new_n1093), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1119), .B1(new_n1123), .B2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1079), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1127), .ZN(new_n1130));
  NOR3_X1   g705(.A1(new_n1129), .A2(KEYINPUT119), .A3(new_n1130), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1118), .B1(new_n1128), .B2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g707(.A(KEYINPUT51), .B1(new_n1113), .B2(G168), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1055), .B1(new_n1113), .B2(G168), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT124), .ZN(new_n1136));
  INV_X1    g711(.A(G168), .ZN(new_n1137));
  AOI211_X1 g712(.A(new_n1137), .B(new_n1101), .C1(new_n1112), .C2(new_n728), .ZN(new_n1138));
  OAI21_X1  g713(.A(KEYINPUT51), .B1(new_n1138), .B2(new_n1055), .ZN(new_n1139));
  AND3_X1   g714(.A1(new_n1135), .A2(new_n1136), .A3(new_n1139), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1136), .B1(new_n1135), .B2(new_n1139), .ZN(new_n1141));
  OAI21_X1  g716(.A(KEYINPUT62), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1135), .A2(new_n1139), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1143), .A2(KEYINPUT124), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT62), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1135), .A2(new_n1139), .A3(new_n1136), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1144), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(G1961), .ZN(new_n1148));
  AND3_X1   g723(.A1(new_n1058), .A2(KEYINPUT121), .A3(new_n1060), .ZN(new_n1149));
  AOI21_X1  g724(.A(KEYINPUT121), .B1(new_n1058), .B2(new_n1060), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1148), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT53), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1152), .B1(new_n1068), .B2(G2078), .ZN(new_n1153));
  AND2_X1   g728(.A1(new_n1151), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n753), .A2(KEYINPUT53), .ZN(new_n1155));
  OR2_X1    g730(.A1(new_n1112), .A2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g731(.A(G301), .B1(new_n1154), .B2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1142), .A2(new_n1147), .A3(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT57), .ZN(new_n1159));
  NAND2_X1  g734(.A1(G299), .A2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n576), .A2(KEYINPUT57), .A3(new_n580), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(G1956), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1097), .A2(new_n1163), .ZN(new_n1164));
  AND3_X1   g739(.A1(new_n1065), .A2(new_n1066), .A3(new_n1067), .ZN(new_n1165));
  XNOR2_X1  g740(.A(KEYINPUT56), .B(G2072), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1162), .A2(new_n1164), .A3(new_n1167), .ZN(new_n1168));
  AND3_X1   g743(.A1(new_n576), .A2(KEYINPUT57), .A3(new_n580), .ZN(new_n1169));
  AOI21_X1  g744(.A(KEYINPUT57), .B1(new_n576), .B2(new_n580), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  AOI21_X1  g746(.A(G1956), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1166), .ZN(new_n1173));
  NOR2_X1   g748(.A1(new_n1068), .A2(new_n1173), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1171), .B1(new_n1172), .B2(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT122), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1164), .A2(new_n1167), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1178), .A2(KEYINPUT122), .A3(new_n1171), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1177), .A2(new_n1179), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n1078), .A2(new_n1028), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1181), .A2(new_n764), .ZN(new_n1182));
  INV_X1    g757(.A(G1348), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1183), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n642), .B1(new_n1182), .B2(new_n1184), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1168), .B1(new_n1180), .B2(new_n1185), .ZN(new_n1186));
  INV_X1    g761(.A(KEYINPUT123), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1175), .A2(new_n1168), .A3(new_n1187), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT61), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1178), .A2(KEYINPUT123), .A3(new_n1171), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1188), .A2(new_n1189), .A3(new_n1190), .ZN(new_n1191));
  NAND4_X1  g766(.A1(new_n1177), .A2(new_n1179), .A3(KEYINPUT61), .A4(new_n1168), .ZN(new_n1192));
  XNOR2_X1  g767(.A(KEYINPUT58), .B(G1341), .ZN(new_n1193));
  OAI22_X1  g768(.A1(new_n1068), .A2(G1996), .B1(new_n1181), .B2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1194), .A2(new_n563), .ZN(new_n1195));
  XNOR2_X1  g770(.A(new_n1195), .B(KEYINPUT59), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1191), .A2(new_n1192), .A3(new_n1196), .ZN(new_n1197));
  NAND3_X1  g772(.A1(new_n1184), .A2(KEYINPUT60), .A3(new_n1182), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1198), .A2(new_n642), .ZN(new_n1199));
  NAND4_X1  g774(.A1(new_n632), .A2(KEYINPUT60), .A3(new_n1182), .A4(new_n1184), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1184), .A2(new_n1182), .ZN(new_n1201));
  INV_X1    g776(.A(KEYINPUT60), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  AND3_X1   g778(.A1(new_n1199), .A2(new_n1200), .A3(new_n1203), .ZN(new_n1204));
  OAI21_X1  g779(.A(new_n1186), .B1(new_n1197), .B2(new_n1204), .ZN(new_n1205));
  AND4_X1   g780(.A1(G301), .A2(new_n1156), .A3(new_n1153), .A4(new_n1151), .ZN(new_n1206));
  INV_X1    g781(.A(G171), .ZN(new_n1207));
  NAND4_X1  g782(.A1(new_n468), .A2(KEYINPUT53), .A3(G40), .A4(new_n753), .ZN(new_n1208));
  OAI21_X1  g783(.A(G2105), .B1(new_n470), .B2(KEYINPUT125), .ZN(new_n1209));
  AOI21_X1  g784(.A(new_n1209), .B1(KEYINPUT125), .B2(new_n470), .ZN(new_n1210));
  NOR2_X1   g785(.A1(new_n1208), .A2(new_n1210), .ZN(new_n1211));
  NAND3_X1  g786(.A1(new_n1027), .A2(new_n1067), .A3(new_n1211), .ZN(new_n1212));
  AND2_X1   g787(.A1(new_n1212), .A2(new_n1153), .ZN(new_n1213));
  AOI21_X1  g788(.A(new_n1207), .B1(new_n1213), .B2(new_n1151), .ZN(new_n1214));
  OAI21_X1  g789(.A(KEYINPUT54), .B1(new_n1206), .B2(new_n1214), .ZN(new_n1215));
  NAND3_X1  g790(.A1(new_n1213), .A2(G301), .A3(new_n1151), .ZN(new_n1216));
  INV_X1    g791(.A(KEYINPUT54), .ZN(new_n1217));
  NAND2_X1  g792(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  OAI21_X1  g793(.A(new_n1215), .B1(new_n1157), .B2(new_n1218), .ZN(new_n1219));
  OAI211_X1 g794(.A(new_n1205), .B(new_n1219), .C1(new_n1141), .C2(new_n1140), .ZN(new_n1220));
  NAND2_X1  g795(.A1(new_n1158), .A2(new_n1220), .ZN(new_n1221));
  NOR2_X1   g796(.A1(new_n1094), .A2(new_n1099), .ZN(new_n1222));
  AOI21_X1  g797(.A(new_n1132), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1223));
  XOR2_X1   g798(.A(G290), .B(G1986), .Z(new_n1224));
  OAI21_X1  g799(.A(new_n1038), .B1(new_n1030), .B2(new_n1224), .ZN(new_n1225));
  OAI21_X1  g800(.A(new_n1054), .B1(new_n1223), .B2(new_n1225), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g801(.A1(G229), .A2(new_n458), .A3(G401), .A4(G227), .ZN(new_n1228));
  OAI211_X1 g802(.A(new_n934), .B(new_n1228), .C1(new_n1019), .C2(new_n1020), .ZN(G225));
  INV_X1    g803(.A(G225), .ZN(G308));
endmodule


