

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U551 ( .A1(n716), .A2(n715), .ZN(n725) );
  XNOR2_X2 U552 ( .A(n671), .B(KEYINPUT64), .ZN(n704) );
  INV_X1 U553 ( .A(KEYINPUT30), .ZN(n707) );
  INV_X1 U554 ( .A(KEYINPUT31), .ZN(n713) );
  INV_X1 U555 ( .A(KEYINPUT94), .ZN(n717) );
  NOR2_X1 U556 ( .A1(G1966), .A2(n764), .ZN(n719) );
  INV_X1 U557 ( .A(KEYINPUT97), .ZN(n755) );
  NOR2_X1 U558 ( .A1(G164), .A2(G1384), .ZN(n771) );
  NOR2_X1 U559 ( .A1(n597), .A2(n596), .ZN(n598) );
  AND2_X2 U560 ( .A1(n530), .A2(G2104), .ZN(n872) );
  NOR2_X1 U561 ( .A1(G651), .A2(n639), .ZN(n649) );
  XOR2_X1 U562 ( .A(KEYINPUT1), .B(n521), .Z(n642) );
  NOR2_X1 U563 ( .A1(n539), .A2(n538), .ZN(G160) );
  NOR2_X1 U564 ( .A1(G651), .A2(G543), .ZN(n644) );
  NAND2_X1 U565 ( .A1(n644), .A2(G89), .ZN(n515) );
  XNOR2_X1 U566 ( .A(n515), .B(KEYINPUT4), .ZN(n518) );
  INV_X1 U567 ( .A(G651), .ZN(n520) );
  XOR2_X1 U568 ( .A(G543), .B(KEYINPUT0), .Z(n516) );
  XNOR2_X1 U569 ( .A(KEYINPUT68), .B(n516), .ZN(n639) );
  NOR2_X1 U570 ( .A1(n520), .A2(n639), .ZN(n643) );
  NAND2_X1 U571 ( .A1(G76), .A2(n643), .ZN(n517) );
  NAND2_X1 U572 ( .A1(n518), .A2(n517), .ZN(n519) );
  XNOR2_X1 U573 ( .A(n519), .B(KEYINPUT5), .ZN(n526) );
  NOR2_X1 U574 ( .A1(G543), .A2(n520), .ZN(n521) );
  NAND2_X1 U575 ( .A1(G63), .A2(n642), .ZN(n523) );
  NAND2_X1 U576 ( .A1(G51), .A2(n649), .ZN(n522) );
  NAND2_X1 U577 ( .A1(n523), .A2(n522), .ZN(n524) );
  XOR2_X1 U578 ( .A(KEYINPUT6), .B(n524), .Z(n525) );
  NAND2_X1 U579 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U580 ( .A(n527), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U581 ( .A(KEYINPUT66), .B(KEYINPUT23), .Z(n529) );
  INV_X1 U582 ( .A(G2105), .ZN(n530) );
  NAND2_X1 U583 ( .A1(G101), .A2(n872), .ZN(n528) );
  XNOR2_X1 U584 ( .A(n529), .B(n528), .ZN(n533) );
  NOR2_X1 U585 ( .A1(G2104), .A2(n530), .ZN(n563) );
  NAND2_X1 U586 ( .A1(G125), .A2(n563), .ZN(n531) );
  XOR2_X1 U587 ( .A(KEYINPUT65), .B(n531), .Z(n532) );
  NAND2_X1 U588 ( .A1(n533), .A2(n532), .ZN(n539) );
  XNOR2_X1 U589 ( .A(KEYINPUT17), .B(KEYINPUT67), .ZN(n535) );
  NOR2_X1 U590 ( .A1(G2104), .A2(G2105), .ZN(n534) );
  XNOR2_X2 U591 ( .A(n535), .B(n534), .ZN(n871) );
  NAND2_X1 U592 ( .A1(G137), .A2(n871), .ZN(n537) );
  AND2_X1 U593 ( .A1(G2104), .A2(G2105), .ZN(n875) );
  NAND2_X1 U594 ( .A1(G113), .A2(n875), .ZN(n536) );
  NAND2_X1 U595 ( .A1(n537), .A2(n536), .ZN(n538) );
  NAND2_X1 U596 ( .A1(G138), .A2(n871), .ZN(n541) );
  NAND2_X1 U597 ( .A1(G102), .A2(n872), .ZN(n540) );
  NAND2_X1 U598 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U599 ( .A(n542), .B(KEYINPUT82), .ZN(n546) );
  NAND2_X1 U600 ( .A1(G114), .A2(n875), .ZN(n544) );
  NAND2_X1 U601 ( .A1(G126), .A2(n563), .ZN(n543) );
  NAND2_X1 U602 ( .A1(n544), .A2(n543), .ZN(n545) );
  NOR2_X1 U603 ( .A1(n546), .A2(n545), .ZN(G164) );
  XNOR2_X1 U604 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  INV_X1 U605 ( .A(G82), .ZN(G220) );
  INV_X1 U606 ( .A(G132), .ZN(G219) );
  XNOR2_X1 U607 ( .A(KEYINPUT71), .B(G57), .ZN(G237) );
  NOR2_X1 U608 ( .A1(G220), .A2(G219), .ZN(n547) );
  XOR2_X1 U609 ( .A(KEYINPUT22), .B(n547), .Z(n548) );
  NOR2_X1 U610 ( .A1(G218), .A2(n548), .ZN(n549) );
  NAND2_X1 U611 ( .A1(G96), .A2(n549), .ZN(n915) );
  NAND2_X1 U612 ( .A1(n915), .A2(G2106), .ZN(n553) );
  NAND2_X1 U613 ( .A1(G108), .A2(G120), .ZN(n550) );
  NOR2_X1 U614 ( .A1(G237), .A2(n550), .ZN(n551) );
  NAND2_X1 U615 ( .A1(G69), .A2(n551), .ZN(n916) );
  NAND2_X1 U616 ( .A1(n916), .A2(G567), .ZN(n552) );
  AND2_X1 U617 ( .A1(n553), .A2(n552), .ZN(G319) );
  NAND2_X1 U618 ( .A1(G64), .A2(n642), .ZN(n555) );
  NAND2_X1 U619 ( .A1(G52), .A2(n649), .ZN(n554) );
  NAND2_X1 U620 ( .A1(n555), .A2(n554), .ZN(n560) );
  NAND2_X1 U621 ( .A1(G77), .A2(n643), .ZN(n557) );
  NAND2_X1 U622 ( .A1(G90), .A2(n644), .ZN(n556) );
  NAND2_X1 U623 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U624 ( .A(KEYINPUT9), .B(n558), .Z(n559) );
  NOR2_X1 U625 ( .A1(n560), .A2(n559), .ZN(G171) );
  AND2_X1 U626 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U627 ( .A1(G135), .A2(n871), .ZN(n562) );
  NAND2_X1 U628 ( .A1(G111), .A2(n875), .ZN(n561) );
  NAND2_X1 U629 ( .A1(n562), .A2(n561), .ZN(n567) );
  INV_X1 U630 ( .A(n563), .ZN(n564) );
  INV_X1 U631 ( .A(n564), .ZN(n876) );
  NAND2_X1 U632 ( .A1(n876), .A2(G123), .ZN(n565) );
  XOR2_X1 U633 ( .A(KEYINPUT18), .B(n565), .Z(n566) );
  NOR2_X1 U634 ( .A1(n567), .A2(n566), .ZN(n569) );
  NAND2_X1 U635 ( .A1(n872), .A2(G99), .ZN(n568) );
  NAND2_X1 U636 ( .A1(n569), .A2(n568), .ZN(n918) );
  XNOR2_X1 U637 ( .A(G2096), .B(n918), .ZN(n570) );
  OR2_X1 U638 ( .A1(G2100), .A2(n570), .ZN(G156) );
  NAND2_X1 U639 ( .A1(G75), .A2(n643), .ZN(n572) );
  NAND2_X1 U640 ( .A1(G88), .A2(n644), .ZN(n571) );
  NAND2_X1 U641 ( .A1(n572), .A2(n571), .ZN(n576) );
  NAND2_X1 U642 ( .A1(G62), .A2(n642), .ZN(n574) );
  NAND2_X1 U643 ( .A1(G50), .A2(n649), .ZN(n573) );
  NAND2_X1 U644 ( .A1(n574), .A2(n573), .ZN(n575) );
  NOR2_X1 U645 ( .A1(n576), .A2(n575), .ZN(G166) );
  XOR2_X1 U646 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U647 ( .A1(G7), .A2(G661), .ZN(n577) );
  XNOR2_X1 U648 ( .A(n577), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U649 ( .A(G223), .ZN(n819) );
  NAND2_X1 U650 ( .A1(n819), .A2(G567), .ZN(n578) );
  XOR2_X1 U651 ( .A(KEYINPUT11), .B(n578), .Z(G234) );
  NAND2_X1 U652 ( .A1(G56), .A2(n642), .ZN(n579) );
  XOR2_X1 U653 ( .A(KEYINPUT14), .B(n579), .Z(n586) );
  NAND2_X1 U654 ( .A1(n644), .A2(G81), .ZN(n580) );
  XOR2_X1 U655 ( .A(KEYINPUT12), .B(n580), .Z(n583) );
  NAND2_X1 U656 ( .A1(n643), .A2(G68), .ZN(n581) );
  XOR2_X1 U657 ( .A(KEYINPUT72), .B(n581), .Z(n582) );
  NOR2_X1 U658 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U659 ( .A(n584), .B(KEYINPUT13), .ZN(n585) );
  NOR2_X1 U660 ( .A1(n586), .A2(n585), .ZN(n588) );
  NAND2_X1 U661 ( .A1(n649), .A2(G43), .ZN(n587) );
  NAND2_X1 U662 ( .A1(n588), .A2(n587), .ZN(n971) );
  INV_X1 U663 ( .A(G860), .ZN(n618) );
  OR2_X1 U664 ( .A1(n971), .A2(n618), .ZN(G153) );
  INV_X1 U665 ( .A(G171), .ZN(G301) );
  NAND2_X1 U666 ( .A1(G868), .A2(G301), .ZN(n600) );
  NAND2_X1 U667 ( .A1(G79), .A2(n643), .ZN(n590) );
  NAND2_X1 U668 ( .A1(G54), .A2(n649), .ZN(n589) );
  NAND2_X1 U669 ( .A1(n590), .A2(n589), .ZN(n597) );
  NAND2_X1 U670 ( .A1(n642), .A2(G66), .ZN(n591) );
  XNOR2_X1 U671 ( .A(KEYINPUT73), .B(n591), .ZN(n594) );
  NAND2_X1 U672 ( .A1(n644), .A2(G92), .ZN(n592) );
  XOR2_X1 U673 ( .A(KEYINPUT74), .B(n592), .Z(n593) );
  NOR2_X1 U674 ( .A1(n594), .A2(n593), .ZN(n595) );
  XNOR2_X1 U675 ( .A(n595), .B(KEYINPUT75), .ZN(n596) );
  XOR2_X1 U676 ( .A(KEYINPUT15), .B(n598), .Z(n986) );
  OR2_X1 U677 ( .A1(n986), .A2(G868), .ZN(n599) );
  NAND2_X1 U678 ( .A1(n600), .A2(n599), .ZN(G284) );
  NAND2_X1 U679 ( .A1(n644), .A2(G91), .ZN(n601) );
  XOR2_X1 U680 ( .A(KEYINPUT69), .B(n601), .Z(n603) );
  NAND2_X1 U681 ( .A1(n643), .A2(G78), .ZN(n602) );
  NAND2_X1 U682 ( .A1(n603), .A2(n602), .ZN(n604) );
  XOR2_X1 U683 ( .A(KEYINPUT70), .B(n604), .Z(n608) );
  NAND2_X1 U684 ( .A1(G65), .A2(n642), .ZN(n606) );
  NAND2_X1 U685 ( .A1(G53), .A2(n649), .ZN(n605) );
  AND2_X1 U686 ( .A1(n606), .A2(n605), .ZN(n607) );
  NAND2_X1 U687 ( .A1(n608), .A2(n607), .ZN(G299) );
  INV_X1 U688 ( .A(G868), .ZN(n609) );
  NOR2_X1 U689 ( .A1(G286), .A2(n609), .ZN(n611) );
  NOR2_X1 U690 ( .A1(G868), .A2(G299), .ZN(n610) );
  NOR2_X1 U691 ( .A1(n611), .A2(n610), .ZN(G297) );
  NAND2_X1 U692 ( .A1(n618), .A2(G559), .ZN(n612) );
  NAND2_X1 U693 ( .A1(n612), .A2(n986), .ZN(n613) );
  XNOR2_X1 U694 ( .A(n613), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U695 ( .A1(G868), .A2(n971), .ZN(n616) );
  NAND2_X1 U696 ( .A1(G868), .A2(n986), .ZN(n614) );
  NOR2_X1 U697 ( .A1(G559), .A2(n614), .ZN(n615) );
  NOR2_X1 U698 ( .A1(n616), .A2(n615), .ZN(G282) );
  NAND2_X1 U699 ( .A1(G559), .A2(n986), .ZN(n617) );
  XOR2_X1 U700 ( .A(n971), .B(n617), .Z(n658) );
  NAND2_X1 U701 ( .A1(n618), .A2(n658), .ZN(n626) );
  NAND2_X1 U702 ( .A1(G67), .A2(n642), .ZN(n620) );
  NAND2_X1 U703 ( .A1(G55), .A2(n649), .ZN(n619) );
  NAND2_X1 U704 ( .A1(n620), .A2(n619), .ZN(n621) );
  XNOR2_X1 U705 ( .A(KEYINPUT76), .B(n621), .ZN(n625) );
  NAND2_X1 U706 ( .A1(G80), .A2(n643), .ZN(n623) );
  NAND2_X1 U707 ( .A1(G93), .A2(n644), .ZN(n622) );
  NAND2_X1 U708 ( .A1(n623), .A2(n622), .ZN(n624) );
  NOR2_X1 U709 ( .A1(n625), .A2(n624), .ZN(n660) );
  XOR2_X1 U710 ( .A(n626), .B(n660), .Z(G145) );
  NAND2_X1 U711 ( .A1(G61), .A2(n642), .ZN(n628) );
  NAND2_X1 U712 ( .A1(G86), .A2(n644), .ZN(n627) );
  NAND2_X1 U713 ( .A1(n628), .A2(n627), .ZN(n629) );
  XNOR2_X1 U714 ( .A(KEYINPUT77), .B(n629), .ZN(n635) );
  NAND2_X1 U715 ( .A1(G73), .A2(n643), .ZN(n630) );
  XOR2_X1 U716 ( .A(KEYINPUT2), .B(n630), .Z(n633) );
  NAND2_X1 U717 ( .A1(n649), .A2(G48), .ZN(n631) );
  XOR2_X1 U718 ( .A(KEYINPUT78), .B(n631), .Z(n632) );
  NOR2_X1 U719 ( .A1(n633), .A2(n632), .ZN(n634) );
  NAND2_X1 U720 ( .A1(n635), .A2(n634), .ZN(G305) );
  NAND2_X1 U721 ( .A1(G49), .A2(n649), .ZN(n637) );
  NAND2_X1 U722 ( .A1(G74), .A2(G651), .ZN(n636) );
  NAND2_X1 U723 ( .A1(n637), .A2(n636), .ZN(n638) );
  NOR2_X1 U724 ( .A1(n642), .A2(n638), .ZN(n641) );
  NAND2_X1 U725 ( .A1(G87), .A2(n639), .ZN(n640) );
  NAND2_X1 U726 ( .A1(n641), .A2(n640), .ZN(G288) );
  AND2_X1 U727 ( .A1(n642), .A2(G60), .ZN(n648) );
  NAND2_X1 U728 ( .A1(G72), .A2(n643), .ZN(n646) );
  NAND2_X1 U729 ( .A1(G85), .A2(n644), .ZN(n645) );
  NAND2_X1 U730 ( .A1(n646), .A2(n645), .ZN(n647) );
  NOR2_X1 U731 ( .A1(n648), .A2(n647), .ZN(n651) );
  NAND2_X1 U732 ( .A1(n649), .A2(G47), .ZN(n650) );
  NAND2_X1 U733 ( .A1(n651), .A2(n650), .ZN(G290) );
  XNOR2_X1 U734 ( .A(KEYINPUT79), .B(G305), .ZN(n652) );
  XNOR2_X1 U735 ( .A(n652), .B(G288), .ZN(n653) );
  XNOR2_X1 U736 ( .A(KEYINPUT19), .B(n653), .ZN(n655) );
  XNOR2_X1 U737 ( .A(G290), .B(G166), .ZN(n654) );
  XNOR2_X1 U738 ( .A(n655), .B(n654), .ZN(n656) );
  XOR2_X1 U739 ( .A(n660), .B(n656), .Z(n657) );
  XNOR2_X1 U740 ( .A(G299), .B(n657), .ZN(n846) );
  XNOR2_X1 U741 ( .A(n658), .B(n846), .ZN(n659) );
  NAND2_X1 U742 ( .A1(n659), .A2(G868), .ZN(n662) );
  OR2_X1 U743 ( .A1(G868), .A2(n660), .ZN(n661) );
  NAND2_X1 U744 ( .A1(n662), .A2(n661), .ZN(G295) );
  NAND2_X1 U745 ( .A1(G2084), .A2(G2078), .ZN(n663) );
  XOR2_X1 U746 ( .A(KEYINPUT20), .B(n663), .Z(n664) );
  NAND2_X1 U747 ( .A1(G2090), .A2(n664), .ZN(n665) );
  XNOR2_X1 U748 ( .A(KEYINPUT21), .B(n665), .ZN(n666) );
  NAND2_X1 U749 ( .A1(n666), .A2(G2072), .ZN(G158) );
  NAND2_X1 U750 ( .A1(G661), .A2(G483), .ZN(n667) );
  XOR2_X1 U751 ( .A(KEYINPUT80), .B(n667), .Z(n668) );
  NAND2_X1 U752 ( .A1(n668), .A2(G319), .ZN(n669) );
  XNOR2_X1 U753 ( .A(n669), .B(KEYINPUT81), .ZN(n823) );
  NAND2_X1 U754 ( .A1(n823), .A2(G36), .ZN(G176) );
  INV_X1 U755 ( .A(G166), .ZN(G303) );
  NAND2_X1 U756 ( .A1(G160), .A2(G40), .ZN(n770) );
  XOR2_X1 U757 ( .A(KEYINPUT86), .B(n770), .Z(n670) );
  NAND2_X1 U758 ( .A1(n670), .A2(n771), .ZN(n671) );
  NAND2_X1 U759 ( .A1(n704), .A2(G8), .ZN(n672) );
  XNOR2_X1 U760 ( .A(n672), .B(KEYINPUT87), .ZN(n758) );
  INV_X1 U761 ( .A(n758), .ZN(n764) );
  XOR2_X1 U762 ( .A(G1996), .B(KEYINPUT92), .Z(n944) );
  NOR2_X1 U763 ( .A1(n704), .A2(n944), .ZN(n673) );
  XOR2_X1 U764 ( .A(n673), .B(KEYINPUT26), .Z(n675) );
  NAND2_X1 U765 ( .A1(n704), .A2(G1341), .ZN(n674) );
  NAND2_X1 U766 ( .A1(n675), .A2(n674), .ZN(n686) );
  INV_X1 U767 ( .A(n704), .ZN(n699) );
  NAND2_X1 U768 ( .A1(G2067), .A2(n699), .ZN(n677) );
  NAND2_X1 U769 ( .A1(n704), .A2(G1348), .ZN(n676) );
  NAND2_X1 U770 ( .A1(n677), .A2(n676), .ZN(n679) );
  OR2_X1 U771 ( .A1(n971), .A2(n679), .ZN(n678) );
  NOR2_X1 U772 ( .A1(n686), .A2(n678), .ZN(n682) );
  INV_X1 U773 ( .A(n679), .ZN(n680) );
  AND2_X1 U774 ( .A1(n680), .A2(n986), .ZN(n681) );
  NOR2_X1 U775 ( .A1(n682), .A2(n681), .ZN(n691) );
  NAND2_X1 U776 ( .A1(G2072), .A2(n699), .ZN(n683) );
  XOR2_X1 U777 ( .A(KEYINPUT27), .B(n683), .Z(n685) );
  NAND2_X1 U778 ( .A1(n704), .A2(G1956), .ZN(n684) );
  NAND2_X1 U779 ( .A1(n685), .A2(n684), .ZN(n693) );
  NOR2_X1 U780 ( .A1(n693), .A2(G299), .ZN(n689) );
  NOR2_X1 U781 ( .A1(n971), .A2(n686), .ZN(n687) );
  AND2_X1 U782 ( .A1(n986), .A2(n687), .ZN(n688) );
  NOR2_X1 U783 ( .A1(n689), .A2(n688), .ZN(n690) );
  NAND2_X1 U784 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U785 ( .A(n692), .B(KEYINPUT93), .ZN(n697) );
  NAND2_X1 U786 ( .A1(n693), .A2(G299), .ZN(n694) );
  XNOR2_X1 U787 ( .A(n694), .B(KEYINPUT91), .ZN(n695) );
  XNOR2_X1 U788 ( .A(n695), .B(KEYINPUT28), .ZN(n696) );
  NOR2_X1 U789 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U790 ( .A(n698), .B(KEYINPUT29), .ZN(n703) );
  XNOR2_X1 U791 ( .A(G2078), .B(KEYINPUT25), .ZN(n945) );
  NAND2_X1 U792 ( .A1(n699), .A2(n945), .ZN(n701) );
  XOR2_X1 U793 ( .A(G1961), .B(KEYINPUT90), .Z(n1012) );
  NAND2_X1 U794 ( .A1(n704), .A2(n1012), .ZN(n700) );
  NAND2_X1 U795 ( .A1(n701), .A2(n700), .ZN(n710) );
  NAND2_X1 U796 ( .A1(G171), .A2(n710), .ZN(n702) );
  NAND2_X1 U797 ( .A1(n703), .A2(n702), .ZN(n716) );
  NOR2_X1 U798 ( .A1(n704), .A2(G2084), .ZN(n705) );
  XNOR2_X1 U799 ( .A(KEYINPUT89), .B(n705), .ZN(n720) );
  NAND2_X1 U800 ( .A1(G8), .A2(n720), .ZN(n706) );
  NOR2_X1 U801 ( .A1(n719), .A2(n706), .ZN(n708) );
  XNOR2_X1 U802 ( .A(n708), .B(n707), .ZN(n709) );
  NOR2_X1 U803 ( .A1(n709), .A2(G168), .ZN(n712) );
  NOR2_X1 U804 ( .A1(G171), .A2(n710), .ZN(n711) );
  NOR2_X1 U805 ( .A1(n712), .A2(n711), .ZN(n714) );
  XNOR2_X1 U806 ( .A(n714), .B(n713), .ZN(n715) );
  XNOR2_X1 U807 ( .A(n725), .B(n717), .ZN(n718) );
  NOR2_X1 U808 ( .A1(n719), .A2(n718), .ZN(n723) );
  INV_X1 U809 ( .A(n720), .ZN(n721) );
  NAND2_X1 U810 ( .A1(G8), .A2(n721), .ZN(n722) );
  NAND2_X1 U811 ( .A1(n723), .A2(n722), .ZN(n736) );
  AND2_X1 U812 ( .A1(G286), .A2(G8), .ZN(n724) );
  NAND2_X1 U813 ( .A1(n725), .A2(n724), .ZN(n733) );
  INV_X1 U814 ( .A(G8), .ZN(n731) );
  NOR2_X1 U815 ( .A1(G1971), .A2(n764), .ZN(n727) );
  NOR2_X1 U816 ( .A1(n704), .A2(G2090), .ZN(n726) );
  NOR2_X1 U817 ( .A1(n727), .A2(n726), .ZN(n728) );
  XOR2_X1 U818 ( .A(KEYINPUT95), .B(n728), .Z(n729) );
  NAND2_X1 U819 ( .A1(n729), .A2(G303), .ZN(n730) );
  OR2_X1 U820 ( .A1(n731), .A2(n730), .ZN(n732) );
  AND2_X1 U821 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U822 ( .A(KEYINPUT32), .B(n734), .ZN(n735) );
  NAND2_X1 U823 ( .A1(n736), .A2(n735), .ZN(n763) );
  INV_X1 U824 ( .A(n763), .ZN(n746) );
  NOR2_X1 U825 ( .A1(G1976), .A2(G288), .ZN(n739) );
  INV_X1 U826 ( .A(n739), .ZN(n738) );
  INV_X1 U827 ( .A(G1971), .ZN(n1004) );
  NAND2_X1 U828 ( .A1(G166), .A2(n1004), .ZN(n737) );
  NAND2_X1 U829 ( .A1(n738), .A2(n737), .ZN(n982) );
  XNOR2_X1 U830 ( .A(G1981), .B(G305), .ZN(n969) );
  INV_X1 U831 ( .A(KEYINPUT33), .ZN(n742) );
  NAND2_X1 U832 ( .A1(n758), .A2(n739), .ZN(n740) );
  NOR2_X1 U833 ( .A1(n742), .A2(n740), .ZN(n741) );
  XNOR2_X1 U834 ( .A(n741), .B(KEYINPUT96), .ZN(n748) );
  OR2_X1 U835 ( .A1(n748), .A2(n742), .ZN(n743) );
  OR2_X1 U836 ( .A1(n969), .A2(n743), .ZN(n752) );
  INV_X1 U837 ( .A(n752), .ZN(n744) );
  OR2_X1 U838 ( .A1(n982), .A2(n744), .ZN(n745) );
  NOR2_X1 U839 ( .A1(n746), .A2(n745), .ZN(n754) );
  NAND2_X1 U840 ( .A1(G1976), .A2(G288), .ZN(n975) );
  INV_X1 U841 ( .A(n975), .ZN(n747) );
  OR2_X1 U842 ( .A1(n747), .A2(n764), .ZN(n749) );
  OR2_X1 U843 ( .A1(n749), .A2(n748), .ZN(n750) );
  OR2_X1 U844 ( .A1(n750), .A2(n969), .ZN(n751) );
  AND2_X1 U845 ( .A1(n752), .A2(n751), .ZN(n753) );
  NOR2_X1 U846 ( .A1(n754), .A2(n753), .ZN(n756) );
  XNOR2_X1 U847 ( .A(n756), .B(n755), .ZN(n769) );
  NOR2_X1 U848 ( .A1(G1981), .A2(G305), .ZN(n757) );
  XNOR2_X1 U849 ( .A(n757), .B(KEYINPUT24), .ZN(n759) );
  NAND2_X1 U850 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U851 ( .A(n760), .B(KEYINPUT88), .ZN(n767) );
  NOR2_X1 U852 ( .A1(G2090), .A2(G303), .ZN(n761) );
  NAND2_X1 U853 ( .A1(G8), .A2(n761), .ZN(n762) );
  NAND2_X1 U854 ( .A1(n763), .A2(n762), .ZN(n765) );
  NAND2_X1 U855 ( .A1(n765), .A2(n764), .ZN(n766) );
  NAND2_X1 U856 ( .A1(n767), .A2(n766), .ZN(n768) );
  NOR2_X1 U857 ( .A1(n769), .A2(n768), .ZN(n791) );
  NOR2_X1 U858 ( .A1(n771), .A2(n770), .ZN(n814) );
  XOR2_X1 U859 ( .A(KEYINPUT84), .B(KEYINPUT38), .Z(n773) );
  NAND2_X1 U860 ( .A1(G105), .A2(n872), .ZN(n772) );
  XNOR2_X1 U861 ( .A(n773), .B(n772), .ZN(n777) );
  NAND2_X1 U862 ( .A1(G141), .A2(n871), .ZN(n775) );
  NAND2_X1 U863 ( .A1(G117), .A2(n875), .ZN(n774) );
  NAND2_X1 U864 ( .A1(n775), .A2(n774), .ZN(n776) );
  NOR2_X1 U865 ( .A1(n777), .A2(n776), .ZN(n779) );
  NAND2_X1 U866 ( .A1(n876), .A2(G129), .ZN(n778) );
  NAND2_X1 U867 ( .A1(n779), .A2(n778), .ZN(n884) );
  NAND2_X1 U868 ( .A1(G1996), .A2(n884), .ZN(n787) );
  NAND2_X1 U869 ( .A1(G131), .A2(n871), .ZN(n781) );
  NAND2_X1 U870 ( .A1(G107), .A2(n875), .ZN(n780) );
  NAND2_X1 U871 ( .A1(n781), .A2(n780), .ZN(n785) );
  NAND2_X1 U872 ( .A1(G95), .A2(n872), .ZN(n783) );
  NAND2_X1 U873 ( .A1(G119), .A2(n876), .ZN(n782) );
  NAND2_X1 U874 ( .A1(n783), .A2(n782), .ZN(n784) );
  OR2_X1 U875 ( .A1(n785), .A2(n784), .ZN(n888) );
  NAND2_X1 U876 ( .A1(G1991), .A2(n888), .ZN(n786) );
  NAND2_X1 U877 ( .A1(n787), .A2(n786), .ZN(n927) );
  NAND2_X1 U878 ( .A1(n814), .A2(n927), .ZN(n806) );
  XOR2_X1 U879 ( .A(n806), .B(KEYINPUT85), .Z(n789) );
  XNOR2_X1 U880 ( .A(G1986), .B(G290), .ZN(n977) );
  NAND2_X1 U881 ( .A1(n977), .A2(n814), .ZN(n788) );
  NAND2_X1 U882 ( .A1(n789), .A2(n788), .ZN(n790) );
  NOR2_X1 U883 ( .A1(n791), .A2(n790), .ZN(n802) );
  XNOR2_X1 U884 ( .A(G2067), .B(KEYINPUT37), .ZN(n812) );
  NAND2_X1 U885 ( .A1(n871), .A2(G140), .ZN(n792) );
  XOR2_X1 U886 ( .A(KEYINPUT83), .B(n792), .Z(n794) );
  NAND2_X1 U887 ( .A1(n872), .A2(G104), .ZN(n793) );
  NAND2_X1 U888 ( .A1(n794), .A2(n793), .ZN(n795) );
  XNOR2_X1 U889 ( .A(KEYINPUT34), .B(n795), .ZN(n800) );
  NAND2_X1 U890 ( .A1(G116), .A2(n875), .ZN(n797) );
  NAND2_X1 U891 ( .A1(G128), .A2(n876), .ZN(n796) );
  NAND2_X1 U892 ( .A1(n797), .A2(n796), .ZN(n798) );
  XOR2_X1 U893 ( .A(KEYINPUT35), .B(n798), .Z(n799) );
  NOR2_X1 U894 ( .A1(n800), .A2(n799), .ZN(n801) );
  XNOR2_X1 U895 ( .A(KEYINPUT36), .B(n801), .ZN(n894) );
  NOR2_X1 U896 ( .A1(n812), .A2(n894), .ZN(n939) );
  NAND2_X1 U897 ( .A1(n814), .A2(n939), .ZN(n810) );
  NAND2_X1 U898 ( .A1(n802), .A2(n810), .ZN(n817) );
  NOR2_X1 U899 ( .A1(G1996), .A2(n884), .ZN(n803) );
  XOR2_X1 U900 ( .A(KEYINPUT98), .B(n803), .Z(n922) );
  NOR2_X1 U901 ( .A1(G1986), .A2(G290), .ZN(n804) );
  XNOR2_X1 U902 ( .A(KEYINPUT99), .B(n804), .ZN(n805) );
  OR2_X1 U903 ( .A1(n888), .A2(G1991), .ZN(n919) );
  NAND2_X1 U904 ( .A1(n805), .A2(n919), .ZN(n807) );
  NAND2_X1 U905 ( .A1(n807), .A2(n806), .ZN(n808) );
  NAND2_X1 U906 ( .A1(n922), .A2(n808), .ZN(n809) );
  XOR2_X1 U907 ( .A(KEYINPUT39), .B(n809), .Z(n811) );
  NAND2_X1 U908 ( .A1(n811), .A2(n810), .ZN(n813) );
  NAND2_X1 U909 ( .A1(n812), .A2(n894), .ZN(n936) );
  NAND2_X1 U910 ( .A1(n813), .A2(n936), .ZN(n815) );
  NAND2_X1 U911 ( .A1(n815), .A2(n814), .ZN(n816) );
  NAND2_X1 U912 ( .A1(n817), .A2(n816), .ZN(n818) );
  XNOR2_X1 U913 ( .A(n818), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U914 ( .A1(n819), .A2(G2106), .ZN(n820) );
  XNOR2_X1 U915 ( .A(n820), .B(KEYINPUT102), .ZN(G217) );
  AND2_X1 U916 ( .A1(G15), .A2(G2), .ZN(n821) );
  NAND2_X1 U917 ( .A1(G661), .A2(n821), .ZN(G259) );
  NAND2_X1 U918 ( .A1(G3), .A2(G1), .ZN(n822) );
  NAND2_X1 U919 ( .A1(n823), .A2(n822), .ZN(G188) );
  XOR2_X1 U920 ( .A(KEYINPUT42), .B(G2090), .Z(n825) );
  XNOR2_X1 U921 ( .A(G2084), .B(G2078), .ZN(n824) );
  XNOR2_X1 U922 ( .A(n825), .B(n824), .ZN(n826) );
  XOR2_X1 U923 ( .A(n826), .B(G2100), .Z(n828) );
  XNOR2_X1 U924 ( .A(G2067), .B(G2072), .ZN(n827) );
  XNOR2_X1 U925 ( .A(n828), .B(n827), .ZN(n832) );
  XOR2_X1 U926 ( .A(G2096), .B(KEYINPUT43), .Z(n830) );
  XNOR2_X1 U927 ( .A(KEYINPUT103), .B(G2678), .ZN(n829) );
  XNOR2_X1 U928 ( .A(n830), .B(n829), .ZN(n831) );
  XOR2_X1 U929 ( .A(n832), .B(n831), .Z(G227) );
  XOR2_X1 U930 ( .A(KEYINPUT105), .B(G1981), .Z(n834) );
  XNOR2_X1 U931 ( .A(G1996), .B(G1991), .ZN(n833) );
  XNOR2_X1 U932 ( .A(n834), .B(n833), .ZN(n835) );
  XOR2_X1 U933 ( .A(n835), .B(KEYINPUT41), .Z(n837) );
  XNOR2_X1 U934 ( .A(G1956), .B(G1976), .ZN(n836) );
  XNOR2_X1 U935 ( .A(n837), .B(n836), .ZN(n841) );
  XOR2_X1 U936 ( .A(G1971), .B(G1961), .Z(n839) );
  XNOR2_X1 U937 ( .A(G1986), .B(G1966), .ZN(n838) );
  XNOR2_X1 U938 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U939 ( .A(n841), .B(n840), .Z(n843) );
  XNOR2_X1 U940 ( .A(KEYINPUT104), .B(G2474), .ZN(n842) );
  XNOR2_X1 U941 ( .A(n843), .B(n842), .ZN(G229) );
  XNOR2_X1 U942 ( .A(n971), .B(KEYINPUT115), .ZN(n845) );
  XNOR2_X1 U943 ( .A(G171), .B(n986), .ZN(n844) );
  XNOR2_X1 U944 ( .A(n845), .B(n844), .ZN(n848) );
  XOR2_X1 U945 ( .A(G286), .B(n846), .Z(n847) );
  XNOR2_X1 U946 ( .A(n848), .B(n847), .ZN(n849) );
  NOR2_X1 U947 ( .A1(G37), .A2(n849), .ZN(G397) );
  NAND2_X1 U948 ( .A1(n876), .A2(G124), .ZN(n850) );
  XNOR2_X1 U949 ( .A(n850), .B(KEYINPUT44), .ZN(n852) );
  NAND2_X1 U950 ( .A1(G136), .A2(n871), .ZN(n851) );
  NAND2_X1 U951 ( .A1(n852), .A2(n851), .ZN(n853) );
  XOR2_X1 U952 ( .A(KEYINPUT106), .B(n853), .Z(n855) );
  NAND2_X1 U953 ( .A1(n875), .A2(G112), .ZN(n854) );
  NAND2_X1 U954 ( .A1(n855), .A2(n854), .ZN(n858) );
  NAND2_X1 U955 ( .A1(G100), .A2(n872), .ZN(n856) );
  XNOR2_X1 U956 ( .A(KEYINPUT107), .B(n856), .ZN(n857) );
  NOR2_X1 U957 ( .A1(n858), .A2(n857), .ZN(G162) );
  XNOR2_X1 U958 ( .A(KEYINPUT109), .B(KEYINPUT110), .ZN(n863) );
  NAND2_X1 U959 ( .A1(G142), .A2(n871), .ZN(n860) );
  NAND2_X1 U960 ( .A1(G106), .A2(n872), .ZN(n859) );
  NAND2_X1 U961 ( .A1(n860), .A2(n859), .ZN(n861) );
  XNOR2_X1 U962 ( .A(n861), .B(KEYINPUT45), .ZN(n862) );
  XNOR2_X1 U963 ( .A(n863), .B(n862), .ZN(n868) );
  NAND2_X1 U964 ( .A1(n875), .A2(G118), .ZN(n864) );
  XNOR2_X1 U965 ( .A(n864), .B(KEYINPUT108), .ZN(n866) );
  NAND2_X1 U966 ( .A1(G130), .A2(n876), .ZN(n865) );
  NAND2_X1 U967 ( .A1(n866), .A2(n865), .ZN(n867) );
  NOR2_X1 U968 ( .A1(n868), .A2(n867), .ZN(n893) );
  XOR2_X1 U969 ( .A(KEYINPUT48), .B(KEYINPUT113), .Z(n870) );
  XNOR2_X1 U970 ( .A(G162), .B(KEYINPUT46), .ZN(n869) );
  XNOR2_X1 U971 ( .A(n870), .B(n869), .ZN(n887) );
  NAND2_X1 U972 ( .A1(G139), .A2(n871), .ZN(n874) );
  NAND2_X1 U973 ( .A1(G103), .A2(n872), .ZN(n873) );
  NAND2_X1 U974 ( .A1(n874), .A2(n873), .ZN(n883) );
  XNOR2_X1 U975 ( .A(KEYINPUT47), .B(KEYINPUT112), .ZN(n881) );
  NAND2_X1 U976 ( .A1(n875), .A2(G115), .ZN(n879) );
  NAND2_X1 U977 ( .A1(n876), .A2(G127), .ZN(n877) );
  XOR2_X1 U978 ( .A(KEYINPUT111), .B(n877), .Z(n878) );
  NAND2_X1 U979 ( .A1(n879), .A2(n878), .ZN(n880) );
  XOR2_X1 U980 ( .A(n881), .B(n880), .Z(n882) );
  NOR2_X1 U981 ( .A1(n883), .A2(n882), .ZN(n930) );
  XNOR2_X1 U982 ( .A(n930), .B(n884), .ZN(n885) );
  XNOR2_X1 U983 ( .A(n885), .B(n918), .ZN(n886) );
  XOR2_X1 U984 ( .A(n887), .B(n886), .Z(n890) );
  XOR2_X1 U985 ( .A(G160), .B(n888), .Z(n889) );
  XNOR2_X1 U986 ( .A(n890), .B(n889), .ZN(n891) );
  XNOR2_X1 U987 ( .A(G164), .B(n891), .ZN(n892) );
  XNOR2_X1 U988 ( .A(n893), .B(n892), .ZN(n895) );
  XOR2_X1 U989 ( .A(n895), .B(n894), .Z(n896) );
  NOR2_X1 U990 ( .A1(G37), .A2(n896), .ZN(n897) );
  XNOR2_X1 U991 ( .A(KEYINPUT114), .B(n897), .ZN(G395) );
  XNOR2_X1 U992 ( .A(KEYINPUT116), .B(KEYINPUT49), .ZN(n899) );
  NOR2_X1 U993 ( .A1(G227), .A2(G229), .ZN(n898) );
  XNOR2_X1 U994 ( .A(n899), .B(n898), .ZN(n912) );
  XNOR2_X1 U995 ( .A(G2454), .B(G2443), .ZN(n909) );
  XOR2_X1 U996 ( .A(KEYINPUT100), .B(G2430), .Z(n901) );
  XNOR2_X1 U997 ( .A(G2446), .B(KEYINPUT101), .ZN(n900) );
  XNOR2_X1 U998 ( .A(n901), .B(n900), .ZN(n905) );
  XOR2_X1 U999 ( .A(G2451), .B(G2427), .Z(n903) );
  XNOR2_X1 U1000 ( .A(G1348), .B(G1341), .ZN(n902) );
  XNOR2_X1 U1001 ( .A(n903), .B(n902), .ZN(n904) );
  XOR2_X1 U1002 ( .A(n905), .B(n904), .Z(n907) );
  XNOR2_X1 U1003 ( .A(G2435), .B(G2438), .ZN(n906) );
  XNOR2_X1 U1004 ( .A(n907), .B(n906), .ZN(n908) );
  XNOR2_X1 U1005 ( .A(n909), .B(n908), .ZN(n910) );
  NAND2_X1 U1006 ( .A1(n910), .A2(G14), .ZN(n917) );
  NAND2_X1 U1007 ( .A1(G319), .A2(n917), .ZN(n911) );
  NOR2_X1 U1008 ( .A1(n912), .A2(n911), .ZN(n914) );
  NOR2_X1 U1009 ( .A1(G397), .A2(G395), .ZN(n913) );
  NAND2_X1 U1010 ( .A1(n914), .A2(n913), .ZN(G225) );
  XNOR2_X1 U1011 ( .A(KEYINPUT117), .B(G225), .ZN(G308) );
  INV_X1 U1013 ( .A(G120), .ZN(G236) );
  INV_X1 U1014 ( .A(G108), .ZN(G238) );
  INV_X1 U1015 ( .A(G96), .ZN(G221) );
  INV_X1 U1016 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1017 ( .A1(n916), .A2(n915), .ZN(G325) );
  INV_X1 U1018 ( .A(G325), .ZN(G261) );
  INV_X1 U1019 ( .A(n917), .ZN(G401) );
  NAND2_X1 U1020 ( .A1(n919), .A2(n918), .ZN(n925) );
  XNOR2_X1 U1021 ( .A(G2090), .B(G162), .ZN(n920) );
  XNOR2_X1 U1022 ( .A(n920), .B(KEYINPUT118), .ZN(n921) );
  NAND2_X1 U1023 ( .A1(n922), .A2(n921), .ZN(n923) );
  XOR2_X1 U1024 ( .A(KEYINPUT51), .B(n923), .Z(n924) );
  NOR2_X1 U1025 ( .A1(n925), .A2(n924), .ZN(n929) );
  XOR2_X1 U1026 ( .A(G160), .B(G2084), .Z(n926) );
  NOR2_X1 U1027 ( .A1(n927), .A2(n926), .ZN(n928) );
  NAND2_X1 U1028 ( .A1(n929), .A2(n928), .ZN(n935) );
  XOR2_X1 U1029 ( .A(G2072), .B(n930), .Z(n932) );
  XOR2_X1 U1030 ( .A(G164), .B(G2078), .Z(n931) );
  NOR2_X1 U1031 ( .A1(n932), .A2(n931), .ZN(n933) );
  XOR2_X1 U1032 ( .A(KEYINPUT50), .B(n933), .Z(n934) );
  NOR2_X1 U1033 ( .A1(n935), .A2(n934), .ZN(n937) );
  NAND2_X1 U1034 ( .A1(n937), .A2(n936), .ZN(n938) );
  NOR2_X1 U1035 ( .A1(n939), .A2(n938), .ZN(n940) );
  XOR2_X1 U1036 ( .A(KEYINPUT52), .B(n940), .Z(n941) );
  NOR2_X1 U1037 ( .A1(KEYINPUT55), .A2(n941), .ZN(n942) );
  XNOR2_X1 U1038 ( .A(KEYINPUT119), .B(n942), .ZN(n943) );
  NAND2_X1 U1039 ( .A1(n943), .A2(G29), .ZN(n1025) );
  XOR2_X1 U1040 ( .A(n944), .B(G32), .Z(n947) );
  XOR2_X1 U1041 ( .A(n945), .B(G27), .Z(n946) );
  NOR2_X1 U1042 ( .A1(n947), .A2(n946), .ZN(n955) );
  XNOR2_X1 U1043 ( .A(G2067), .B(G26), .ZN(n949) );
  XNOR2_X1 U1044 ( .A(G33), .B(G2072), .ZN(n948) );
  NOR2_X1 U1045 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1046 ( .A1(G28), .A2(n950), .ZN(n953) );
  XOR2_X1 U1047 ( .A(KEYINPUT121), .B(G1991), .Z(n951) );
  XNOR2_X1 U1048 ( .A(G25), .B(n951), .ZN(n952) );
  NOR2_X1 U1049 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1050 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1051 ( .A(n956), .B(KEYINPUT53), .ZN(n957) );
  XNOR2_X1 U1052 ( .A(KEYINPUT122), .B(n957), .ZN(n960) );
  XOR2_X1 U1053 ( .A(G2090), .B(KEYINPUT120), .Z(n958) );
  XNOR2_X1 U1054 ( .A(G35), .B(n958), .ZN(n959) );
  NAND2_X1 U1055 ( .A1(n960), .A2(n959), .ZN(n963) );
  XNOR2_X1 U1056 ( .A(G34), .B(G2084), .ZN(n961) );
  XNOR2_X1 U1057 ( .A(KEYINPUT54), .B(n961), .ZN(n962) );
  NOR2_X1 U1058 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1059 ( .A(KEYINPUT55), .B(n964), .ZN(n966) );
  INV_X1 U1060 ( .A(G29), .ZN(n965) );
  NAND2_X1 U1061 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1062 ( .A1(n967), .A2(G11), .ZN(n1023) );
  XNOR2_X1 U1063 ( .A(G16), .B(KEYINPUT56), .ZN(n992) );
  XOR2_X1 U1064 ( .A(G168), .B(G1966), .Z(n968) );
  NOR2_X1 U1065 ( .A1(n969), .A2(n968), .ZN(n970) );
  XOR2_X1 U1066 ( .A(KEYINPUT57), .B(n970), .Z(n990) );
  XNOR2_X1 U1067 ( .A(G301), .B(G1961), .ZN(n973) );
  XNOR2_X1 U1068 ( .A(n971), .B(G1341), .ZN(n972) );
  NOR2_X1 U1069 ( .A1(n973), .A2(n972), .ZN(n985) );
  NAND2_X1 U1070 ( .A1(G1971), .A2(G303), .ZN(n974) );
  NAND2_X1 U1071 ( .A1(n975), .A2(n974), .ZN(n976) );
  NOR2_X1 U1072 ( .A1(n977), .A2(n976), .ZN(n980) );
  XNOR2_X1 U1073 ( .A(G1956), .B(KEYINPUT123), .ZN(n978) );
  XNOR2_X1 U1074 ( .A(n978), .B(G299), .ZN(n979) );
  NAND2_X1 U1075 ( .A1(n980), .A2(n979), .ZN(n981) );
  NOR2_X1 U1076 ( .A1(n982), .A2(n981), .ZN(n983) );
  XNOR2_X1 U1077 ( .A(n983), .B(KEYINPUT124), .ZN(n984) );
  NAND2_X1 U1078 ( .A1(n985), .A2(n984), .ZN(n988) );
  XOR2_X1 U1079 ( .A(G1348), .B(n986), .Z(n987) );
  NOR2_X1 U1080 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1081 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1082 ( .A1(n992), .A2(n991), .ZN(n1021) );
  INV_X1 U1083 ( .A(G16), .ZN(n1019) );
  XOR2_X1 U1084 ( .A(KEYINPUT126), .B(G4), .Z(n994) );
  XNOR2_X1 U1085 ( .A(G1348), .B(KEYINPUT59), .ZN(n993) );
  XNOR2_X1 U1086 ( .A(n994), .B(n993), .ZN(n997) );
  XOR2_X1 U1087 ( .A(KEYINPUT125), .B(G1341), .Z(n995) );
  XNOR2_X1 U1088 ( .A(G19), .B(n995), .ZN(n996) );
  NOR2_X1 U1089 ( .A1(n997), .A2(n996), .ZN(n1001) );
  XNOR2_X1 U1090 ( .A(G1956), .B(G20), .ZN(n999) );
  XNOR2_X1 U1091 ( .A(G6), .B(G1981), .ZN(n998) );
  NOR2_X1 U1092 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1093 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1094 ( .A(n1002), .B(KEYINPUT127), .ZN(n1003) );
  XNOR2_X1 U1095 ( .A(KEYINPUT60), .B(n1003), .ZN(n1011) );
  XOR2_X1 U1096 ( .A(G1986), .B(G24), .Z(n1006) );
  XNOR2_X1 U1097 ( .A(n1004), .B(G22), .ZN(n1005) );
  NAND2_X1 U1098 ( .A1(n1006), .A2(n1005), .ZN(n1008) );
  XNOR2_X1 U1099 ( .A(G23), .B(G1976), .ZN(n1007) );
  NOR2_X1 U1100 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1101 ( .A(KEYINPUT58), .B(n1009), .ZN(n1010) );
  NAND2_X1 U1102 ( .A1(n1011), .A2(n1010), .ZN(n1016) );
  XOR2_X1 U1103 ( .A(G1966), .B(G21), .Z(n1014) );
  XNOR2_X1 U1104 ( .A(n1012), .B(G5), .ZN(n1013) );
  NAND2_X1 U1105 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NOR2_X1 U1106 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1107 ( .A(KEYINPUT61), .B(n1017), .ZN(n1018) );
  NAND2_X1 U1108 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1109 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NOR2_X1 U1110 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1111 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XOR2_X1 U1112 ( .A(KEYINPUT62), .B(n1026), .Z(G311) );
  INV_X1 U1113 ( .A(G311), .ZN(G150) );
endmodule

