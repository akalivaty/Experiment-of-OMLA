

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764;

  AND2_X1 U368 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U369 ( .A(n606), .B(KEYINPUT103), .ZN(n683) );
  OR2_X1 U370 ( .A1(n542), .A2(n545), .ZN(n541) );
  XNOR2_X1 U371 ( .A(n612), .B(n442), .ZN(n597) );
  AND2_X1 U372 ( .A1(n408), .A2(n407), .ZN(n406) );
  XNOR2_X1 U373 ( .A(n737), .B(n437), .ZN(n671) );
  BUF_X1 U374 ( .A(G113), .Z(n347) );
  XNOR2_X1 U375 ( .A(n506), .B(n465), .ZN(n750) );
  XNOR2_X1 U376 ( .A(G110), .B(KEYINPUT16), .ZN(n430) );
  INV_X1 U377 ( .A(G146), .ZN(n401) );
  INV_X2 U378 ( .A(G953), .ZN(n742) );
  XNOR2_X2 U379 ( .A(n346), .B(KEYINPUT69), .ZN(n599) );
  NAND2_X1 U380 ( .A1(n579), .A2(n578), .ZN(n346) );
  NAND2_X2 U381 ( .A1(n415), .A2(n414), .ZN(n423) );
  BUF_X2 U382 ( .A(n693), .Z(n371) );
  NAND2_X2 U383 ( .A1(n348), .A2(n602), .ZN(n529) );
  XNOR2_X2 U384 ( .A(n499), .B(n498), .ZN(n348) );
  XNOR2_X1 U385 ( .A(G137), .B(n347), .ZN(n486) );
  NOR2_X1 U386 ( .A1(G953), .A2(G237), .ZN(n509) );
  XOR2_X1 U387 ( .A(n648), .B(n647), .Z(n349) );
  AND2_X2 U388 ( .A1(n416), .A2(n418), .ZN(n415) );
  XNOR2_X2 U389 ( .A(n453), .B(n452), .ZN(n523) );
  NOR2_X1 U390 ( .A1(n710), .A2(n707), .ZN(n592) );
  AND2_X1 U391 ( .A1(n390), .A2(n389), .ZN(n388) );
  NAND2_X1 U392 ( .A1(n413), .A2(n556), .ZN(n661) );
  AND2_X1 U393 ( .A1(n652), .A2(n393), .ZN(n355) );
  AND2_X1 U394 ( .A1(n557), .A2(n691), .ZN(n555) );
  XNOR2_X1 U395 ( .A(n550), .B(n549), .ZN(n557) );
  NAND2_X1 U396 ( .A1(n532), .A2(n533), .ZN(n372) );
  NAND2_X1 U397 ( .A1(n557), .A2(n350), .ZN(n652) );
  AND2_X1 U398 ( .A1(n691), .A2(n552), .ZN(n350) );
  OR2_X1 U399 ( .A1(n637), .A2(n417), .ZN(n414) );
  BUF_X1 U400 ( .A(n662), .Z(n351) );
  XNOR2_X2 U401 ( .A(n751), .B(G146), .ZN(n491) );
  OR2_X1 U402 ( .A1(n538), .A2(n537), .ZN(n673) );
  XNOR2_X2 U403 ( .A(n463), .B(n400), .ZN(n506) );
  BUF_X1 U404 ( .A(n548), .Z(n533) );
  XNOR2_X2 U405 ( .A(n436), .B(n435), .ZN(n737) );
  OR2_X2 U406 ( .A1(n648), .A2(G902), .ZN(n397) );
  XNOR2_X2 U407 ( .A(n523), .B(n454), .ZN(n751) );
  NAND2_X1 U408 ( .A1(n661), .A2(n655), .ZN(n562) );
  XNOR2_X1 U409 ( .A(KEYINPUT4), .B(G131), .ZN(n454) );
  INV_X1 U410 ( .A(KEYINPUT10), .ZN(n400) );
  XNOR2_X1 U411 ( .A(n481), .B(n480), .ZN(n693) );
  INV_X1 U412 ( .A(KEYINPUT100), .ZN(n394) );
  INV_X1 U413 ( .A(n544), .ZN(n391) );
  NOR2_X1 U414 ( .A1(n761), .A2(n763), .ZN(n596) );
  INV_X1 U415 ( .A(KEYINPUT11), .ZN(n378) );
  XOR2_X1 U416 ( .A(KEYINPUT95), .B(KEYINPUT12), .Z(n501) );
  XNOR2_X1 U417 ( .A(G902), .B(KEYINPUT15), .ZN(n635) );
  NOR2_X1 U418 ( .A1(n635), .A2(KEYINPUT64), .ZN(n422) );
  NAND2_X1 U419 ( .A1(n411), .A2(n421), .ZN(n420) );
  NAND2_X1 U420 ( .A1(n636), .A2(KEYINPUT2), .ZN(n421) );
  OR2_X1 U421 ( .A1(n641), .A2(G902), .ZN(n492) );
  XNOR2_X1 U422 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U423 ( .A(n491), .B(n461), .ZN(n648) );
  XNOR2_X1 U424 ( .A(G107), .B(G104), .ZN(n457) );
  XNOR2_X1 U425 ( .A(n581), .B(n580), .ZN(n625) );
  XNOR2_X1 U426 ( .A(n476), .B(n475), .ZN(n663) );
  XNOR2_X1 U427 ( .A(n750), .B(n468), .ZN(n476) );
  NAND2_X1 U428 ( .A1(n709), .A2(n394), .ZN(n393) );
  NOR2_X1 U429 ( .A1(n618), .A2(n617), .ZN(n619) );
  NAND2_X1 U430 ( .A1(n384), .A2(n387), .ZN(n383) );
  AND2_X1 U431 ( .A1(n386), .A2(n385), .ZN(n384) );
  NAND2_X1 U432 ( .A1(G237), .A2(G234), .ZN(n443) );
  XNOR2_X1 U433 ( .A(n504), .B(n377), .ZN(n505) );
  XNOR2_X1 U434 ( .A(n503), .B(n378), .ZN(n377) );
  XNOR2_X1 U435 ( .A(KEYINPUT93), .B(KEYINPUT94), .ZN(n500) );
  XNOR2_X1 U436 ( .A(G140), .B(G122), .ZN(n507) );
  XOR2_X1 U437 ( .A(G131), .B(G143), .Z(n508) );
  XNOR2_X1 U438 ( .A(G101), .B(G110), .ZN(n456) );
  XNOR2_X1 U439 ( .A(KEYINPUT66), .B(G140), .ZN(n459) );
  XNOR2_X1 U440 ( .A(KEYINPUT4), .B(KEYINPUT83), .ZN(n427) );
  INV_X1 U441 ( .A(G237), .ZN(n438) );
  AND2_X1 U442 ( .A1(n409), .A2(n381), .ZN(n407) );
  XNOR2_X1 U443 ( .A(n369), .B(n571), .ZN(n577) );
  NAND2_X1 U444 ( .A1(n697), .A2(n381), .ZN(n369) );
  NAND2_X1 U445 ( .A1(n411), .A2(n439), .ZN(n409) );
  NAND2_X1 U446 ( .A1(n399), .A2(n398), .ZN(n690) );
  INV_X1 U447 ( .A(n694), .ZN(n398) );
  INV_X1 U448 ( .A(n693), .ZN(n399) );
  XOR2_X1 U449 ( .A(KEYINPUT71), .B(KEYINPUT88), .Z(n467) );
  XNOR2_X1 U450 ( .A(KEYINPUT76), .B(KEYINPUT89), .ZN(n470) );
  INV_X1 U451 ( .A(G134), .ZN(n452) );
  NAND2_X1 U452 ( .A1(KEYINPUT64), .A2(n725), .ZN(n417) );
  NAND2_X1 U453 ( .A1(n420), .A2(n419), .ZN(n418) );
  NAND2_X1 U454 ( .A1(n635), .A2(n636), .ZN(n419) );
  AND2_X1 U455 ( .A1(n683), .A2(n611), .ZN(n629) );
  INV_X1 U456 ( .A(KEYINPUT1), .ZN(n396) );
  XNOR2_X1 U457 ( .A(n583), .B(n582), .ZN(n761) );
  NOR2_X1 U458 ( .A1(n625), .A2(n606), .ZN(n583) );
  XNOR2_X1 U459 ( .A(n555), .B(KEYINPUT102), .ZN(n413) );
  INV_X1 U460 ( .A(KEYINPUT122), .ZN(n374) );
  INV_X1 U461 ( .A(KEYINPUT60), .ZN(n365) );
  INV_X1 U462 ( .A(KEYINPUT56), .ZN(n367) );
  OR2_X1 U463 ( .A1(n411), .A2(n439), .ZN(n352) );
  AND2_X1 U464 ( .A1(n655), .A2(n560), .ZN(n353) );
  NOR2_X1 U465 ( .A1(n713), .A2(n719), .ZN(n354) );
  AND2_X1 U466 ( .A1(n661), .A2(n353), .ZN(n356) );
  AND2_X1 U467 ( .A1(n543), .A2(KEYINPUT100), .ZN(n357) );
  NOR2_X1 U468 ( .A1(n559), .A2(n558), .ZN(n358) );
  AND2_X1 U469 ( .A1(n408), .A2(n409), .ZN(n359) );
  XOR2_X1 U470 ( .A(n451), .B(KEYINPUT0), .Z(n360) );
  INV_X1 U471 ( .A(n635), .ZN(n411) );
  XOR2_X1 U472 ( .A(n666), .B(KEYINPUT59), .Z(n361) );
  XOR2_X1 U473 ( .A(n671), .B(n670), .Z(n362) );
  XOR2_X1 U474 ( .A(n641), .B(n640), .Z(n363) );
  AND2_X1 U475 ( .A1(n394), .A2(KEYINPUT101), .ZN(n364) );
  XNOR2_X1 U476 ( .A(n649), .B(n349), .ZN(n650) );
  XNOR2_X1 U477 ( .A(n642), .B(n363), .ZN(n645) );
  INV_X1 U478 ( .A(n626), .ZN(n381) );
  XNOR2_X1 U479 ( .A(n366), .B(n365), .ZN(G60) );
  NAND2_X1 U480 ( .A1(n379), .A2(n644), .ZN(n366) );
  XNOR2_X1 U481 ( .A(n368), .B(n367), .ZN(G51) );
  NAND2_X1 U482 ( .A1(n380), .A2(n644), .ZN(n368) );
  NAND2_X1 U483 ( .A1(n406), .A2(n410), .ZN(n373) );
  NAND2_X1 U484 ( .A1(n392), .A2(KEYINPUT101), .ZN(n390) );
  NAND2_X1 U485 ( .A1(n355), .A2(n395), .ZN(n392) );
  XNOR2_X2 U486 ( .A(n531), .B(KEYINPUT92), .ZN(n702) );
  NAND2_X1 U487 ( .A1(n370), .A2(n553), .ZN(n554) );
  NAND2_X1 U488 ( .A1(n388), .A2(n383), .ZN(n370) );
  XNOR2_X2 U489 ( .A(n372), .B(n534), .ZN(n656) );
  NOR2_X1 U490 ( .A1(n622), .A2(n621), .ZN(n624) );
  XNOR2_X2 U491 ( .A(n373), .B(n441), .ZN(n612) );
  XNOR2_X1 U492 ( .A(n375), .B(n374), .ZN(G66) );
  NAND2_X1 U493 ( .A1(n665), .A2(n644), .ZN(n375) );
  XNOR2_X2 U494 ( .A(n376), .B(n360), .ZN(n548) );
  NOR2_X2 U495 ( .A1(n597), .A2(n450), .ZN(n376) );
  NOR2_X1 U496 ( .A1(n634), .A2(n633), .ZN(n752) );
  XNOR2_X1 U497 ( .A(n513), .B(n512), .ZN(n666) );
  XNOR2_X1 U498 ( .A(n667), .B(n361), .ZN(n379) );
  XNOR2_X1 U499 ( .A(n672), .B(n362), .ZN(n380) );
  INV_X1 U500 ( .A(KEYINPUT101), .ZN(n385) );
  NAND2_X1 U501 ( .A1(n391), .A2(n394), .ZN(n386) );
  INV_X1 U502 ( .A(n392), .ZN(n387) );
  NAND2_X1 U503 ( .A1(n391), .A2(n364), .ZN(n389) );
  NAND2_X1 U504 ( .A1(n544), .A2(n357), .ZN(n395) );
  XNOR2_X2 U505 ( .A(n589), .B(n396), .ZN(n627) );
  XNOR2_X2 U506 ( .A(n397), .B(n462), .ZN(n589) );
  XNOR2_X2 U507 ( .A(n401), .B(G125), .ZN(n463) );
  NAND2_X1 U508 ( .A1(n402), .A2(n356), .ZN(n404) );
  NAND2_X1 U509 ( .A1(n403), .A2(n405), .ZN(n402) );
  INV_X1 U510 ( .A(n662), .ZN(n403) );
  NAND2_X1 U511 ( .A1(n404), .A2(n563), .ZN(n565) );
  INV_X1 U512 ( .A(KEYINPUT44), .ZN(n405) );
  XNOR2_X2 U513 ( .A(n529), .B(KEYINPUT35), .ZN(n662) );
  NAND2_X1 U514 ( .A1(n410), .A2(n359), .ZN(n631) );
  OR2_X2 U515 ( .A1(n671), .A2(n352), .ZN(n408) );
  NAND2_X1 U516 ( .A1(n671), .A2(n439), .ZN(n410) );
  NOR2_X2 U517 ( .A1(n724), .A2(n725), .ZN(n638) );
  XNOR2_X2 U518 ( .A(n412), .B(KEYINPUT32), .ZN(n655) );
  NAND2_X1 U519 ( .A1(n557), .A2(n358), .ZN(n412) );
  NAND2_X1 U520 ( .A1(n637), .A2(n422), .ZN(n416) );
  NOR2_X4 U521 ( .A1(n423), .A2(n638), .ZN(n732) );
  INV_X1 U522 ( .A(KEYINPUT46), .ZN(n595) );
  BUF_X1 U523 ( .A(n502), .Z(n503) );
  INV_X1 U524 ( .A(n584), .ZN(n576) );
  INV_X1 U525 ( .A(KEYINPUT48), .ZN(n623) );
  AND2_X1 U526 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U527 ( .A(n491), .B(n490), .ZN(n641) );
  INV_X1 U528 ( .A(KEYINPUT64), .ZN(n636) );
  INV_X1 U529 ( .A(n736), .ZN(n644) );
  NAND2_X1 U530 ( .A1(n742), .A2(G224), .ZN(n425) );
  XNOR2_X1 U531 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n424) );
  XNOR2_X1 U532 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U533 ( .A(n426), .B(n463), .ZN(n429) );
  XNOR2_X2 U534 ( .A(G143), .B(G128), .ZN(n453) );
  XNOR2_X1 U535 ( .A(n453), .B(n427), .ZN(n428) );
  XNOR2_X1 U536 ( .A(n429), .B(n428), .ZN(n437) );
  XNOR2_X2 U537 ( .A(G104), .B(G113), .ZN(n502) );
  XNOR2_X1 U538 ( .A(n502), .B(n430), .ZN(n432) );
  INV_X1 U539 ( .A(G107), .ZN(n431) );
  XNOR2_X1 U540 ( .A(n431), .B(G122), .ZN(n516) );
  XNOR2_X1 U541 ( .A(n432), .B(n516), .ZN(n436) );
  XNOR2_X1 U542 ( .A(G101), .B(G116), .ZN(n434) );
  XNOR2_X1 U543 ( .A(KEYINPUT3), .B(G119), .ZN(n433) );
  XNOR2_X1 U544 ( .A(n434), .B(n433), .ZN(n489) );
  INV_X1 U545 ( .A(n489), .ZN(n435) );
  INV_X1 U546 ( .A(G902), .ZN(n526) );
  NAND2_X1 U547 ( .A1(n526), .A2(n438), .ZN(n440) );
  NAND2_X1 U548 ( .A1(n440), .A2(G210), .ZN(n439) );
  AND2_X1 U549 ( .A1(n440), .A2(G214), .ZN(n626) );
  INV_X1 U550 ( .A(KEYINPUT80), .ZN(n441) );
  XNOR2_X1 U551 ( .A(KEYINPUT70), .B(KEYINPUT19), .ZN(n442) );
  XNOR2_X1 U552 ( .A(n443), .B(KEYINPUT84), .ZN(n444) );
  XNOR2_X1 U553 ( .A(KEYINPUT14), .B(n444), .ZN(n445) );
  NAND2_X1 U554 ( .A1(G952), .A2(n445), .ZN(n717) );
  NOR2_X1 U555 ( .A1(n717), .A2(G953), .ZN(n574) );
  INV_X1 U556 ( .A(n574), .ZN(n449) );
  NAND2_X1 U557 ( .A1(n445), .A2(G902), .ZN(n446) );
  XNOR2_X1 U558 ( .A(n446), .B(KEYINPUT85), .ZN(n572) );
  NOR2_X1 U559 ( .A1(G898), .A2(n742), .ZN(n738) );
  NAND2_X1 U560 ( .A1(n572), .A2(n738), .ZN(n447) );
  XNOR2_X1 U561 ( .A(n447), .B(KEYINPUT86), .ZN(n448) );
  AND2_X1 U562 ( .A1(n449), .A2(n448), .ZN(n450) );
  INV_X1 U563 ( .A(KEYINPUT82), .ZN(n451) );
  XNOR2_X1 U564 ( .A(n548), .B(KEYINPUT87), .ZN(n538) );
  NAND2_X1 U565 ( .A1(n742), .A2(G227), .ZN(n455) );
  XNOR2_X1 U566 ( .A(n456), .B(n455), .ZN(n458) );
  XNOR2_X1 U567 ( .A(n458), .B(n457), .ZN(n460) );
  XNOR2_X1 U568 ( .A(n459), .B(G137), .ZN(n464) );
  XNOR2_X1 U569 ( .A(n460), .B(n464), .ZN(n461) );
  INV_X1 U570 ( .A(G469), .ZN(n462) );
  INV_X1 U571 ( .A(n464), .ZN(n465) );
  XNOR2_X1 U572 ( .A(G128), .B(KEYINPUT23), .ZN(n466) );
  XNOR2_X1 U573 ( .A(n467), .B(n466), .ZN(n468) );
  NAND2_X1 U574 ( .A1(G234), .A2(n742), .ZN(n469) );
  XOR2_X1 U575 ( .A(KEYINPUT8), .B(n469), .Z(n517) );
  AND2_X1 U576 ( .A1(n517), .A2(G221), .ZN(n474) );
  XOR2_X1 U577 ( .A(G119), .B(G110), .Z(n471) );
  XNOR2_X1 U578 ( .A(n471), .B(n470), .ZN(n472) );
  XOR2_X1 U579 ( .A(n472), .B(KEYINPUT24), .Z(n473) );
  XNOR2_X1 U580 ( .A(n474), .B(n473), .ZN(n475) );
  NAND2_X1 U581 ( .A1(n663), .A2(n526), .ZN(n481) );
  NAND2_X1 U582 ( .A1(n635), .A2(G234), .ZN(n478) );
  XNOR2_X1 U583 ( .A(KEYINPUT90), .B(KEYINPUT20), .ZN(n477) );
  XNOR2_X1 U584 ( .A(n478), .B(n477), .ZN(n482) );
  NAND2_X1 U585 ( .A1(G217), .A2(n482), .ZN(n479) );
  XNOR2_X1 U586 ( .A(n479), .B(KEYINPUT25), .ZN(n480) );
  NAND2_X1 U587 ( .A1(n482), .A2(G221), .ZN(n483) );
  XNOR2_X1 U588 ( .A(n483), .B(KEYINPUT21), .ZN(n694) );
  INV_X1 U589 ( .A(n690), .ZN(n484) );
  AND2_X2 U590 ( .A1(n627), .A2(n484), .ZN(n530) );
  NAND2_X1 U591 ( .A1(n509), .A2(G210), .ZN(n485) );
  XNOR2_X1 U592 ( .A(n485), .B(KEYINPUT5), .ZN(n487) );
  XNOR2_X1 U593 ( .A(n487), .B(n486), .ZN(n488) );
  XOR2_X1 U594 ( .A(n488), .B(n489), .Z(n490) );
  XNOR2_X2 U595 ( .A(n492), .B(G472), .ZN(n697) );
  XNOR2_X1 U596 ( .A(n697), .B(KEYINPUT6), .ZN(n608) );
  INV_X1 U597 ( .A(n608), .ZN(n493) );
  NAND2_X1 U598 ( .A1(n530), .A2(n493), .ZN(n495) );
  XNOR2_X1 U599 ( .A(KEYINPUT67), .B(KEYINPUT33), .ZN(n494) );
  XNOR2_X1 U600 ( .A(n495), .B(n494), .ZN(n719) );
  OR2_X2 U601 ( .A1(n538), .A2(n719), .ZN(n499) );
  XNOR2_X1 U602 ( .A(KEYINPUT72), .B(KEYINPUT34), .ZN(n497) );
  INV_X1 U603 ( .A(KEYINPUT68), .ZN(n496) );
  XNOR2_X1 U604 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U605 ( .A(n501), .B(n500), .ZN(n504) );
  XOR2_X1 U606 ( .A(n506), .B(n505), .Z(n513) );
  XNOR2_X1 U607 ( .A(n508), .B(n507), .ZN(n511) );
  NAND2_X1 U608 ( .A1(n509), .A2(G214), .ZN(n510) );
  NAND2_X1 U609 ( .A1(n666), .A2(n526), .ZN(n515) );
  XOR2_X1 U610 ( .A(KEYINPUT13), .B(G475), .Z(n514) );
  XNOR2_X1 U611 ( .A(n515), .B(n514), .ZN(n546) );
  XOR2_X1 U612 ( .A(n516), .B(KEYINPUT98), .Z(n519) );
  NAND2_X1 U613 ( .A1(G217), .A2(n517), .ZN(n518) );
  XNOR2_X1 U614 ( .A(n519), .B(n518), .ZN(n525) );
  XOR2_X1 U615 ( .A(KEYINPUT9), .B(KEYINPUT97), .Z(n521) );
  XNOR2_X1 U616 ( .A(G116), .B(KEYINPUT7), .ZN(n520) );
  XNOR2_X1 U617 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U618 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U619 ( .A(n525), .B(n524), .ZN(n734) );
  NAND2_X1 U620 ( .A1(n734), .A2(n526), .ZN(n527) );
  XNOR2_X1 U621 ( .A(n527), .B(G478), .ZN(n545) );
  AND2_X1 U622 ( .A1(n546), .A2(n545), .ZN(n602) );
  NAND2_X1 U623 ( .A1(n662), .A2(KEYINPUT44), .ZN(n553) );
  NAND2_X1 U624 ( .A1(n530), .A2(n697), .ZN(n531) );
  INV_X1 U625 ( .A(n702), .ZN(n532) );
  INV_X1 U626 ( .A(KEYINPUT31), .ZN(n534) );
  NOR2_X1 U627 ( .A1(n690), .A2(n589), .ZN(n536) );
  INV_X1 U628 ( .A(KEYINPUT91), .ZN(n535) );
  XNOR2_X1 U629 ( .A(n536), .B(n535), .ZN(n579) );
  INV_X1 U630 ( .A(n697), .ZN(n586) );
  NAND2_X1 U631 ( .A1(n579), .A2(n586), .ZN(n537) );
  NAND2_X1 U632 ( .A1(n656), .A2(n673), .ZN(n544) );
  INV_X1 U633 ( .A(KEYINPUT96), .ZN(n539) );
  XNOR2_X1 U634 ( .A(n546), .B(n539), .ZN(n542) );
  INV_X1 U635 ( .A(KEYINPUT99), .ZN(n540) );
  XNOR2_X2 U636 ( .A(n541), .B(n540), .ZN(n606) );
  NAND2_X1 U637 ( .A1(n542), .A2(n545), .ZN(n677) );
  AND2_X1 U638 ( .A1(n606), .A2(n677), .ZN(n709) );
  INV_X1 U639 ( .A(n709), .ZN(n543) );
  OR2_X1 U640 ( .A1(n546), .A2(n545), .ZN(n707) );
  NOR2_X1 U641 ( .A1(n707), .A2(n694), .ZN(n547) );
  NAND2_X1 U642 ( .A1(n548), .A2(n547), .ZN(n550) );
  INV_X1 U643 ( .A(KEYINPUT22), .ZN(n549) );
  INV_X1 U644 ( .A(n627), .ZN(n691) );
  INV_X1 U645 ( .A(n371), .ZN(n551) );
  AND2_X1 U646 ( .A1(n608), .A2(n551), .ZN(n552) );
  XNOR2_X1 U647 ( .A(n554), .B(KEYINPUT79), .ZN(n567) );
  AND2_X1 U648 ( .A1(n586), .A2(n371), .ZN(n556) );
  XNOR2_X1 U649 ( .A(n608), .B(KEYINPUT73), .ZN(n559) );
  NAND2_X1 U650 ( .A1(n627), .A2(n371), .ZN(n558) );
  INV_X1 U651 ( .A(KEYINPUT65), .ZN(n560) );
  NAND2_X1 U652 ( .A1(n560), .A2(KEYINPUT44), .ZN(n561) );
  NAND2_X1 U653 ( .A1(n562), .A2(n561), .ZN(n563) );
  NAND2_X1 U654 ( .A1(n405), .A2(KEYINPUT65), .ZN(n564) );
  NAND2_X1 U655 ( .A1(n567), .A2(n566), .ZN(n570) );
  INV_X1 U656 ( .A(KEYINPUT77), .ZN(n568) );
  XNOR2_X1 U657 ( .A(n568), .B(KEYINPUT45), .ZN(n569) );
  XNOR2_X1 U658 ( .A(n570), .B(n569), .ZN(n741) );
  XNOR2_X1 U659 ( .A(KEYINPUT30), .B(KEYINPUT105), .ZN(n571) );
  NAND2_X1 U660 ( .A1(G953), .A2(n572), .ZN(n573) );
  NOR2_X1 U661 ( .A1(G900), .A2(n573), .ZN(n575) );
  NOR2_X1 U662 ( .A1(n575), .A2(n574), .ZN(n584) );
  XNOR2_X1 U663 ( .A(n631), .B(KEYINPUT38), .ZN(n705) );
  NAND2_X1 U664 ( .A1(n599), .A2(n705), .ZN(n581) );
  XOR2_X1 U665 ( .A(KEYINPUT78), .B(KEYINPUT39), .Z(n580) );
  XNOR2_X1 U666 ( .A(KEYINPUT108), .B(KEYINPUT40), .ZN(n582) );
  NOR2_X1 U667 ( .A1(n584), .A2(n694), .ZN(n585) );
  NAND2_X1 U668 ( .A1(n371), .A2(n585), .ZN(n607) );
  OR2_X1 U669 ( .A1(n607), .A2(n586), .ZN(n588) );
  INV_X1 U670 ( .A(KEYINPUT28), .ZN(n587) );
  XNOR2_X1 U671 ( .A(n588), .B(n587), .ZN(n591) );
  XNOR2_X1 U672 ( .A(n589), .B(KEYINPUT107), .ZN(n590) );
  NAND2_X1 U673 ( .A1(n591), .A2(n590), .ZN(n598) );
  NAND2_X1 U674 ( .A1(n705), .A2(n381), .ZN(n710) );
  XNOR2_X1 U675 ( .A(KEYINPUT41), .B(n592), .ZN(n720) );
  OR2_X1 U676 ( .A1(n598), .A2(n720), .ZN(n593) );
  XNOR2_X1 U677 ( .A(n593), .B(KEYINPUT42), .ZN(n594) );
  XNOR2_X1 U678 ( .A(KEYINPUT109), .B(n594), .ZN(n763) );
  XNOR2_X1 U679 ( .A(n596), .B(n595), .ZN(n622) );
  OR2_X1 U680 ( .A1(n597), .A2(n598), .ZN(n678) );
  OR2_X1 U681 ( .A1(n709), .A2(n678), .ZN(n616) );
  NAND2_X1 U682 ( .A1(n616), .A2(KEYINPUT47), .ZN(n604) );
  INV_X1 U683 ( .A(n599), .ZN(n600) );
  NOR2_X1 U684 ( .A1(n631), .A2(n600), .ZN(n601) );
  NAND2_X1 U685 ( .A1(n602), .A2(n601), .ZN(n603) );
  XNOR2_X1 U686 ( .A(n603), .B(KEYINPUT106), .ZN(n762) );
  NAND2_X1 U687 ( .A1(n604), .A2(n762), .ZN(n605) );
  XNOR2_X1 U688 ( .A(n605), .B(KEYINPUT75), .ZN(n620) );
  OR2_X1 U689 ( .A1(n608), .A2(n607), .ZN(n610) );
  INV_X1 U690 ( .A(KEYINPUT104), .ZN(n609) );
  XNOR2_X1 U691 ( .A(n610), .B(n609), .ZN(n611) );
  NAND2_X1 U692 ( .A1(n629), .A2(n612), .ZN(n614) );
  XOR2_X1 U693 ( .A(KEYINPUT36), .B(KEYINPUT110), .Z(n613) );
  XNOR2_X1 U694 ( .A(n614), .B(n613), .ZN(n615) );
  NAND2_X1 U695 ( .A1(n615), .A2(n627), .ZN(n687) );
  INV_X1 U696 ( .A(n687), .ZN(n618) );
  NOR2_X1 U697 ( .A1(n616), .A2(KEYINPUT47), .ZN(n617) );
  NAND2_X1 U698 ( .A1(n620), .A2(n619), .ZN(n621) );
  XNOR2_X1 U699 ( .A(n624), .B(n623), .ZN(n634) );
  NOR2_X1 U700 ( .A1(n625), .A2(n677), .ZN(n689) );
  NOR2_X1 U701 ( .A1(n627), .A2(n626), .ZN(n628) );
  NAND2_X1 U702 ( .A1(n629), .A2(n628), .ZN(n630) );
  XNOR2_X1 U703 ( .A(n630), .B(KEYINPUT43), .ZN(n632) );
  AND2_X1 U704 ( .A1(n632), .A2(n631), .ZN(n659) );
  OR2_X1 U705 ( .A1(n689), .A2(n659), .ZN(n633) );
  AND2_X2 U706 ( .A1(n741), .A2(n752), .ZN(n637) );
  INV_X1 U707 ( .A(n637), .ZN(n724) );
  INV_X1 U708 ( .A(KEYINPUT2), .ZN(n725) );
  NAND2_X1 U709 ( .A1(n732), .A2(G472), .ZN(n642) );
  XOR2_X1 U710 ( .A(KEYINPUT111), .B(KEYINPUT112), .Z(n639) );
  XNOR2_X1 U711 ( .A(n639), .B(KEYINPUT62), .ZN(n640) );
  INV_X1 U712 ( .A(G952), .ZN(n643) );
  AND2_X1 U713 ( .A1(n643), .A2(G953), .ZN(n736) );
  NAND2_X1 U714 ( .A1(n645), .A2(n644), .ZN(n646) );
  XNOR2_X1 U715 ( .A(n646), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U716 ( .A1(n732), .A2(G469), .ZN(n649) );
  XOR2_X1 U717 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n647) );
  NAND2_X1 U718 ( .A1(n650), .A2(n644), .ZN(n651) );
  XNOR2_X1 U719 ( .A(n651), .B(KEYINPUT121), .ZN(G54) );
  XNOR2_X1 U720 ( .A(n652), .B(G101), .ZN(G3) );
  INV_X1 U721 ( .A(n683), .ZN(n657) );
  NOR2_X1 U722 ( .A1(n657), .A2(n673), .ZN(n653) );
  XOR2_X1 U723 ( .A(G104), .B(n653), .Z(G6) );
  NOR2_X1 U724 ( .A1(n656), .A2(n677), .ZN(n654) );
  XOR2_X1 U725 ( .A(G116), .B(n654), .Z(G18) );
  XNOR2_X1 U726 ( .A(n655), .B(G119), .ZN(G21) );
  NOR2_X1 U727 ( .A1(n657), .A2(n656), .ZN(n658) );
  XOR2_X1 U728 ( .A(n347), .B(n658), .Z(G15) );
  XOR2_X1 U729 ( .A(G140), .B(n659), .Z(G42) );
  XOR2_X1 U730 ( .A(G110), .B(KEYINPUT113), .Z(n660) );
  XNOR2_X1 U731 ( .A(n661), .B(n660), .ZN(G12) );
  XOR2_X1 U732 ( .A(G122), .B(n351), .Z(G24) );
  NAND2_X1 U733 ( .A1(n732), .A2(G217), .ZN(n664) );
  XNOR2_X1 U734 ( .A(n664), .B(n663), .ZN(n665) );
  NAND2_X1 U735 ( .A1(n732), .A2(G475), .ZN(n667) );
  NAND2_X1 U736 ( .A1(n732), .A2(G210), .ZN(n672) );
  XOR2_X1 U737 ( .A(KEYINPUT55), .B(KEYINPUT81), .Z(n669) );
  XNOR2_X1 U738 ( .A(KEYINPUT54), .B(KEYINPUT120), .ZN(n668) );
  XOR2_X1 U739 ( .A(n669), .B(n668), .Z(n670) );
  NOR2_X1 U740 ( .A1(n673), .A2(n677), .ZN(n675) );
  XNOR2_X1 U741 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n674) );
  XNOR2_X1 U742 ( .A(n675), .B(n674), .ZN(n676) );
  XNOR2_X1 U743 ( .A(G107), .B(n676), .ZN(G9) );
  XOR2_X1 U744 ( .A(G128), .B(KEYINPUT29), .Z(n681) );
  INV_X1 U745 ( .A(n677), .ZN(n679) );
  INV_X1 U746 ( .A(n678), .ZN(n682) );
  NAND2_X1 U747 ( .A1(n679), .A2(n682), .ZN(n680) );
  XNOR2_X1 U748 ( .A(n681), .B(n680), .ZN(G30) );
  NAND2_X1 U749 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X1 U750 ( .A(n684), .B(KEYINPUT114), .ZN(n685) );
  XNOR2_X1 U751 ( .A(G146), .B(n685), .ZN(G48) );
  INV_X1 U752 ( .A(G125), .ZN(n686) );
  XNOR2_X1 U753 ( .A(n687), .B(n686), .ZN(n688) );
  XNOR2_X1 U754 ( .A(n688), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U755 ( .A(G134), .B(n689), .Z(G36) );
  NAND2_X1 U756 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U757 ( .A(n692), .B(KEYINPUT50), .ZN(n700) );
  XOR2_X1 U758 ( .A(KEYINPUT115), .B(KEYINPUT49), .Z(n696) );
  NAND2_X1 U759 ( .A1(n694), .A2(n371), .ZN(n695) );
  XNOR2_X1 U760 ( .A(n696), .B(n695), .ZN(n698) );
  NOR2_X1 U761 ( .A1(n698), .A2(n697), .ZN(n699) );
  NAND2_X1 U762 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U763 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U764 ( .A(KEYINPUT51), .B(n703), .ZN(n704) );
  NOR2_X1 U765 ( .A1(n704), .A2(n720), .ZN(n714) );
  NOR2_X1 U766 ( .A1(n705), .A2(n381), .ZN(n706) );
  NOR2_X1 U767 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U768 ( .A(n708), .B(KEYINPUT116), .ZN(n712) );
  NOR2_X1 U769 ( .A1(n710), .A2(n709), .ZN(n711) );
  NOR2_X1 U770 ( .A1(n712), .A2(n711), .ZN(n713) );
  NOR2_X1 U771 ( .A1(n714), .A2(n354), .ZN(n715) );
  XNOR2_X1 U772 ( .A(n715), .B(KEYINPUT52), .ZN(n716) );
  NOR2_X1 U773 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U774 ( .A(n718), .B(KEYINPUT117), .ZN(n722) );
  OR2_X1 U775 ( .A1(n720), .A2(n719), .ZN(n721) );
  NAND2_X1 U776 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U777 ( .A(KEYINPUT118), .B(n723), .ZN(n728) );
  NAND2_X1 U778 ( .A1(n724), .A2(KEYINPUT74), .ZN(n726) );
  XNOR2_X1 U779 ( .A(n726), .B(n725), .ZN(n727) );
  NOR2_X1 U780 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U781 ( .A(n729), .B(KEYINPUT119), .ZN(n730) );
  NOR2_X1 U782 ( .A1(G953), .A2(n730), .ZN(n731) );
  XNOR2_X1 U783 ( .A(KEYINPUT53), .B(n731), .ZN(G75) );
  NAND2_X1 U784 ( .A1(n732), .A2(G478), .ZN(n733) );
  XOR2_X1 U785 ( .A(n734), .B(n733), .Z(n735) );
  NOR2_X1 U786 ( .A1(n736), .A2(n735), .ZN(G63) );
  XOR2_X1 U787 ( .A(KEYINPUT123), .B(n737), .Z(n739) );
  NOR2_X1 U788 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U789 ( .A(KEYINPUT124), .B(n740), .ZN(n749) );
  BUF_X1 U790 ( .A(n741), .Z(n743) );
  NAND2_X1 U791 ( .A1(n743), .A2(n742), .ZN(n747) );
  NAND2_X1 U792 ( .A1(G953), .A2(G224), .ZN(n744) );
  XNOR2_X1 U793 ( .A(n744), .B(KEYINPUT61), .ZN(n745) );
  NAND2_X1 U794 ( .A1(n745), .A2(G898), .ZN(n746) );
  NAND2_X1 U795 ( .A1(n747), .A2(n746), .ZN(n748) );
  XNOR2_X1 U796 ( .A(n749), .B(n748), .ZN(G69) );
  XOR2_X1 U797 ( .A(n751), .B(n750), .Z(n755) );
  XNOR2_X1 U798 ( .A(n752), .B(n755), .ZN(n753) );
  NOR2_X1 U799 ( .A1(G953), .A2(n753), .ZN(n754) );
  XNOR2_X1 U800 ( .A(n754), .B(KEYINPUT125), .ZN(n760) );
  XNOR2_X1 U801 ( .A(n755), .B(G227), .ZN(n756) );
  NAND2_X1 U802 ( .A1(n756), .A2(G900), .ZN(n757) );
  XNOR2_X1 U803 ( .A(KEYINPUT126), .B(n757), .ZN(n758) );
  NAND2_X1 U804 ( .A1(n758), .A2(G953), .ZN(n759) );
  NAND2_X1 U805 ( .A1(n760), .A2(n759), .ZN(G72) );
  XOR2_X1 U806 ( .A(n761), .B(G131), .Z(G33) );
  XNOR2_X1 U807 ( .A(G143), .B(n762), .ZN(G45) );
  XNOR2_X1 U808 ( .A(G137), .B(KEYINPUT127), .ZN(n764) );
  XNOR2_X1 U809 ( .A(n764), .B(n763), .ZN(G39) );
endmodule

