//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 0 1 0 1 1 1 1 1 0 1 1 1 1 1 0 1 0 1 1 0 0 1 0 0 0 0 1 0 0 0 0 1 1 0 0 0 0 0 0 0 1 1 0 0 1 0 0 0 1 0 0 0 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:53 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n444, new_n448, new_n450, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n571, new_n572, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n581, new_n582,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n608, new_n609, new_n610, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n637, new_n639, new_n640,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT64), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  AND2_X1   g018(.A1(G2072), .A2(G2078), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  NAND2_X1  g022(.A1(G94), .A2(G452), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT65), .ZN(G173));
  NAND2_X1  g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g026(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g027(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT2), .Z(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI22_X1  g034(.A1(new_n455), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT66), .Z(G319));
  INV_X1    g036(.A(G137), .ZN(new_n462));
  OR2_X1    g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  AND2_X1   g040(.A1(KEYINPUT67), .A2(G2105), .ZN(new_n466));
  NOR2_X1   g041(.A1(KEYINPUT67), .A2(G2105), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  AND2_X1   g044(.A1(new_n469), .A2(G2104), .ZN(new_n470));
  AOI22_X1  g045(.A1(new_n465), .A2(new_n468), .B1(G101), .B2(new_n470), .ZN(new_n471));
  XNOR2_X1  g046(.A(KEYINPUT67), .B(G2105), .ZN(new_n472));
  INV_X1    g047(.A(G125), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n473), .B1(new_n463), .B2(new_n464), .ZN(new_n474));
  AND2_X1   g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n472), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n471), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G160));
  AND3_X1   g053(.A1(new_n463), .A2(KEYINPUT68), .A3(new_n464), .ZN(new_n479));
  AOI21_X1  g054(.A(KEYINPUT68), .B1(new_n463), .B2(new_n464), .ZN(new_n480));
  OAI21_X1  g055(.A(new_n472), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(G124), .ZN(new_n482));
  NOR2_X1   g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  XOR2_X1   g058(.A(new_n483), .B(KEYINPUT69), .Z(new_n484));
  OAI21_X1  g059(.A(G2104), .B1(new_n468), .B2(G112), .ZN(new_n485));
  OAI22_X1  g060(.A1(new_n481), .A2(new_n482), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n469), .B1(new_n479), .B2(new_n480), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n486), .B1(G136), .B2(new_n488), .ZN(G162));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n490));
  OR2_X1    g065(.A1(new_n490), .A2(KEYINPUT71), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(new_n492));
  AND2_X1   g067(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n493));
  NOR2_X1   g068(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n494));
  OAI21_X1  g069(.A(G138), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n492), .B1(new_n495), .B2(new_n472), .ZN(new_n496));
  XNOR2_X1  g071(.A(KEYINPUT3), .B(G2104), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n468), .A2(new_n497), .A3(G138), .A4(new_n491), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n469), .A2(G114), .ZN(new_n500));
  OAI21_X1  g075(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n501));
  OAI21_X1  g076(.A(KEYINPUT70), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  OR2_X1    g077(.A1(G102), .A2(G2105), .ZN(new_n503));
  INV_X1    g078(.A(G114), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(G2105), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT70), .ZN(new_n506));
  NAND4_X1  g081(.A1(new_n503), .A2(new_n505), .A3(new_n506), .A4(G2104), .ZN(new_n507));
  AND2_X1   g082(.A1(G126), .A2(G2105), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n502), .A2(new_n507), .B1(new_n497), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n499), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(G164));
  INV_X1    g086(.A(G543), .ZN(new_n512));
  OAI21_X1  g087(.A(KEYINPUT73), .B1(new_n512), .B2(KEYINPUT5), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT73), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT5), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n514), .A2(new_n515), .A3(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n513), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(KEYINPUT72), .A2(G651), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT6), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g095(.A1(KEYINPUT72), .A2(KEYINPUT6), .A3(G651), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n512), .A2(KEYINPUT5), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n517), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(KEYINPUT74), .ZN(new_n525));
  AOI22_X1  g100(.A1(new_n513), .A2(new_n516), .B1(KEYINPUT5), .B2(new_n512), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT74), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n526), .A2(new_n527), .A3(new_n522), .ZN(new_n528));
  AND2_X1   g103(.A1(new_n525), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(G88), .ZN(new_n530));
  NAND2_X1  g105(.A1(G75), .A2(G543), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n531), .B(KEYINPUT75), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n517), .A2(new_n523), .ZN(new_n533));
  INV_X1    g108(.A(G62), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n512), .B1(new_n520), .B2(new_n521), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n535), .A2(G651), .B1(G50), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n530), .A2(new_n537), .ZN(G303));
  INV_X1    g113(.A(G303), .ZN(G166));
  NAND2_X1  g114(.A1(new_n533), .A2(KEYINPUT76), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT76), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n526), .A2(new_n541), .ZN(new_n542));
  NAND4_X1  g117(.A1(new_n540), .A2(G63), .A3(new_n542), .A4(G651), .ZN(new_n543));
  NAND3_X1  g118(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n544));
  OR2_X1    g119(.A1(new_n544), .A2(KEYINPUT7), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n544), .A2(KEYINPUT7), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n536), .A2(G51), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  AND2_X1   g122(.A1(new_n543), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n529), .A2(G89), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n548), .A2(new_n549), .ZN(G286));
  INV_X1    g125(.A(G286), .ZN(G168));
  INV_X1    g126(.A(G651), .ZN(new_n552));
  NAND2_X1  g127(.A1(G77), .A2(G543), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n540), .A2(new_n542), .ZN(new_n554));
  INV_X1    g129(.A(G64), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  AOI21_X1  g131(.A(new_n552), .B1(new_n556), .B2(KEYINPUT77), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n557), .B1(KEYINPUT77), .B2(new_n556), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n529), .A2(G90), .B1(G52), .B2(new_n536), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n558), .A2(new_n559), .ZN(G301));
  INV_X1    g135(.A(G301), .ZN(G171));
  XNOR2_X1  g136(.A(KEYINPUT78), .B(G81), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n529), .A2(new_n562), .B1(G43), .B2(new_n536), .ZN(new_n563));
  AND3_X1   g138(.A1(new_n540), .A2(G56), .A3(new_n542), .ZN(new_n564));
  AND2_X1   g139(.A1(G68), .A2(G543), .ZN(new_n565));
  OAI21_X1  g140(.A(G651), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n563), .A2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G860), .ZN(G153));
  NAND4_X1  g144(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g145(.A1(G1), .A2(G3), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n571), .B(KEYINPUT8), .ZN(new_n572));
  NAND4_X1  g147(.A1(G319), .A2(G483), .A3(G661), .A4(new_n572), .ZN(G188));
  NAND2_X1  g148(.A1(new_n536), .A2(G53), .ZN(new_n574));
  XOR2_X1   g149(.A(new_n574), .B(KEYINPUT9), .Z(new_n575));
  AOI21_X1  g150(.A(new_n575), .B1(G91), .B2(new_n529), .ZN(new_n576));
  AND2_X1   g151(.A1(new_n526), .A2(KEYINPUT79), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n526), .A2(KEYINPUT79), .ZN(new_n578));
  OAI21_X1  g153(.A(G65), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(G78), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n579), .B1(new_n580), .B2(new_n512), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n581), .A2(G651), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n576), .A2(new_n582), .ZN(G299));
  NAND2_X1  g158(.A1(new_n536), .A2(G49), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n585), .B1(new_n529), .B2(G87), .ZN(new_n586));
  AOI21_X1  g161(.A(G74), .B1(new_n540), .B2(new_n542), .ZN(new_n587));
  NOR3_X1   g162(.A1(new_n587), .A2(KEYINPUT80), .A3(new_n552), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT80), .ZN(new_n589));
  INV_X1    g164(.A(G74), .ZN(new_n590));
  AND3_X1   g165(.A1(new_n517), .A2(new_n541), .A3(new_n523), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n541), .B1(new_n517), .B2(new_n523), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n590), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n589), .B1(new_n593), .B2(G651), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n586), .B1(new_n588), .B2(new_n594), .ZN(G288));
  NAND3_X1  g170(.A1(new_n525), .A2(G86), .A3(new_n528), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n536), .A2(G48), .ZN(new_n597));
  AND2_X1   g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT81), .ZN(new_n599));
  AND2_X1   g174(.A1(G73), .A2(G543), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n600), .B1(new_n526), .B2(G61), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n599), .B1(new_n601), .B2(new_n552), .ZN(new_n602));
  AND3_X1   g177(.A1(new_n517), .A2(G61), .A3(new_n523), .ZN(new_n603));
  OAI211_X1 g178(.A(KEYINPUT81), .B(G651), .C1(new_n603), .C2(new_n600), .ZN(new_n604));
  AND3_X1   g179(.A1(new_n602), .A2(new_n604), .A3(KEYINPUT82), .ZN(new_n605));
  AOI21_X1  g180(.A(KEYINPUT82), .B1(new_n602), .B2(new_n604), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n598), .B1(new_n605), .B2(new_n606), .ZN(G305));
  AOI22_X1  g182(.A1(new_n529), .A2(G85), .B1(G47), .B2(new_n536), .ZN(new_n608));
  AND3_X1   g183(.A1(new_n540), .A2(G60), .A3(new_n542), .ZN(new_n609));
  AND2_X1   g184(.A1(G72), .A2(G543), .ZN(new_n610));
  OAI21_X1  g185(.A(G651), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n608), .A2(new_n611), .ZN(G290));
  NAND2_X1  g187(.A1(G301), .A2(G868), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT83), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n536), .A2(G54), .ZN(new_n615));
  OAI21_X1  g190(.A(G66), .B1(new_n577), .B2(new_n578), .ZN(new_n616));
  NAND2_X1  g191(.A1(G79), .A2(G543), .ZN(new_n617));
  AND2_X1   g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  OAI211_X1 g193(.A(new_n614), .B(new_n615), .C1(new_n618), .C2(new_n552), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n552), .B1(new_n616), .B2(new_n617), .ZN(new_n620));
  INV_X1    g195(.A(new_n615), .ZN(new_n621));
  OAI21_X1  g196(.A(KEYINPUT83), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n619), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n529), .A2(G92), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(KEYINPUT10), .Z(new_n625));
  NAND2_X1  g200(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  INV_X1    g201(.A(new_n626), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n613), .B1(new_n627), .B2(G868), .ZN(G284));
  OAI21_X1  g203(.A(new_n613), .B1(new_n627), .B2(G868), .ZN(G321));
  NAND2_X1  g204(.A1(G286), .A2(G868), .ZN(new_n630));
  NOR2_X1   g205(.A1(new_n630), .A2(KEYINPUT84), .ZN(new_n631));
  AND2_X1   g206(.A1(new_n630), .A2(KEYINPUT84), .ZN(new_n632));
  INV_X1    g207(.A(G868), .ZN(new_n633));
  NAND2_X1  g208(.A1(G299), .A2(new_n633), .ZN(new_n634));
  AOI21_X1  g209(.A(new_n631), .B1(new_n632), .B2(new_n634), .ZN(G297));
  AOI21_X1  g210(.A(new_n631), .B1(new_n632), .B2(new_n634), .ZN(G280));
  INV_X1    g211(.A(G559), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n627), .B1(new_n637), .B2(G860), .ZN(G148));
  NAND2_X1  g213(.A1(new_n627), .A2(new_n637), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n639), .A2(G868), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n640), .B1(G868), .B2(new_n568), .ZN(G323));
  XNOR2_X1  g216(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OAI221_X1 g217(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n468), .C2(G111), .ZN(new_n643));
  INV_X1    g218(.A(G135), .ZN(new_n644));
  INV_X1    g219(.A(G123), .ZN(new_n645));
  OAI221_X1 g220(.A(new_n643), .B1(new_n487), .B2(new_n644), .C1(new_n645), .C2(new_n481), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT85), .ZN(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(new_n648));
  OR2_X1    g223(.A1(new_n648), .A2(G2096), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n648), .A2(G2096), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n497), .A2(new_n470), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT12), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT13), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(G2100), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n649), .A2(new_n650), .A3(new_n654), .ZN(G156));
  XNOR2_X1  g230(.A(G2427), .B(G2438), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(G2430), .ZN(new_n657));
  XNOR2_X1  g232(.A(KEYINPUT15), .B(G2435), .ZN(new_n658));
  OR2_X1    g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n657), .A2(new_n658), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n659), .A2(KEYINPUT14), .A3(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2451), .B(G2454), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT16), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n661), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2443), .B(G2446), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1341), .B(G1348), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT86), .ZN(new_n669));
  OAI211_X1 g244(.A(new_n669), .B(G14), .C1(new_n667), .C2(new_n666), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(G401));
  XOR2_X1   g246(.A(G2084), .B(G2090), .Z(new_n672));
  XNOR2_X1  g247(.A(G2067), .B(G2678), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n673), .B(KEYINPUT87), .Z(new_n674));
  NOR2_X1   g249(.A1(G2072), .A2(G2078), .ZN(new_n675));
  OR2_X1    g250(.A1(new_n444), .A2(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(new_n677));
  AOI21_X1  g252(.A(new_n672), .B1(new_n674), .B2(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n676), .B(KEYINPUT17), .Z(new_n679));
  OAI21_X1  g254(.A(new_n678), .B1(new_n674), .B2(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(new_n680), .B(KEYINPUT88), .Z(new_n681));
  NAND3_X1  g256(.A1(new_n676), .A2(new_n672), .A3(new_n673), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT18), .ZN(new_n683));
  AND2_X1   g258(.A1(new_n674), .A2(new_n672), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n683), .B1(new_n684), .B2(new_n679), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n681), .A2(new_n685), .ZN(new_n686));
  XOR2_X1   g261(.A(G2096), .B(G2100), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(G227));
  XOR2_X1   g263(.A(G1971), .B(G1976), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT19), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1956), .B(G2474), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1961), .B(G1966), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  AND2_X1   g268(.A1(new_n691), .A2(new_n692), .ZN(new_n694));
  NOR3_X1   g269(.A1(new_n690), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n690), .A2(new_n693), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT89), .B(KEYINPUT20), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  AOI211_X1 g273(.A(new_n695), .B(new_n698), .C1(new_n690), .C2(new_n694), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT90), .ZN(new_n700));
  XOR2_X1   g275(.A(G1981), .B(G1986), .Z(new_n701));
  XNOR2_X1  g276(.A(G1991), .B(G1996), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  XOR2_X1   g278(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n700), .B(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(G229));
  MUX2_X1   g282(.A(G6), .B(G305), .S(G16), .Z(new_n708));
  XOR2_X1   g283(.A(KEYINPUT32), .B(G1981), .Z(new_n709));
  XOR2_X1   g284(.A(new_n708), .B(new_n709), .Z(new_n710));
  INV_X1    g285(.A(G16), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(G22), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(G166), .B2(new_n711), .ZN(new_n713));
  INV_X1    g288(.A(G1971), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n711), .A2(G23), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n525), .A2(new_n528), .ZN(new_n717));
  INV_X1    g292(.A(G87), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n584), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  OAI21_X1  g294(.A(KEYINPUT80), .B1(new_n587), .B2(new_n552), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n593), .A2(new_n589), .A3(G651), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n719), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n716), .B1(new_n722), .B2(new_n711), .ZN(new_n723));
  XOR2_X1   g298(.A(KEYINPUT33), .B(G1976), .Z(new_n724));
  NAND2_X1  g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  OR2_X1    g300(.A1(new_n723), .A2(new_n724), .ZN(new_n726));
  NAND3_X1  g301(.A1(new_n715), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  OR3_X1    g302(.A1(new_n710), .A2(KEYINPUT34), .A3(new_n727), .ZN(new_n728));
  OAI21_X1  g303(.A(KEYINPUT34), .B1(new_n710), .B2(new_n727), .ZN(new_n729));
  INV_X1    g304(.A(G29), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n730), .A2(G25), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n488), .A2(G131), .ZN(new_n732));
  INV_X1    g307(.A(new_n481), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n733), .A2(G119), .ZN(new_n734));
  OAI221_X1 g309(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n468), .C2(G107), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n732), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(new_n736), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n731), .B1(new_n737), .B2(new_n730), .ZN(new_n738));
  XOR2_X1   g313(.A(KEYINPUT35), .B(G1991), .Z(new_n739));
  XOR2_X1   g314(.A(new_n738), .B(new_n739), .Z(new_n740));
  MUX2_X1   g315(.A(G24), .B(G290), .S(G16), .Z(new_n741));
  AND2_X1   g316(.A1(new_n741), .A2(G1986), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n741), .A2(G1986), .ZN(new_n743));
  NOR3_X1   g318(.A1(new_n740), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  AND3_X1   g319(.A1(new_n728), .A2(new_n729), .A3(new_n744), .ZN(new_n745));
  XNOR2_X1  g320(.A(KEYINPUT91), .B(KEYINPUT36), .ZN(new_n746));
  AND2_X1   g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n745), .A2(new_n746), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n730), .A2(G27), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G164), .B2(new_n730), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(G2078), .ZN(new_n752));
  XNOR2_X1  g327(.A(KEYINPUT31), .B(G11), .ZN(new_n753));
  INV_X1    g328(.A(KEYINPUT30), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n754), .A2(G28), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT97), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n730), .B1(new_n754), .B2(G28), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n753), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT24), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n730), .B1(new_n759), .B2(G34), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(new_n759), .B2(G34), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(G160), .B2(G29), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n758), .B1(new_n762), .B2(G2084), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n488), .A2(G141), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n733), .A2(G129), .ZN(new_n765));
  NAND3_X1  g340(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n766));
  INV_X1    g341(.A(KEYINPUT26), .ZN(new_n767));
  OR2_X1    g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n766), .A2(new_n767), .ZN(new_n769));
  AOI22_X1  g344(.A1(new_n768), .A2(new_n769), .B1(G105), .B2(new_n470), .ZN(new_n770));
  NAND3_X1  g345(.A1(new_n764), .A2(new_n765), .A3(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(new_n771), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n772), .A2(new_n730), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(new_n730), .B2(G32), .ZN(new_n774));
  XNOR2_X1  g349(.A(KEYINPUT27), .B(G1996), .ZN(new_n775));
  OAI221_X1 g350(.A(new_n763), .B1(G2084), .B2(new_n762), .C1(new_n774), .C2(new_n775), .ZN(new_n776));
  AOI211_X1 g351(.A(new_n752), .B(new_n776), .C1(G29), .C2(new_n647), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n711), .A2(G20), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT23), .ZN(new_n779));
  INV_X1    g354(.A(G299), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n779), .B1(new_n780), .B2(new_n711), .ZN(new_n781));
  INV_X1    g356(.A(G1956), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  AOI22_X1  g358(.A1(new_n497), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n784), .A2(new_n468), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(KEYINPUT95), .Z(new_n786));
  NAND2_X1  g361(.A1(new_n488), .A2(G139), .ZN(new_n787));
  NAND3_X1  g362(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(KEYINPUT25), .Z(new_n789));
  NAND3_X1  g364(.A1(new_n786), .A2(new_n787), .A3(new_n789), .ZN(new_n790));
  MUX2_X1   g365(.A(G33), .B(new_n790), .S(G29), .Z(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(G2072), .Z(new_n792));
  NAND2_X1  g367(.A1(new_n730), .A2(G35), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G162), .B2(new_n730), .ZN(new_n794));
  XOR2_X1   g369(.A(KEYINPUT29), .B(G2090), .Z(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NAND4_X1  g371(.A1(new_n777), .A2(new_n783), .A3(new_n792), .A4(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n711), .A2(G21), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(G168), .B2(new_n711), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(G1966), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n774), .A2(new_n775), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT96), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n711), .A2(G19), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(new_n568), .B2(new_n711), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(G1341), .ZN(new_n805));
  NOR4_X1   g380(.A1(new_n797), .A2(new_n800), .A3(new_n802), .A4(new_n805), .ZN(new_n806));
  NOR2_X1   g381(.A1(G4), .A2(G16), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT92), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(new_n626), .B2(new_n711), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(G1348), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n730), .A2(G26), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(KEYINPUT28), .Z(new_n812));
  OAI221_X1 g387(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n468), .C2(G116), .ZN(new_n813));
  INV_X1    g388(.A(G140), .ZN(new_n814));
  INV_X1    g389(.A(G128), .ZN(new_n815));
  OAI221_X1 g390(.A(new_n813), .B1(new_n487), .B2(new_n814), .C1(new_n815), .C2(new_n481), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT93), .ZN(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n812), .B1(new_n818), .B2(G29), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT94), .ZN(new_n820));
  INV_X1    g395(.A(G2067), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n711), .A2(G5), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n823), .B1(G171), .B2(new_n711), .ZN(new_n824));
  INV_X1    g399(.A(G1961), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  NAND4_X1  g401(.A1(new_n806), .A2(new_n810), .A3(new_n822), .A4(new_n826), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n749), .A2(new_n827), .ZN(G311));
  INV_X1    g403(.A(G311), .ZN(G150));
  NOR2_X1   g404(.A1(new_n626), .A2(new_n637), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT38), .ZN(new_n831));
  INV_X1    g406(.A(G67), .ZN(new_n832));
  INV_X1    g407(.A(G80), .ZN(new_n833));
  OAI22_X1  g408(.A1(new_n554), .A2(new_n832), .B1(new_n833), .B2(new_n512), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n834), .A2(KEYINPUT98), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT98), .ZN(new_n836));
  OAI221_X1 g411(.A(new_n836), .B1(new_n833), .B2(new_n512), .C1(new_n554), .C2(new_n832), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n835), .A2(G651), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n838), .A2(KEYINPUT99), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT99), .ZN(new_n840));
  NAND4_X1  g415(.A1(new_n835), .A2(new_n840), .A3(new_n837), .A4(G651), .ZN(new_n841));
  AOI22_X1  g416(.A1(new_n529), .A2(G93), .B1(G55), .B2(new_n536), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n839), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n843), .A2(new_n567), .ZN(new_n844));
  INV_X1    g419(.A(new_n842), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n845), .B1(new_n838), .B2(KEYINPUT99), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n568), .B1(new_n846), .B2(new_n841), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n844), .A2(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n831), .B(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT39), .ZN(new_n850));
  AOI21_X1  g425(.A(G860), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n851), .B1(new_n850), .B2(new_n849), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n843), .A2(G860), .ZN(new_n853));
  XOR2_X1   g428(.A(new_n853), .B(KEYINPUT37), .Z(new_n854));
  NAND2_X1  g429(.A1(new_n852), .A2(new_n854), .ZN(G145));
  NAND2_X1  g430(.A1(new_n818), .A2(new_n510), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n817), .A2(G164), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n858), .A2(new_n772), .ZN(new_n859));
  OR2_X1    g434(.A1(new_n790), .A2(KEYINPUT100), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n856), .A2(new_n771), .A3(new_n857), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n862), .A2(KEYINPUT100), .A3(new_n790), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n790), .A2(KEYINPUT100), .ZN(new_n864));
  NAND4_X1  g439(.A1(new_n859), .A2(new_n864), .A3(new_n860), .A4(new_n861), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  XOR2_X1   g441(.A(new_n736), .B(KEYINPUT101), .Z(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(new_n652), .ZN(new_n868));
  OAI221_X1 g443(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n468), .C2(G118), .ZN(new_n869));
  INV_X1    g444(.A(G142), .ZN(new_n870));
  INV_X1    g445(.A(G130), .ZN(new_n871));
  OAI221_X1 g446(.A(new_n869), .B1(new_n487), .B2(new_n870), .C1(new_n871), .C2(new_n481), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n868), .B(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n866), .A2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n873), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n875), .A2(new_n863), .A3(new_n865), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n647), .B(G160), .ZN(new_n878));
  XOR2_X1   g453(.A(new_n878), .B(G162), .Z(new_n879));
  AOI21_X1  g454(.A(G37), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(new_n879), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n874), .A2(new_n876), .A3(new_n881), .ZN(new_n882));
  AND3_X1   g457(.A1(new_n880), .A2(KEYINPUT40), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(KEYINPUT40), .B1(new_n880), .B2(new_n882), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n883), .A2(new_n884), .ZN(G395));
  NAND2_X1  g460(.A1(new_n843), .A2(new_n633), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n848), .B(new_n639), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n627), .A2(new_n780), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n780), .B1(new_n623), .B2(new_n625), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n888), .A2(KEYINPUT41), .A3(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT41), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n626), .A2(G299), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n892), .B1(new_n893), .B2(new_n889), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n891), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n887), .A2(new_n895), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n893), .A2(new_n889), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n896), .B1(new_n897), .B2(new_n887), .ZN(new_n898));
  XNOR2_X1  g473(.A(G305), .B(G166), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n722), .B(G290), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT102), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n899), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n900), .A2(new_n901), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n902), .B(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(KEYINPUT103), .B(KEYINPUT42), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n904), .B(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n898), .B(new_n906), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n886), .B1(new_n907), .B2(new_n633), .ZN(G295));
  OAI21_X1  g483(.A(new_n886), .B1(new_n907), .B2(new_n633), .ZN(G331));
  NAND2_X1  g484(.A1(G301), .A2(G168), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n558), .A2(G286), .A3(new_n559), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n912), .B1(new_n844), .B2(new_n847), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n843), .A2(new_n567), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n846), .A2(new_n568), .A3(new_n841), .ZN(new_n915));
  NAND4_X1  g490(.A1(new_n914), .A2(new_n915), .A3(new_n911), .A4(new_n910), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n913), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(new_n897), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n891), .A2(new_n913), .A3(new_n894), .A4(new_n916), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(new_n904), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n918), .A2(new_n904), .A3(new_n919), .ZN(new_n923));
  INV_X1    g498(.A(G37), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n922), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(KEYINPUT43), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT104), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT43), .ZN(new_n928));
  NAND4_X1  g503(.A1(new_n922), .A2(new_n923), .A3(new_n928), .A4(new_n924), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n926), .A2(new_n927), .A3(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT44), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n925), .A2(KEYINPUT104), .A3(KEYINPUT43), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n926), .A2(KEYINPUT44), .A3(new_n929), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(G397));
  XNOR2_X1  g510(.A(new_n817), .B(new_n821), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n936), .B1(G1996), .B2(new_n771), .ZN(new_n937));
  INV_X1    g512(.A(G1384), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n510), .A2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT45), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT105), .ZN(new_n942));
  INV_X1    g517(.A(G40), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n942), .B1(new_n477), .B2(new_n943), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n471), .A2(new_n476), .A3(KEYINPUT105), .A4(G40), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n941), .A2(new_n946), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n947), .B(KEYINPUT107), .ZN(new_n948));
  INV_X1    g523(.A(new_n947), .ZN(new_n949));
  OR2_X1    g524(.A1(new_n949), .A2(G1996), .ZN(new_n950));
  OAI22_X1  g525(.A1(new_n937), .A2(new_n948), .B1(new_n771), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n737), .A2(new_n739), .ZN(new_n952));
  OR2_X1    g527(.A1(new_n737), .A2(new_n739), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n948), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  OR2_X1    g529(.A1(new_n951), .A2(new_n954), .ZN(new_n955));
  NOR2_X1   g530(.A1(G290), .A2(G1986), .ZN(new_n956));
  XNOR2_X1  g531(.A(new_n956), .B(KEYINPUT106), .ZN(new_n957));
  NAND2_X1  g532(.A1(G290), .A2(G1986), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n949), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n955), .A2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT54), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT117), .ZN(new_n962));
  AOI21_X1  g537(.A(KEYINPUT108), .B1(new_n510), .B2(new_n938), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT108), .ZN(new_n964));
  AOI211_X1 g539(.A(new_n964), .B(G1384), .C1(new_n499), .C2(new_n509), .ZN(new_n965));
  NOR3_X1   g540(.A1(new_n963), .A2(new_n965), .A3(KEYINPUT50), .ZN(new_n966));
  AOI21_X1  g541(.A(G1384), .B1(new_n499), .B2(new_n509), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT50), .ZN(new_n968));
  OAI211_X1 g543(.A(new_n944), .B(new_n945), .C1(new_n967), .C2(new_n968), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n962), .B1(new_n966), .B2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(new_n969), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n939), .A2(new_n964), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n967), .A2(KEYINPUT108), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n972), .A2(new_n968), .A3(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n971), .A2(new_n974), .A3(KEYINPUT117), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n970), .A2(new_n975), .A3(new_n825), .ZN(new_n976));
  OR2_X1    g551(.A1(new_n976), .A2(KEYINPUT124), .ZN(new_n977));
  INV_X1    g552(.A(new_n946), .ZN(new_n978));
  INV_X1    g553(.A(G2078), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n967), .A2(KEYINPUT45), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n978), .A2(new_n979), .A3(new_n941), .A4(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT53), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n976), .A2(KEYINPUT124), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n477), .A2(new_n943), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n982), .A2(G2078), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n941), .A2(new_n985), .A3(new_n980), .A4(new_n986), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n977), .A2(new_n983), .A3(new_n984), .A4(new_n987), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n988), .A2(G171), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n980), .A2(new_n944), .A3(new_n945), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n972), .A2(new_n973), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n990), .B1(new_n991), .B2(new_n940), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(new_n986), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n976), .A2(new_n983), .A3(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(G171), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT123), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n994), .A2(KEYINPUT123), .A3(G171), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n961), .B1(new_n989), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n988), .A2(G171), .ZN(new_n1001));
  OAI211_X1 g576(.A(new_n1001), .B(KEYINPUT54), .C1(G171), .C2(new_n994), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n966), .A2(new_n969), .ZN(new_n1003));
  INV_X1    g578(.A(G2090), .ZN(new_n1004));
  AND3_X1   g579(.A1(new_n980), .A2(new_n944), .A3(new_n945), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(new_n941), .ZN(new_n1006));
  AOI22_X1  g581(.A1(new_n1003), .A2(new_n1004), .B1(new_n1006), .B2(new_n714), .ZN(new_n1007));
  NAND2_X1  g582(.A1(G303), .A2(G8), .ZN(new_n1008));
  XNOR2_X1  g583(.A(KEYINPUT109), .B(KEYINPUT55), .ZN(new_n1009));
  XNOR2_X1  g584(.A(new_n1008), .B(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(G8), .ZN(new_n1011));
  NOR3_X1   g586(.A1(new_n1007), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(G1981), .ZN(new_n1014));
  OAI211_X1 g589(.A(new_n1014), .B(new_n598), .C1(new_n605), .C2(new_n606), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n602), .A2(new_n604), .A3(new_n596), .A4(new_n597), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(G1981), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT49), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1015), .A2(KEYINPUT49), .A3(new_n1017), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n963), .A2(new_n965), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1011), .B1(new_n1022), .B2(new_n978), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1020), .A2(new_n1021), .A3(new_n1023), .ZN(new_n1024));
  OAI211_X1 g599(.A(new_n586), .B(G1976), .C1(new_n588), .C2(new_n594), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n972), .A2(new_n944), .A3(new_n945), .A4(new_n973), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1025), .A2(new_n1026), .A3(G8), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT52), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1028), .B1(new_n722), .B2(G1976), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1028), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1013), .A2(new_n1024), .A3(new_n1032), .ZN(new_n1033));
  OAI21_X1  g608(.A(KEYINPUT50), .B1(new_n963), .B2(new_n965), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1034), .A2(KEYINPUT112), .A3(new_n978), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n967), .A2(new_n968), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g612(.A(KEYINPUT112), .B1(new_n1034), .B2(new_n978), .ZN(new_n1038));
  OAI21_X1  g613(.A(KEYINPUT113), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT112), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n968), .B1(new_n972), .B2(new_n973), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1040), .B1(new_n1041), .B2(new_n946), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT113), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n1042), .A2(new_n1043), .A3(new_n1036), .A4(new_n1035), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1039), .A2(new_n1004), .A3(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1006), .A2(new_n714), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(G8), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1033), .B1(new_n1048), .B2(new_n1010), .ZN(new_n1049));
  NOR3_X1   g624(.A1(new_n966), .A2(G2084), .A3(new_n969), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n940), .B1(new_n963), .B2(new_n965), .ZN(new_n1051));
  AOI21_X1  g626(.A(G1966), .B1(new_n1005), .B2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(G8), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(G286), .A2(G8), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1053), .A2(KEYINPUT51), .A3(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT51), .ZN(new_n1056));
  INV_X1    g631(.A(G1966), .ZN(new_n1057));
  AOI21_X1  g632(.A(KEYINPUT45), .B1(new_n972), .B2(new_n973), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1057), .B1(new_n1058), .B2(new_n990), .ZN(new_n1059));
  INV_X1    g634(.A(G2084), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n971), .A2(new_n974), .A3(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1062));
  OAI211_X1 g637(.A(new_n1056), .B(G8), .C1(new_n1062), .C2(G286), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT122), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1054), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1064), .B1(new_n1062), .B2(new_n1065), .ZN(new_n1066));
  AOI211_X1 g641(.A(KEYINPUT122), .B(new_n1054), .C1(new_n1059), .C2(new_n1061), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n1055), .B(new_n1063), .C1(new_n1066), .C2(new_n1067), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1000), .A2(new_n1002), .A3(new_n1049), .A4(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT61), .ZN(new_n1070));
  INV_X1    g645(.A(new_n941), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1071), .A2(new_n990), .ZN(new_n1072));
  XNOR2_X1  g647(.A(KEYINPUT56), .B(G2072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1042), .A2(new_n1036), .A3(new_n1035), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1075), .B1(new_n1076), .B2(new_n782), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT57), .ZN(new_n1078));
  XNOR2_X1  g653(.A(G299), .B(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(KEYINPUT116), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n782), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1081));
  AND4_X1   g656(.A1(KEYINPUT116), .A2(new_n1081), .A3(new_n1079), .A4(new_n1074), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g658(.A(KEYINPUT119), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1081), .A2(new_n1074), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT119), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1079), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1085), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1084), .A2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1070), .B1(new_n1083), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(KEYINPUT120), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT120), .ZN(new_n1092));
  OAI211_X1 g667(.A(new_n1092), .B(new_n1070), .C1(new_n1083), .C2(new_n1089), .ZN(new_n1093));
  INV_X1    g668(.A(G1348), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n970), .A2(new_n975), .A3(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1026), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(new_n821), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n626), .A2(KEYINPUT121), .ZN(new_n1100));
  OR2_X1    g675(.A1(new_n626), .A2(KEYINPUT121), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1099), .A2(KEYINPUT60), .A3(new_n1100), .A4(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT60), .ZN(new_n1103));
  OAI211_X1 g678(.A(KEYINPUT121), .B(new_n626), .C1(new_n1098), .C2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1098), .A2(new_n1103), .ZN(new_n1105));
  AND3_X1   g680(.A1(new_n1102), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1006), .A2(G1996), .ZN(new_n1107));
  XOR2_X1   g682(.A(KEYINPUT118), .B(KEYINPUT58), .Z(new_n1108));
  XNOR2_X1  g683(.A(new_n1108), .B(G1341), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1096), .A2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n568), .B1(new_n1107), .B2(new_n1110), .ZN(new_n1111));
  XNOR2_X1  g686(.A(new_n1111), .B(KEYINPUT59), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1113));
  OAI21_X1  g688(.A(KEYINPUT61), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1112), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1106), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1091), .A2(new_n1093), .A3(new_n1116), .ZN(new_n1117));
  OAI22_X1  g692(.A1(new_n1099), .A2(new_n626), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1118), .B1(new_n1080), .B2(new_n1082), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1069), .B1(new_n1117), .B2(new_n1119), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1065), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(KEYINPUT122), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1062), .A2(new_n1064), .A3(new_n1065), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT62), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1124), .A2(new_n1125), .A3(new_n1055), .A4(new_n1063), .ZN(new_n1126));
  AND2_X1   g701(.A1(new_n999), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1068), .A2(KEYINPUT62), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1127), .A2(new_n1049), .A3(KEYINPUT125), .A4(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT125), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1128), .A2(new_n999), .A3(new_n1126), .ZN(new_n1131));
  AND3_X1   g706(.A1(new_n1015), .A2(KEYINPUT49), .A3(new_n1017), .ZN(new_n1132));
  AOI21_X1  g707(.A(KEYINPUT49), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1023), .ZN(new_n1134));
  NOR3_X1   g709(.A1(new_n1132), .A2(new_n1133), .A3(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(G1976), .ZN(new_n1136));
  AOI21_X1  g711(.A(KEYINPUT52), .B1(G288), .B2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1137), .A2(new_n1023), .A3(new_n1025), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1027), .A2(KEYINPUT52), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NOR3_X1   g715(.A1(new_n1012), .A2(new_n1135), .A3(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1011), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1010), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1141), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1130), .B1(new_n1131), .B2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1129), .A2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT110), .ZN(new_n1147));
  NOR3_X1   g722(.A1(new_n1135), .A2(new_n1140), .A3(new_n1147), .ZN(new_n1148));
  AOI21_X1  g723(.A(KEYINPUT110), .B1(new_n1032), .B2(new_n1024), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1012), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  XOR2_X1   g725(.A(new_n1023), .B(KEYINPUT111), .Z(new_n1151));
  NOR3_X1   g726(.A1(new_n1135), .A2(G1976), .A3(G288), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1015), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1151), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1150), .A2(new_n1154), .ZN(new_n1155));
  OAI21_X1  g730(.A(KEYINPUT114), .B1(new_n1007), .B2(new_n1011), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n971), .A2(new_n974), .ZN(new_n1157));
  OAI22_X1  g732(.A1(new_n1157), .A2(G2090), .B1(new_n1072), .B2(G1971), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT114), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1158), .A2(new_n1159), .A3(G8), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1156), .A2(new_n1010), .A3(new_n1160), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1161), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT115), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  OAI211_X1 g739(.A(new_n1161), .B(KEYINPUT115), .C1(new_n1148), .C2(new_n1149), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT63), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1062), .A2(G8), .A3(G168), .ZN(new_n1167));
  NOR3_X1   g742(.A1(new_n1012), .A2(new_n1166), .A3(new_n1167), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1164), .A2(new_n1165), .A3(new_n1168), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1166), .B1(new_n1144), .B2(new_n1167), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1155), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1146), .A2(new_n1171), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n960), .B1(new_n1120), .B2(new_n1172), .ZN(new_n1173));
  XNOR2_X1  g748(.A(new_n950), .B(KEYINPUT46), .ZN(new_n1174));
  INV_X1    g749(.A(new_n948), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1175), .B1(new_n936), .B2(new_n771), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1174), .A2(new_n1176), .ZN(new_n1177));
  XNOR2_X1  g752(.A(new_n1177), .B(KEYINPUT47), .ZN(new_n1178));
  NOR2_X1   g753(.A1(new_n957), .A2(new_n949), .ZN(new_n1179));
  XNOR2_X1  g754(.A(new_n1179), .B(KEYINPUT48), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1178), .B1(new_n955), .B2(new_n1180), .ZN(new_n1181));
  OAI22_X1  g756(.A1(new_n951), .A2(new_n952), .B1(G2067), .B2(new_n818), .ZN(new_n1182));
  XOR2_X1   g757(.A(new_n1182), .B(KEYINPUT126), .Z(new_n1183));
  AOI21_X1  g758(.A(new_n1181), .B1(new_n1183), .B2(new_n1175), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1173), .A2(new_n1184), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g760(.A(new_n460), .ZN(new_n1187));
  OR2_X1    g761(.A1(G227), .A2(new_n1187), .ZN(new_n1188));
  OR2_X1    g762(.A1(new_n1188), .A2(KEYINPUT127), .ZN(new_n1189));
  NAND2_X1  g763(.A1(new_n1188), .A2(KEYINPUT127), .ZN(new_n1190));
  NAND4_X1  g764(.A1(new_n1189), .A2(new_n670), .A3(new_n706), .A4(new_n1190), .ZN(new_n1191));
  AOI21_X1  g765(.A(new_n1191), .B1(new_n880), .B2(new_n882), .ZN(new_n1192));
  AND3_X1   g766(.A1(new_n1192), .A2(new_n932), .A3(new_n930), .ZN(G308));
  NAND3_X1  g767(.A1(new_n1192), .A2(new_n930), .A3(new_n932), .ZN(G225));
endmodule


