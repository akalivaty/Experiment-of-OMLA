//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 1 0 1 1 1 1 0 1 1 0 1 0 1 0 1 1 1 0 0 1 1 0 0 0 0 0 1 1 1 1 0 1 1 1 1 1 1 1 1 0 1 0 0 1 0 0 1 1 1 0 1 1 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:34 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n699,
    new_n700, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n715,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n729, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n904, new_n905,
    new_n906, new_n907, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  INV_X1    g002(.A(G146), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G143), .ZN(new_n190));
  INV_X1    g004(.A(G143), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G146), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n190), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G128), .ZN(new_n194));
  OR2_X1    g008(.A1(new_n194), .A2(KEYINPUT1), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n193), .A2(new_n195), .ZN(new_n196));
  OAI211_X1 g010(.A(new_n191), .B(G146), .C1(new_n194), .C2(KEYINPUT1), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n194), .A2(new_n189), .A3(G143), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n196), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT74), .ZN(new_n201));
  INV_X1    g015(.A(G107), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n201), .B1(new_n202), .B2(G104), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(G104), .ZN(new_n204));
  INV_X1    g018(.A(G104), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n205), .A2(KEYINPUT74), .A3(G107), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n203), .A2(new_n204), .A3(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G101), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT76), .ZN(new_n209));
  INV_X1    g023(.A(G101), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n205), .A2(G107), .ZN(new_n211));
  AND3_X1   g025(.A1(new_n202), .A2(KEYINPUT3), .A3(G104), .ZN(new_n212));
  AOI21_X1  g026(.A(KEYINPUT3), .B1(new_n202), .B2(G104), .ZN(new_n213));
  OAI211_X1 g027(.A(new_n210), .B(new_n211), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  AND3_X1   g028(.A1(new_n208), .A2(new_n209), .A3(new_n214), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n209), .B1(new_n208), .B2(new_n214), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n200), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(new_n199), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(KEYINPUT75), .ZN(new_n219));
  INV_X1    g033(.A(new_n196), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT75), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n199), .A2(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n219), .A2(new_n220), .A3(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n223), .A2(new_n214), .A3(new_n208), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n217), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT11), .ZN(new_n226));
  INV_X1    g040(.A(G134), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n226), .B1(new_n227), .B2(G137), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(G137), .ZN(new_n229));
  INV_X1    g043(.A(G137), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n230), .A2(KEYINPUT11), .A3(G134), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n228), .A2(new_n229), .A3(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(G131), .ZN(new_n233));
  INV_X1    g047(.A(G131), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n228), .A2(new_n231), .A3(new_n234), .A4(new_n229), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  AOI21_X1  g050(.A(KEYINPUT12), .B1(new_n225), .B2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT12), .ZN(new_n238));
  INV_X1    g052(.A(new_n236), .ZN(new_n239));
  AOI211_X1 g053(.A(new_n238), .B(new_n239), .C1(new_n217), .C2(new_n224), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n237), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT3), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n242), .B1(new_n205), .B2(G107), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n202), .A2(KEYINPUT3), .A3(G104), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(new_n211), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G101), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT73), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n247), .A2(new_n248), .A3(KEYINPUT4), .A4(new_n214), .ZN(new_n249));
  INV_X1    g063(.A(new_n214), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n210), .B1(new_n245), .B2(new_n211), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n252));
  NOR3_X1   g066(.A1(new_n250), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n246), .A2(new_n252), .A3(G101), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(KEYINPUT73), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n249), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  NAND4_X1  g070(.A1(new_n190), .A2(new_n192), .A3(KEYINPUT0), .A4(G128), .ZN(new_n257));
  AND2_X1   g071(.A1(new_n190), .A2(new_n192), .ZN(new_n258));
  XNOR2_X1  g072(.A(KEYINPUT0), .B(G128), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n257), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n256), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT10), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n224), .A2(new_n263), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n215), .A2(new_n216), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n220), .A2(new_n218), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n265), .A2(KEYINPUT10), .A3(new_n266), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n262), .A2(new_n239), .A3(new_n264), .A4(new_n267), .ZN(new_n268));
  XNOR2_X1  g082(.A(G110), .B(G140), .ZN(new_n269));
  INV_X1    g083(.A(G953), .ZN(new_n270));
  AND2_X1   g084(.A1(new_n270), .A2(G227), .ZN(new_n271));
  XOR2_X1   g085(.A(new_n269), .B(new_n271), .Z(new_n272));
  NAND2_X1  g086(.A1(new_n268), .A2(new_n272), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n241), .A2(new_n273), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n262), .A2(new_n264), .A3(new_n267), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(new_n236), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n272), .B1(new_n276), .B2(new_n268), .ZN(new_n277));
  OAI211_X1 g091(.A(new_n187), .B(new_n188), .C1(new_n274), .C2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(G469), .A2(G902), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n268), .B1(new_n237), .B2(new_n240), .ZN(new_n280));
  INV_X1    g094(.A(new_n272), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n276), .A2(new_n268), .A3(new_n272), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n282), .A2(G469), .A3(new_n283), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n278), .A2(new_n279), .A3(new_n284), .ZN(new_n285));
  XOR2_X1   g099(.A(KEYINPUT9), .B(G234), .Z(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  OAI21_X1  g101(.A(G221), .B1(new_n287), .B2(G902), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n285), .A2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT77), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n285), .A2(KEYINPUT77), .A3(new_n288), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(G217), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n294), .B1(G234), .B2(new_n188), .ZN(new_n295));
  OR2_X1    g109(.A1(KEYINPUT69), .A2(KEYINPUT23), .ZN(new_n296));
  NAND2_X1  g110(.A1(KEYINPUT69), .A2(KEYINPUT23), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n296), .A2(G119), .A3(new_n194), .A4(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n194), .A2(G119), .ZN(new_n299));
  INV_X1    g113(.A(G119), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(G128), .ZN(new_n301));
  AND2_X1   g115(.A1(KEYINPUT69), .A2(KEYINPUT23), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n299), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n298), .A2(new_n303), .A3(G110), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT70), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND4_X1  g120(.A1(new_n298), .A2(new_n303), .A3(KEYINPUT70), .A4(G110), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(G140), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(G125), .ZN(new_n310));
  INV_X1    g124(.A(G125), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(G140), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT16), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NOR3_X1   g129(.A1(new_n311), .A2(KEYINPUT16), .A3(G140), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n189), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  XNOR2_X1  g131(.A(G125), .B(G140), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n316), .B1(new_n318), .B2(KEYINPUT16), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G146), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n317), .A2(new_n320), .ZN(new_n321));
  AND2_X1   g135(.A1(new_n299), .A2(new_n301), .ZN(new_n322));
  XOR2_X1   g136(.A(KEYINPUT24), .B(G110), .Z(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n308), .A2(new_n321), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(G221), .A2(G234), .ZN(new_n326));
  OAI21_X1  g140(.A(KEYINPUT22), .B1(new_n326), .B2(G953), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT22), .ZN(new_n328));
  NAND4_X1  g142(.A1(new_n328), .A2(new_n270), .A3(G221), .A4(G234), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n327), .A2(new_n329), .A3(G137), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  AOI21_X1  g145(.A(G137), .B1(new_n327), .B2(new_n329), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  AND2_X1   g147(.A1(new_n298), .A2(new_n303), .ZN(new_n334));
  OAI22_X1  g148(.A1(new_n334), .A2(G110), .B1(new_n322), .B2(new_n323), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n313), .A2(G146), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n336), .B1(new_n319), .B2(G146), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  AND3_X1   g152(.A1(new_n325), .A2(new_n333), .A3(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT71), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n340), .B1(new_n331), .B2(new_n332), .ZN(new_n341));
  INV_X1    g155(.A(new_n332), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n342), .A2(KEYINPUT71), .A3(new_n330), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n344), .B1(new_n325), .B2(new_n338), .ZN(new_n345));
  OAI21_X1  g159(.A(KEYINPUT72), .B1(new_n339), .B2(new_n345), .ZN(new_n346));
  AOI22_X1  g160(.A1(new_n306), .A2(new_n307), .B1(new_n322), .B2(new_n323), .ZN(new_n347));
  AOI22_X1  g161(.A1(new_n347), .A2(new_n321), .B1(new_n335), .B2(new_n337), .ZN(new_n348));
  AOI21_X1  g162(.A(KEYINPUT72), .B1(new_n348), .B2(new_n333), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n346), .A2(new_n350), .A3(new_n188), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT25), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n325), .A2(new_n338), .A3(new_n333), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n354), .B1(new_n348), .B2(new_n344), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n349), .B1(new_n355), .B2(KEYINPUT72), .ZN(new_n356));
  AOI21_X1  g170(.A(KEYINPUT25), .B1(new_n356), .B2(new_n188), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n295), .B1(new_n353), .B2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n356), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n295), .A2(G902), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n358), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT30), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n230), .A2(G134), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n227), .A2(G137), .ZN(new_n365));
  OAI21_X1  g179(.A(G131), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n235), .A2(new_n366), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n367), .A2(KEYINPUT64), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT64), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n369), .B1(new_n235), .B2(new_n366), .ZN(new_n370));
  NOR3_X1   g184(.A1(new_n368), .A2(new_n200), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n261), .A2(new_n236), .ZN(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n363), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT65), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n372), .A2(new_n375), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n200), .A2(new_n367), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n261), .A2(new_n236), .A3(KEYINPUT65), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n376), .A2(KEYINPUT30), .A3(new_n378), .A4(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n300), .A2(G116), .ZN(new_n381));
  INV_X1    g195(.A(G116), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(G119), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  XOR2_X1   g199(.A(KEYINPUT2), .B(G113), .Z(new_n386));
  OR2_X1    g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n385), .A2(new_n386), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n374), .A2(new_n380), .A3(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(G237), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n391), .A2(new_n270), .A3(G210), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT27), .ZN(new_n393));
  XNOR2_X1  g207(.A(new_n392), .B(new_n393), .ZN(new_n394));
  XNOR2_X1  g208(.A(new_n394), .B(KEYINPUT26), .ZN(new_n395));
  XNOR2_X1  g209(.A(new_n395), .B(new_n210), .ZN(new_n396));
  INV_X1    g210(.A(new_n389), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n376), .A2(new_n397), .A3(new_n378), .A4(new_n379), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n390), .A2(new_n396), .A3(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT31), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND4_X1  g215(.A1(new_n390), .A2(new_n396), .A3(KEYINPUT31), .A4(new_n398), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  OR2_X1    g217(.A1(new_n395), .A2(G101), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n395), .A2(G101), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT66), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n396), .A2(KEYINPUT66), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NOR3_X1   g224(.A1(new_n373), .A2(new_n389), .A3(new_n377), .ZN(new_n411));
  OR2_X1    g225(.A1(new_n411), .A2(KEYINPUT28), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n389), .B1(new_n371), .B2(new_n373), .ZN(new_n413));
  AND2_X1   g227(.A1(new_n413), .A2(new_n398), .ZN(new_n414));
  XNOR2_X1  g228(.A(KEYINPUT67), .B(KEYINPUT28), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n412), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n410), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n403), .A2(new_n417), .ZN(new_n418));
  NOR2_X1   g232(.A1(G472), .A2(G902), .ZN(new_n419));
  AOI21_X1  g233(.A(KEYINPUT32), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  AOI22_X1  g234(.A1(new_n401), .A2(new_n402), .B1(new_n410), .B2(new_n416), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT32), .ZN(new_n422));
  INV_X1    g236(.A(new_n419), .ZN(new_n423));
  NOR3_X1   g237(.A1(new_n421), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n420), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n376), .A2(new_n378), .A3(new_n379), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(new_n389), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n427), .A2(KEYINPUT68), .A3(new_n398), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT68), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n426), .A2(new_n429), .A3(new_n389), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n428), .A2(KEYINPUT28), .A3(new_n430), .ZN(new_n431));
  NAND4_X1  g245(.A1(new_n431), .A2(KEYINPUT29), .A3(new_n396), .A4(new_n412), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT29), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n433), .B1(new_n410), .B2(new_n416), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n396), .B1(new_n390), .B2(new_n398), .ZN(new_n435));
  OAI211_X1 g249(.A(new_n432), .B(new_n188), .C1(new_n434), .C2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(G472), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n362), .B1(new_n425), .B2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(G478), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n439), .A2(KEYINPUT15), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n194), .A2(G143), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT13), .ZN(new_n443));
  OAI21_X1  g257(.A(KEYINPUT86), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT86), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n441), .A2(new_n445), .A3(KEYINPUT13), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n194), .A2(G143), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n444), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n441), .A2(KEYINPUT13), .ZN(new_n449));
  OAI21_X1  g263(.A(G134), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  AND2_X1   g264(.A1(new_n442), .A2(new_n447), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(new_n227), .ZN(new_n452));
  INV_X1    g266(.A(G122), .ZN(new_n453));
  OR2_X1    g267(.A1(new_n453), .A2(KEYINPUT85), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(KEYINPUT85), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n382), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n453), .A2(G116), .ZN(new_n457));
  OAI21_X1  g271(.A(G107), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  NOR3_X1   g273(.A1(new_n456), .A2(G107), .A3(new_n457), .ZN(new_n460));
  OAI211_X1 g274(.A(new_n450), .B(new_n452), .C1(new_n459), .C2(new_n460), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n451), .B(new_n227), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n456), .A2(new_n457), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n463), .B1(KEYINPUT14), .B2(new_n202), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT14), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n456), .A2(new_n465), .ZN(new_n466));
  OAI211_X1 g280(.A(new_n462), .B(new_n464), .C1(new_n458), .C2(new_n466), .ZN(new_n467));
  NOR3_X1   g281(.A1(new_n287), .A2(new_n294), .A3(G953), .ZN(new_n468));
  AND3_X1   g282(.A1(new_n461), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n468), .B1(new_n461), .B2(new_n467), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n188), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT87), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n440), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n471), .A2(new_n472), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n461), .A2(new_n467), .ZN(new_n475));
  INV_X1    g289(.A(new_n468), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n461), .A2(new_n467), .A3(new_n468), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n479), .A2(KEYINPUT87), .A3(new_n188), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n474), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n473), .B1(new_n481), .B2(new_n440), .ZN(new_n482));
  INV_X1    g296(.A(G475), .ZN(new_n483));
  INV_X1    g297(.A(new_n321), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n391), .A2(new_n270), .A3(G214), .ZN(new_n485));
  XNOR2_X1  g299(.A(new_n485), .B(new_n191), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n486), .A2(KEYINPUT17), .A3(G131), .ZN(new_n487));
  OAI21_X1  g301(.A(KEYINPUT82), .B1(new_n486), .B2(G131), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n486), .A2(G131), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n485), .B(G143), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT82), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n490), .A2(new_n491), .A3(new_n234), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n488), .A2(new_n489), .A3(new_n492), .ZN(new_n493));
  OAI211_X1 g307(.A(new_n484), .B(new_n487), .C1(new_n493), .C2(KEYINPUT17), .ZN(new_n494));
  XNOR2_X1  g308(.A(G113), .B(G122), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n495), .B(new_n205), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT18), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n490), .B1(new_n497), .B2(new_n234), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n318), .A2(new_n189), .ZN(new_n499));
  OAI221_X1 g313(.A(new_n498), .B1(new_n336), .B2(new_n499), .C1(new_n489), .C2(new_n497), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n494), .A2(new_n496), .A3(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  XNOR2_X1  g316(.A(new_n318), .B(KEYINPUT19), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(new_n189), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n493), .A2(new_n320), .A3(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n496), .B1(new_n505), .B2(new_n500), .ZN(new_n506));
  OAI211_X1 g320(.A(new_n483), .B(new_n188), .C1(new_n502), .C2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n506), .ZN(new_n508));
  AOI21_X1  g322(.A(KEYINPUT83), .B1(new_n508), .B2(new_n501), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n507), .B1(KEYINPUT20), .B2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT83), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n511), .B1(new_n502), .B2(new_n506), .ZN(new_n512));
  AOI21_X1  g326(.A(G475), .B1(new_n508), .B2(new_n501), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT20), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n512), .A2(new_n513), .A3(new_n514), .A4(new_n188), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n510), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n270), .A2(G952), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n517), .B1(G234), .B2(G237), .ZN(new_n518));
  XOR2_X1   g332(.A(KEYINPUT21), .B(G898), .Z(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(G234), .A2(G237), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n521), .A2(G902), .A3(G953), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n518), .B1(new_n520), .B2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n496), .B1(new_n494), .B2(new_n500), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n188), .B1(new_n502), .B2(new_n526), .ZN(new_n527));
  XOR2_X1   g341(.A(KEYINPUT84), .B(G475), .Z(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n482), .A2(new_n516), .A3(new_n525), .A4(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT88), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  AOI22_X1  g347(.A1(new_n510), .A2(new_n515), .B1(new_n527), .B2(new_n529), .ZN(new_n534));
  NAND4_X1  g348(.A1(new_n534), .A2(KEYINPUT88), .A3(new_n525), .A4(new_n482), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT6), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT5), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n384), .A2(new_n538), .ZN(new_n539));
  OAI21_X1  g353(.A(G113), .B1(new_n381), .B2(KEYINPUT5), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n388), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NOR3_X1   g355(.A1(new_n215), .A2(new_n216), .A3(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n542), .B1(new_n256), .B2(new_n389), .ZN(new_n543));
  XOR2_X1   g357(.A(G110), .B(G122), .Z(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n545), .A2(KEYINPUT78), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n537), .B1(new_n543), .B2(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n247), .A2(KEYINPUT4), .A3(new_n214), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n549), .A2(KEYINPUT73), .A3(new_n254), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n397), .B1(new_n550), .B2(new_n249), .ZN(new_n551));
  OAI211_X1 g365(.A(KEYINPUT6), .B(new_n546), .C1(new_n551), .C2(new_n542), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n543), .A2(new_n545), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n548), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n260), .A2(G125), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n555), .B1(new_n266), .B2(G125), .ZN(new_n556));
  INV_X1    g370(.A(G224), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n557), .A2(G953), .ZN(new_n558));
  XNOR2_X1  g372(.A(new_n556), .B(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n554), .A2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT80), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n556), .B1(new_n561), .B2(new_n558), .ZN(new_n562));
  OAI21_X1  g376(.A(KEYINPUT7), .B1(new_n557), .B2(G953), .ZN(new_n563));
  XNOR2_X1  g377(.A(new_n562), .B(new_n563), .ZN(new_n564));
  XOR2_X1   g378(.A(new_n544), .B(KEYINPUT8), .Z(new_n565));
  OAI22_X1  g379(.A1(new_n540), .A2(KEYINPUT79), .B1(new_n384), .B2(new_n538), .ZN(new_n566));
  AND2_X1   g380(.A1(new_n540), .A2(KEYINPUT79), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n388), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NOR3_X1   g382(.A1(new_n568), .A2(new_n215), .A3(new_n216), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n208), .A2(new_n214), .ZN(new_n570));
  AND2_X1   g384(.A1(new_n541), .A2(new_n570), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n565), .B1(new_n569), .B2(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n564), .A2(new_n553), .A3(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n560), .A2(new_n188), .A3(new_n573), .ZN(new_n574));
  OAI21_X1  g388(.A(G210), .B1(G237), .B2(G902), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  NAND4_X1  g391(.A1(new_n560), .A2(new_n188), .A3(new_n575), .A4(new_n573), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n577), .A2(KEYINPUT81), .A3(new_n578), .ZN(new_n579));
  OAI21_X1  g393(.A(G214), .B1(G237), .B2(G902), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT81), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n574), .A2(new_n581), .A3(new_n576), .ZN(new_n582));
  AND3_X1   g396(.A1(new_n579), .A2(new_n580), .A3(new_n582), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n293), .A2(new_n438), .A3(new_n536), .A4(new_n583), .ZN(new_n584));
  XNOR2_X1  g398(.A(new_n584), .B(G101), .ZN(G3));
  OAI21_X1  g399(.A(G472), .B1(new_n421), .B2(G902), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n418), .A2(new_n419), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AOI211_X1 g402(.A(new_n362), .B(new_n588), .C1(new_n291), .C2(new_n292), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n516), .A2(new_n530), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT33), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n479), .A2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT89), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n479), .A2(KEYINPUT89), .A3(new_n591), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT90), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n591), .B1(new_n469), .B2(new_n596), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n470), .B1(KEYINPUT90), .B2(new_n478), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n439), .A2(G902), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n594), .A2(new_n595), .A3(new_n599), .A4(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n471), .A2(new_n439), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n590), .A2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n580), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n606), .B1(new_n577), .B2(new_n578), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n605), .A2(new_n525), .A3(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n589), .A2(new_n609), .ZN(new_n610));
  XOR2_X1   g424(.A(new_n610), .B(KEYINPUT91), .Z(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(KEYINPUT34), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n612), .B(new_n205), .ZN(G6));
  NAND2_X1  g427(.A1(new_n607), .A2(new_n525), .ZN(new_n614));
  INV_X1    g428(.A(new_n482), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n507), .A2(new_n514), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n513), .A2(KEYINPUT20), .A3(new_n188), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n616), .A2(new_n530), .A3(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n615), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n614), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n589), .A2(new_n621), .ZN(new_n622));
  XOR2_X1   g436(.A(KEYINPUT35), .B(G107), .Z(new_n623));
  XNOR2_X1  g437(.A(new_n622), .B(new_n623), .ZN(G9));
  INV_X1    g438(.A(KEYINPUT92), .ZN(new_n625));
  AOI21_X1  g439(.A(KEYINPUT36), .B1(new_n341), .B2(new_n343), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n348), .B(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n627), .A2(new_n361), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n358), .A2(new_n625), .A3(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n295), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n351), .A2(new_n352), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n356), .A2(KEYINPUT25), .A3(new_n188), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n631), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  OAI21_X1  g448(.A(KEYINPUT92), .B1(new_n634), .B2(new_n628), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n630), .A2(new_n635), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n636), .B1(new_n533), .B2(new_n535), .ZN(new_n637));
  INV_X1    g451(.A(new_n588), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n637), .A2(new_n293), .A3(new_n583), .A4(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(KEYINPUT93), .ZN(new_n640));
  XNOR2_X1  g454(.A(KEYINPUT37), .B(G110), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(G12));
  AOI21_X1  g456(.A(new_n636), .B1(new_n425), .B2(new_n437), .ZN(new_n643));
  XOR2_X1   g457(.A(new_n518), .B(KEYINPUT94), .Z(new_n644));
  INV_X1    g458(.A(G900), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n644), .B1(new_n645), .B2(new_n523), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n620), .A2(new_n646), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n643), .A2(new_n293), .A3(new_n607), .A4(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(G128), .ZN(G30));
  NAND2_X1  g463(.A1(new_n579), .A2(new_n582), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(KEYINPUT95), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(KEYINPUT38), .ZN(new_n652));
  AND3_X1   g466(.A1(new_n410), .A2(new_n430), .A3(new_n428), .ZN(new_n653));
  INV_X1    g467(.A(new_n399), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n188), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(G472), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n425), .A2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n652), .A2(new_n658), .ZN(new_n659));
  NOR3_X1   g473(.A1(new_n534), .A2(new_n482), .A3(new_n606), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(new_n636), .ZN(new_n661));
  XOR2_X1   g475(.A(new_n661), .B(KEYINPUT96), .Z(new_n662));
  XOR2_X1   g476(.A(new_n646), .B(KEYINPUT39), .Z(new_n663));
  NAND2_X1  g477(.A1(new_n293), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(KEYINPUT97), .ZN(new_n665));
  INV_X1    g479(.A(KEYINPUT40), .ZN(new_n666));
  AND2_X1   g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n665), .A2(new_n666), .ZN(new_n668));
  OAI211_X1 g482(.A(new_n659), .B(new_n662), .C1(new_n667), .C2(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(G143), .ZN(G45));
  AND2_X1   g484(.A1(new_n643), .A2(new_n293), .ZN(new_n671));
  INV_X1    g485(.A(new_n607), .ZN(new_n672));
  INV_X1    g486(.A(new_n646), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n590), .A2(new_n603), .A3(new_n673), .ZN(new_n674));
  OAI21_X1  g488(.A(KEYINPUT98), .B1(new_n672), .B2(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(new_n674), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT98), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n676), .A2(new_n677), .A3(new_n607), .ZN(new_n678));
  AND3_X1   g492(.A1(new_n671), .A2(new_n675), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(new_n189), .ZN(G48));
  INV_X1    g494(.A(new_n420), .ZN(new_n681));
  INV_X1    g495(.A(new_n424), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n681), .A2(new_n682), .A3(new_n437), .ZN(new_n683));
  INV_X1    g497(.A(new_n362), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(new_n274), .ZN(new_n686));
  INV_X1    g500(.A(new_n277), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n187), .B1(new_n688), .B2(new_n188), .ZN(new_n689));
  INV_X1    g503(.A(new_n278), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n288), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n685), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(new_n609), .ZN(new_n694));
  XNOR2_X1  g508(.A(KEYINPUT41), .B(G113), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(G15));
  NAND2_X1  g510(.A1(new_n693), .A2(new_n621), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G116), .ZN(G18));
  NOR2_X1   g512(.A1(new_n692), .A2(new_n672), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n699), .A2(new_n683), .A3(new_n637), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G119), .ZN(G21));
  AOI211_X1 g515(.A(new_n408), .B(new_n409), .C1(new_n431), .C2(new_n412), .ZN(new_n702));
  INV_X1    g516(.A(new_n403), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n419), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(new_n586), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n705), .A2(new_n362), .ZN(new_n706));
  INV_X1    g520(.A(new_n288), .ZN(new_n707));
  NOR3_X1   g521(.A1(new_n689), .A2(new_n690), .A3(new_n707), .ZN(new_n708));
  AND3_X1   g522(.A1(new_n706), .A2(new_n525), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n577), .A2(new_n578), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n660), .A2(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n709), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G122), .ZN(G24));
  NOR3_X1   g528(.A1(new_n636), .A2(new_n674), .A3(new_n705), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n699), .A2(new_n715), .ZN(new_n716));
  XOR2_X1   g530(.A(KEYINPUT99), .B(G125), .Z(new_n717));
  XNOR2_X1  g531(.A(new_n716), .B(new_n717), .ZN(G27));
  INV_X1    g532(.A(new_n289), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n606), .B1(new_n579), .B2(new_n582), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n438), .A2(new_n719), .A3(new_n676), .A4(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT100), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n722), .A2(KEYINPUT42), .ZN(new_n723));
  AND2_X1   g537(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n722), .A2(KEYINPUT42), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n723), .B1(new_n721), .B2(new_n725), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(new_n234), .ZN(G33));
  NAND4_X1  g542(.A1(new_n438), .A2(new_n719), .A3(new_n647), .A4(new_n720), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G134), .ZN(G36));
  NAND2_X1  g544(.A1(new_n603), .A2(new_n534), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT43), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n731), .B(new_n732), .ZN(new_n733));
  AND4_X1   g547(.A1(new_n588), .A2(new_n733), .A3(new_n635), .A4(new_n630), .ZN(new_n734));
  OR2_X1    g548(.A1(new_n734), .A2(KEYINPUT44), .ZN(new_n735));
  INV_X1    g549(.A(new_n720), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n736), .B1(new_n734), .B2(KEYINPUT44), .ZN(new_n737));
  AND2_X1   g551(.A1(new_n282), .A2(new_n283), .ZN(new_n738));
  OAI21_X1  g552(.A(G469), .B1(new_n738), .B2(KEYINPUT45), .ZN(new_n739));
  OR2_X1    g553(.A1(new_n739), .A2(KEYINPUT101), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n738), .A2(KEYINPUT45), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n739), .A2(KEYINPUT101), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n740), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(new_n279), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT46), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n690), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n743), .A2(KEYINPUT46), .A3(new_n279), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n707), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n735), .A2(new_n737), .A3(new_n663), .A4(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(KEYINPUT102), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G137), .ZN(G39));
  INV_X1    g565(.A(KEYINPUT47), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n748), .B(new_n752), .ZN(new_n753));
  NOR4_X1   g567(.A1(new_n736), .A2(new_n683), .A3(new_n684), .A4(new_n674), .ZN(new_n754));
  XOR2_X1   g568(.A(new_n754), .B(KEYINPUT103), .Z(new_n755));
  OR2_X1    g569(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G140), .ZN(G42));
  INV_X1    g571(.A(new_n691), .ZN(new_n758));
  OR2_X1    g572(.A1(new_n758), .A2(KEYINPUT49), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(KEYINPUT49), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n362), .A2(new_n606), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n759), .A2(new_n760), .A3(new_n288), .A4(new_n761), .ZN(new_n762));
  NOR3_X1   g576(.A1(new_n762), .A2(new_n657), .A3(new_n731), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n652), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n636), .A2(new_n705), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(new_n676), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n720), .A2(new_n719), .ZN(new_n767));
  OAI21_X1  g581(.A(KEYINPUT107), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT107), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n715), .A2(new_n769), .A3(new_n719), .A4(new_n720), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  OAI211_X1 g585(.A(new_n771), .B(new_n729), .C1(new_n724), .C2(new_n726), .ZN(new_n772));
  NOR3_X1   g586(.A1(new_n736), .A2(new_n615), .A3(new_n646), .ZN(new_n773));
  AND3_X1   g587(.A1(new_n773), .A2(new_n671), .A3(new_n619), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  AOI22_X1  g589(.A1(new_n693), .A2(new_n609), .B1(new_n709), .B2(new_n712), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT104), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n776), .A2(new_n700), .A3(new_n777), .A4(new_n697), .ZN(new_n778));
  INV_X1    g592(.A(new_n621), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n438), .A2(new_n708), .ZN(new_n780));
  INV_X1    g594(.A(new_n637), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n683), .A2(new_n708), .A3(new_n607), .ZN(new_n782));
  OAI22_X1  g596(.A1(new_n779), .A2(new_n780), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n706), .A2(new_n525), .A3(new_n708), .ZN(new_n784));
  OAI22_X1  g598(.A1(new_n780), .A2(new_n608), .B1(new_n784), .B2(new_n711), .ZN(new_n785));
  OAI21_X1  g599(.A(KEYINPUT104), .B1(new_n783), .B2(new_n785), .ZN(new_n786));
  AND2_X1   g600(.A1(new_n778), .A2(new_n786), .ZN(new_n787));
  NOR3_X1   g601(.A1(new_n588), .A2(new_n362), .A3(new_n524), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n293), .A2(new_n583), .A3(new_n605), .A4(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT105), .ZN(new_n790));
  AND3_X1   g604(.A1(new_n584), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n790), .B1(new_n584), .B2(new_n789), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n590), .A2(new_n482), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n293), .A2(new_n583), .A3(new_n794), .A4(new_n788), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n639), .A2(new_n795), .ZN(new_n796));
  AOI21_X1  g610(.A(KEYINPUT106), .B1(new_n793), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n584), .A2(new_n789), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n798), .A2(KEYINPUT105), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n584), .A2(new_n789), .A3(new_n790), .ZN(new_n800));
  AND4_X1   g614(.A1(KEYINPUT106), .A2(new_n799), .A3(new_n796), .A4(new_n800), .ZN(new_n801));
  OAI211_X1 g615(.A(new_n775), .B(new_n787), .C1(new_n797), .C2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT108), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n793), .A2(KEYINPUT106), .A3(new_n796), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n799), .A2(new_n796), .A3(new_n800), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT106), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n805), .A2(new_n808), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n809), .A2(KEYINPUT108), .A3(new_n775), .A4(new_n787), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n648), .A2(new_n716), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n679), .A2(new_n811), .ZN(new_n812));
  NOR3_X1   g626(.A1(new_n634), .A2(new_n628), .A3(new_n646), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n712), .A2(new_n719), .A3(new_n657), .A4(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT52), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  AND2_X1   g631(.A1(new_n814), .A2(KEYINPUT52), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n812), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n804), .A2(new_n810), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n821), .A2(KEYINPUT53), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT109), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n811), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n648), .A2(new_n716), .A3(KEYINPUT109), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n679), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(new_n818), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT110), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n826), .A2(KEYINPUT110), .A3(new_n818), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n831), .A2(new_n817), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT53), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n832), .A2(new_n833), .A3(new_n804), .A4(new_n810), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n822), .A2(new_n834), .A3(KEYINPUT54), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n821), .A2(new_n833), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT54), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n776), .A2(new_n697), .A3(new_n700), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT111), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n833), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  OR2_X1    g654(.A1(new_n838), .A2(new_n839), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n809), .A2(new_n775), .A3(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n832), .A2(new_n840), .A3(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n836), .A2(new_n837), .A3(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT112), .ZN(new_n845));
  AND3_X1   g659(.A1(new_n835), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n845), .B1(new_n835), .B2(new_n844), .ZN(new_n847));
  AND2_X1   g661(.A1(new_n733), .A2(new_n644), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n848), .A2(new_n706), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n652), .A2(new_n849), .A3(new_n606), .A4(new_n708), .ZN(new_n850));
  XNOR2_X1  g664(.A(new_n850), .B(KEYINPUT50), .ZN(new_n851));
  INV_X1    g665(.A(new_n851), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n736), .A2(new_n692), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n848), .A2(new_n853), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n854), .A2(new_n636), .A3(new_n705), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n853), .A2(new_n684), .A3(new_n518), .A4(new_n658), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n856), .A2(new_n590), .A3(new_n603), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  OR2_X1    g672(.A1(new_n858), .A2(KEYINPUT113), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(KEYINPUT113), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n852), .A2(KEYINPUT114), .A3(new_n859), .A4(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT114), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n859), .A2(new_n860), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n862), .B1(new_n863), .B2(new_n851), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n753), .B1(new_n288), .B2(new_n758), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n865), .A2(new_n720), .A3(new_n849), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n861), .A2(new_n864), .A3(KEYINPUT51), .A4(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n849), .A2(new_n607), .A3(new_n708), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n866), .A2(new_n852), .A3(new_n858), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT51), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n854), .A2(new_n685), .ZN(new_n872));
  AND2_X1   g686(.A1(new_n872), .A2(KEYINPUT48), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n872), .A2(KEYINPUT48), .ZN(new_n874));
  XOR2_X1   g688(.A(new_n517), .B(KEYINPUT115), .Z(new_n875));
  OAI21_X1  g689(.A(new_n875), .B1(new_n856), .B2(new_n604), .ZN(new_n876));
  NOR3_X1   g690(.A1(new_n873), .A2(new_n874), .A3(new_n876), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n867), .A2(new_n868), .A3(new_n871), .A4(new_n877), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n846), .A2(new_n847), .A3(new_n878), .ZN(new_n879));
  NOR2_X1   g693(.A1(G952), .A2(G953), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n764), .B1(new_n879), .B2(new_n880), .ZN(G75));
  INV_X1    g695(.A(KEYINPUT56), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n836), .A2(new_n843), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n883), .A2(G902), .ZN(new_n884));
  INV_X1    g698(.A(G210), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n882), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n554), .B(new_n559), .ZN(new_n887));
  XOR2_X1   g701(.A(new_n887), .B(KEYINPUT55), .Z(new_n888));
  OAI21_X1  g702(.A(new_n888), .B1(KEYINPUT116), .B2(KEYINPUT56), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n886), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n270), .A2(G952), .ZN(new_n891));
  INV_X1    g705(.A(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(new_n889), .ZN(new_n893));
  OAI211_X1 g707(.A(new_n882), .B(new_n893), .C1(new_n884), .C2(new_n885), .ZN(new_n894));
  AND3_X1   g708(.A1(new_n890), .A2(new_n892), .A3(new_n894), .ZN(G51));
  XOR2_X1   g709(.A(new_n279), .B(KEYINPUT57), .Z(new_n896));
  INV_X1    g710(.A(new_n844), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n837), .B1(new_n836), .B2(new_n843), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n896), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n688), .B(KEYINPUT117), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  OR2_X1    g715(.A1(new_n884), .A2(new_n743), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n891), .B1(new_n901), .B2(new_n902), .ZN(G54));
  NAND4_X1  g717(.A1(new_n883), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n502), .A2(new_n506), .ZN(new_n905));
  AND2_X1   g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n904), .A2(new_n905), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n906), .A2(new_n907), .A3(new_n891), .ZN(G60));
  NAND3_X1  g722(.A1(new_n594), .A2(new_n599), .A3(new_n595), .ZN(new_n909));
  NAND2_X1  g723(.A1(G478), .A2(G902), .ZN(new_n910));
  XOR2_X1   g724(.A(new_n910), .B(KEYINPUT59), .Z(new_n911));
  NOR2_X1   g725(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n912), .B1(new_n897), .B2(new_n898), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(new_n892), .ZN(new_n914));
  INV_X1    g728(.A(new_n911), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n915), .B1(new_n846), .B2(new_n847), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n914), .B1(new_n916), .B2(new_n909), .ZN(G63));
  INV_X1    g731(.A(KEYINPUT61), .ZN(new_n918));
  AND2_X1   g732(.A1(new_n832), .A2(new_n840), .ZN(new_n919));
  AOI22_X1  g733(.A1(new_n919), .A2(new_n842), .B1(new_n833), .B2(new_n821), .ZN(new_n920));
  NAND2_X1  g734(.A1(G217), .A2(G902), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(KEYINPUT60), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n359), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(new_n892), .ZN(new_n924));
  INV_X1    g738(.A(new_n922), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n883), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n926), .A2(new_n627), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n918), .B1(new_n924), .B2(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n891), .B1(new_n926), .B2(new_n359), .ZN(new_n929));
  OAI211_X1 g743(.A(new_n929), .B(KEYINPUT61), .C1(new_n627), .C2(new_n926), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n928), .A2(new_n930), .ZN(G66));
  NAND2_X1  g745(.A1(new_n809), .A2(new_n787), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(new_n270), .ZN(new_n933));
  OAI21_X1  g747(.A(G953), .B1(new_n520), .B2(new_n557), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(new_n554), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n936), .B1(G898), .B2(new_n270), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n935), .B(new_n937), .ZN(G69));
  NAND2_X1  g752(.A1(new_n374), .A2(new_n380), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n939), .B(KEYINPUT120), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(new_n503), .ZN(new_n941));
  XNOR2_X1  g755(.A(KEYINPUT118), .B(KEYINPUT119), .ZN(new_n942));
  XOR2_X1   g756(.A(new_n941), .B(new_n942), .Z(new_n943));
  INV_X1    g757(.A(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n270), .B1(new_n944), .B2(KEYINPUT124), .ZN(new_n945));
  NAND2_X1  g759(.A1(G227), .A2(G900), .ZN(new_n946));
  AND2_X1   g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n438), .B1(new_n605), .B2(new_n794), .ZN(new_n949));
  OR3_X1    g763(.A1(new_n665), .A2(new_n736), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n749), .A2(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT121), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n951), .B(new_n952), .ZN(new_n953));
  AOI21_X1  g767(.A(KEYINPUT62), .B1(new_n669), .B2(new_n826), .ZN(new_n954));
  AND3_X1   g768(.A1(new_n669), .A2(KEYINPUT62), .A3(new_n826), .ZN(new_n955));
  OAI211_X1 g769(.A(new_n953), .B(new_n756), .C1(new_n954), .C2(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n944), .B1(new_n956), .B2(new_n270), .ZN(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n270), .A2(G900), .ZN(new_n959));
  NAND4_X1  g773(.A1(new_n748), .A2(new_n438), .A3(new_n663), .A4(new_n712), .ZN(new_n960));
  OAI211_X1 g774(.A(new_n960), .B(new_n729), .C1(new_n724), .C2(new_n726), .ZN(new_n961));
  INV_X1    g775(.A(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(KEYINPUT122), .ZN(new_n963));
  AND3_X1   g777(.A1(new_n749), .A2(new_n963), .A3(new_n826), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n963), .B1(new_n749), .B2(new_n826), .ZN(new_n965));
  OAI211_X1 g779(.A(new_n756), .B(new_n962), .C1(new_n964), .C2(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n959), .B1(new_n966), .B2(new_n270), .ZN(new_n967));
  OR2_X1    g781(.A1(new_n967), .A2(KEYINPUT123), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n967), .A2(KEYINPUT123), .ZN(new_n969));
  AND2_X1   g783(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  OAI211_X1 g784(.A(new_n948), .B(new_n958), .C1(new_n970), .C2(new_n943), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n943), .B1(new_n968), .B2(new_n969), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n947), .B1(new_n972), .B2(new_n957), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n971), .A2(new_n973), .ZN(G72));
  NAND2_X1  g788(.A1(G472), .A2(G902), .ZN(new_n975));
  XOR2_X1   g789(.A(new_n975), .B(KEYINPUT63), .Z(new_n976));
  XOR2_X1   g790(.A(new_n976), .B(KEYINPUT125), .Z(new_n977));
  OAI21_X1  g791(.A(new_n977), .B1(new_n966), .B2(new_n932), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n390), .A2(new_n398), .ZN(new_n979));
  XOR2_X1   g793(.A(new_n979), .B(KEYINPUT126), .Z(new_n980));
  NAND3_X1  g794(.A1(new_n978), .A2(new_n406), .A3(new_n980), .ZN(new_n981));
  AND2_X1   g795(.A1(new_n981), .A2(new_n892), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n977), .B1(new_n956), .B2(new_n932), .ZN(new_n983));
  INV_X1    g797(.A(new_n980), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n983), .A2(new_n396), .A3(new_n984), .ZN(new_n985));
  OR2_X1    g799(.A1(new_n654), .A2(new_n435), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n822), .A2(new_n834), .A3(new_n976), .A4(new_n986), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n982), .A2(new_n985), .A3(new_n987), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n988), .A2(KEYINPUT127), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT127), .ZN(new_n990));
  NAND4_X1  g804(.A1(new_n982), .A2(new_n985), .A3(new_n990), .A4(new_n987), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n989), .A2(new_n991), .ZN(G57));
endmodule


