

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590;

  XOR2_X2 U321 ( .A(n463), .B(KEYINPUT41), .Z(n574) );
  XOR2_X1 U322 ( .A(G99GAT), .B(G85GAT), .Z(n441) );
  INV_X1 U323 ( .A(KEYINPUT117), .ZN(n460) );
  AND2_X1 U324 ( .A1(n380), .A2(n379), .ZN(n381) );
  NOR2_X1 U325 ( .A1(n529), .A2(n378), .ZN(n379) );
  XNOR2_X1 U326 ( .A(G211GAT), .B(KEYINPUT89), .ZN(n340) );
  XOR2_X1 U327 ( .A(n452), .B(n451), .Z(n581) );
  INV_X1 U328 ( .A(n544), .ZN(n536) );
  INV_X1 U329 ( .A(n543), .ZN(n378) );
  NOR2_X1 U330 ( .A1(n489), .A2(n543), .ZN(n578) );
  AND2_X1 U331 ( .A1(G228GAT), .A2(G233GAT), .ZN(n289) );
  XOR2_X1 U332 ( .A(n354), .B(n353), .Z(n290) );
  XNOR2_X1 U333 ( .A(n425), .B(n289), .ZN(n349) );
  XNOR2_X1 U334 ( .A(KEYINPUT75), .B(KEYINPUT31), .ZN(n436) );
  XNOR2_X1 U335 ( .A(n350), .B(n349), .ZN(n352) );
  XNOR2_X1 U336 ( .A(n437), .B(n436), .ZN(n440) );
  INV_X1 U337 ( .A(KEYINPUT10), .ZN(n396) );
  XNOR2_X1 U338 ( .A(n355), .B(n290), .ZN(n359) );
  XNOR2_X1 U339 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U340 ( .A(n397), .B(n396), .ZN(n402) );
  XNOR2_X1 U341 ( .A(n359), .B(n358), .ZN(n487) );
  XNOR2_X1 U342 ( .A(n447), .B(n446), .ZN(n450) );
  XNOR2_X1 U343 ( .A(n402), .B(n401), .ZN(n406) );
  XOR2_X1 U344 ( .A(n554), .B(n413), .Z(n588) );
  XNOR2_X1 U345 ( .A(n361), .B(KEYINPUT67), .ZN(n544) );
  XOR2_X1 U346 ( .A(n412), .B(n411), .Z(n554) );
  INV_X1 U347 ( .A(G43GAT), .ZN(n482) );
  XNOR2_X1 U348 ( .A(n476), .B(G197GAT), .ZN(n477) );
  XNOR2_X1 U349 ( .A(n482), .B(KEYINPUT40), .ZN(n483) );
  XNOR2_X1 U350 ( .A(n478), .B(n477), .ZN(G1352GAT) );
  XNOR2_X1 U351 ( .A(n484), .B(n483), .ZN(G1330GAT) );
  XOR2_X1 U352 ( .A(G85GAT), .B(G120GAT), .Z(n292) );
  XNOR2_X1 U353 ( .A(G29GAT), .B(G134GAT), .ZN(n291) );
  XNOR2_X1 U354 ( .A(n292), .B(n291), .ZN(n296) );
  XOR2_X1 U355 ( .A(G57GAT), .B(G148GAT), .Z(n294) );
  XNOR2_X1 U356 ( .A(G141GAT), .B(G1GAT), .ZN(n293) );
  XNOR2_X1 U357 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U358 ( .A(n296), .B(n295), .Z(n301) );
  XOR2_X1 U359 ( .A(KEYINPUT93), .B(KEYINPUT92), .Z(n298) );
  NAND2_X1 U360 ( .A1(G225GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U361 ( .A(n298), .B(n297), .ZN(n299) );
  XNOR2_X1 U362 ( .A(KEYINPUT91), .B(n299), .ZN(n300) );
  XNOR2_X1 U363 ( .A(n301), .B(n300), .ZN(n305) );
  XOR2_X1 U364 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n303) );
  XNOR2_X1 U365 ( .A(KEYINPUT4), .B(KEYINPUT5), .ZN(n302) );
  XNOR2_X1 U366 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U367 ( .A(n305), .B(n304), .Z(n311) );
  XOR2_X1 U368 ( .A(G127GAT), .B(KEYINPUT0), .Z(n307) );
  XNOR2_X1 U369 ( .A(G113GAT), .B(KEYINPUT81), .ZN(n306) );
  XNOR2_X1 U370 ( .A(n307), .B(n306), .ZN(n367) );
  XOR2_X1 U371 ( .A(G155GAT), .B(KEYINPUT2), .Z(n309) );
  XNOR2_X1 U372 ( .A(G162GAT), .B(KEYINPUT3), .ZN(n308) );
  XNOR2_X1 U373 ( .A(n309), .B(n308), .ZN(n356) );
  XNOR2_X1 U374 ( .A(n367), .B(n356), .ZN(n310) );
  XOR2_X1 U375 ( .A(n311), .B(n310), .Z(n541) );
  INV_X1 U376 ( .A(n541), .ZN(n529) );
  XNOR2_X1 U377 ( .A(KEYINPUT37), .B(KEYINPUT105), .ZN(n416) );
  XOR2_X1 U378 ( .A(G78GAT), .B(G155GAT), .Z(n313) );
  XNOR2_X1 U379 ( .A(G8GAT), .B(G211GAT), .ZN(n312) );
  XNOR2_X1 U380 ( .A(n313), .B(n312), .ZN(n317) );
  XOR2_X1 U381 ( .A(KEYINPUT12), .B(KEYINPUT79), .Z(n315) );
  XNOR2_X1 U382 ( .A(G64GAT), .B(KEYINPUT15), .ZN(n314) );
  XNOR2_X1 U383 ( .A(n315), .B(n314), .ZN(n316) );
  XNOR2_X1 U384 ( .A(n317), .B(n316), .ZN(n328) );
  XOR2_X1 U385 ( .A(G15GAT), .B(G1GAT), .Z(n421) );
  XOR2_X1 U386 ( .A(G71GAT), .B(G127GAT), .Z(n319) );
  XNOR2_X1 U387 ( .A(G22GAT), .B(G183GAT), .ZN(n318) );
  XNOR2_X1 U388 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U389 ( .A(n421), .B(n320), .Z(n322) );
  NAND2_X1 U390 ( .A1(G231GAT), .A2(G233GAT), .ZN(n321) );
  XNOR2_X1 U391 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U392 ( .A(n323), .B(KEYINPUT80), .Z(n326) );
  XNOR2_X1 U393 ( .A(G57GAT), .B(KEYINPUT74), .ZN(n324) );
  XNOR2_X1 U394 ( .A(n324), .B(KEYINPUT13), .ZN(n434) );
  XNOR2_X1 U395 ( .A(n434), .B(KEYINPUT14), .ZN(n325) );
  XNOR2_X1 U396 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U397 ( .A(n328), .B(n327), .Z(n585) );
  INV_X1 U398 ( .A(n585), .ZN(n577) );
  XOR2_X1 U399 ( .A(G169GAT), .B(G8GAT), .Z(n422) );
  XOR2_X1 U400 ( .A(G64GAT), .B(G92GAT), .Z(n330) );
  XNOR2_X1 U401 ( .A(G176GAT), .B(G204GAT), .ZN(n329) );
  XNOR2_X1 U402 ( .A(n330), .B(n329), .ZN(n435) );
  XOR2_X1 U403 ( .A(n422), .B(n435), .Z(n332) );
  NAND2_X1 U404 ( .A1(G226GAT), .A2(G233GAT), .ZN(n331) );
  XNOR2_X1 U405 ( .A(n332), .B(n331), .ZN(n336) );
  XOR2_X1 U406 ( .A(KEYINPUT94), .B(KEYINPUT95), .Z(n334) );
  XNOR2_X1 U407 ( .A(G36GAT), .B(G190GAT), .ZN(n333) );
  XNOR2_X1 U408 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U409 ( .A(n336), .B(n335), .Z(n345) );
  XOR2_X1 U410 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n338) );
  XNOR2_X1 U411 ( .A(KEYINPUT85), .B(G183GAT), .ZN(n337) );
  XNOR2_X1 U412 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U413 ( .A(KEYINPUT17), .B(n339), .Z(n375) );
  XNOR2_X1 U414 ( .A(n340), .B(KEYINPUT21), .ZN(n341) );
  XOR2_X1 U415 ( .A(n341), .B(KEYINPUT90), .Z(n343) );
  XNOR2_X1 U416 ( .A(G197GAT), .B(G218GAT), .ZN(n342) );
  XNOR2_X1 U417 ( .A(n343), .B(n342), .ZN(n357) );
  XNOR2_X1 U418 ( .A(n375), .B(n357), .ZN(n344) );
  XNOR2_X1 U419 ( .A(n345), .B(n344), .ZN(n531) );
  XNOR2_X1 U420 ( .A(n531), .B(KEYINPUT96), .ZN(n346) );
  XNOR2_X1 U421 ( .A(n346), .B(KEYINPUT27), .ZN(n540) );
  XOR2_X1 U422 ( .A(KEYINPUT88), .B(KEYINPUT87), .Z(n348) );
  XNOR2_X1 U423 ( .A(G50GAT), .B(KEYINPUT22), .ZN(n347) );
  XNOR2_X1 U424 ( .A(n348), .B(n347), .ZN(n350) );
  XOR2_X1 U425 ( .A(G141GAT), .B(G22GAT), .Z(n425) );
  XNOR2_X1 U426 ( .A(G106GAT), .B(G78GAT), .ZN(n351) );
  XNOR2_X1 U427 ( .A(n351), .B(G148GAT), .ZN(n448) );
  XOR2_X1 U428 ( .A(n352), .B(n448), .Z(n355) );
  XOR2_X1 U429 ( .A(KEYINPUT86), .B(KEYINPUT23), .Z(n354) );
  XNOR2_X1 U430 ( .A(G204GAT), .B(KEYINPUT24), .ZN(n353) );
  XNOR2_X1 U431 ( .A(n357), .B(n356), .ZN(n358) );
  INV_X1 U432 ( .A(KEYINPUT28), .ZN(n360) );
  XNOR2_X1 U433 ( .A(n487), .B(n360), .ZN(n361) );
  NOR2_X1 U434 ( .A1(n540), .A2(n544), .ZN(n380) );
  XOR2_X1 U435 ( .A(KEYINPUT65), .B(G99GAT), .Z(n363) );
  XNOR2_X1 U436 ( .A(G43GAT), .B(G15GAT), .ZN(n362) );
  XNOR2_X1 U437 ( .A(n363), .B(n362), .ZN(n364) );
  XOR2_X1 U438 ( .A(n364), .B(G176GAT), .Z(n366) );
  XOR2_X1 U439 ( .A(G120GAT), .B(G71GAT), .Z(n437) );
  XNOR2_X1 U440 ( .A(G169GAT), .B(n437), .ZN(n365) );
  XNOR2_X1 U441 ( .A(n366), .B(n365), .ZN(n371) );
  XOR2_X1 U442 ( .A(G190GAT), .B(G134GAT), .Z(n398) );
  XOR2_X1 U443 ( .A(n367), .B(n398), .Z(n369) );
  NAND2_X1 U444 ( .A1(G227GAT), .A2(G233GAT), .ZN(n368) );
  XNOR2_X1 U445 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U446 ( .A(n371), .B(n370), .Z(n377) );
  XOR2_X1 U447 ( .A(KEYINPUT83), .B(KEYINPUT82), .Z(n373) );
  XNOR2_X1 U448 ( .A(KEYINPUT84), .B(KEYINPUT20), .ZN(n372) );
  XNOR2_X1 U449 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U450 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U451 ( .A(n377), .B(n376), .ZN(n543) );
  XNOR2_X1 U452 ( .A(n381), .B(KEYINPUT97), .ZN(n391) );
  NAND2_X1 U453 ( .A1(n487), .A2(n543), .ZN(n382) );
  XNOR2_X1 U454 ( .A(n382), .B(KEYINPUT98), .ZN(n383) );
  XNOR2_X1 U455 ( .A(KEYINPUT26), .B(n383), .ZN(n559) );
  NOR2_X1 U456 ( .A1(n540), .A2(n559), .ZN(n384) );
  XNOR2_X1 U457 ( .A(KEYINPUT99), .B(n384), .ZN(n388) );
  NOR2_X1 U458 ( .A1(n543), .A2(n531), .ZN(n385) );
  NOR2_X1 U459 ( .A1(n487), .A2(n385), .ZN(n386) );
  XNOR2_X1 U460 ( .A(KEYINPUT25), .B(n386), .ZN(n387) );
  NAND2_X1 U461 ( .A1(n388), .A2(n387), .ZN(n389) );
  NAND2_X1 U462 ( .A1(n529), .A2(n389), .ZN(n390) );
  NAND2_X1 U463 ( .A1(n391), .A2(n390), .ZN(n392) );
  XOR2_X1 U464 ( .A(KEYINPUT100), .B(n392), .Z(n499) );
  NOR2_X1 U465 ( .A1(n577), .A2(n499), .ZN(n414) );
  XOR2_X1 U466 ( .A(KEYINPUT76), .B(G92GAT), .Z(n394) );
  XNOR2_X1 U467 ( .A(G162GAT), .B(G106GAT), .ZN(n393) );
  XNOR2_X1 U468 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U469 ( .A(G218GAT), .B(n395), .ZN(n397) );
  XOR2_X1 U470 ( .A(KEYINPUT78), .B(KEYINPUT77), .Z(n400) );
  XNOR2_X1 U471 ( .A(n398), .B(n441), .ZN(n399) );
  XNOR2_X1 U472 ( .A(n400), .B(n399), .ZN(n401) );
  XOR2_X1 U473 ( .A(KEYINPUT66), .B(KEYINPUT11), .Z(n404) );
  NAND2_X1 U474 ( .A1(G232GAT), .A2(G233GAT), .ZN(n403) );
  XNOR2_X1 U475 ( .A(n404), .B(n403), .ZN(n405) );
  XOR2_X1 U476 ( .A(n406), .B(n405), .Z(n412) );
  XNOR2_X1 U477 ( .A(G36GAT), .B(KEYINPUT7), .ZN(n407) );
  XNOR2_X1 U478 ( .A(n407), .B(G29GAT), .ZN(n408) );
  XOR2_X1 U479 ( .A(n408), .B(KEYINPUT8), .Z(n410) );
  XNOR2_X1 U480 ( .A(G43GAT), .B(G50GAT), .ZN(n409) );
  XNOR2_X1 U481 ( .A(n410), .B(n409), .ZN(n420) );
  XNOR2_X1 U482 ( .A(n420), .B(KEYINPUT9), .ZN(n411) );
  XOR2_X1 U483 ( .A(KEYINPUT36), .B(KEYINPUT104), .Z(n413) );
  NAND2_X1 U484 ( .A1(n414), .A2(n588), .ZN(n415) );
  XOR2_X1 U485 ( .A(n416), .B(n415), .Z(n528) );
  XOR2_X1 U486 ( .A(KEYINPUT71), .B(KEYINPUT30), .Z(n418) );
  XNOR2_X1 U487 ( .A(KEYINPUT68), .B(KEYINPUT29), .ZN(n417) );
  XNOR2_X1 U488 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U489 ( .A(n420), .B(n419), .ZN(n433) );
  XOR2_X1 U490 ( .A(G197GAT), .B(G113GAT), .Z(n424) );
  XNOR2_X1 U491 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U492 ( .A(n424), .B(n423), .ZN(n426) );
  XOR2_X1 U493 ( .A(n426), .B(n425), .Z(n431) );
  XOR2_X1 U494 ( .A(KEYINPUT69), .B(KEYINPUT72), .Z(n428) );
  NAND2_X1 U495 ( .A1(G229GAT), .A2(G233GAT), .ZN(n427) );
  XNOR2_X1 U496 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U497 ( .A(KEYINPUT70), .B(n429), .ZN(n430) );
  XNOR2_X1 U498 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U499 ( .A(n433), .B(n432), .ZN(n560) );
  XNOR2_X1 U500 ( .A(n560), .B(KEYINPUT73), .ZN(n546) );
  XNOR2_X1 U501 ( .A(n435), .B(n434), .ZN(n452) );
  INV_X1 U502 ( .A(n441), .ZN(n439) );
  INV_X1 U503 ( .A(n440), .ZN(n438) );
  NAND2_X1 U504 ( .A1(n439), .A2(n438), .ZN(n443) );
  NAND2_X1 U505 ( .A1(n441), .A2(n440), .ZN(n442) );
  NAND2_X1 U506 ( .A1(n443), .A2(n442), .ZN(n447) );
  AND2_X1 U507 ( .A1(G230GAT), .A2(G233GAT), .ZN(n445) );
  INV_X1 U508 ( .A(KEYINPUT33), .ZN(n444) );
  XNOR2_X1 U509 ( .A(n448), .B(KEYINPUT32), .ZN(n449) );
  XNOR2_X1 U510 ( .A(n450), .B(n449), .ZN(n451) );
  AND2_X1 U511 ( .A1(n546), .A2(n581), .ZN(n500) );
  AND2_X1 U512 ( .A1(n528), .A2(n500), .ZN(n453) );
  XOR2_X1 U513 ( .A(KEYINPUT38), .B(n453), .Z(n511) );
  NOR2_X1 U514 ( .A1(n529), .A2(n511), .ZN(n455) );
  XNOR2_X1 U515 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n454) );
  XNOR2_X1 U516 ( .A(n455), .B(n454), .ZN(G1328GAT) );
  XOR2_X1 U517 ( .A(KEYINPUT45), .B(KEYINPUT116), .Z(n457) );
  NAND2_X1 U518 ( .A1(n577), .A2(n588), .ZN(n456) );
  XNOR2_X1 U519 ( .A(n457), .B(n456), .ZN(n458) );
  NAND2_X1 U520 ( .A1(n458), .A2(n581), .ZN(n459) );
  NOR2_X1 U521 ( .A1(n546), .A2(n459), .ZN(n461) );
  XNOR2_X1 U522 ( .A(n461), .B(n460), .ZN(n471) );
  INV_X1 U523 ( .A(KEYINPUT64), .ZN(n462) );
  XNOR2_X1 U524 ( .A(n581), .B(n462), .ZN(n463) );
  INV_X1 U525 ( .A(n574), .ZN(n564) );
  NOR2_X1 U526 ( .A1(n564), .A2(n560), .ZN(n464) );
  XNOR2_X1 U527 ( .A(n464), .B(KEYINPUT114), .ZN(n465) );
  XNOR2_X1 U528 ( .A(KEYINPUT46), .B(n465), .ZN(n467) );
  INV_X1 U529 ( .A(n554), .ZN(n569) );
  OR2_X1 U530 ( .A1(n577), .A2(n554), .ZN(n466) );
  OR2_X1 U531 ( .A1(n467), .A2(n466), .ZN(n469) );
  XOR2_X1 U532 ( .A(KEYINPUT115), .B(KEYINPUT47), .Z(n468) );
  XNOR2_X1 U533 ( .A(n469), .B(n468), .ZN(n470) );
  NOR2_X1 U534 ( .A1(n471), .A2(n470), .ZN(n472) );
  XNOR2_X1 U535 ( .A(KEYINPUT48), .B(n472), .ZN(n539) );
  NOR2_X1 U536 ( .A1(n531), .A2(n539), .ZN(n473) );
  XNOR2_X1 U537 ( .A(n473), .B(KEYINPUT54), .ZN(n485) );
  NOR2_X1 U538 ( .A1(n559), .A2(n541), .ZN(n474) );
  AND2_X1 U539 ( .A1(n485), .A2(n474), .ZN(n475) );
  XOR2_X1 U540 ( .A(KEYINPUT127), .B(n475), .Z(n587) );
  INV_X1 U541 ( .A(n587), .ZN(n584) );
  NOR2_X1 U542 ( .A1(n584), .A2(n560), .ZN(n478) );
  XNOR2_X1 U543 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n476) );
  NOR2_X1 U544 ( .A1(n531), .A2(n511), .ZN(n481) );
  INV_X1 U545 ( .A(G36GAT), .ZN(n479) );
  XNOR2_X1 U546 ( .A(n479), .B(KEYINPUT106), .ZN(n480) );
  XNOR2_X1 U547 ( .A(n481), .B(n480), .ZN(G1329GAT) );
  NOR2_X1 U548 ( .A1(n543), .A2(n511), .ZN(n484) );
  NAND2_X1 U549 ( .A1(n485), .A2(n529), .ZN(n486) );
  NOR2_X1 U550 ( .A1(n487), .A2(n486), .ZN(n488) );
  XNOR2_X1 U551 ( .A(n488), .B(KEYINPUT55), .ZN(n489) );
  NAND2_X1 U552 ( .A1(n578), .A2(n554), .ZN(n493) );
  XOR2_X1 U553 ( .A(KEYINPUT58), .B(KEYINPUT126), .Z(n491) );
  INV_X1 U554 ( .A(G190GAT), .ZN(n490) );
  XNOR2_X1 U555 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U556 ( .A(n493), .B(n492), .ZN(G1351GAT) );
  NAND2_X1 U557 ( .A1(n578), .A2(n546), .ZN(n496) );
  XOR2_X1 U558 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n494) );
  XNOR2_X1 U559 ( .A(n494), .B(G169GAT), .ZN(n495) );
  XNOR2_X1 U560 ( .A(n496), .B(n495), .ZN(G1348GAT) );
  NOR2_X1 U561 ( .A1(n554), .A2(n585), .ZN(n497) );
  XOR2_X1 U562 ( .A(KEYINPUT16), .B(n497), .Z(n498) );
  NOR2_X1 U563 ( .A1(n499), .A2(n498), .ZN(n516) );
  NAND2_X1 U564 ( .A1(n500), .A2(n516), .ZN(n509) );
  NOR2_X1 U565 ( .A1(n529), .A2(n509), .ZN(n502) );
  XNOR2_X1 U566 ( .A(KEYINPUT34), .B(KEYINPUT101), .ZN(n501) );
  XNOR2_X1 U567 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U568 ( .A(G1GAT), .B(n503), .ZN(G1324GAT) );
  NOR2_X1 U569 ( .A1(n531), .A2(n509), .ZN(n504) );
  XOR2_X1 U570 ( .A(G8GAT), .B(n504), .Z(G1325GAT) );
  NOR2_X1 U571 ( .A1(n509), .A2(n543), .ZN(n508) );
  XOR2_X1 U572 ( .A(KEYINPUT102), .B(KEYINPUT103), .Z(n506) );
  XNOR2_X1 U573 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n505) );
  XNOR2_X1 U574 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U575 ( .A(n508), .B(n507), .ZN(G1326GAT) );
  NOR2_X1 U576 ( .A1(n536), .A2(n509), .ZN(n510) );
  XOR2_X1 U577 ( .A(G22GAT), .B(n510), .Z(G1327GAT) );
  NOR2_X1 U578 ( .A1(n536), .A2(n511), .ZN(n512) );
  XOR2_X1 U579 ( .A(G50GAT), .B(n512), .Z(G1331GAT) );
  XOR2_X1 U580 ( .A(KEYINPUT109), .B(KEYINPUT42), .Z(n514) );
  XNOR2_X1 U581 ( .A(G57GAT), .B(KEYINPUT108), .ZN(n513) );
  XNOR2_X1 U582 ( .A(n514), .B(n513), .ZN(n518) );
  NAND2_X1 U583 ( .A1(n574), .A2(n560), .ZN(n515) );
  XNOR2_X1 U584 ( .A(KEYINPUT107), .B(n515), .ZN(n527) );
  NAND2_X1 U585 ( .A1(n527), .A2(n516), .ZN(n523) );
  NOR2_X1 U586 ( .A1(n529), .A2(n523), .ZN(n517) );
  XOR2_X1 U587 ( .A(n518), .B(n517), .Z(G1332GAT) );
  NOR2_X1 U588 ( .A1(n531), .A2(n523), .ZN(n519) );
  XOR2_X1 U589 ( .A(KEYINPUT110), .B(n519), .Z(n520) );
  XNOR2_X1 U590 ( .A(G64GAT), .B(n520), .ZN(G1333GAT) );
  NOR2_X1 U591 ( .A1(n543), .A2(n523), .ZN(n522) );
  XNOR2_X1 U592 ( .A(G71GAT), .B(KEYINPUT111), .ZN(n521) );
  XNOR2_X1 U593 ( .A(n522), .B(n521), .ZN(G1334GAT) );
  NOR2_X1 U594 ( .A1(n536), .A2(n523), .ZN(n525) );
  XNOR2_X1 U595 ( .A(KEYINPUT112), .B(KEYINPUT43), .ZN(n524) );
  XNOR2_X1 U596 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U597 ( .A(G78GAT), .B(n526), .ZN(G1335GAT) );
  NAND2_X1 U598 ( .A1(n528), .A2(n527), .ZN(n535) );
  NOR2_X1 U599 ( .A1(n529), .A2(n535), .ZN(n530) );
  XOR2_X1 U600 ( .A(G85GAT), .B(n530), .Z(G1336GAT) );
  NOR2_X1 U601 ( .A1(n531), .A2(n535), .ZN(n532) );
  XOR2_X1 U602 ( .A(G92GAT), .B(n532), .Z(G1337GAT) );
  NOR2_X1 U603 ( .A1(n543), .A2(n535), .ZN(n534) );
  XNOR2_X1 U604 ( .A(G99GAT), .B(KEYINPUT113), .ZN(n533) );
  XNOR2_X1 U605 ( .A(n534), .B(n533), .ZN(G1338GAT) );
  NOR2_X1 U606 ( .A1(n536), .A2(n535), .ZN(n537) );
  XOR2_X1 U607 ( .A(KEYINPUT44), .B(n537), .Z(n538) );
  XNOR2_X1 U608 ( .A(G106GAT), .B(n538), .ZN(G1339GAT) );
  XOR2_X1 U609 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n548) );
  NOR2_X1 U610 ( .A1(n540), .A2(n539), .ZN(n542) );
  NAND2_X1 U611 ( .A1(n542), .A2(n541), .ZN(n558) );
  OR2_X1 U612 ( .A1(n544), .A2(n543), .ZN(n545) );
  NOR2_X1 U613 ( .A1(n558), .A2(n545), .ZN(n555) );
  NAND2_X1 U614 ( .A1(n555), .A2(n546), .ZN(n547) );
  XNOR2_X1 U615 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U616 ( .A(G113GAT), .B(n549), .ZN(G1340GAT) );
  XOR2_X1 U617 ( .A(G120GAT), .B(KEYINPUT49), .Z(n551) );
  NAND2_X1 U618 ( .A1(n555), .A2(n574), .ZN(n550) );
  XNOR2_X1 U619 ( .A(n551), .B(n550), .ZN(G1341GAT) );
  NAND2_X1 U620 ( .A1(n555), .A2(n577), .ZN(n552) );
  XNOR2_X1 U621 ( .A(n552), .B(KEYINPUT50), .ZN(n553) );
  XNOR2_X1 U622 ( .A(G127GAT), .B(n553), .ZN(G1342GAT) );
  XOR2_X1 U623 ( .A(G134GAT), .B(KEYINPUT51), .Z(n557) );
  NAND2_X1 U624 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U625 ( .A(n557), .B(n556), .ZN(G1343GAT) );
  OR2_X1 U626 ( .A1(n559), .A2(n558), .ZN(n568) );
  NOR2_X1 U627 ( .A1(n560), .A2(n568), .ZN(n561) );
  XOR2_X1 U628 ( .A(G141GAT), .B(n561), .Z(G1344GAT) );
  XOR2_X1 U629 ( .A(KEYINPUT52), .B(KEYINPUT120), .Z(n563) );
  XNOR2_X1 U630 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n562) );
  XNOR2_X1 U631 ( .A(n563), .B(n562), .ZN(n566) );
  NOR2_X1 U632 ( .A1(n564), .A2(n568), .ZN(n565) );
  XOR2_X1 U633 ( .A(n566), .B(n565), .Z(G1345GAT) );
  NOR2_X1 U634 ( .A1(n585), .A2(n568), .ZN(n567) );
  XOR2_X1 U635 ( .A(G155GAT), .B(n567), .Z(G1346GAT) );
  NOR2_X1 U636 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U637 ( .A(G162GAT), .B(n570), .Z(G1347GAT) );
  XOR2_X1 U638 ( .A(KEYINPUT57), .B(KEYINPUT124), .Z(n572) );
  XNOR2_X1 U639 ( .A(G176GAT), .B(KEYINPUT123), .ZN(n571) );
  XNOR2_X1 U640 ( .A(n572), .B(n571), .ZN(n573) );
  XOR2_X1 U641 ( .A(KEYINPUT56), .B(n573), .Z(n576) );
  NAND2_X1 U642 ( .A1(n574), .A2(n578), .ZN(n575) );
  XNOR2_X1 U643 ( .A(n576), .B(n575), .ZN(G1349GAT) );
  XOR2_X1 U644 ( .A(G183GAT), .B(KEYINPUT125), .Z(n580) );
  NAND2_X1 U645 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U646 ( .A(n580), .B(n579), .ZN(G1350GAT) );
  NOR2_X1 U647 ( .A1(n584), .A2(n581), .ZN(n583) );
  XNOR2_X1 U648 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n582) );
  XNOR2_X1 U649 ( .A(n583), .B(n582), .ZN(G1353GAT) );
  NOR2_X1 U650 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U651 ( .A(G211GAT), .B(n586), .Z(G1354GAT) );
  NAND2_X1 U652 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U653 ( .A(n589), .B(KEYINPUT62), .ZN(n590) );
  XNOR2_X1 U654 ( .A(G218GAT), .B(n590), .ZN(G1355GAT) );
endmodule

