//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 0 0 1 0 0 0 1 1 0 1 0 1 1 1 0 0 0 1 0 0 1 0 1 0 1 1 1 1 1 0 1 1 1 0 1 0 1 0 0 0 1 0 0 1 1 1 0 0 1 1 1 1 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:59 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n449, new_n450, new_n452, new_n455,
    new_n456, new_n457, new_n458, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n574, new_n575, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n592, new_n593, new_n594, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n624, new_n627, new_n628, new_n630, new_n631, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n846, new_n847, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n965, new_n966,
    new_n967, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1209;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT65), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT66), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g022(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT68), .ZN(new_n449));
  AND2_X1   g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n449), .B(new_n450), .ZN(G223));
  NAND2_X1  g026(.A1(new_n450), .A2(G567), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT69), .Z(G234));
  NAND2_X1  g028(.A1(new_n450), .A2(G2106), .ZN(G217));
  NOR4_X1   g029(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT2), .Z(new_n456));
  NOR4_X1   g031(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n456), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  AOI22_X1  g035(.A1(new_n456), .A2(G2106), .B1(G567), .B2(new_n458), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT70), .ZN(new_n467));
  AND3_X1   g042(.A1(new_n464), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n467), .B1(new_n464), .B2(new_n466), .ZN(new_n469));
  OAI21_X1  g044(.A(G125), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n462), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  AND3_X1   g047(.A1(KEYINPUT71), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(KEYINPUT3), .B1(KEYINPUT71), .B2(G2104), .ZN(new_n474));
  OAI211_X1 g049(.A(G137), .B(new_n462), .C1(new_n473), .C2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n463), .A2(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G101), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n475), .A2(KEYINPUT72), .A3(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  AOI21_X1  g054(.A(KEYINPUT72), .B1(new_n475), .B2(new_n477), .ZN(new_n480));
  NOR3_X1   g055(.A1(new_n472), .A2(new_n479), .A3(new_n480), .ZN(G160));
  OAI21_X1  g056(.A(new_n462), .B1(new_n473), .B2(new_n474), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G136), .ZN(new_n484));
  OAI21_X1  g059(.A(G2105), .B1(new_n473), .B2(new_n474), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G124), .ZN(new_n487));
  NOR2_X1   g062(.A1(G100), .A2(G2105), .ZN(new_n488));
  XOR2_X1   g063(.A(new_n488), .B(KEYINPUT73), .Z(new_n489));
  OAI21_X1  g064(.A(G2104), .B1(new_n462), .B2(G112), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n484), .B(new_n487), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  XOR2_X1   g066(.A(new_n491), .B(KEYINPUT74), .Z(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G162));
  OAI21_X1  g068(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT75), .ZN(new_n496));
  INV_X1    g071(.A(G114), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n496), .B1(new_n497), .B2(G2105), .ZN(new_n498));
  NOR3_X1   g073(.A1(new_n462), .A2(KEYINPUT75), .A3(G114), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n495), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(G126), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n500), .B1(new_n501), .B2(new_n485), .ZN(new_n502));
  INV_X1    g077(.A(G138), .ZN(new_n503));
  NOR3_X1   g078(.A1(new_n503), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n504), .B1(new_n468), .B2(new_n469), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT76), .ZN(new_n506));
  OAI211_X1 g081(.A(G138), .B(new_n462), .C1(new_n473), .C2(new_n474), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n505), .A2(new_n506), .B1(KEYINPUT4), .B2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(new_n504), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n465), .A2(G2104), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n511));
  OAI21_X1  g086(.A(KEYINPUT70), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n464), .A2(new_n466), .A3(new_n467), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n509), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(KEYINPUT76), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n502), .B1(new_n508), .B2(new_n515), .ZN(G164));
  OR2_X1    g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(KEYINPUT6), .A2(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AND2_X1   g094(.A1(G50), .A2(G543), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n519), .A2(KEYINPUT77), .A3(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(new_n521), .ZN(new_n522));
  AOI21_X1  g097(.A(KEYINPUT77), .B1(new_n519), .B2(new_n520), .ZN(new_n523));
  INV_X1    g098(.A(G543), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n524), .A2(KEYINPUT5), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT5), .ZN(new_n526));
  OAI21_X1  g101(.A(KEYINPUT78), .B1(new_n526), .B2(G543), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT78), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n528), .A2(new_n524), .A3(KEYINPUT5), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n525), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(new_n519), .ZN(new_n531));
  XNOR2_X1  g106(.A(KEYINPUT79), .B(G88), .ZN(new_n532));
  OAI22_X1  g107(.A1(new_n522), .A2(new_n523), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n530), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n534));
  INV_X1    g109(.A(G651), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n533), .A2(new_n536), .ZN(G166));
  INV_X1    g112(.A(new_n531), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G89), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n517), .A2(KEYINPUT80), .A3(new_n518), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT80), .ZN(new_n541));
  AND2_X1   g116(.A1(KEYINPUT6), .A2(G651), .ZN(new_n542));
  NOR2_X1   g117(.A1(KEYINPUT6), .A2(G651), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  AND3_X1   g119(.A1(new_n540), .A2(new_n544), .A3(G543), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G51), .ZN(new_n546));
  NAND3_X1  g121(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT7), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n530), .A2(G63), .A3(G651), .ZN(new_n549));
  NAND4_X1  g124(.A1(new_n539), .A2(new_n546), .A3(new_n548), .A4(new_n549), .ZN(G286));
  INV_X1    g125(.A(G286), .ZN(G168));
  AOI22_X1  g126(.A1(new_n530), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n552), .A2(new_n535), .ZN(new_n553));
  INV_X1    g128(.A(G90), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n540), .A2(new_n544), .A3(G543), .ZN(new_n555));
  INV_X1    g130(.A(G52), .ZN(new_n556));
  OAI22_X1  g131(.A1(new_n531), .A2(new_n554), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n553), .A2(new_n557), .ZN(G171));
  NAND2_X1  g133(.A1(G68), .A2(G543), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n527), .A2(new_n529), .ZN(new_n560));
  INV_X1    g135(.A(new_n525), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(G56), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n559), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G651), .ZN(new_n565));
  NAND4_X1  g140(.A1(new_n540), .A2(new_n544), .A3(G43), .A4(G543), .ZN(new_n566));
  NAND4_X1  g141(.A1(new_n560), .A2(G81), .A3(new_n561), .A4(new_n519), .ZN(new_n567));
  AND3_X1   g142(.A1(new_n566), .A2(new_n567), .A3(KEYINPUT81), .ZN(new_n568));
  AOI21_X1  g143(.A(KEYINPUT81), .B1(new_n566), .B2(new_n567), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n565), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(G860), .ZN(G153));
  NAND4_X1  g147(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g148(.A1(G1), .A2(G3), .ZN(new_n574));
  XNOR2_X1  g149(.A(new_n574), .B(KEYINPUT8), .ZN(new_n575));
  NAND4_X1  g150(.A1(G319), .A2(G483), .A3(G661), .A4(new_n575), .ZN(G188));
  NAND4_X1  g151(.A1(new_n540), .A2(new_n544), .A3(G53), .A4(G543), .ZN(new_n577));
  AOI21_X1  g152(.A(KEYINPUT83), .B1(KEYINPUT82), .B2(KEYINPUT9), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n538), .A2(G91), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n578), .B1(KEYINPUT83), .B2(KEYINPUT9), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n545), .A2(G53), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n530), .A2(G65), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT85), .ZN(new_n583));
  NAND2_X1  g158(.A1(G78), .A2(G543), .ZN(new_n584));
  XOR2_X1   g159(.A(new_n584), .B(KEYINPUT84), .Z(new_n585));
  NAND3_X1  g160(.A1(new_n582), .A2(new_n583), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n586), .A2(G651), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n583), .B1(new_n582), .B2(new_n585), .ZN(new_n588));
  OAI211_X1 g163(.A(new_n579), .B(new_n581), .C1(new_n587), .C2(new_n588), .ZN(G299));
  INV_X1    g164(.A(G171), .ZN(G301));
  INV_X1    g165(.A(G166), .ZN(G303));
  NAND2_X1  g166(.A1(new_n545), .A2(G49), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n530), .A2(G87), .A3(new_n519), .ZN(new_n593));
  OAI21_X1  g168(.A(G651), .B1(new_n530), .B2(G74), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(G288));
  NAND2_X1  g170(.A1(new_n530), .A2(G61), .ZN(new_n596));
  NAND2_X1  g171(.A1(G73), .A2(G543), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n535), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n560), .A2(G86), .A3(new_n561), .ZN(new_n599));
  NAND2_X1  g174(.A1(G48), .A2(G543), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n599), .A2(new_n600), .B1(new_n517), .B2(new_n518), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(new_n602), .ZN(G305));
  AOI22_X1  g178(.A1(new_n538), .A2(G85), .B1(new_n545), .B2(G47), .ZN(new_n604));
  AND2_X1   g179(.A1(new_n530), .A2(G60), .ZN(new_n605));
  AND2_X1   g180(.A1(G72), .A2(G543), .ZN(new_n606));
  OAI211_X1 g181(.A(KEYINPUT86), .B(G651), .C1(new_n605), .C2(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT86), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n606), .B1(new_n530), .B2(G60), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n609), .B2(new_n535), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n604), .A2(new_n607), .A3(new_n610), .ZN(G290));
  NAND3_X1  g186(.A1(new_n530), .A2(G92), .A3(new_n519), .ZN(new_n612));
  INV_X1    g187(.A(KEYINPUT10), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n612), .B(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(G79), .A2(G543), .ZN(new_n615));
  INV_X1    g190(.A(G66), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n562), .B2(new_n616), .ZN(new_n617));
  AOI22_X1  g192(.A1(new_n617), .A2(G651), .B1(G54), .B2(new_n545), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n614), .A2(new_n618), .ZN(new_n619));
  INV_X1    g194(.A(G868), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n621), .B1(new_n620), .B2(G171), .ZN(G321));
  XOR2_X1   g197(.A(G321), .B(KEYINPUT87), .Z(G284));
  NAND2_X1  g198(.A1(G299), .A2(new_n620), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n624), .B1(new_n620), .B2(G168), .ZN(G297));
  OAI21_X1  g200(.A(new_n624), .B1(new_n620), .B2(G168), .ZN(G280));
  INV_X1    g201(.A(new_n619), .ZN(new_n627));
  XNOR2_X1  g202(.A(KEYINPUT88), .B(G559), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n627), .B1(G860), .B2(new_n628), .ZN(G148));
  NAND2_X1  g204(.A1(new_n627), .A2(new_n628), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n630), .A2(G868), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n631), .B1(G868), .B2(new_n571), .ZN(G323));
  XNOR2_X1  g207(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g208(.A1(new_n512), .A2(new_n513), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n634), .A2(new_n476), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT12), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT89), .B(KEYINPUT13), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(G2100), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n636), .B(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n483), .A2(G135), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n486), .A2(G123), .ZN(new_n641));
  NOR2_X1   g216(.A1(new_n462), .A2(G111), .ZN(new_n642));
  OAI21_X1  g217(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n643));
  OAI211_X1 g218(.A(new_n640), .B(new_n641), .C1(new_n642), .C2(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT90), .B(G2096), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n639), .A2(new_n646), .ZN(G156));
  XNOR2_X1  g222(.A(G2427), .B(G2438), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G2430), .ZN(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT15), .B(G2435), .ZN(new_n650));
  OR2_X1    g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n649), .A2(new_n650), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n651), .A2(KEYINPUT14), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2451), .B(G2454), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT16), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n653), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2443), .B(G2446), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1341), .B(G1348), .ZN(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n656), .A2(new_n657), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n658), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT91), .ZN(new_n663));
  INV_X1    g238(.A(G14), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n658), .A2(new_n661), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n664), .B1(new_n665), .B2(new_n659), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(G401));
  XOR2_X1   g243(.A(KEYINPUT92), .B(KEYINPUT18), .Z(new_n669));
  XOR2_X1   g244(.A(G2084), .B(G2090), .Z(new_n670));
  XNOR2_X1  g245(.A(G2067), .B(G2678), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  AND2_X1   g247(.A1(new_n672), .A2(KEYINPUT17), .ZN(new_n673));
  OR2_X1    g248(.A1(new_n670), .A2(new_n671), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n669), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(G2072), .B(G2078), .Z(new_n676));
  AOI21_X1  g251(.A(new_n676), .B1(new_n672), .B2(new_n669), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n675), .B(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(G2096), .B(G2100), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT93), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n678), .B(new_n680), .ZN(G227));
  XOR2_X1   g256(.A(G1991), .B(G1996), .Z(new_n682));
  XOR2_X1   g257(.A(G1971), .B(G1976), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT19), .ZN(new_n684));
  XOR2_X1   g259(.A(G1956), .B(G2474), .Z(new_n685));
  XOR2_X1   g260(.A(G1961), .B(G1966), .Z(new_n686));
  AND2_X1   g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT95), .ZN(new_n689));
  XOR2_X1   g264(.A(KEYINPUT94), .B(KEYINPUT20), .Z(new_n690));
  OR2_X1    g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n689), .A2(new_n690), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n685), .A2(new_n686), .ZN(new_n693));
  NOR3_X1   g268(.A1(new_n684), .A2(new_n687), .A3(new_n693), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n694), .B1(new_n684), .B2(new_n693), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n691), .A2(new_n692), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n696), .A2(new_n698), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n682), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(G1981), .B(G1986), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  NOR3_X1   g280(.A1(new_n700), .A2(new_n701), .A3(new_n682), .ZN(new_n706));
  OR3_X1    g281(.A1(new_n703), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n705), .B1(new_n703), .B2(new_n706), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(G229));
  XOR2_X1   g285(.A(KEYINPUT96), .B(G29), .Z(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n712), .A2(G35), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n713), .B1(G162), .B2(new_n712), .ZN(new_n714));
  XOR2_X1   g289(.A(new_n714), .B(KEYINPUT29), .Z(new_n715));
  INV_X1    g290(.A(G2090), .ZN(new_n716));
  AND2_X1   g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(G16), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(G19), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(new_n571), .B2(new_n718), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(G1341), .Z(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(new_n715), .B2(new_n716), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n711), .A2(G26), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(KEYINPUT28), .Z(new_n724));
  OR2_X1    g299(.A1(G104), .A2(G2105), .ZN(new_n725));
  OAI211_X1 g300(.A(new_n725), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT105), .ZN(new_n727));
  INV_X1    g302(.A(G140), .ZN(new_n728));
  OAI21_X1  g303(.A(KEYINPUT104), .B1(new_n482), .B2(new_n728), .ZN(new_n729));
  OR3_X1    g304(.A1(new_n482), .A2(KEYINPUT104), .A3(new_n728), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n486), .A2(G128), .ZN(new_n731));
  NAND4_X1  g306(.A1(new_n727), .A2(new_n729), .A3(new_n730), .A4(new_n731), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n724), .B1(new_n732), .B2(G29), .ZN(new_n733));
  INV_X1    g308(.A(G2067), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n733), .B(new_n734), .ZN(new_n735));
  XOR2_X1   g310(.A(KEYINPUT31), .B(G11), .Z(new_n736));
  INV_X1    g311(.A(G28), .ZN(new_n737));
  OR2_X1    g312(.A1(new_n737), .A2(KEYINPUT30), .ZN(new_n738));
  AOI21_X1  g313(.A(G29), .B1(new_n737), .B2(KEYINPUT30), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n736), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n718), .A2(G5), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(G171), .B2(new_n718), .ZN(new_n742));
  OAI221_X1 g317(.A(new_n740), .B1(new_n644), .B2(new_n711), .C1(new_n742), .C2(G1961), .ZN(new_n743));
  OR2_X1    g318(.A1(new_n735), .A2(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(KEYINPUT24), .ZN(new_n745));
  OR2_X1    g320(.A1(new_n745), .A2(G34), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n745), .A2(G34), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n711), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(G160), .ZN(new_n749));
  INV_X1    g324(.A(G29), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n748), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(G2084), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  NOR4_X1   g328(.A1(new_n717), .A2(new_n722), .A3(new_n744), .A4(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n750), .A2(G32), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n483), .A2(G141), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n486), .A2(G129), .ZN(new_n757));
  NAND3_X1  g332(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT26), .ZN(new_n759));
  OR2_X1    g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n758), .A2(new_n759), .ZN(new_n761));
  AOI22_X1  g336(.A1(new_n760), .A2(new_n761), .B1(G105), .B2(new_n476), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n756), .A2(new_n757), .A3(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(new_n763), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n755), .B1(new_n764), .B2(new_n750), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT27), .ZN(new_n766));
  INV_X1    g341(.A(G1996), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  XNOR2_X1  g343(.A(KEYINPUT108), .B(G1956), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n718), .A2(G20), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT23), .Z(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(G299), .B2(G16), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n768), .B1(new_n769), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n718), .A2(G4), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(new_n627), .B2(new_n718), .ZN(new_n775));
  XOR2_X1   g350(.A(KEYINPUT103), .B(G1348), .Z(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n742), .A2(G1961), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n750), .A2(G33), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n780));
  INV_X1    g355(.A(KEYINPUT25), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(G139), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n782), .B1(new_n783), .B2(new_n482), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n634), .A2(G127), .ZN(new_n785));
  INV_X1    g360(.A(G115), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n785), .B1(new_n786), .B2(new_n463), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n784), .B1(new_n787), .B2(G2105), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n779), .B1(new_n788), .B2(new_n750), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(G2072), .Z(new_n790));
  NAND4_X1  g365(.A1(new_n773), .A2(new_n777), .A3(new_n778), .A4(new_n790), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n712), .A2(G27), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(G164), .B2(new_n712), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(G2078), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n718), .A2(G21), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(G168), .B2(new_n718), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(KEYINPUT106), .Z(new_n797));
  OAI22_X1  g372(.A1(new_n797), .A2(G1966), .B1(new_n769), .B2(new_n772), .ZN(new_n798));
  NOR3_X1   g373(.A1(new_n791), .A2(new_n794), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n797), .A2(G1966), .ZN(new_n800));
  XOR2_X1   g375(.A(new_n800), .B(KEYINPUT107), .Z(new_n801));
  NAND3_X1  g376(.A1(new_n754), .A2(new_n799), .A3(new_n801), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n712), .A2(G25), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n483), .A2(G131), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n486), .A2(G119), .ZN(new_n805));
  OR2_X1    g380(.A1(G95), .A2(G2105), .ZN(new_n806));
  OAI211_X1 g381(.A(new_n806), .B(G2104), .C1(G107), .C2(new_n462), .ZN(new_n807));
  AND3_X1   g382(.A1(new_n804), .A2(new_n805), .A3(new_n807), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n803), .B1(new_n808), .B2(new_n712), .ZN(new_n809));
  XOR2_X1   g384(.A(new_n809), .B(KEYINPUT97), .Z(new_n810));
  XOR2_X1   g385(.A(KEYINPUT35), .B(G1991), .Z(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT98), .ZN(new_n813));
  AND2_X1   g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n812), .A2(new_n813), .ZN(new_n815));
  MUX2_X1   g390(.A(G24), .B(G290), .S(G16), .Z(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(G1986), .ZN(new_n817));
  NOR3_X1   g392(.A1(new_n814), .A2(new_n815), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n718), .A2(G6), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n819), .B1(new_n602), .B2(new_n718), .ZN(new_n820));
  XOR2_X1   g395(.A(new_n820), .B(KEYINPUT100), .Z(new_n821));
  XNOR2_X1  g396(.A(KEYINPUT32), .B(G1981), .ZN(new_n822));
  INV_X1    g397(.A(new_n822), .ZN(new_n823));
  OR2_X1    g398(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n821), .A2(new_n823), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n718), .A2(G22), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(G166), .B2(new_n718), .ZN(new_n827));
  INV_X1    g402(.A(G1971), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n718), .A2(G23), .ZN(new_n830));
  INV_X1    g405(.A(G288), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n830), .B1(new_n831), .B2(new_n718), .ZN(new_n832));
  XNOR2_X1  g407(.A(KEYINPUT33), .B(G1976), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT101), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n832), .B(new_n834), .ZN(new_n835));
  NAND4_X1  g410(.A1(new_n824), .A2(new_n825), .A3(new_n829), .A4(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(KEYINPUT99), .B(KEYINPUT34), .ZN(new_n837));
  OR2_X1    g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n836), .A2(new_n837), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n818), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  XOR2_X1   g415(.A(KEYINPUT102), .B(KEYINPUT36), .Z(new_n841));
  NOR2_X1   g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n840), .A2(new_n841), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n802), .B1(new_n843), .B2(new_n844), .ZN(G311));
  AND2_X1   g420(.A1(new_n799), .A2(new_n801), .ZN(new_n846));
  INV_X1    g421(.A(new_n844), .ZN(new_n847));
  OAI211_X1 g422(.A(new_n754), .B(new_n846), .C1(new_n847), .C2(new_n842), .ZN(G150));
  NAND2_X1  g423(.A1(new_n627), .A2(G559), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(KEYINPUT38), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n530), .A2(G67), .ZN(new_n851));
  NAND2_X1  g426(.A1(G80), .A2(G543), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n535), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND4_X1  g428(.A1(new_n560), .A2(G93), .A3(new_n561), .A4(new_n519), .ZN(new_n854));
  INV_X1    g429(.A(G55), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n854), .B1(new_n555), .B2(new_n855), .ZN(new_n856));
  OR2_X1    g431(.A1(new_n853), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n570), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n566), .A2(new_n567), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT81), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n566), .A2(new_n567), .A3(KEYINPUT81), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n853), .A2(new_n856), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n863), .A2(new_n565), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n858), .A2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n850), .B(new_n867), .ZN(new_n868));
  OR2_X1    g443(.A1(new_n868), .A2(KEYINPUT39), .ZN(new_n869));
  INV_X1    g444(.A(G860), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n868), .A2(KEYINPUT39), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n869), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n864), .A2(new_n870), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(KEYINPUT37), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n872), .A2(new_n874), .ZN(G145));
  OR2_X1    g450(.A1(G106), .A2(G2105), .ZN(new_n876));
  OAI211_X1 g451(.A(new_n876), .B(G2104), .C1(G118), .C2(new_n462), .ZN(new_n877));
  INV_X1    g452(.A(G142), .ZN(new_n878));
  INV_X1    g453(.A(G130), .ZN(new_n879));
  OAI221_X1 g454(.A(new_n877), .B1(new_n482), .B2(new_n878), .C1(new_n879), .C2(new_n485), .ZN(new_n880));
  OR2_X1    g455(.A1(new_n880), .A2(KEYINPUT109), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(KEYINPUT109), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  XOR2_X1   g458(.A(new_n635), .B(KEYINPUT12), .Z(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n636), .A2(new_n881), .A3(new_n882), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n808), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n885), .A2(new_n886), .A3(new_n808), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT110), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n889), .A2(KEYINPUT110), .A3(new_n890), .ZN(new_n894));
  INV_X1    g469(.A(new_n732), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n895), .A2(G164), .ZN(new_n896));
  INV_X1    g471(.A(new_n502), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n507), .A2(KEYINPUT4), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n898), .B1(new_n514), .B2(KEYINPUT76), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n505), .A2(new_n506), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n897), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(new_n732), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n896), .A2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n788), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n896), .A2(new_n788), .A3(new_n902), .ZN(new_n906));
  AND3_X1   g481(.A1(new_n905), .A2(new_n763), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n763), .B1(new_n905), .B2(new_n906), .ZN(new_n908));
  OAI211_X1 g483(.A(new_n893), .B(new_n894), .C1(new_n907), .C2(new_n908), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n907), .A2(new_n908), .ZN(new_n910));
  AOI21_X1  g485(.A(KEYINPUT110), .B1(new_n889), .B2(new_n890), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  XOR2_X1   g487(.A(G160), .B(new_n644), .Z(new_n913));
  XNOR2_X1  g488(.A(new_n913), .B(new_n492), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n909), .A2(new_n912), .A3(new_n914), .ZN(new_n915));
  XNOR2_X1  g490(.A(KEYINPUT111), .B(G37), .ZN(new_n916));
  AND2_X1   g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT112), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n909), .A2(new_n912), .ZN(new_n919));
  INV_X1    g494(.A(new_n914), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n918), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  AOI211_X1 g496(.A(KEYINPUT112), .B(new_n914), .C1(new_n909), .C2(new_n912), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n917), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  XNOR2_X1  g498(.A(KEYINPUT113), .B(KEYINPUT40), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n923), .B(new_n924), .ZN(G395));
  NAND4_X1  g500(.A1(new_n831), .A2(new_n607), .A3(new_n610), .A4(new_n604), .ZN(new_n926));
  NAND2_X1  g501(.A1(G290), .A2(G288), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT114), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n926), .A2(new_n927), .A3(KEYINPUT114), .ZN(new_n931));
  XNOR2_X1  g506(.A(G166), .B(new_n602), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n930), .A2(new_n931), .A3(new_n933), .ZN(new_n934));
  NAND4_X1  g509(.A1(new_n932), .A2(KEYINPUT114), .A3(new_n927), .A4(new_n926), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  XOR2_X1   g511(.A(KEYINPUT115), .B(KEYINPUT42), .Z(new_n937));
  AND2_X1   g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n936), .A2(new_n937), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  XNOR2_X1  g515(.A(new_n866), .B(new_n630), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n538), .A2(G91), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n577), .A2(new_n578), .ZN(new_n943));
  AND3_X1   g518(.A1(new_n942), .A2(new_n581), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n582), .A2(new_n585), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(KEYINPUT85), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n946), .A2(G651), .A3(new_n586), .ZN(new_n947));
  NAND4_X1  g522(.A1(new_n944), .A2(new_n947), .A3(new_n614), .A4(new_n618), .ZN(new_n948));
  NAND2_X1  g523(.A1(G299), .A2(new_n619), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(KEYINPUT41), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT41), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n948), .A2(new_n949), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  OR2_X1    g529(.A1(new_n941), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n941), .A2(new_n950), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n940), .A2(new_n957), .ZN(new_n958));
  OAI211_X1 g533(.A(new_n956), .B(new_n955), .C1(new_n938), .C2(new_n939), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n620), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(new_n960), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n864), .A2(G868), .ZN(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n961), .A2(new_n963), .ZN(G295));
  INV_X1    g539(.A(KEYINPUT116), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n961), .A2(new_n965), .A3(new_n963), .ZN(new_n966));
  OAI21_X1  g541(.A(KEYINPUT116), .B1(new_n960), .B2(new_n962), .ZN(new_n967));
  AND2_X1   g542(.A1(new_n966), .A2(new_n967), .ZN(G331));
  INV_X1    g543(.A(new_n916), .ZN(new_n969));
  INV_X1    g544(.A(new_n950), .ZN(new_n970));
  AND3_X1   g545(.A1(new_n858), .A2(new_n865), .A3(G301), .ZN(new_n971));
  AOI21_X1  g546(.A(G301), .B1(new_n858), .B2(new_n865), .ZN(new_n972));
  NOR3_X1   g547(.A1(new_n971), .A2(new_n972), .A3(G286), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n570), .A2(new_n857), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n864), .B1(new_n863), .B2(new_n565), .ZN(new_n975));
  OAI21_X1  g550(.A(G171), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n858), .A2(new_n865), .A3(G301), .ZN(new_n977));
  AOI21_X1  g552(.A(G168), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n970), .B1(new_n973), .B2(new_n978), .ZN(new_n979));
  OAI21_X1  g554(.A(G286), .B1(new_n971), .B2(new_n972), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n976), .A2(G168), .A3(new_n977), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n954), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n979), .A2(new_n982), .ZN(new_n983));
  OAI21_X1  g558(.A(KEYINPUT118), .B1(new_n983), .B2(new_n936), .ZN(new_n984));
  AND2_X1   g559(.A1(new_n934), .A2(new_n935), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT118), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n985), .A2(new_n979), .A3(new_n982), .A4(new_n986), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n969), .B1(new_n984), .B2(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n950), .B1(new_n980), .B2(new_n981), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n973), .A2(new_n978), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT119), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n953), .A2(new_n991), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n948), .A2(new_n949), .A3(KEYINPUT119), .A4(new_n952), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n992), .A2(new_n951), .A3(new_n993), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n989), .B1(new_n990), .B2(new_n994), .ZN(new_n995));
  OAI21_X1  g570(.A(KEYINPUT120), .B1(new_n995), .B2(new_n985), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT120), .ZN(new_n997));
  AND3_X1   g572(.A1(new_n994), .A2(new_n981), .A3(new_n980), .ZN(new_n998));
  OAI211_X1 g573(.A(new_n997), .B(new_n936), .C1(new_n998), .C2(new_n989), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n996), .A2(new_n999), .ZN(new_n1000));
  AND3_X1   g575(.A1(new_n988), .A2(new_n1000), .A3(KEYINPUT43), .ZN(new_n1001));
  AOI21_X1  g576(.A(G37), .B1(new_n984), .B2(new_n987), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT117), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n985), .B1(new_n983), .B2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n1004), .B1(new_n1003), .B2(new_n983), .ZN(new_n1005));
  AOI21_X1  g580(.A(KEYINPUT43), .B1(new_n1002), .B2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g581(.A(KEYINPUT44), .B1(new_n1001), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT44), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT43), .ZN(new_n1009));
  AND3_X1   g584(.A1(new_n988), .A2(new_n1000), .A3(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1009), .B1(new_n1002), .B2(new_n1005), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1008), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1007), .A2(new_n1012), .ZN(G397));
  INV_X1    g588(.A(KEYINPUT57), .ZN(new_n1014));
  XNOR2_X1  g589(.A(G299), .B(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(G125), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1016), .B1(new_n512), .B2(new_n513), .ZN(new_n1017));
  INV_X1    g592(.A(new_n471), .ZN(new_n1018));
  OAI21_X1  g593(.A(G2105), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(new_n480), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n1019), .A2(new_n1020), .A3(G40), .A4(new_n478), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT45), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1022), .A2(G1384), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1021), .B1(new_n901), .B2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1022), .B1(G164), .B2(G1384), .ZN(new_n1025));
  XNOR2_X1  g600(.A(KEYINPUT56), .B(G2072), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1024), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  NOR2_X1   g602(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n901), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1021), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT50), .ZN(new_n1032));
  INV_X1    g607(.A(G1384), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1032), .B1(new_n901), .B2(new_n1033), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1031), .A2(new_n1034), .ZN(new_n1035));
  OAI211_X1 g610(.A(new_n1015), .B(new_n1027), .C1(new_n1035), .C2(G1956), .ZN(new_n1036));
  NOR4_X1   g611(.A1(G164), .A2(new_n1021), .A3(G1384), .A4(G2067), .ZN(new_n1037));
  INV_X1    g612(.A(new_n776), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1021), .B1(new_n901), .B2(new_n1028), .ZN(new_n1039));
  OAI21_X1  g614(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1038), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  OAI211_X1 g616(.A(new_n1036), .B(new_n627), .C1(new_n1037), .C2(new_n1041), .ZN(new_n1042));
  XNOR2_X1  g617(.A(G299), .B(KEYINPUT57), .ZN(new_n1043));
  AND3_X1   g618(.A1(new_n1024), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1044));
  AOI21_X1  g619(.A(G1956), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1043), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  AND2_X1   g621(.A1(new_n1042), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT60), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1048), .B1(new_n1041), .B2(new_n1037), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1037), .B1(new_n776), .B2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n619), .B1(new_n1051), .B2(KEYINPUT60), .ZN(new_n1052));
  NOR4_X1   g627(.A1(new_n1041), .A2(new_n1037), .A3(new_n1048), .A4(new_n627), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1049), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  XNOR2_X1  g629(.A(KEYINPUT125), .B(KEYINPUT59), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1024), .A2(new_n1025), .A3(new_n767), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n505), .A2(new_n506), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n515), .A2(new_n1057), .A3(new_n898), .ZN(new_n1058));
  AOI21_X1  g633(.A(G1384), .B1(new_n1058), .B2(new_n897), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(new_n1030), .ZN(new_n1060));
  XOR2_X1   g635(.A(KEYINPUT58), .B(G1341), .Z(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  AOI211_X1 g637(.A(new_n570), .B(new_n1055), .C1(new_n1056), .C2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1056), .A2(new_n1062), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(new_n571), .ZN(new_n1065));
  NOR2_X1   g640(.A1(KEYINPUT125), .A2(KEYINPUT59), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1063), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1046), .A2(new_n1036), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT61), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1054), .A2(new_n1067), .A3(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1046), .A2(new_n1036), .A3(KEYINPUT61), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(KEYINPUT126), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT126), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1046), .A2(new_n1036), .A3(new_n1074), .A4(KEYINPUT61), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1047), .B1(new_n1071), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1023), .ZN(new_n1078));
  OAI211_X1 g653(.A(G40), .B(G160), .C1(G164), .C2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(KEYINPUT45), .B1(new_n901), .B2(new_n1033), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n828), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1039), .A2(new_n1040), .A3(new_n716), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(G8), .ZN(new_n1084));
  XNOR2_X1  g659(.A(KEYINPUT122), .B(KEYINPUT55), .ZN(new_n1085));
  OAI211_X1 g660(.A(G8), .B(new_n1085), .C1(new_n533), .C2(new_n536), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(G303), .A2(G8), .ZN(new_n1088));
  NAND2_X1  g663(.A1(KEYINPUT122), .A2(KEYINPUT55), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1087), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1084), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(G8), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1092), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1090), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT49), .ZN(new_n1096));
  INV_X1    g671(.A(G1981), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n596), .A2(new_n597), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(G651), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n599), .A2(new_n600), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(new_n519), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1097), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1102));
  NOR3_X1   g677(.A1(new_n598), .A2(new_n601), .A3(G1981), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1096), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n602), .A2(new_n1097), .ZN(new_n1105));
  OAI21_X1  g680(.A(G1981), .B1(new_n598), .B2(new_n601), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1105), .A2(KEYINPUT49), .A3(new_n1106), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1060), .A2(new_n1104), .A3(new_n1107), .A4(G8), .ZN(new_n1108));
  INV_X1    g683(.A(G1976), .ZN(new_n1109));
  NOR2_X1   g684(.A1(G288), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(KEYINPUT52), .B1(G288), .B2(new_n1109), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1060), .A2(G8), .A3(new_n1111), .A4(new_n1112), .ZN(new_n1113));
  AOI211_X1 g688(.A(new_n1092), .B(new_n1110), .C1(new_n1059), .C2(new_n1030), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT52), .ZN(new_n1115));
  OAI211_X1 g690(.A(new_n1108), .B(new_n1113), .C1(new_n1114), .C2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1116), .ZN(new_n1117));
  AND3_X1   g692(.A1(new_n1091), .A2(new_n1095), .A3(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(G1966), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1119), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1039), .A2(new_n1040), .A3(new_n752), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1120), .A2(G168), .A3(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(G8), .ZN(new_n1123));
  AOI21_X1  g698(.A(G168), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1124));
  OAI21_X1  g699(.A(KEYINPUT51), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT51), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1122), .A2(new_n1126), .A3(G8), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1125), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(G2078), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1024), .A2(new_n1025), .A3(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT53), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(G1961), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1050), .A2(new_n1133), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1024), .A2(new_n1025), .A3(KEYINPUT53), .A4(new_n1129), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1132), .A2(new_n1134), .A3(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1136), .A2(G171), .ZN(new_n1137));
  AND2_X1   g712(.A1(new_n1130), .A2(KEYINPUT127), .ZN(new_n1138));
  OAI21_X1  g713(.A(KEYINPUT53), .B1(new_n1130), .B2(KEYINPUT127), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1134), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1132), .A2(G301), .ZN(new_n1141));
  OAI211_X1 g716(.A(new_n1137), .B(KEYINPUT54), .C1(new_n1140), .C2(new_n1141), .ZN(new_n1142));
  AND3_X1   g717(.A1(new_n1118), .A2(new_n1128), .A3(new_n1142), .ZN(new_n1143));
  AND4_X1   g718(.A1(G301), .A2(new_n1132), .A3(new_n1134), .A4(new_n1135), .ZN(new_n1144));
  OAI211_X1 g719(.A(new_n1132), .B(new_n1134), .C1(new_n1138), .C2(new_n1139), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1144), .B1(new_n1145), .B2(G171), .ZN(new_n1146));
  OR2_X1    g721(.A1(new_n1146), .A2(KEYINPUT54), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1077), .A2(new_n1143), .A3(new_n1147), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1092), .B1(new_n1059), .B2(new_n1030), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1149), .ZN(new_n1150));
  NOR2_X1   g725(.A1(G288), .A2(G1976), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1103), .B1(new_n1108), .B2(new_n1151), .ZN(new_n1152));
  OAI22_X1  g727(.A1(new_n1095), .A2(new_n1116), .B1(new_n1150), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT62), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1154), .B1(new_n1125), .B2(new_n1127), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1116), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1156), .A2(new_n1091), .A3(new_n1145), .A4(G171), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1125), .A2(new_n1154), .A3(new_n1127), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1153), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  AOI211_X1 g735(.A(new_n1092), .B(G286), .C1(new_n1120), .C2(new_n1121), .ZN(new_n1161));
  NAND4_X1  g736(.A1(new_n1091), .A2(new_n1095), .A3(new_n1117), .A4(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT63), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT123), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1162), .A2(KEYINPUT123), .A3(new_n1163), .ZN(new_n1167));
  AND2_X1   g742(.A1(new_n1161), .A2(KEYINPUT63), .ZN(new_n1168));
  AND2_X1   g743(.A1(new_n1093), .A2(KEYINPUT124), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1090), .B1(new_n1093), .B2(KEYINPUT124), .ZN(new_n1170));
  OAI211_X1 g745(.A(new_n1168), .B(new_n1156), .C1(new_n1169), .C2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1166), .A2(new_n1167), .A3(new_n1171), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1148), .A2(new_n1160), .A3(new_n1172), .ZN(new_n1173));
  NOR2_X1   g748(.A1(new_n1025), .A2(new_n1021), .ZN(new_n1174));
  XNOR2_X1  g749(.A(new_n732), .B(G2067), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  XNOR2_X1  g751(.A(new_n1176), .B(KEYINPUT121), .ZN(new_n1177));
  XNOR2_X1  g752(.A(new_n763), .B(G1996), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1177), .B1(new_n1174), .B2(new_n1178), .ZN(new_n1179));
  NOR2_X1   g754(.A1(new_n808), .A2(new_n811), .ZN(new_n1180));
  AND2_X1   g755(.A1(new_n808), .A2(new_n811), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1174), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1179), .A2(new_n1182), .ZN(new_n1183));
  XNOR2_X1  g758(.A(G290), .B(G1986), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1183), .B1(new_n1174), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1173), .A2(new_n1185), .ZN(new_n1186));
  INV_X1    g761(.A(new_n1174), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1179), .A2(new_n1181), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n895), .A2(new_n734), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n1187), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  NOR3_X1   g765(.A1(new_n1187), .A2(G1986), .A3(G290), .ZN(new_n1191));
  XNOR2_X1  g766(.A(new_n1191), .B(KEYINPUT48), .ZN(new_n1192));
  NOR2_X1   g767(.A1(new_n1183), .A2(new_n1192), .ZN(new_n1193));
  OR3_X1    g768(.A1(new_n1187), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1194));
  OAI21_X1  g769(.A(KEYINPUT46), .B1(new_n1187), .B2(G1996), .ZN(new_n1195));
  OR2_X1    g770(.A1(new_n1175), .A2(new_n763), .ZN(new_n1196));
  AOI22_X1  g771(.A1(new_n1194), .A2(new_n1195), .B1(new_n1196), .B2(new_n1174), .ZN(new_n1197));
  XNOR2_X1  g772(.A(new_n1197), .B(KEYINPUT47), .ZN(new_n1198));
  NOR3_X1   g773(.A1(new_n1190), .A2(new_n1193), .A3(new_n1198), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1186), .A2(new_n1199), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g775(.A(G319), .ZN(new_n1202));
  AOI211_X1 g776(.A(new_n1202), .B(G227), .C1(new_n663), .C2(new_n666), .ZN(new_n1203));
  NAND3_X1  g777(.A1(new_n923), .A2(new_n709), .A3(new_n1203), .ZN(new_n1204));
  NAND2_X1  g778(.A1(new_n1002), .A2(new_n1005), .ZN(new_n1205));
  NAND2_X1  g779(.A1(new_n1205), .A2(KEYINPUT43), .ZN(new_n1206));
  NAND3_X1  g780(.A1(new_n988), .A2(new_n1000), .A3(new_n1009), .ZN(new_n1207));
  AOI21_X1  g781(.A(new_n1204), .B1(new_n1206), .B2(new_n1207), .ZN(G308));
  NAND2_X1  g782(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1209));
  NAND4_X1  g783(.A1(new_n1209), .A2(new_n709), .A3(new_n923), .A4(new_n1203), .ZN(G225));
endmodule


