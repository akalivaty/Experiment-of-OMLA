

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X2 U554 ( .A1(n535), .A2(G2104), .ZN(n869) );
  OR2_X1 U555 ( .A1(G299), .A2(n714), .ZN(n711) );
  NOR2_X1 U556 ( .A1(G651), .A2(G543), .ZN(n651) );
  AND2_X1 U557 ( .A1(n725), .A2(n521), .ZN(n520) );
  XNOR2_X1 U558 ( .A(KEYINPUT91), .B(n724), .ZN(n521) );
  NOR2_X2 U559 ( .A1(n589), .A2(n588), .ZN(n932) );
  NOR2_X2 U560 ( .A1(n576), .A2(n575), .ZN(G160) );
  XOR2_X1 U561 ( .A(G543), .B(KEYINPUT0), .Z(n522) );
  AND2_X1 U562 ( .A1(n538), .A2(n537), .ZN(n523) );
  INV_X1 U563 ( .A(KEYINPUT64), .ZN(n689) );
  INV_X1 U564 ( .A(KEYINPUT94), .ZN(n697) );
  NOR2_X1 U565 ( .A1(G164), .A2(G1384), .ZN(n765) );
  NOR2_X1 U566 ( .A1(G651), .A2(n632), .ZN(n655) );
  NOR2_X1 U567 ( .A1(n527), .A2(n632), .ZN(n650) );
  XNOR2_X1 U568 ( .A(n534), .B(KEYINPUT83), .ZN(n539) );
  AND2_X1 U569 ( .A1(n539), .A2(n523), .ZN(G164) );
  INV_X1 U570 ( .A(G651), .ZN(n527) );
  NOR2_X1 U571 ( .A1(G543), .A2(n527), .ZN(n524) );
  XOR2_X1 U572 ( .A(KEYINPUT1), .B(n524), .Z(n654) );
  NAND2_X1 U573 ( .A1(G65), .A2(n654), .ZN(n526) );
  XNOR2_X1 U574 ( .A(KEYINPUT66), .B(n522), .ZN(n632) );
  NAND2_X1 U575 ( .A1(G53), .A2(n655), .ZN(n525) );
  NAND2_X1 U576 ( .A1(n526), .A2(n525), .ZN(n531) );
  NAND2_X1 U577 ( .A1(G78), .A2(n650), .ZN(n529) );
  NAND2_X1 U578 ( .A1(G91), .A2(n651), .ZN(n528) );
  NAND2_X1 U579 ( .A1(n529), .A2(n528), .ZN(n530) );
  OR2_X1 U580 ( .A1(n531), .A2(n530), .ZN(G299) );
  AND2_X1 U581 ( .A1(G2105), .A2(G2104), .ZN(n873) );
  NAND2_X1 U582 ( .A1(G114), .A2(n873), .ZN(n533) );
  INV_X1 U583 ( .A(G2105), .ZN(n535) );
  NOR2_X2 U584 ( .A1(G2104), .A2(n535), .ZN(n874) );
  NAND2_X1 U585 ( .A1(G126), .A2(n874), .ZN(n532) );
  NAND2_X1 U586 ( .A1(n533), .A2(n532), .ZN(n534) );
  NAND2_X1 U587 ( .A1(G102), .A2(n869), .ZN(n538) );
  OR2_X1 U588 ( .A1(G2105), .A2(G2104), .ZN(n536) );
  XNOR2_X2 U589 ( .A(n536), .B(KEYINPUT17), .ZN(n870) );
  NAND2_X1 U590 ( .A1(n870), .A2(G138), .ZN(n537) );
  XOR2_X1 U591 ( .A(G2446), .B(G2451), .Z(n541) );
  XNOR2_X1 U592 ( .A(G2454), .B(KEYINPUT107), .ZN(n540) );
  XNOR2_X1 U593 ( .A(n541), .B(n540), .ZN(n548) );
  XOR2_X1 U594 ( .A(G2438), .B(G2430), .Z(n543) );
  XNOR2_X1 U595 ( .A(G2435), .B(G2443), .ZN(n542) );
  XNOR2_X1 U596 ( .A(n543), .B(n542), .ZN(n544) );
  XOR2_X1 U597 ( .A(n544), .B(G2427), .Z(n546) );
  XNOR2_X1 U598 ( .A(G1348), .B(G1341), .ZN(n545) );
  XNOR2_X1 U599 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U600 ( .A(n548), .B(n547), .ZN(n549) );
  AND2_X1 U601 ( .A1(n549), .A2(G14), .ZN(G401) );
  AND2_X1 U602 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U603 ( .A(G132), .ZN(G219) );
  INV_X1 U604 ( .A(G57), .ZN(G237) );
  NAND2_X1 U605 ( .A1(G64), .A2(n654), .ZN(n551) );
  NAND2_X1 U606 ( .A1(G52), .A2(n655), .ZN(n550) );
  NAND2_X1 U607 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U608 ( .A(KEYINPUT68), .B(n552), .ZN(n557) );
  NAND2_X1 U609 ( .A1(G77), .A2(n650), .ZN(n554) );
  NAND2_X1 U610 ( .A1(G90), .A2(n651), .ZN(n553) );
  NAND2_X1 U611 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U612 ( .A(KEYINPUT9), .B(n555), .Z(n556) );
  NOR2_X1 U613 ( .A1(n557), .A2(n556), .ZN(G171) );
  NAND2_X1 U614 ( .A1(G63), .A2(n654), .ZN(n559) );
  NAND2_X1 U615 ( .A1(G51), .A2(n655), .ZN(n558) );
  NAND2_X1 U616 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U617 ( .A(KEYINPUT6), .B(n560), .ZN(n566) );
  NAND2_X1 U618 ( .A1(n651), .A2(G89), .ZN(n561) );
  XNOR2_X1 U619 ( .A(n561), .B(KEYINPUT4), .ZN(n563) );
  NAND2_X1 U620 ( .A1(G76), .A2(n650), .ZN(n562) );
  NAND2_X1 U621 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U622 ( .A(n564), .B(KEYINPUT5), .Z(n565) );
  NOR2_X1 U623 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U624 ( .A(KEYINPUT73), .B(n567), .Z(n568) );
  XOR2_X1 U625 ( .A(KEYINPUT7), .B(n568), .Z(G168) );
  XOR2_X1 U626 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U627 ( .A1(G101), .A2(n869), .ZN(n569) );
  XOR2_X1 U628 ( .A(KEYINPUT23), .B(n569), .Z(n572) );
  NAND2_X1 U629 ( .A1(G113), .A2(n873), .ZN(n570) );
  XOR2_X1 U630 ( .A(KEYINPUT65), .B(n570), .Z(n571) );
  NAND2_X1 U631 ( .A1(n572), .A2(n571), .ZN(n576) );
  NAND2_X1 U632 ( .A1(G137), .A2(n870), .ZN(n574) );
  NAND2_X1 U633 ( .A1(G125), .A2(n874), .ZN(n573) );
  NAND2_X1 U634 ( .A1(n574), .A2(n573), .ZN(n575) );
  NAND2_X1 U635 ( .A1(G7), .A2(G661), .ZN(n577) );
  XNOR2_X1 U636 ( .A(n577), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U637 ( .A(G223), .ZN(n843) );
  NAND2_X1 U638 ( .A1(n843), .A2(G567), .ZN(n578) );
  XOR2_X1 U639 ( .A(KEYINPUT11), .B(n578), .Z(G234) );
  NAND2_X1 U640 ( .A1(G56), .A2(n654), .ZN(n579) );
  XNOR2_X1 U641 ( .A(n579), .B(KEYINPUT70), .ZN(n580) );
  XNOR2_X1 U642 ( .A(n580), .B(KEYINPUT14), .ZN(n582) );
  NAND2_X1 U643 ( .A1(G43), .A2(n655), .ZN(n581) );
  NAND2_X1 U644 ( .A1(n582), .A2(n581), .ZN(n589) );
  NAND2_X1 U645 ( .A1(G68), .A2(n650), .ZN(n585) );
  NAND2_X1 U646 ( .A1(n651), .A2(G81), .ZN(n583) );
  XNOR2_X1 U647 ( .A(n583), .B(KEYINPUT12), .ZN(n584) );
  NAND2_X1 U648 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U649 ( .A(n586), .B(KEYINPUT13), .ZN(n587) );
  XNOR2_X1 U650 ( .A(KEYINPUT71), .B(n587), .ZN(n588) );
  NAND2_X1 U651 ( .A1(G860), .A2(n932), .ZN(n590) );
  XNOR2_X1 U652 ( .A(n590), .B(KEYINPUT72), .ZN(G153) );
  INV_X1 U653 ( .A(G171), .ZN(G301) );
  NAND2_X1 U654 ( .A1(G868), .A2(G301), .ZN(n599) );
  NAND2_X1 U655 ( .A1(G79), .A2(n650), .ZN(n592) );
  NAND2_X1 U656 ( .A1(G92), .A2(n651), .ZN(n591) );
  NAND2_X1 U657 ( .A1(n592), .A2(n591), .ZN(n596) );
  NAND2_X1 U658 ( .A1(G66), .A2(n654), .ZN(n594) );
  NAND2_X1 U659 ( .A1(G54), .A2(n655), .ZN(n593) );
  NAND2_X1 U660 ( .A1(n594), .A2(n593), .ZN(n595) );
  NOR2_X1 U661 ( .A1(n596), .A2(n595), .ZN(n597) );
  XNOR2_X1 U662 ( .A(n597), .B(KEYINPUT15), .ZN(n941) );
  INV_X1 U663 ( .A(G868), .ZN(n669) );
  NAND2_X1 U664 ( .A1(n941), .A2(n669), .ZN(n598) );
  NAND2_X1 U665 ( .A1(n599), .A2(n598), .ZN(G284) );
  NOR2_X1 U666 ( .A1(G868), .A2(G299), .ZN(n601) );
  NOR2_X1 U667 ( .A1(G286), .A2(n669), .ZN(n600) );
  NOR2_X1 U668 ( .A1(n601), .A2(n600), .ZN(G297) );
  INV_X1 U669 ( .A(G860), .ZN(n602) );
  NAND2_X1 U670 ( .A1(n602), .A2(G559), .ZN(n603) );
  INV_X1 U671 ( .A(n941), .ZN(n624) );
  NAND2_X1 U672 ( .A1(n603), .A2(n624), .ZN(n604) );
  XNOR2_X1 U673 ( .A(n604), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U674 ( .A1(n624), .A2(G868), .ZN(n605) );
  NOR2_X1 U675 ( .A1(G559), .A2(n605), .ZN(n607) );
  AND2_X1 U676 ( .A1(n669), .A2(n932), .ZN(n606) );
  NOR2_X1 U677 ( .A1(n607), .A2(n606), .ZN(G282) );
  XNOR2_X1 U678 ( .A(G2100), .B(KEYINPUT75), .ZN(n617) );
  NAND2_X1 U679 ( .A1(G123), .A2(n874), .ZN(n608) );
  XNOR2_X1 U680 ( .A(n608), .B(KEYINPUT18), .ZN(n615) );
  NAND2_X1 U681 ( .A1(G111), .A2(n873), .ZN(n610) );
  NAND2_X1 U682 ( .A1(G135), .A2(n870), .ZN(n609) );
  NAND2_X1 U683 ( .A1(n610), .A2(n609), .ZN(n613) );
  NAND2_X1 U684 ( .A1(n869), .A2(G99), .ZN(n611) );
  XOR2_X1 U685 ( .A(KEYINPUT74), .B(n611), .Z(n612) );
  NOR2_X1 U686 ( .A1(n613), .A2(n612), .ZN(n614) );
  NAND2_X1 U687 ( .A1(n615), .A2(n614), .ZN(n868) );
  INV_X1 U688 ( .A(n868), .ZN(n1000) );
  XNOR2_X1 U689 ( .A(n1000), .B(G2096), .ZN(n616) );
  NAND2_X1 U690 ( .A1(n617), .A2(n616), .ZN(G156) );
  NAND2_X1 U691 ( .A1(G67), .A2(n654), .ZN(n619) );
  NAND2_X1 U692 ( .A1(G55), .A2(n655), .ZN(n618) );
  NAND2_X1 U693 ( .A1(n619), .A2(n618), .ZN(n623) );
  NAND2_X1 U694 ( .A1(G80), .A2(n650), .ZN(n621) );
  NAND2_X1 U695 ( .A1(G93), .A2(n651), .ZN(n620) );
  NAND2_X1 U696 ( .A1(n621), .A2(n620), .ZN(n622) );
  OR2_X1 U697 ( .A1(n623), .A2(n622), .ZN(n670) );
  XOR2_X1 U698 ( .A(n932), .B(KEYINPUT76), .Z(n626) );
  NAND2_X1 U699 ( .A1(G559), .A2(n624), .ZN(n625) );
  XNOR2_X1 U700 ( .A(n626), .B(n625), .ZN(n667) );
  NOR2_X1 U701 ( .A1(n667), .A2(G860), .ZN(n627) );
  XOR2_X1 U702 ( .A(KEYINPUT77), .B(n627), .Z(n628) );
  XOR2_X1 U703 ( .A(n670), .B(n628), .Z(G145) );
  NAND2_X1 U704 ( .A1(G49), .A2(n655), .ZN(n630) );
  NAND2_X1 U705 ( .A1(G74), .A2(G651), .ZN(n629) );
  NAND2_X1 U706 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U707 ( .A1(n654), .A2(n631), .ZN(n634) );
  NAND2_X1 U708 ( .A1(G87), .A2(n632), .ZN(n633) );
  NAND2_X1 U709 ( .A1(n634), .A2(n633), .ZN(G288) );
  NAND2_X1 U710 ( .A1(G47), .A2(n655), .ZN(n636) );
  NAND2_X1 U711 ( .A1(G85), .A2(n651), .ZN(n635) );
  NAND2_X1 U712 ( .A1(n636), .A2(n635), .ZN(n639) );
  NAND2_X1 U713 ( .A1(G72), .A2(n650), .ZN(n637) );
  XNOR2_X1 U714 ( .A(KEYINPUT67), .B(n637), .ZN(n638) );
  NOR2_X1 U715 ( .A1(n639), .A2(n638), .ZN(n641) );
  NAND2_X1 U716 ( .A1(n654), .A2(G60), .ZN(n640) );
  NAND2_X1 U717 ( .A1(n641), .A2(n640), .ZN(G290) );
  NAND2_X1 U718 ( .A1(G86), .A2(n651), .ZN(n648) );
  NAND2_X1 U719 ( .A1(G61), .A2(n654), .ZN(n643) );
  NAND2_X1 U720 ( .A1(G48), .A2(n655), .ZN(n642) );
  NAND2_X1 U721 ( .A1(n643), .A2(n642), .ZN(n646) );
  NAND2_X1 U722 ( .A1(n650), .A2(G73), .ZN(n644) );
  XOR2_X1 U723 ( .A(KEYINPUT2), .B(n644), .Z(n645) );
  NOR2_X1 U724 ( .A1(n646), .A2(n645), .ZN(n647) );
  NAND2_X1 U725 ( .A1(n648), .A2(n647), .ZN(n649) );
  XNOR2_X1 U726 ( .A(n649), .B(KEYINPUT78), .ZN(G305) );
  NAND2_X1 U727 ( .A1(G75), .A2(n650), .ZN(n653) );
  NAND2_X1 U728 ( .A1(G88), .A2(n651), .ZN(n652) );
  NAND2_X1 U729 ( .A1(n653), .A2(n652), .ZN(n659) );
  NAND2_X1 U730 ( .A1(G62), .A2(n654), .ZN(n657) );
  NAND2_X1 U731 ( .A1(G50), .A2(n655), .ZN(n656) );
  NAND2_X1 U732 ( .A1(n657), .A2(n656), .ZN(n658) );
  NOR2_X1 U733 ( .A1(n659), .A2(n658), .ZN(G166) );
  INV_X1 U734 ( .A(G166), .ZN(G303) );
  XNOR2_X1 U735 ( .A(KEYINPUT79), .B(KEYINPUT80), .ZN(n661) );
  XNOR2_X1 U736 ( .A(G288), .B(KEYINPUT19), .ZN(n660) );
  XNOR2_X1 U737 ( .A(n661), .B(n660), .ZN(n662) );
  XOR2_X1 U738 ( .A(n670), .B(n662), .Z(n664) );
  XNOR2_X1 U739 ( .A(G290), .B(G305), .ZN(n663) );
  XNOR2_X1 U740 ( .A(n664), .B(n663), .ZN(n665) );
  XNOR2_X1 U741 ( .A(n665), .B(G303), .ZN(n666) );
  XNOR2_X1 U742 ( .A(n666), .B(G299), .ZN(n893) );
  XOR2_X1 U743 ( .A(n893), .B(n667), .Z(n668) );
  NOR2_X1 U744 ( .A1(n669), .A2(n668), .ZN(n672) );
  NOR2_X1 U745 ( .A1(G868), .A2(n670), .ZN(n671) );
  NOR2_X1 U746 ( .A1(n672), .A2(n671), .ZN(G295) );
  NAND2_X1 U747 ( .A1(G2078), .A2(G2084), .ZN(n673) );
  XNOR2_X1 U748 ( .A(n673), .B(KEYINPUT81), .ZN(n674) );
  XNOR2_X1 U749 ( .A(n674), .B(KEYINPUT20), .ZN(n675) );
  NAND2_X1 U750 ( .A1(n675), .A2(G2090), .ZN(n676) );
  XNOR2_X1 U751 ( .A(KEYINPUT21), .B(n676), .ZN(n677) );
  NAND2_X1 U752 ( .A1(n677), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U753 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U754 ( .A(KEYINPUT69), .B(G82), .ZN(G220) );
  NAND2_X1 U755 ( .A1(G120), .A2(G69), .ZN(n678) );
  NOR2_X1 U756 ( .A1(G237), .A2(n678), .ZN(n679) );
  NAND2_X1 U757 ( .A1(G108), .A2(n679), .ZN(n850) );
  NAND2_X1 U758 ( .A1(n850), .A2(G567), .ZN(n685) );
  NOR2_X1 U759 ( .A1(G219), .A2(G220), .ZN(n680) );
  XOR2_X1 U760 ( .A(KEYINPUT22), .B(n680), .Z(n681) );
  NOR2_X1 U761 ( .A1(G218), .A2(n681), .ZN(n682) );
  NAND2_X1 U762 ( .A1(G96), .A2(n682), .ZN(n849) );
  NAND2_X1 U763 ( .A1(G2106), .A2(n849), .ZN(n683) );
  XNOR2_X1 U764 ( .A(KEYINPUT82), .B(n683), .ZN(n684) );
  NAND2_X1 U765 ( .A1(n685), .A2(n684), .ZN(n923) );
  NAND2_X1 U766 ( .A1(G483), .A2(G661), .ZN(n686) );
  NOR2_X1 U767 ( .A1(n923), .A2(n686), .ZN(n848) );
  NAND2_X1 U768 ( .A1(n848), .A2(G36), .ZN(G176) );
  NAND2_X1 U769 ( .A1(G160), .A2(G40), .ZN(n688) );
  INV_X1 U770 ( .A(KEYINPUT84), .ZN(n687) );
  XNOR2_X1 U771 ( .A(n688), .B(n687), .ZN(n764) );
  NAND2_X1 U772 ( .A1(n764), .A2(n765), .ZN(n692) );
  XNOR2_X1 U773 ( .A(n692), .B(n689), .ZN(n690) );
  NAND2_X1 U774 ( .A1(n690), .A2(G1996), .ZN(n691) );
  XNOR2_X1 U775 ( .A(n691), .B(KEYINPUT26), .ZN(n694) );
  XNOR2_X2 U776 ( .A(n692), .B(KEYINPUT64), .ZN(n738) );
  NAND2_X1 U777 ( .A1(G1341), .A2(n738), .ZN(n693) );
  NAND2_X1 U778 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U779 ( .A(n695), .B(KEYINPUT93), .ZN(n696) );
  NAND2_X1 U780 ( .A1(n696), .A2(n932), .ZN(n703) );
  NOR2_X1 U781 ( .A1(n941), .A2(n703), .ZN(n698) );
  XNOR2_X1 U782 ( .A(n698), .B(n697), .ZN(n702) );
  NAND2_X1 U783 ( .A1(n738), .A2(G1348), .ZN(n700) );
  INV_X1 U784 ( .A(n738), .ZN(n720) );
  XOR2_X1 U785 ( .A(KEYINPUT89), .B(n720), .Z(n706) );
  NAND2_X1 U786 ( .A1(G2067), .A2(n706), .ZN(n699) );
  NAND2_X1 U787 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U788 ( .A1(n702), .A2(n701), .ZN(n705) );
  NAND2_X1 U789 ( .A1(n941), .A2(n703), .ZN(n704) );
  NAND2_X1 U790 ( .A1(n705), .A2(n704), .ZN(n712) );
  INV_X1 U791 ( .A(n706), .ZN(n719) );
  INV_X1 U792 ( .A(G2072), .ZN(n976) );
  NOR2_X1 U793 ( .A1(n719), .A2(n976), .ZN(n708) );
  XNOR2_X1 U794 ( .A(KEYINPUT27), .B(KEYINPUT92), .ZN(n707) );
  XNOR2_X1 U795 ( .A(n708), .B(n707), .ZN(n710) );
  NAND2_X1 U796 ( .A1(n719), .A2(G1956), .ZN(n709) );
  NAND2_X1 U797 ( .A1(n710), .A2(n709), .ZN(n714) );
  NAND2_X1 U798 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U799 ( .A(KEYINPUT95), .B(n713), .ZN(n717) );
  NAND2_X1 U800 ( .A1(G299), .A2(n714), .ZN(n715) );
  XOR2_X1 U801 ( .A(KEYINPUT28), .B(n715), .Z(n716) );
  NOR2_X1 U802 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U803 ( .A(n718), .B(KEYINPUT29), .ZN(n725) );
  XOR2_X1 U804 ( .A(G2078), .B(KEYINPUT25), .Z(n983) );
  NOR2_X1 U805 ( .A1(n719), .A2(n983), .ZN(n722) );
  NOR2_X1 U806 ( .A1(G1961), .A2(n720), .ZN(n721) );
  NOR2_X1 U807 ( .A1(n722), .A2(n721), .ZN(n723) );
  XOR2_X1 U808 ( .A(KEYINPUT90), .B(n723), .Z(n730) );
  AND2_X1 U809 ( .A1(G171), .A2(n730), .ZN(n724) );
  NAND2_X1 U810 ( .A1(n738), .A2(G8), .ZN(n804) );
  NOR2_X1 U811 ( .A1(G1966), .A2(n804), .ZN(n752) );
  NOR2_X1 U812 ( .A1(n738), .A2(G2084), .ZN(n750) );
  NOR2_X1 U813 ( .A1(n752), .A2(n750), .ZN(n726) );
  NAND2_X1 U814 ( .A1(G8), .A2(n726), .ZN(n727) );
  XNOR2_X1 U815 ( .A(KEYINPUT30), .B(n727), .ZN(n728) );
  XNOR2_X1 U816 ( .A(n728), .B(KEYINPUT96), .ZN(n729) );
  NOR2_X1 U817 ( .A1(G168), .A2(n729), .ZN(n732) );
  NOR2_X1 U818 ( .A1(G171), .A2(n730), .ZN(n731) );
  NOR2_X1 U819 ( .A1(n732), .A2(n731), .ZN(n733) );
  XOR2_X1 U820 ( .A(KEYINPUT31), .B(n733), .Z(n734) );
  XNOR2_X1 U821 ( .A(n734), .B(KEYINPUT97), .ZN(n735) );
  NOR2_X1 U822 ( .A1(n520), .A2(n735), .ZN(n736) );
  XNOR2_X1 U823 ( .A(n736), .B(KEYINPUT98), .ZN(n751) );
  INV_X1 U824 ( .A(n751), .ZN(n737) );
  NAND2_X1 U825 ( .A1(n737), .A2(G286), .ZN(n746) );
  INV_X1 U826 ( .A(G8), .ZN(n744) );
  NOR2_X1 U827 ( .A1(n738), .A2(G2090), .ZN(n739) );
  XNOR2_X1 U828 ( .A(KEYINPUT99), .B(n739), .ZN(n742) );
  NOR2_X1 U829 ( .A1(G1971), .A2(n804), .ZN(n740) );
  NOR2_X1 U830 ( .A1(G166), .A2(n740), .ZN(n741) );
  NAND2_X1 U831 ( .A1(n742), .A2(n741), .ZN(n743) );
  OR2_X1 U832 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U833 ( .A1(n746), .A2(n745), .ZN(n749) );
  XOR2_X1 U834 ( .A(KEYINPUT32), .B(KEYINPUT101), .Z(n747) );
  XOR2_X1 U835 ( .A(KEYINPUT100), .B(n747), .Z(n748) );
  XNOR2_X1 U836 ( .A(n749), .B(n748), .ZN(n809) );
  NAND2_X1 U837 ( .A1(n750), .A2(G8), .ZN(n754) );
  NOR2_X1 U838 ( .A1(n752), .A2(n751), .ZN(n753) );
  NAND2_X1 U839 ( .A1(n754), .A2(n753), .ZN(n807) );
  NAND2_X1 U840 ( .A1(n809), .A2(n807), .ZN(n763) );
  NAND2_X1 U841 ( .A1(G8), .A2(G166), .ZN(n755) );
  NOR2_X1 U842 ( .A1(G2090), .A2(n755), .ZN(n756) );
  XNOR2_X1 U843 ( .A(n756), .B(KEYINPUT103), .ZN(n761) );
  NOR2_X1 U844 ( .A1(G1981), .A2(G305), .ZN(n757) );
  XOR2_X1 U845 ( .A(n757), .B(KEYINPUT24), .Z(n758) );
  NOR2_X1 U846 ( .A1(n804), .A2(n758), .ZN(n759) );
  XNOR2_X1 U847 ( .A(n759), .B(KEYINPUT88), .ZN(n796) );
  INV_X1 U848 ( .A(n796), .ZN(n760) );
  AND2_X1 U849 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U850 ( .A1(n763), .A2(n762), .ZN(n799) );
  INV_X1 U851 ( .A(n765), .ZN(n766) );
  NAND2_X1 U852 ( .A1(n764), .A2(n766), .ZN(n794) );
  INV_X1 U853 ( .A(n794), .ZN(n838) );
  XNOR2_X1 U854 ( .A(KEYINPUT37), .B(G2067), .ZN(n836) );
  NAND2_X1 U855 ( .A1(G104), .A2(n869), .ZN(n768) );
  NAND2_X1 U856 ( .A1(G140), .A2(n870), .ZN(n767) );
  NAND2_X1 U857 ( .A1(n768), .A2(n767), .ZN(n769) );
  XNOR2_X1 U858 ( .A(KEYINPUT34), .B(n769), .ZN(n775) );
  NAND2_X1 U859 ( .A1(G116), .A2(n873), .ZN(n771) );
  NAND2_X1 U860 ( .A1(G128), .A2(n874), .ZN(n770) );
  NAND2_X1 U861 ( .A1(n771), .A2(n770), .ZN(n772) );
  XNOR2_X1 U862 ( .A(KEYINPUT85), .B(n772), .ZN(n773) );
  XNOR2_X1 U863 ( .A(KEYINPUT35), .B(n773), .ZN(n774) );
  NOR2_X1 U864 ( .A1(n775), .A2(n774), .ZN(n776) );
  XNOR2_X1 U865 ( .A(KEYINPUT36), .B(n776), .ZN(n883) );
  NOR2_X1 U866 ( .A1(n836), .A2(n883), .ZN(n999) );
  NAND2_X1 U867 ( .A1(n838), .A2(n999), .ZN(n834) );
  NAND2_X1 U868 ( .A1(G117), .A2(n873), .ZN(n778) );
  NAND2_X1 U869 ( .A1(G129), .A2(n874), .ZN(n777) );
  NAND2_X1 U870 ( .A1(n778), .A2(n777), .ZN(n779) );
  XNOR2_X1 U871 ( .A(KEYINPUT86), .B(n779), .ZN(n783) );
  NAND2_X1 U872 ( .A1(G105), .A2(n869), .ZN(n780) );
  XNOR2_X1 U873 ( .A(n780), .B(KEYINPUT38), .ZN(n781) );
  XNOR2_X1 U874 ( .A(n781), .B(KEYINPUT87), .ZN(n782) );
  NOR2_X1 U875 ( .A1(n783), .A2(n782), .ZN(n785) );
  NAND2_X1 U876 ( .A1(n870), .A2(G141), .ZN(n784) );
  NAND2_X1 U877 ( .A1(n785), .A2(n784), .ZN(n865) );
  AND2_X1 U878 ( .A1(n865), .A2(G1996), .ZN(n793) );
  NAND2_X1 U879 ( .A1(G95), .A2(n869), .ZN(n787) );
  NAND2_X1 U880 ( .A1(G131), .A2(n870), .ZN(n786) );
  NAND2_X1 U881 ( .A1(n787), .A2(n786), .ZN(n791) );
  NAND2_X1 U882 ( .A1(G107), .A2(n873), .ZN(n789) );
  NAND2_X1 U883 ( .A1(G119), .A2(n874), .ZN(n788) );
  NAND2_X1 U884 ( .A1(n789), .A2(n788), .ZN(n790) );
  OR2_X1 U885 ( .A1(n791), .A2(n790), .ZN(n886) );
  AND2_X1 U886 ( .A1(n886), .A2(G1991), .ZN(n792) );
  NOR2_X1 U887 ( .A1(n793), .A2(n792), .ZN(n996) );
  NOR2_X1 U888 ( .A1(n996), .A2(n794), .ZN(n830) );
  INV_X1 U889 ( .A(n830), .ZN(n795) );
  NAND2_X1 U890 ( .A1(n834), .A2(n795), .ZN(n818) );
  NOR2_X1 U891 ( .A1(n796), .A2(n804), .ZN(n797) );
  NOR2_X1 U892 ( .A1(n818), .A2(n797), .ZN(n798) );
  NAND2_X1 U893 ( .A1(n799), .A2(n798), .ZN(n823) );
  INV_X1 U894 ( .A(n804), .ZN(n801) );
  NAND2_X1 U895 ( .A1(G288), .A2(G1976), .ZN(n800) );
  XNOR2_X1 U896 ( .A(n800), .B(KEYINPUT102), .ZN(n940) );
  AND2_X1 U897 ( .A1(n801), .A2(n940), .ZN(n802) );
  NOR2_X1 U898 ( .A1(KEYINPUT33), .A2(n802), .ZN(n806) );
  NOR2_X1 U899 ( .A1(G1976), .A2(G288), .ZN(n812) );
  NAND2_X1 U900 ( .A1(n812), .A2(KEYINPUT33), .ZN(n803) );
  NOR2_X1 U901 ( .A1(n804), .A2(n803), .ZN(n805) );
  NOR2_X1 U902 ( .A1(n806), .A2(n805), .ZN(n810) );
  AND2_X1 U903 ( .A1(n807), .A2(n810), .ZN(n808) );
  NAND2_X1 U904 ( .A1(n809), .A2(n808), .ZN(n817) );
  INV_X1 U905 ( .A(n810), .ZN(n815) );
  NOR2_X1 U906 ( .A1(G1971), .A2(G303), .ZN(n811) );
  NOR2_X1 U907 ( .A1(n812), .A2(n811), .ZN(n939) );
  INV_X1 U908 ( .A(KEYINPUT33), .ZN(n813) );
  AND2_X1 U909 ( .A1(n939), .A2(n813), .ZN(n814) );
  OR2_X1 U910 ( .A1(n815), .A2(n814), .ZN(n816) );
  NAND2_X1 U911 ( .A1(n817), .A2(n816), .ZN(n821) );
  XOR2_X1 U912 ( .A(G1981), .B(G305), .Z(n929) );
  INV_X1 U913 ( .A(n818), .ZN(n819) );
  AND2_X1 U914 ( .A1(n929), .A2(n819), .ZN(n820) );
  NAND2_X1 U915 ( .A1(n821), .A2(n820), .ZN(n822) );
  NAND2_X1 U916 ( .A1(n823), .A2(n822), .ZN(n825) );
  XNOR2_X1 U917 ( .A(G1986), .B(G290), .ZN(n926) );
  NAND2_X1 U918 ( .A1(n926), .A2(n838), .ZN(n824) );
  NAND2_X1 U919 ( .A1(n825), .A2(n824), .ZN(n841) );
  XOR2_X1 U920 ( .A(KEYINPUT106), .B(KEYINPUT39), .Z(n826) );
  XNOR2_X1 U921 ( .A(KEYINPUT105), .B(n826), .ZN(n833) );
  NOR2_X1 U922 ( .A1(G1996), .A2(n865), .ZN(n1011) );
  NOR2_X1 U923 ( .A1(G1991), .A2(n886), .ZN(n1001) );
  NOR2_X1 U924 ( .A1(G1986), .A2(G290), .ZN(n827) );
  XNOR2_X1 U925 ( .A(KEYINPUT104), .B(n827), .ZN(n828) );
  NOR2_X1 U926 ( .A1(n1001), .A2(n828), .ZN(n829) );
  NOR2_X1 U927 ( .A1(n830), .A2(n829), .ZN(n831) );
  NOR2_X1 U928 ( .A1(n1011), .A2(n831), .ZN(n832) );
  XNOR2_X1 U929 ( .A(n833), .B(n832), .ZN(n835) );
  NAND2_X1 U930 ( .A1(n835), .A2(n834), .ZN(n837) );
  NAND2_X1 U931 ( .A1(n836), .A2(n883), .ZN(n1017) );
  NAND2_X1 U932 ( .A1(n837), .A2(n1017), .ZN(n839) );
  NAND2_X1 U933 ( .A1(n839), .A2(n838), .ZN(n840) );
  NAND2_X1 U934 ( .A1(n841), .A2(n840), .ZN(n842) );
  XNOR2_X1 U935 ( .A(KEYINPUT40), .B(n842), .ZN(G329) );
  NAND2_X1 U936 ( .A1(G2106), .A2(n843), .ZN(G217) );
  INV_X1 U937 ( .A(G661), .ZN(n845) );
  NAND2_X1 U938 ( .A1(G2), .A2(G15), .ZN(n844) );
  NOR2_X1 U939 ( .A1(n845), .A2(n844), .ZN(n846) );
  XOR2_X1 U940 ( .A(KEYINPUT108), .B(n846), .Z(G259) );
  NAND2_X1 U941 ( .A1(G3), .A2(G1), .ZN(n847) );
  NAND2_X1 U942 ( .A1(n848), .A2(n847), .ZN(G188) );
  XNOR2_X1 U943 ( .A(G69), .B(KEYINPUT109), .ZN(G235) );
  INV_X1 U945 ( .A(G120), .ZN(G236) );
  INV_X1 U946 ( .A(G96), .ZN(G221) );
  NOR2_X1 U947 ( .A1(n850), .A2(n849), .ZN(G325) );
  INV_X1 U948 ( .A(G325), .ZN(G261) );
  NAND2_X1 U949 ( .A1(G124), .A2(n874), .ZN(n851) );
  XNOR2_X1 U950 ( .A(n851), .B(KEYINPUT44), .ZN(n853) );
  NAND2_X1 U951 ( .A1(n869), .A2(G100), .ZN(n852) );
  NAND2_X1 U952 ( .A1(n853), .A2(n852), .ZN(n857) );
  NAND2_X1 U953 ( .A1(G112), .A2(n873), .ZN(n855) );
  NAND2_X1 U954 ( .A1(G136), .A2(n870), .ZN(n854) );
  NAND2_X1 U955 ( .A1(n855), .A2(n854), .ZN(n856) );
  NOR2_X1 U956 ( .A1(n857), .A2(n856), .ZN(G162) );
  NAND2_X1 U957 ( .A1(G118), .A2(n873), .ZN(n859) );
  NAND2_X1 U958 ( .A1(G130), .A2(n874), .ZN(n858) );
  NAND2_X1 U959 ( .A1(n859), .A2(n858), .ZN(n864) );
  NAND2_X1 U960 ( .A1(G106), .A2(n869), .ZN(n861) );
  NAND2_X1 U961 ( .A1(G142), .A2(n870), .ZN(n860) );
  NAND2_X1 U962 ( .A1(n861), .A2(n860), .ZN(n862) );
  XOR2_X1 U963 ( .A(n862), .B(KEYINPUT45), .Z(n863) );
  NOR2_X1 U964 ( .A1(n864), .A2(n863), .ZN(n866) );
  XNOR2_X1 U965 ( .A(n866), .B(n865), .ZN(n867) );
  XNOR2_X1 U966 ( .A(G162), .B(n867), .ZN(n885) );
  XNOR2_X1 U967 ( .A(G160), .B(n868), .ZN(n881) );
  NAND2_X1 U968 ( .A1(G103), .A2(n869), .ZN(n872) );
  NAND2_X1 U969 ( .A1(G139), .A2(n870), .ZN(n871) );
  NAND2_X1 U970 ( .A1(n872), .A2(n871), .ZN(n879) );
  NAND2_X1 U971 ( .A1(G115), .A2(n873), .ZN(n876) );
  NAND2_X1 U972 ( .A1(G127), .A2(n874), .ZN(n875) );
  NAND2_X1 U973 ( .A1(n876), .A2(n875), .ZN(n877) );
  XOR2_X1 U974 ( .A(KEYINPUT47), .B(n877), .Z(n878) );
  NOR2_X1 U975 ( .A1(n879), .A2(n878), .ZN(n880) );
  XNOR2_X1 U976 ( .A(KEYINPUT112), .B(n880), .ZN(n1005) );
  XNOR2_X1 U977 ( .A(n881), .B(n1005), .ZN(n882) );
  XNOR2_X1 U978 ( .A(n883), .B(n882), .ZN(n884) );
  XNOR2_X1 U979 ( .A(n885), .B(n884), .ZN(n891) );
  XOR2_X1 U980 ( .A(KEYINPUT113), .B(KEYINPUT46), .Z(n888) );
  XOR2_X1 U981 ( .A(n886), .B(KEYINPUT48), .Z(n887) );
  XNOR2_X1 U982 ( .A(n888), .B(n887), .ZN(n889) );
  XNOR2_X1 U983 ( .A(G164), .B(n889), .ZN(n890) );
  XNOR2_X1 U984 ( .A(n891), .B(n890), .ZN(n892) );
  NOR2_X1 U985 ( .A1(G37), .A2(n892), .ZN(G395) );
  XNOR2_X1 U986 ( .A(G171), .B(n893), .ZN(n895) );
  XNOR2_X1 U987 ( .A(n941), .B(n932), .ZN(n894) );
  XNOR2_X1 U988 ( .A(n895), .B(n894), .ZN(n896) );
  XNOR2_X1 U989 ( .A(n896), .B(G286), .ZN(n897) );
  NOR2_X1 U990 ( .A1(G37), .A2(n897), .ZN(G397) );
  XOR2_X1 U991 ( .A(G2096), .B(G2100), .Z(n899) );
  XNOR2_X1 U992 ( .A(KEYINPUT42), .B(G2678), .ZN(n898) );
  XNOR2_X1 U993 ( .A(n899), .B(n898), .ZN(n903) );
  XOR2_X1 U994 ( .A(KEYINPUT43), .B(G2072), .Z(n901) );
  XNOR2_X1 U995 ( .A(G2067), .B(G2090), .ZN(n900) );
  XNOR2_X1 U996 ( .A(n901), .B(n900), .ZN(n902) );
  XOR2_X1 U997 ( .A(n903), .B(n902), .Z(n905) );
  XNOR2_X1 U998 ( .A(G2078), .B(G2084), .ZN(n904) );
  XNOR2_X1 U999 ( .A(n905), .B(n904), .ZN(G227) );
  XOR2_X1 U1000 ( .A(KEYINPUT41), .B(G1976), .Z(n907) );
  XNOR2_X1 U1001 ( .A(G1996), .B(G1991), .ZN(n906) );
  XNOR2_X1 U1002 ( .A(n907), .B(n906), .ZN(n908) );
  XOR2_X1 U1003 ( .A(n908), .B(KEYINPUT110), .Z(n910) );
  XNOR2_X1 U1004 ( .A(G1981), .B(G1966), .ZN(n909) );
  XNOR2_X1 U1005 ( .A(n910), .B(n909), .ZN(n914) );
  XOR2_X1 U1006 ( .A(G1961), .B(G1956), .Z(n912) );
  XNOR2_X1 U1007 ( .A(G1986), .B(G1971), .ZN(n911) );
  XNOR2_X1 U1008 ( .A(n912), .B(n911), .ZN(n913) );
  XOR2_X1 U1009 ( .A(n914), .B(n913), .Z(n916) );
  XNOR2_X1 U1010 ( .A(KEYINPUT111), .B(G2474), .ZN(n915) );
  XNOR2_X1 U1011 ( .A(n916), .B(n915), .ZN(G229) );
  NOR2_X1 U1012 ( .A1(G401), .A2(n923), .ZN(n920) );
  NOR2_X1 U1013 ( .A1(G227), .A2(G229), .ZN(n917) );
  XNOR2_X1 U1014 ( .A(KEYINPUT49), .B(n917), .ZN(n918) );
  NOR2_X1 U1015 ( .A1(G397), .A2(n918), .ZN(n919) );
  NAND2_X1 U1016 ( .A1(n920), .A2(n919), .ZN(n921) );
  NOR2_X1 U1017 ( .A1(G395), .A2(n921), .ZN(n922) );
  XOR2_X1 U1018 ( .A(KEYINPUT114), .B(n922), .Z(G225) );
  XNOR2_X1 U1019 ( .A(KEYINPUT115), .B(G225), .ZN(G308) );
  INV_X1 U1020 ( .A(n923), .ZN(G319) );
  INV_X1 U1021 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1022 ( .A(G16), .B(KEYINPUT56), .ZN(n924) );
  XNOR2_X1 U1023 ( .A(n924), .B(KEYINPUT122), .ZN(n947) );
  XNOR2_X1 U1024 ( .A(G1956), .B(G299), .ZN(n925) );
  NOR2_X1 U1025 ( .A1(n926), .A2(n925), .ZN(n928) );
  NAND2_X1 U1026 ( .A1(G1971), .A2(G303), .ZN(n927) );
  NAND2_X1 U1027 ( .A1(n928), .A2(n927), .ZN(n938) );
  XNOR2_X1 U1028 ( .A(G168), .B(G1966), .ZN(n930) );
  NAND2_X1 U1029 ( .A1(n930), .A2(n929), .ZN(n931) );
  XNOR2_X1 U1030 ( .A(n931), .B(KEYINPUT57), .ZN(n936) );
  XOR2_X1 U1031 ( .A(n932), .B(G1341), .Z(n934) );
  XNOR2_X1 U1032 ( .A(G301), .B(G1961), .ZN(n933) );
  NOR2_X1 U1033 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1034 ( .A1(n936), .A2(n935), .ZN(n937) );
  NOR2_X1 U1035 ( .A1(n938), .A2(n937), .ZN(n945) );
  NAND2_X1 U1036 ( .A1(n940), .A2(n939), .ZN(n943) );
  XNOR2_X1 U1037 ( .A(G1348), .B(n941), .ZN(n942) );
  NOR2_X1 U1038 ( .A1(n943), .A2(n942), .ZN(n944) );
  NAND2_X1 U1039 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1040 ( .A1(n947), .A2(n946), .ZN(n1026) );
  XNOR2_X1 U1041 ( .A(G1348), .B(KEYINPUT59), .ZN(n948) );
  XNOR2_X1 U1042 ( .A(n948), .B(G4), .ZN(n952) );
  XNOR2_X1 U1043 ( .A(G1981), .B(G6), .ZN(n950) );
  XNOR2_X1 U1044 ( .A(G1341), .B(G19), .ZN(n949) );
  NOR2_X1 U1045 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1046 ( .A1(n952), .A2(n951), .ZN(n955) );
  XOR2_X1 U1047 ( .A(KEYINPUT123), .B(G1956), .Z(n953) );
  XNOR2_X1 U1048 ( .A(G20), .B(n953), .ZN(n954) );
  NOR2_X1 U1049 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1050 ( .A(KEYINPUT60), .B(n956), .ZN(n957) );
  XNOR2_X1 U1051 ( .A(n957), .B(KEYINPUT124), .ZN(n961) );
  XNOR2_X1 U1052 ( .A(G1961), .B(G5), .ZN(n959) );
  XNOR2_X1 U1053 ( .A(G1966), .B(G21), .ZN(n958) );
  NOR2_X1 U1054 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1055 ( .A1(n961), .A2(n960), .ZN(n968) );
  XNOR2_X1 U1056 ( .A(G1976), .B(G23), .ZN(n963) );
  XNOR2_X1 U1057 ( .A(G1971), .B(G22), .ZN(n962) );
  NOR2_X1 U1058 ( .A1(n963), .A2(n962), .ZN(n965) );
  XOR2_X1 U1059 ( .A(G1986), .B(G24), .Z(n964) );
  NAND2_X1 U1060 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1061 ( .A(KEYINPUT58), .B(n966), .ZN(n967) );
  NOR2_X1 U1062 ( .A1(n968), .A2(n967), .ZN(n969) );
  XOR2_X1 U1063 ( .A(KEYINPUT61), .B(n969), .Z(n970) );
  NOR2_X1 U1064 ( .A1(G16), .A2(n970), .ZN(n971) );
  XNOR2_X1 U1065 ( .A(KEYINPUT125), .B(n971), .ZN(n972) );
  NAND2_X1 U1066 ( .A1(n972), .A2(G11), .ZN(n1024) );
  XOR2_X1 U1067 ( .A(G32), .B(G1996), .Z(n987) );
  XNOR2_X1 U1068 ( .A(KEYINPUT118), .B(G25), .ZN(n973) );
  XOR2_X1 U1069 ( .A(n973), .B(G1991), .Z(n974) );
  NAND2_X1 U1070 ( .A1(n974), .A2(G28), .ZN(n975) );
  XNOR2_X1 U1071 ( .A(n975), .B(KEYINPUT119), .ZN(n982) );
  XNOR2_X1 U1072 ( .A(n976), .B(G33), .ZN(n979) );
  XOR2_X1 U1073 ( .A(G2067), .B(G26), .Z(n977) );
  XNOR2_X1 U1074 ( .A(KEYINPUT120), .B(n977), .ZN(n978) );
  NAND2_X1 U1075 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1076 ( .A(n980), .B(KEYINPUT121), .ZN(n981) );
  NAND2_X1 U1077 ( .A1(n982), .A2(n981), .ZN(n985) );
  XNOR2_X1 U1078 ( .A(G27), .B(n983), .ZN(n984) );
  NOR2_X1 U1079 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1080 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1081 ( .A(n988), .B(KEYINPUT53), .ZN(n991) );
  XOR2_X1 U1082 ( .A(G2084), .B(G34), .Z(n989) );
  XNOR2_X1 U1083 ( .A(KEYINPUT54), .B(n989), .ZN(n990) );
  NAND2_X1 U1084 ( .A1(n991), .A2(n990), .ZN(n993) );
  XNOR2_X1 U1085 ( .A(G35), .B(G2090), .ZN(n992) );
  NOR2_X1 U1086 ( .A1(n993), .A2(n992), .ZN(n994) );
  NOR2_X1 U1087 ( .A1(G29), .A2(n994), .ZN(n995) );
  XNOR2_X1 U1088 ( .A(n995), .B(KEYINPUT55), .ZN(n1022) );
  XNOR2_X1 U1089 ( .A(G160), .B(G2084), .ZN(n997) );
  NAND2_X1 U1090 ( .A1(n997), .A2(n996), .ZN(n998) );
  NOR2_X1 U1091 ( .A1(n999), .A2(n998), .ZN(n1003) );
  NOR2_X1 U1092 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1093 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XNOR2_X1 U1094 ( .A(KEYINPUT116), .B(n1004), .ZN(n1016) );
  XNOR2_X1 U1095 ( .A(G2072), .B(KEYINPUT117), .ZN(n1006) );
  XNOR2_X1 U1096 ( .A(n1006), .B(n1005), .ZN(n1008) );
  XOR2_X1 U1097 ( .A(G164), .B(G2078), .Z(n1007) );
  NOR2_X1 U1098 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1099 ( .A(KEYINPUT50), .B(n1009), .ZN(n1014) );
  XOR2_X1 U1100 ( .A(G2090), .B(G162), .Z(n1010) );
  NOR2_X1 U1101 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XOR2_X1 U1102 ( .A(KEYINPUT51), .B(n1012), .Z(n1013) );
  NAND2_X1 U1103 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NOR2_X1 U1104 ( .A1(n1016), .A2(n1015), .ZN(n1018) );
  NAND2_X1 U1105 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1106 ( .A(KEYINPUT52), .B(n1019), .ZN(n1020) );
  NAND2_X1 U1107 ( .A1(G29), .A2(n1020), .ZN(n1021) );
  NAND2_X1 U1108 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NOR2_X1 U1109 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1110 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1111 ( .A(n1027), .B(KEYINPUT126), .ZN(n1028) );
  XNOR2_X1 U1112 ( .A(KEYINPUT62), .B(n1028), .ZN(G150) );
  INV_X1 U1113 ( .A(G150), .ZN(G311) );
endmodule

