//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 1 0 1 0 0 1 1 1 0 0 0 0 0 1 1 0 0 0 1 0 1 0 1 0 0 0 1 1 1 1 0 0 1 0 1 0 0 0 0 1 1 0 1 1 0 1 0 0 1 0 1 0 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:49 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1232, new_n1233, new_n1234, new_n1235, new_n1237,
    new_n1238, new_n1239, new_n1240, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1306, new_n1307, new_n1308;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n202), .A2(G50), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(new_n206), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g0016(.A(KEYINPUT64), .B(G244), .ZN(new_n217));
  AND2_X1   g0017(.A1(new_n217), .A2(G77), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G107), .A2(G264), .ZN(new_n222));
  NAND4_X1  g0022(.A1(new_n219), .A2(new_n220), .A3(new_n221), .A4(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n208), .B1(new_n218), .B2(new_n223), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n211), .B(new_n216), .C1(KEYINPUT1), .C2(new_n224), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n225), .B1(KEYINPUT1), .B2(new_n224), .ZN(G361));
  XNOR2_X1  g0026(.A(G238), .B(G244), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(G232), .ZN(new_n228));
  XNOR2_X1  g0028(.A(KEYINPUT2), .B(G226), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XOR2_X1   g0030(.A(G264), .B(G270), .Z(new_n231));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n230), .B(new_n233), .ZN(G358));
  XNOR2_X1  g0034(.A(G50), .B(G68), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G58), .B(G77), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n235), .B(new_n236), .Z(new_n237));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XNOR2_X1  g0038(.A(G107), .B(G116), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G351));
  XNOR2_X1  g0041(.A(KEYINPUT15), .B(G87), .ZN(new_n242));
  INV_X1    g0042(.A(new_n242), .ZN(new_n243));
  INV_X1    g0043(.A(G33), .ZN(new_n244));
  NOR2_X1   g0044(.A1(new_n244), .A2(G20), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  INV_X1    g0046(.A(G77), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n206), .A2(new_n244), .ZN(new_n248));
  INV_X1    g0048(.A(G58), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(KEYINPUT8), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT8), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G58), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  OAI221_X1 g0054(.A(new_n246), .B1(new_n206), .B2(new_n247), .C1(new_n248), .C2(new_n254), .ZN(new_n255));
  NAND3_X1  g0055(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(new_n214), .ZN(new_n257));
  AND2_X1   g0057(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n259), .A2(new_n214), .A3(new_n256), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n205), .A2(G20), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G77), .ZN(new_n262));
  OAI22_X1  g0062(.A1(new_n260), .A2(new_n262), .B1(G77), .B2(new_n259), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n258), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT65), .ZN(new_n266));
  AND2_X1   g0066(.A1(G33), .A2(G41), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n266), .B1(new_n267), .B2(new_n214), .ZN(new_n268));
  NAND2_X1  g0068(.A1(G33), .A2(G41), .ZN(new_n269));
  NAND4_X1  g0069(.A1(new_n269), .A2(KEYINPUT65), .A3(G1), .A4(G13), .ZN(new_n270));
  AND2_X1   g0070(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n271), .A2(new_n217), .A3(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(new_n272), .ZN(new_n274));
  NAND4_X1  g0074(.A1(new_n268), .A2(new_n274), .A3(G274), .A4(new_n270), .ZN(new_n275));
  AND2_X1   g0075(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G179), .ZN(new_n277));
  OR2_X1    g0077(.A1(KEYINPUT3), .A2(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(KEYINPUT3), .A2(G33), .ZN(new_n279));
  AOI21_X1  g0079(.A(G1698), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G232), .ZN(new_n281));
  XNOR2_X1  g0081(.A(KEYINPUT3), .B(G33), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n282), .A2(G238), .A3(G1698), .ZN(new_n283));
  INV_X1    g0083(.A(G107), .ZN(new_n284));
  OAI211_X1 g0084(.A(new_n281), .B(new_n283), .C1(new_n284), .C2(new_n282), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n267), .A2(new_n214), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n276), .A2(new_n277), .A3(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n276), .A2(new_n287), .ZN(new_n289));
  INV_X1    g0089(.A(G169), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n265), .A2(new_n288), .A3(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G200), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n293), .B1(new_n276), .B2(new_n287), .ZN(new_n294));
  INV_X1    g0094(.A(G190), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n264), .B1(new_n289), .B2(new_n295), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n292), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  XOR2_X1   g0097(.A(new_n297), .B(KEYINPUT66), .Z(new_n298));
  NAND2_X1  g0098(.A1(new_n280), .A2(G222), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n282), .A2(G223), .A3(G1698), .ZN(new_n300));
  OAI211_X1 g0100(.A(new_n299), .B(new_n300), .C1(new_n247), .C2(new_n282), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(new_n286), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n271), .A2(G226), .A3(new_n272), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n302), .A2(new_n275), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(G200), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n261), .A2(G50), .ZN(new_n306));
  OAI22_X1  g0106(.A1(new_n260), .A2(new_n306), .B1(G50), .B2(new_n259), .ZN(new_n307));
  INV_X1    g0107(.A(G150), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n248), .A2(new_n308), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n309), .B1(new_n245), .B2(new_n253), .ZN(new_n310));
  OAI21_X1  g0110(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n307), .B1(new_n312), .B2(new_n257), .ZN(new_n313));
  OR2_X1    g0113(.A1(new_n313), .A2(KEYINPUT9), .ZN(new_n314));
  NAND4_X1  g0114(.A1(new_n302), .A2(G190), .A3(new_n275), .A4(new_n303), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n313), .A2(KEYINPUT9), .ZN(new_n316));
  NAND4_X1  g0116(.A1(new_n305), .A2(new_n314), .A3(new_n315), .A4(new_n316), .ZN(new_n317));
  XNOR2_X1  g0117(.A(new_n317), .B(KEYINPUT10), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n313), .B1(new_n304), .B2(new_n290), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n319), .B1(G179), .B2(new_n304), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n245), .A2(G77), .ZN(new_n323));
  INV_X1    g0123(.A(G50), .ZN(new_n324));
  OAI221_X1 g0124(.A(new_n323), .B1(new_n206), .B2(G68), .C1(new_n324), .C2(new_n248), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n325), .A2(KEYINPUT11), .A3(new_n257), .ZN(new_n326));
  INV_X1    g0126(.A(new_n259), .ZN(new_n327));
  INV_X1    g0127(.A(G68), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  XNOR2_X1  g0129(.A(new_n329), .B(KEYINPUT12), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n261), .A2(G68), .ZN(new_n331));
  OAI211_X1 g0131(.A(new_n326), .B(new_n330), .C1(new_n260), .C2(new_n331), .ZN(new_n332));
  AOI21_X1  g0132(.A(KEYINPUT11), .B1(new_n325), .B2(new_n257), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(G232), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(G1698), .ZN(new_n337));
  AND2_X1   g0137(.A1(KEYINPUT3), .A2(G33), .ZN(new_n338));
  NOR2_X1   g0138(.A1(KEYINPUT3), .A2(G33), .ZN(new_n339));
  OAI221_X1 g0139(.A(new_n337), .B1(G226), .B2(G1698), .C1(new_n338), .C2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(G97), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n244), .A2(new_n342), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n286), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT13), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n268), .A2(G238), .A3(new_n270), .A4(new_n272), .ZN(new_n346));
  NAND4_X1  g0146(.A1(new_n344), .A2(new_n345), .A3(new_n275), .A4(new_n346), .ZN(new_n347));
  NOR2_X1   g0147(.A1(G226), .A2(G1698), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n348), .B1(new_n336), .B2(G1698), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n343), .B1(new_n349), .B2(new_n282), .ZN(new_n350));
  INV_X1    g0150(.A(new_n286), .ZN(new_n351));
  OAI211_X1 g0151(.A(new_n275), .B(new_n346), .C1(new_n350), .C2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(KEYINPUT13), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n347), .A2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT67), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(KEYINPUT14), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n354), .A2(G169), .A3(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n347), .A2(G179), .A3(new_n353), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n356), .B1(new_n354), .B2(G169), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n335), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n354), .A2(G200), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n334), .B(new_n362), .C1(new_n295), .C2(new_n354), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n253), .A2(new_n261), .ZN(new_n366));
  OAI22_X1  g0166(.A1(new_n366), .A2(new_n260), .B1(new_n259), .B2(new_n253), .ZN(new_n367));
  XNOR2_X1  g0167(.A(new_n367), .B(KEYINPUT69), .ZN(new_n368));
  INV_X1    g0168(.A(new_n257), .ZN(new_n369));
  AND2_X1   g0169(.A1(G58), .A2(G68), .ZN(new_n370));
  OAI21_X1  g0170(.A(G20), .B1(new_n370), .B2(new_n201), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n206), .A2(new_n244), .A3(G159), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT68), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n371), .A2(KEYINPUT68), .A3(new_n372), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n338), .A2(new_n339), .ZN(new_n378));
  AOI21_X1  g0178(.A(KEYINPUT7), .B1(new_n378), .B2(new_n206), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT7), .ZN(new_n380));
  NOR4_X1   g0180(.A1(new_n338), .A2(new_n339), .A3(new_n380), .A4(G20), .ZN(new_n381));
  OAI21_X1  g0181(.A(G68), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n377), .A2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT16), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n369), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n377), .A2(new_n382), .A3(KEYINPUT16), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n368), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n268), .A2(G232), .A3(new_n270), .A4(new_n272), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n275), .A2(new_n388), .ZN(new_n389));
  OR2_X1    g0189(.A1(G223), .A2(G1698), .ZN(new_n390));
  INV_X1    g0190(.A(G226), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(G1698), .ZN(new_n392));
  OAI211_X1 g0192(.A(new_n390), .B(new_n392), .C1(new_n338), .C2(new_n339), .ZN(new_n393));
  NAND2_X1  g0193(.A1(G33), .A2(G87), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n351), .B1(new_n395), .B2(KEYINPUT70), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT70), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n393), .A2(new_n397), .A3(new_n394), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n389), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(new_n277), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n400), .B1(G169), .B2(new_n399), .ZN(new_n401));
  OAI21_X1  g0201(.A(KEYINPUT18), .B1(new_n387), .B2(new_n401), .ZN(new_n402));
  AND3_X1   g0202(.A1(new_n371), .A2(KEYINPUT68), .A3(new_n372), .ZN(new_n403));
  AOI21_X1  g0203(.A(KEYINPUT68), .B1(new_n371), .B2(new_n372), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n380), .B1(new_n282), .B2(G20), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n378), .A2(KEYINPUT7), .A3(new_n206), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n328), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n384), .B1(new_n405), .B2(new_n408), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n409), .A2(new_n257), .A3(new_n386), .ZN(new_n410));
  INV_X1    g0210(.A(new_n368), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n399), .A2(G190), .ZN(new_n412));
  AND3_X1   g0212(.A1(new_n393), .A2(new_n397), .A3(new_n394), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n397), .B1(new_n393), .B2(new_n394), .ZN(new_n414));
  NOR3_X1   g0214(.A1(new_n413), .A2(new_n414), .A3(new_n351), .ZN(new_n415));
  OAI21_X1  g0215(.A(G200), .B1(new_n415), .B2(new_n389), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n410), .A2(new_n411), .A3(new_n412), .A4(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT17), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NOR3_X1   g0219(.A1(new_n415), .A2(new_n295), .A3(new_n389), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n395), .A2(KEYINPUT70), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n421), .A2(new_n286), .A3(new_n398), .ZN(new_n422));
  INV_X1    g0222(.A(new_n389), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n293), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n420), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n387), .A2(new_n425), .A3(KEYINPUT17), .ZN(new_n426));
  AOI21_X1  g0226(.A(G169), .B1(new_n422), .B2(new_n423), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n427), .B1(new_n277), .B2(new_n399), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n410), .A2(new_n411), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT18), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n402), .A2(new_n419), .A3(new_n426), .A4(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n298), .A2(new_n322), .A3(new_n365), .A4(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(G33), .A2(G283), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n435), .B(new_n206), .C1(G33), .C2(new_n342), .ZN(new_n436));
  INV_X1    g0236(.A(G116), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(G20), .ZN(new_n438));
  AND3_X1   g0238(.A1(new_n257), .A2(KEYINPUT74), .A3(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(KEYINPUT74), .B1(new_n257), .B2(new_n438), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n436), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT20), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  OAI211_X1 g0243(.A(KEYINPUT20), .B(new_n436), .C1(new_n439), .C2(new_n440), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n205), .A2(G33), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n259), .A2(new_n446), .A3(new_n214), .A4(new_n256), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(G116), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n259), .A2(new_n437), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n445), .A2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(G303), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n278), .A2(new_n452), .A3(new_n279), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(new_n286), .ZN(new_n454));
  INV_X1    g0254(.A(G257), .ZN(new_n455));
  INV_X1    g0255(.A(G1698), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(G264), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(G1698), .ZN(new_n459));
  AOI22_X1  g0259(.A1(new_n457), .A2(new_n459), .B1(new_n278), .B2(new_n279), .ZN(new_n460));
  OAI21_X1  g0260(.A(KEYINPUT73), .B1(new_n454), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n457), .A2(new_n459), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(new_n282), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT73), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n463), .A2(new_n464), .A3(new_n286), .A4(new_n453), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n205), .A2(G45), .ZN(new_n466));
  OR2_X1    g0266(.A1(KEYINPUT5), .A2(G41), .ZN(new_n467));
  NAND2_X1  g0267(.A1(KEYINPUT5), .A2(G41), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n466), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n469), .A2(G274), .A3(new_n268), .A4(new_n270), .ZN(new_n470));
  AND2_X1   g0270(.A1(KEYINPUT5), .A2(G41), .ZN(new_n471));
  NOR2_X1   g0271(.A1(KEYINPUT5), .A2(G41), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n205), .B(G45), .C1(new_n471), .C2(new_n472), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n473), .A2(new_n268), .A3(G270), .A4(new_n270), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n461), .A2(new_n465), .A3(new_n470), .A4(new_n474), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n451), .A2(KEYINPUT76), .A3(G169), .A4(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT21), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT76), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n443), .A2(new_n444), .B1(new_n448), .B2(new_n449), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n475), .A2(G169), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n478), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n476), .A2(new_n477), .A3(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n475), .A2(KEYINPUT21), .A3(G169), .ZN(new_n483));
  AND2_X1   g0283(.A1(new_n470), .A2(new_n474), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n484), .A2(G179), .A3(new_n465), .A4(new_n461), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(new_n451), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT75), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n486), .A2(KEYINPUT75), .A3(new_n451), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n475), .A2(G200), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n479), .B(new_n491), .C1(new_n295), .C2(new_n475), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n482), .A2(new_n489), .A3(new_n490), .A4(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(G250), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(new_n456), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n455), .A2(G1698), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n495), .B(new_n496), .C1(new_n338), .C2(new_n339), .ZN(new_n497));
  NAND2_X1  g0297(.A1(G33), .A2(G294), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(KEYINPUT79), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT79), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n497), .A2(new_n501), .A3(new_n498), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n500), .A2(new_n286), .A3(new_n502), .ZN(new_n503));
  AND4_X1   g0303(.A1(G264), .A2(new_n473), .A3(new_n268), .A4(new_n270), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n503), .A2(new_n470), .A3(new_n505), .ZN(new_n506));
  OAI21_X1  g0306(.A(KEYINPUT80), .B1(new_n506), .B2(G190), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n293), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n351), .B1(new_n499), .B2(KEYINPUT79), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n504), .B1(new_n509), .B2(new_n502), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT80), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n510), .A2(new_n511), .A3(new_n295), .A4(new_n470), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n507), .A2(new_n508), .A3(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(G13), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n514), .A2(G1), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n206), .A2(G107), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT78), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n517), .A2(new_n518), .A3(KEYINPUT25), .ZN(new_n519));
  OR2_X1    g0319(.A1(new_n518), .A2(KEYINPUT25), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n518), .A2(KEYINPUT25), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n520), .A2(new_n515), .A3(new_n516), .A4(new_n521), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n519), .B(new_n522), .C1(new_n284), .C2(new_n447), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n206), .B(G87), .C1(new_n338), .C2(new_n339), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(KEYINPUT22), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT22), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n282), .A2(new_n526), .A3(new_n206), .A4(G87), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  AND3_X1   g0328(.A1(new_n284), .A2(KEYINPUT23), .A3(G20), .ZN(new_n529));
  AOI21_X1  g0329(.A(KEYINPUT23), .B1(new_n284), .B2(G20), .ZN(new_n530));
  NAND2_X1  g0330(.A1(G33), .A2(G116), .ZN(new_n531));
  OAI22_X1  g0331(.A1(new_n529), .A2(new_n530), .B1(G20), .B2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n528), .A2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT77), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n532), .B1(new_n525), .B2(new_n527), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(KEYINPUT77), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n536), .A2(KEYINPUT24), .A3(new_n538), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n537), .A2(KEYINPUT77), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT24), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n369), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n523), .B1(new_n539), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n513), .A2(new_n543), .ZN(new_n544));
  OAI211_X1 g0344(.A(G250), .B(G1698), .C1(new_n338), .C2(new_n339), .ZN(new_n545));
  OAI211_X1 g0345(.A(G244), .B(new_n456), .C1(new_n338), .C2(new_n339), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT4), .ZN(new_n547));
  OAI211_X1 g0347(.A(new_n435), .B(new_n545), .C1(new_n546), .C2(new_n547), .ZN(new_n548));
  AOI21_X1  g0348(.A(KEYINPUT4), .B1(new_n280), .B2(G244), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n286), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n473), .A2(new_n268), .A3(G257), .A4(new_n270), .ZN(new_n551));
  AND2_X1   g0351(.A1(new_n470), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(new_n290), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT6), .ZN(new_n555));
  AND2_X1   g0355(.A1(G97), .A2(G107), .ZN(new_n556));
  NOR2_X1   g0356(.A1(G97), .A2(G107), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n555), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n284), .A2(KEYINPUT6), .A3(G97), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(G20), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n206), .A2(new_n244), .A3(G77), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n284), .B1(new_n406), .B2(new_n407), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n257), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n327), .A2(new_n342), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n566), .B1(new_n447), .B2(new_n342), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n550), .A2(new_n552), .A3(new_n277), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n554), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  OAI21_X1  g0371(.A(G107), .B1(new_n379), .B2(new_n381), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n248), .A2(new_n247), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n573), .B1(new_n560), .B2(G20), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n567), .B1(new_n575), .B2(new_n257), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n550), .A2(new_n552), .A3(G190), .ZN(new_n577));
  AND2_X1   g0377(.A1(new_n550), .A2(new_n552), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n576), .B(new_n577), .C1(new_n578), .C2(new_n293), .ZN(new_n579));
  AND2_X1   g0379(.A1(new_n571), .A2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(new_n531), .ZN(new_n581));
  AND2_X1   g0381(.A1(G244), .A2(G1698), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n581), .B1(new_n282), .B2(new_n582), .ZN(new_n583));
  OAI211_X1 g0383(.A(G238), .B(new_n456), .C1(new_n338), .C2(new_n339), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n351), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(G45), .ZN(new_n586));
  OR3_X1    g0386(.A1(new_n586), .A2(G1), .A3(G274), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n466), .A2(new_n494), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n268), .A2(new_n587), .A3(new_n270), .A4(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(new_n589), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n290), .B1(new_n585), .B2(new_n590), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n582), .B1(new_n338), .B2(new_n339), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n584), .A2(new_n531), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(new_n286), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n594), .A2(new_n277), .A3(new_n589), .ZN(new_n595));
  AND2_X1   g0395(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n206), .B(G68), .C1(new_n338), .C2(new_n339), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(KEYINPUT72), .ZN(new_n598));
  XOR2_X1   g0398(.A(KEYINPUT71), .B(KEYINPUT19), .Z(new_n599));
  NAND2_X1  g0399(.A1(new_n245), .A2(G97), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT72), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n282), .A2(new_n602), .A3(new_n206), .A4(G68), .ZN(new_n603));
  XNOR2_X1  g0403(.A(KEYINPUT71), .B(KEYINPUT19), .ZN(new_n604));
  INV_X1    g0404(.A(G87), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n605), .A2(new_n342), .A3(new_n284), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n206), .B1(new_n244), .B2(new_n342), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n604), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n598), .A2(new_n601), .A3(new_n603), .A4(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n257), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n243), .A2(new_n259), .ZN(new_n611));
  INV_X1    g0411(.A(new_n611), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n610), .B(new_n612), .C1(new_n242), .C2(new_n447), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n447), .A2(new_n605), .ZN(new_n614));
  AOI211_X1 g0414(.A(new_n611), .B(new_n614), .C1(new_n609), .C2(new_n257), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n293), .B1(new_n585), .B2(new_n590), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n594), .A2(new_n295), .A3(new_n589), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  AOI22_X1  g0418(.A1(new_n596), .A2(new_n613), .B1(new_n615), .B2(new_n618), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n544), .A2(new_n580), .A3(new_n619), .ZN(new_n620));
  AOI21_X1  g0420(.A(G169), .B1(new_n510), .B2(new_n470), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n506), .A2(G179), .ZN(new_n622));
  NOR3_X1   g0422(.A1(new_n543), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  NOR4_X1   g0423(.A1(new_n434), .A2(new_n493), .A3(new_n620), .A4(new_n623), .ZN(G372));
  INV_X1    g0424(.A(new_n434), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n447), .A2(new_n242), .ZN(new_n626));
  AOI211_X1 g0426(.A(new_n611), .B(new_n626), .C1(new_n609), .C2(new_n257), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n591), .A2(new_n595), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT26), .ZN(new_n630));
  AND2_X1   g0430(.A1(new_n616), .A2(new_n617), .ZN(new_n631));
  INV_X1    g0431(.A(new_n614), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n610), .A2(new_n612), .A3(new_n632), .ZN(new_n633));
  OAI22_X1  g0433(.A1(new_n631), .A2(new_n633), .B1(new_n627), .B2(new_n628), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n630), .B1(new_n634), .B2(new_n571), .ZN(new_n635));
  AND3_X1   g0435(.A1(new_n550), .A2(new_n552), .A3(new_n277), .ZN(new_n636));
  AOI21_X1  g0436(.A(G169), .B1(new_n550), .B2(new_n552), .ZN(new_n637));
  NOR3_X1   g0437(.A1(new_n636), .A2(new_n576), .A3(new_n637), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n619), .A2(new_n638), .A3(KEYINPUT26), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n629), .B1(new_n635), .B2(new_n639), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n622), .A2(new_n621), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n534), .A2(new_n535), .A3(new_n541), .ZN(new_n642));
  OAI21_X1  g0442(.A(KEYINPUT24), .B1(new_n537), .B2(KEYINPUT77), .ZN(new_n643));
  AOI211_X1 g0443(.A(new_n535), .B(new_n532), .C1(new_n525), .C2(new_n527), .ZN(new_n644));
  OAI211_X1 g0444(.A(new_n642), .B(new_n257), .C1(new_n643), .C2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n523), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n641), .A2(new_n647), .ZN(new_n648));
  AND3_X1   g0448(.A1(new_n482), .A2(new_n648), .A3(new_n487), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n640), .B1(new_n649), .B2(new_n620), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n625), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g0451(.A(new_n651), .B(KEYINPUT81), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n402), .A2(new_n431), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n361), .A2(new_n292), .ZN(new_n654));
  AND3_X1   g0454(.A1(new_n419), .A2(new_n363), .A3(new_n426), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n653), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n318), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n320), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  OR2_X1    g0458(.A1(new_n652), .A2(new_n658), .ZN(G369));
  NAND2_X1  g0459(.A1(new_n515), .A2(new_n206), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n660), .A2(KEYINPUT27), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT82), .ZN(new_n662));
  XNOR2_X1  g0462(.A(new_n661), .B(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(G213), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n664), .B1(new_n660), .B2(KEYINPUT27), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  XNOR2_X1  g0467(.A(KEYINPUT83), .B(G343), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(new_n451), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n670), .B1(new_n482), .B2(new_n487), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT84), .ZN(new_n672));
  OR2_X1    g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  AND4_X1   g0473(.A1(new_n482), .A2(new_n489), .A3(new_n490), .A4(new_n492), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(new_n670), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n671), .A2(new_n672), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n673), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  XOR2_X1   g0477(.A(new_n677), .B(KEYINPUT85), .Z(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(G330), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  AND2_X1   g0480(.A1(new_n508), .A2(new_n512), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n647), .B1(new_n681), .B2(new_n507), .ZN(new_n682));
  AOI211_X1 g0482(.A(new_n623), .B(new_n682), .C1(new_n647), .C2(new_n669), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n667), .A2(new_n668), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n648), .A2(new_n684), .ZN(new_n685));
  OR2_X1    g0485(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n680), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n482), .A2(new_n489), .A3(new_n490), .ZN(new_n688));
  AND2_X1   g0488(.A1(new_n688), .A2(new_n684), .ZN(new_n689));
  AOI22_X1  g0489(.A1(new_n683), .A2(new_n689), .B1(new_n623), .B2(new_n684), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n687), .A2(new_n690), .ZN(G399));
  INV_X1    g0491(.A(new_n209), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n692), .A2(G41), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n606), .A2(G116), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n694), .A2(G1), .A3(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n696), .B1(new_n212), .B2(new_n694), .ZN(new_n697));
  XNOR2_X1  g0497(.A(new_n697), .B(KEYINPUT28), .ZN(new_n698));
  INV_X1    g0498(.A(new_n629), .ZN(new_n699));
  NOR3_X1   g0499(.A1(new_n634), .A2(new_n571), .A3(new_n630), .ZN(new_n700));
  AOI21_X1  g0500(.A(KEYINPUT26), .B1(new_n619), .B2(new_n638), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n699), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n619), .A2(new_n571), .A3(new_n579), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n682), .A2(new_n703), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n482), .A2(new_n648), .A3(new_n489), .A4(new_n490), .ZN(new_n705));
  AOI22_X1  g0505(.A1(new_n702), .A2(KEYINPUT87), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT87), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n640), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n669), .B1(new_n706), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(KEYINPUT29), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n650), .A2(new_n684), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT29), .ZN(new_n712));
  AOI21_X1  g0512(.A(KEYINPUT88), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n710), .A2(new_n713), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n709), .A2(KEYINPUT88), .A3(KEYINPUT29), .ZN(new_n715));
  AND2_X1   g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n669), .B1(new_n641), .B2(new_n647), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n674), .A2(new_n704), .A3(KEYINPUT86), .A4(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT86), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n717), .A2(new_n544), .A3(new_n580), .A4(new_n619), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n719), .B1(new_n720), .B2(new_n493), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n718), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT30), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n585), .A2(new_n590), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n578), .A2(new_n510), .A3(new_n724), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n723), .B1(new_n725), .B2(new_n485), .ZN(new_n726));
  AND2_X1   g0526(.A1(new_n510), .A2(new_n724), .ZN(new_n727));
  INV_X1    g0527(.A(new_n485), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n727), .A2(new_n728), .A3(KEYINPUT30), .A4(new_n578), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n724), .A2(G179), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n730), .A2(new_n506), .A3(new_n475), .A4(new_n553), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n726), .A2(new_n729), .A3(new_n731), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n732), .A2(KEYINPUT31), .A3(new_n669), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(KEYINPUT31), .B1(new_n732), .B2(new_n669), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n722), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(G330), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n716), .A2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n698), .B1(new_n740), .B2(G1), .ZN(G364));
  NOR2_X1   g0541(.A1(new_n514), .A2(G20), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n205), .B1(new_n742), .B2(G45), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n693), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n680), .A2(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n746), .B1(G330), .B2(new_n678), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n214), .B1(G20), .B2(new_n290), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n206), .A2(new_n277), .ZN(new_n750));
  NOR2_X1   g0550(.A1(G190), .A2(G200), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n206), .A2(G179), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(new_n751), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  AOI22_X1  g0556(.A1(G311), .A2(new_n753), .B1(new_n756), .B2(G329), .ZN(new_n757));
  INV_X1    g0557(.A(G322), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n750), .A2(G190), .A3(new_n293), .ZN(new_n759));
  OAI211_X1 g0559(.A(new_n757), .B(new_n378), .C1(new_n758), .C2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n750), .ZN(new_n761));
  NOR3_X1   g0561(.A1(new_n761), .A2(G190), .A3(new_n293), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  XOR2_X1   g0563(.A(KEYINPUT33), .B(G317), .Z(new_n764));
  NAND3_X1  g0564(.A1(new_n754), .A2(new_n295), .A3(G200), .ZN(new_n765));
  INV_X1    g0565(.A(G283), .ZN(new_n766));
  OAI22_X1  g0566(.A1(new_n763), .A2(new_n764), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NOR3_X1   g0567(.A1(new_n295), .A2(G179), .A3(G200), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(new_n206), .ZN(new_n769));
  INV_X1    g0569(.A(G294), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n750), .A2(G190), .A3(G200), .ZN(new_n771));
  INV_X1    g0571(.A(G326), .ZN(new_n772));
  OAI22_X1  g0572(.A1(new_n769), .A2(new_n770), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NOR3_X1   g0573(.A1(new_n760), .A2(new_n767), .A3(new_n773), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n754), .A2(G190), .A3(G200), .ZN(new_n775));
  INV_X1    g0575(.A(KEYINPUT92), .ZN(new_n776));
  OR2_X1    g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n775), .A2(new_n776), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g0579(.A(new_n779), .B(KEYINPUT94), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n774), .B1(new_n781), .B2(new_n452), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n282), .B1(new_n779), .B2(new_n605), .ZN(new_n783));
  INV_X1    g0583(.A(KEYINPUT93), .ZN(new_n784));
  OR2_X1    g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n759), .ZN(new_n786));
  AOI22_X1  g0586(.A1(new_n786), .A2(G58), .B1(new_n753), .B2(G77), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n787), .B1(new_n328), .B2(new_n763), .ZN(new_n788));
  INV_X1    g0588(.A(KEYINPUT32), .ZN(new_n789));
  INV_X1    g0589(.A(G159), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n789), .B1(new_n755), .B2(new_n790), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n756), .A2(KEYINPUT32), .A3(G159), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n788), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n783), .A2(new_n784), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n765), .A2(new_n284), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n769), .A2(new_n342), .ZN(new_n796));
  INV_X1    g0596(.A(new_n771), .ZN(new_n797));
  AOI211_X1 g0597(.A(new_n795), .B(new_n796), .C1(G50), .C2(new_n797), .ZN(new_n798));
  NAND4_X1  g0598(.A1(new_n785), .A2(new_n793), .A3(new_n794), .A4(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n749), .B1(new_n782), .B2(new_n799), .ZN(new_n800));
  XNOR2_X1  g0600(.A(new_n745), .B(KEYINPUT89), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(G13), .A2(G33), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n804), .A2(G20), .ZN(new_n805));
  XOR2_X1   g0605(.A(new_n805), .B(KEYINPUT91), .Z(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n692), .A2(new_n282), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n809), .B1(new_n586), .B2(new_n213), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n810), .B1(new_n586), .B2(new_n237), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n692), .A2(new_n378), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n812), .A2(G355), .B1(new_n437), .B2(new_n692), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(KEYINPUT90), .ZN(new_n816));
  AOI211_X1 g0616(.A(new_n807), .B(new_n748), .C1(new_n815), .C2(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n814), .A2(KEYINPUT90), .ZN(new_n818));
  AOI211_X1 g0618(.A(new_n800), .B(new_n802), .C1(new_n817), .C2(new_n818), .ZN(new_n819));
  XNOR2_X1  g0619(.A(new_n819), .B(KEYINPUT95), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n820), .B1(new_n678), .B2(new_n806), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n747), .A2(new_n821), .ZN(G396));
  NOR2_X1   g0622(.A1(new_n748), .A2(new_n803), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n802), .B1(new_n247), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n780), .A2(G107), .ZN(new_n825));
  AOI22_X1  g0625(.A1(new_n762), .A2(G283), .B1(G116), .B2(new_n753), .ZN(new_n826));
  XOR2_X1   g0626(.A(new_n826), .B(KEYINPUT96), .Z(new_n827));
  INV_X1    g0627(.A(G311), .ZN(new_n828));
  OAI221_X1 g0628(.A(new_n378), .B1(new_n755), .B2(new_n828), .C1(new_n759), .C2(new_n770), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n765), .A2(new_n605), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n796), .A2(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n831), .B1(new_n452), .B2(new_n771), .ZN(new_n832));
  NOR3_X1   g0632(.A1(new_n827), .A2(new_n829), .A3(new_n832), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n765), .A2(new_n328), .ZN(new_n834));
  INV_X1    g0634(.A(G132), .ZN(new_n835));
  OAI221_X1 g0635(.A(new_n282), .B1(new_n755), .B2(new_n835), .C1(new_n769), .C2(new_n249), .ZN(new_n836));
  AOI211_X1 g0636(.A(new_n834), .B(new_n836), .C1(new_n780), .C2(G50), .ZN(new_n837));
  AOI22_X1  g0637(.A1(new_n786), .A2(G143), .B1(new_n753), .B2(G159), .ZN(new_n838));
  INV_X1    g0638(.A(G137), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n838), .B1(new_n839), .B2(new_n771), .C1(new_n308), .C2(new_n763), .ZN(new_n840));
  XNOR2_X1  g0640(.A(new_n840), .B(KEYINPUT34), .ZN(new_n841));
  AOI22_X1  g0641(.A1(new_n825), .A2(new_n833), .B1(new_n837), .B2(new_n841), .ZN(new_n842));
  NAND4_X1  g0642(.A1(new_n265), .A2(new_n291), .A3(new_n288), .A4(new_n684), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(new_n844));
  OAI22_X1  g0644(.A1(new_n296), .A2(new_n294), .B1(new_n264), .B2(new_n684), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n844), .B1(new_n292), .B2(new_n845), .ZN(new_n846));
  OAI221_X1 g0646(.A(new_n824), .B1(new_n749), .B2(new_n842), .C1(new_n846), .C2(new_n804), .ZN(new_n847));
  INV_X1    g0647(.A(new_n846), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n711), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n650), .A2(new_n684), .A3(new_n846), .ZN(new_n850));
  AND2_X1   g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n745), .B1(new_n852), .B2(new_n738), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n852), .A2(new_n738), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n847), .B1(new_n854), .B2(new_n855), .ZN(G384));
  OR2_X1    g0656(.A1(new_n560), .A2(KEYINPUT35), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n560), .A2(KEYINPUT35), .ZN(new_n858));
  NAND4_X1  g0658(.A1(new_n857), .A2(G116), .A3(new_n215), .A4(new_n858), .ZN(new_n859));
  XOR2_X1   g0659(.A(KEYINPUT97), .B(KEYINPUT36), .Z(new_n860));
  XNOR2_X1  g0660(.A(new_n859), .B(new_n860), .ZN(new_n861));
  OR3_X1    g0661(.A1(new_n212), .A2(new_n247), .A3(new_n370), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n324), .A2(G68), .ZN(new_n863));
  AOI211_X1 g0663(.A(new_n205), .B(G13), .C1(new_n862), .C2(new_n863), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT99), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT98), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n867), .A2(KEYINPUT37), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n417), .B1(new_n387), .B2(new_n666), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n867), .A2(KEYINPUT37), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n871), .B1(new_n387), .B2(new_n401), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n869), .B1(new_n870), .B2(new_n872), .ZN(new_n873));
  AOI22_X1  g0673(.A1(new_n428), .A2(new_n429), .B1(new_n867), .B2(KEYINPUT37), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n429), .A2(new_n667), .ZN(new_n875));
  NAND4_X1  g0675(.A1(new_n874), .A2(new_n417), .A3(new_n875), .A4(new_n868), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n873), .A2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n875), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n432), .A2(new_n878), .ZN(new_n879));
  AND3_X1   g0679(.A1(new_n877), .A2(new_n879), .A3(KEYINPUT38), .ZN(new_n880));
  AOI21_X1  g0680(.A(KEYINPUT38), .B1(new_n877), .B2(new_n879), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n866), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n877), .A2(new_n879), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT38), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n877), .A2(new_n879), .A3(KEYINPUT38), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n885), .A2(KEYINPUT99), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n882), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n669), .A2(new_n335), .ZN(new_n889));
  AND3_X1   g0689(.A1(new_n361), .A2(new_n363), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n889), .B1(new_n361), .B2(new_n363), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n846), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n892), .B1(new_n722), .B2(new_n736), .ZN(new_n893));
  AOI21_X1  g0693(.A(KEYINPUT40), .B1(new_n888), .B2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT40), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n895), .B1(new_n885), .B2(new_n886), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n894), .B1(new_n893), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n732), .A2(new_n669), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT31), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(new_n733), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n901), .B1(new_n721), .B2(new_n718), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n434), .A2(new_n902), .ZN(new_n903));
  OAI21_X1  g0703(.A(G330), .B1(new_n897), .B2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT100), .ZN(new_n905));
  OR2_X1    g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n904), .A2(new_n905), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n897), .A2(new_n903), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n906), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n890), .A2(new_n891), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n910), .B1(new_n850), .B2(new_n843), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n888), .A2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT39), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n913), .B1(new_n880), .B2(new_n881), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n885), .A2(KEYINPUT39), .A3(new_n886), .ZN(new_n915));
  OR2_X1    g0715(.A1(new_n361), .A2(new_n669), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n914), .A2(new_n915), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n653), .A2(new_n666), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n912), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n434), .B1(new_n714), .B2(new_n715), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n922), .A2(new_n658), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n921), .B(new_n923), .ZN(new_n924));
  AND2_X1   g0724(.A1(new_n909), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(KEYINPUT101), .ZN(new_n926));
  OAI221_X1 g0726(.A(new_n926), .B1(new_n205), .B2(new_n742), .C1(new_n924), .C2(new_n909), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n925), .A2(KEYINPUT101), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n865), .B1(new_n927), .B2(new_n928), .ZN(G367));
  NAND2_X1  g0729(.A1(new_n669), .A2(new_n569), .ZN(new_n930));
  AND2_X1   g0730(.A1(new_n580), .A2(new_n930), .ZN(new_n931));
  NOR3_X1   g0731(.A1(new_n930), .A2(new_n636), .A3(new_n637), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT103), .ZN(new_n933));
  OR3_X1    g0733(.A1(new_n931), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n932), .A2(new_n933), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n683), .A2(new_n689), .ZN(new_n937));
  OR2_X1    g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n571), .B1(new_n936), .B2(new_n648), .ZN(new_n939));
  AOI22_X1  g0739(.A1(new_n938), .A2(KEYINPUT42), .B1(new_n939), .B2(new_n684), .ZN(new_n940));
  OR2_X1    g0740(.A1(new_n938), .A2(KEYINPUT42), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n669), .A2(new_n633), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n942), .A2(new_n699), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n943), .A2(KEYINPUT102), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n942), .A2(new_n619), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n943), .A2(KEYINPUT102), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  AOI22_X1  g0749(.A1(new_n940), .A2(new_n941), .B1(KEYINPUT43), .B2(new_n949), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n949), .A2(KEYINPUT43), .ZN(new_n951));
  XOR2_X1   g0751(.A(new_n950), .B(new_n951), .Z(new_n952));
  NOR2_X1   g0752(.A1(new_n687), .A2(new_n936), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n952), .B(new_n953), .ZN(new_n954));
  XOR2_X1   g0754(.A(new_n693), .B(KEYINPUT41), .Z(new_n955));
  OAI21_X1  g0755(.A(new_n937), .B1(new_n686), .B2(new_n689), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n679), .B(new_n956), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n957), .A2(new_n739), .ZN(new_n958));
  INV_X1    g0758(.A(new_n936), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT44), .ZN(new_n960));
  OR3_X1    g0760(.A1(new_n959), .A2(new_n690), .A3(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n960), .B1(new_n959), .B2(new_n690), .ZN(new_n962));
  AND2_X1   g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n959), .A2(new_n690), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n964), .B(KEYINPUT45), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  OR2_X1    g0766(.A1(new_n966), .A2(new_n687), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n687), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n958), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n955), .B1(new_n969), .B2(new_n740), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n954), .B1(new_n970), .B2(new_n744), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n807), .A2(new_n748), .ZN(new_n972));
  OAI221_X1 g0772(.A(new_n972), .B1(new_n209), .B2(new_n242), .C1(new_n233), .C2(new_n809), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(new_n801), .ZN(new_n974));
  XOR2_X1   g0774(.A(new_n974), .B(KEYINPUT104), .Z(new_n975));
  OAI221_X1 g0775(.A(new_n282), .B1(new_n755), .B2(new_n839), .C1(new_n324), .C2(new_n752), .ZN(new_n976));
  OAI22_X1  g0776(.A1(new_n763), .A2(new_n790), .B1(new_n247), .B2(new_n765), .ZN(new_n977));
  AOI211_X1 g0777(.A(new_n976), .B(new_n977), .C1(G143), .C2(new_n797), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n769), .A2(new_n328), .ZN(new_n979));
  INV_X1    g0779(.A(new_n979), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n980), .B1(new_n308), .B2(new_n759), .ZN(new_n981));
  INV_X1    g0781(.A(new_n779), .ZN(new_n982));
  AOI22_X1  g0782(.A1(new_n981), .A2(KEYINPUT109), .B1(new_n982), .B2(G58), .ZN(new_n983));
  OAI211_X1 g0783(.A(new_n978), .B(new_n983), .C1(KEYINPUT109), .C2(new_n981), .ZN(new_n984));
  AOI21_X1  g0784(.A(KEYINPUT46), .B1(new_n982), .B2(G116), .ZN(new_n985));
  XOR2_X1   g0785(.A(new_n985), .B(KEYINPUT107), .Z(new_n986));
  NAND3_X1  g0786(.A1(new_n780), .A2(KEYINPUT46), .A3(G116), .ZN(new_n987));
  INV_X1    g0787(.A(new_n769), .ZN(new_n988));
  AOI22_X1  g0788(.A1(new_n988), .A2(G107), .B1(new_n753), .B2(G283), .ZN(new_n989));
  INV_X1    g0789(.A(G317), .ZN(new_n990));
  OAI221_X1 g0790(.A(new_n378), .B1(new_n755), .B2(new_n990), .C1(new_n342), .C2(new_n765), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n989), .A2(KEYINPUT105), .B1(new_n991), .B2(KEYINPUT108), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n992), .B1(KEYINPUT105), .B2(new_n989), .ZN(new_n993));
  OAI22_X1  g0793(.A1(new_n759), .A2(new_n452), .B1(new_n771), .B2(new_n828), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(KEYINPUT106), .ZN(new_n995));
  AOI22_X1  g0795(.A1(new_n991), .A2(KEYINPUT108), .B1(G294), .B2(new_n762), .ZN(new_n996));
  NAND4_X1  g0796(.A1(new_n987), .A2(new_n993), .A3(new_n995), .A4(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n984), .B1(new_n986), .B2(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT47), .ZN(new_n999));
  OR2_X1    g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n749), .B1(new_n998), .B2(new_n999), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n975), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(new_n949), .B2(new_n806), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n971), .A2(new_n1003), .ZN(G387));
  XOR2_X1   g0804(.A(new_n679), .B(new_n956), .Z(new_n1005));
  NAND2_X1  g0805(.A1(new_n1005), .A2(new_n744), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n378), .B1(new_n755), .B2(new_n772), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(new_n786), .A2(G317), .B1(new_n753), .B2(G303), .ZN(new_n1008));
  OAI221_X1 g0808(.A(new_n1008), .B1(new_n758), .B2(new_n771), .C1(new_n828), .C2(new_n763), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT48), .ZN(new_n1010));
  OR2_X1    g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n982), .A2(G294), .B1(G283), .B2(new_n988), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1011), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1014));
  XOR2_X1   g0814(.A(new_n1014), .B(KEYINPUT49), .Z(new_n1015));
  INV_X1    g0815(.A(new_n765), .ZN(new_n1016));
  AOI211_X1 g0816(.A(new_n1007), .B(new_n1015), .C1(G116), .C2(new_n1016), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(G68), .A2(new_n753), .B1(new_n756), .B2(G150), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n1018), .B(new_n282), .C1(new_n324), .C2(new_n759), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(G159), .A2(new_n797), .B1(new_n1016), .B2(G97), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n1020), .B1(new_n242), .B2(new_n769), .C1(new_n254), .C2(new_n763), .ZN(new_n1021));
  AOI211_X1 g0821(.A(new_n1019), .B(new_n1021), .C1(G77), .C2(new_n982), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n748), .B1(new_n1017), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n695), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n812), .A2(new_n1024), .B1(new_n284), .B2(new_n692), .ZN(new_n1025));
  XOR2_X1   g0825(.A(new_n1025), .B(KEYINPUT110), .Z(new_n1026));
  NOR2_X1   g0826(.A1(new_n230), .A2(new_n586), .ZN(new_n1027));
  AOI21_X1  g0827(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1028));
  AND3_X1   g0828(.A1(new_n253), .A2(KEYINPUT50), .A3(new_n324), .ZN(new_n1029));
  AOI21_X1  g0829(.A(KEYINPUT50), .B1(new_n253), .B2(new_n324), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n695), .B(new_n1028), .C1(new_n1029), .C2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1031), .A2(new_n808), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1026), .B1(new_n1027), .B2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n802), .B1(new_n1033), .B2(new_n972), .ZN(new_n1034));
  OAI211_X1 g0834(.A(new_n1023), .B(new_n1034), .C1(new_n686), .C2(new_n806), .ZN(new_n1035));
  AND2_X1   g0835(.A1(new_n1006), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n958), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1037), .A2(new_n693), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n1005), .A2(new_n740), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1036), .B1(new_n1038), .B2(new_n1039), .ZN(G393));
  OAI21_X1  g0840(.A(new_n972), .B1(new_n342), .B2(new_n209), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n809), .A2(new_n240), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n801), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n759), .A2(new_n828), .B1(new_n771), .B2(new_n990), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT52), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n769), .A2(new_n437), .ZN(new_n1046));
  AOI211_X1 g0846(.A(new_n795), .B(new_n1046), .C1(G303), .C2(new_n762), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n982), .A2(G283), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n378), .B1(new_n752), .B2(new_n770), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1049), .B1(G322), .B2(new_n756), .ZN(new_n1050));
  NAND4_X1  g0850(.A1(new_n1045), .A2(new_n1047), .A3(new_n1048), .A4(new_n1050), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n759), .A2(new_n790), .B1(new_n771), .B2(new_n308), .ZN(new_n1052));
  XOR2_X1   g0852(.A(new_n1052), .B(KEYINPUT111), .Z(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT51), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n769), .A2(new_n247), .ZN(new_n1055));
  AOI211_X1 g0855(.A(new_n830), .B(new_n1055), .C1(G50), .C2(new_n762), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n982), .A2(G68), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n756), .A2(G143), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n378), .B1(new_n753), .B2(new_n253), .ZN(new_n1059));
  NAND4_X1  g0859(.A1(new_n1056), .A2(new_n1057), .A3(new_n1058), .A4(new_n1059), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1051), .B1(new_n1054), .B2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1043), .B1(new_n1061), .B2(new_n748), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1062), .B1(new_n959), .B2(new_n806), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n967), .A2(new_n968), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1063), .B1(new_n1064), .B2(new_n743), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT112), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  OAI211_X1 g0867(.A(KEYINPUT112), .B(new_n1063), .C1(new_n1064), .C2(new_n743), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1064), .A2(new_n1037), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1070), .A2(new_n693), .A3(new_n969), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1069), .A2(new_n1071), .ZN(G390));
  INV_X1    g0872(.A(G330), .ZN(new_n1073));
  NOR4_X1   g0873(.A1(new_n902), .A2(KEYINPUT113), .A3(new_n1073), .A4(new_n892), .ZN(new_n1074));
  INV_X1    g0874(.A(KEYINPUT113), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1075), .B1(new_n893), .B2(G330), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n845), .A2(new_n292), .ZN(new_n1078));
  AND4_X1   g0878(.A1(new_n482), .A2(new_n648), .A3(new_n489), .A4(new_n490), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n1079), .A2(new_n620), .B1(new_n640), .B2(new_n707), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n702), .A2(KEYINPUT87), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n684), .B(new_n1078), .C1(new_n1080), .C2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n843), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n737), .A2(G330), .A3(new_n846), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1083), .B1(new_n1084), .B2(new_n910), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1077), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n893), .A2(G330), .ZN(new_n1087));
  NOR3_X1   g0887(.A1(new_n902), .A2(new_n1073), .A3(new_n848), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n910), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1087), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n850), .A2(new_n843), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1086), .A2(new_n1092), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n738), .A2(new_n434), .ZN(new_n1094));
  NOR3_X1   g0894(.A1(new_n922), .A2(new_n658), .A3(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n916), .B1(new_n880), .B2(new_n881), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n844), .B1(new_n709), .B2(new_n1078), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1098), .B1(new_n1099), .B2(new_n910), .ZN(new_n1100));
  NOR3_X1   g0900(.A1(new_n880), .A2(new_n881), .A3(new_n913), .ZN(new_n1101));
  AOI21_X1  g0901(.A(KEYINPUT39), .B1(new_n885), .B2(new_n886), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n1101), .A2(new_n1102), .B1(new_n911), .B2(new_n917), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1087), .A2(KEYINPUT113), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n893), .A2(new_n1075), .A3(G330), .ZN(new_n1105));
  NAND4_X1  g0905(.A1(new_n1100), .A2(new_n1103), .A3(new_n1104), .A4(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1087), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1091), .A2(new_n1089), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n1108), .A2(new_n916), .B1(new_n914), .B2(new_n915), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1097), .B1(new_n1083), .B2(new_n1089), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1107), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1106), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1096), .A2(new_n1112), .ZN(new_n1113));
  NAND4_X1  g0913(.A1(new_n1093), .A2(new_n1111), .A3(new_n1095), .A4(new_n1106), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1113), .A2(new_n693), .A3(new_n1114), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n1112), .A2(new_n743), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n803), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1117));
  OAI221_X1 g0917(.A(new_n378), .B1(new_n752), .B2(new_n342), .C1(new_n437), .C2(new_n759), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n763), .A2(new_n284), .B1(new_n247), .B2(new_n769), .ZN(new_n1119));
  AOI211_X1 g0919(.A(new_n1118), .B(new_n1119), .C1(G283), .C2(new_n797), .ZN(new_n1120));
  OAI22_X1  g0920(.A1(new_n765), .A2(new_n328), .B1(new_n755), .B2(new_n770), .ZN(new_n1121));
  XNOR2_X1  g0921(.A(new_n1121), .B(KEYINPUT115), .ZN(new_n1122));
  OAI211_X1 g0922(.A(new_n1120), .B(new_n1122), .C1(new_n605), .C2(new_n781), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(KEYINPUT54), .B(G143), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n763), .A2(new_n839), .B1(new_n752), .B2(new_n1124), .ZN(new_n1125));
  XOR2_X1   g0925(.A(new_n1125), .B(KEYINPUT114), .Z(new_n1126));
  NOR2_X1   g0926(.A1(new_n779), .A2(new_n308), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(new_n1127), .B(KEYINPUT53), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n769), .A2(new_n790), .B1(new_n765), .B2(new_n324), .ZN(new_n1129));
  INV_X1    g0929(.A(G125), .ZN(new_n1130));
  OAI221_X1 g0930(.A(new_n282), .B1(new_n755), .B2(new_n1130), .C1(new_n759), .C2(new_n835), .ZN(new_n1131));
  AOI211_X1 g0931(.A(new_n1129), .B(new_n1131), .C1(G128), .C2(new_n797), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1126), .A2(new_n1128), .A3(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n749), .B1(new_n1123), .B2(new_n1133), .ZN(new_n1134));
  AOI211_X1 g0934(.A(new_n802), .B(new_n1134), .C1(new_n254), .C2(new_n823), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1116), .B1(new_n1117), .B2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1115), .A2(new_n1136), .ZN(G378));
  INV_X1    g0937(.A(KEYINPUT57), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(new_n1114), .B2(new_n1095), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT119), .ZN(new_n1140));
  AOI211_X1 g0940(.A(new_n313), .B(new_n666), .C1(new_n318), .C2(new_n320), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n666), .A2(new_n313), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n321), .A2(new_n1142), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  OR3_X1    g0945(.A1(new_n1141), .A2(new_n1143), .A3(new_n1145), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1145), .B1(new_n1141), .B2(new_n1143), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n896), .A2(new_n893), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1149), .A2(G330), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1148), .B1(new_n894), .B2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1073), .B1(new_n896), .B2(new_n893), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1148), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n892), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n737), .A2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1155), .B1(new_n882), .B2(new_n887), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n1152), .B(new_n1153), .C1(new_n1156), .C2(KEYINPUT40), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1151), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1158), .A2(new_n921), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1151), .A2(new_n1157), .A3(new_n920), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1140), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(new_n1140), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1139), .B1(new_n1161), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(KEYINPUT120), .ZN(new_n1165));
  INV_X1    g0965(.A(KEYINPUT120), .ZN(new_n1166));
  OAI211_X1 g0966(.A(new_n1139), .B(new_n1166), .C1(new_n1161), .C2(new_n1163), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n1077), .A2(new_n1085), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1095), .B1(new_n1112), .B2(new_n1168), .ZN(new_n1169));
  AND3_X1   g0969(.A1(new_n1151), .A2(new_n1157), .A3(new_n920), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n920), .B1(new_n1151), .B2(new_n1157), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1169), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n694), .B1(new_n1172), .B2(new_n1138), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1165), .A2(new_n1167), .A3(new_n1173), .ZN(new_n1174));
  OR2_X1    g0974(.A1(new_n282), .A2(G41), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n1175), .B(new_n324), .C1(G33), .C2(G41), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n762), .A2(G97), .B1(new_n797), .B2(G116), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1016), .A2(G58), .ZN(new_n1178));
  AND3_X1   g0978(.A1(new_n1177), .A2(new_n980), .A3(new_n1178), .ZN(new_n1179));
  OAI22_X1  g0979(.A1(new_n759), .A2(new_n284), .B1(new_n752), .B2(new_n242), .ZN(new_n1180));
  AOI211_X1 g0980(.A(new_n1175), .B(new_n1180), .C1(G283), .C2(new_n756), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1179), .B(new_n1181), .C1(new_n247), .C2(new_n779), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1176), .B1(new_n1183), .B2(KEYINPUT58), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n769), .A2(new_n308), .ZN(new_n1185));
  OAI22_X1  g0985(.A1(new_n771), .A2(new_n1130), .B1(new_n752), .B2(new_n839), .ZN(new_n1186));
  AOI211_X1 g0986(.A(new_n1185), .B(new_n1186), .C1(G132), .C2(new_n762), .ZN(new_n1187));
  INV_X1    g0987(.A(G128), .ZN(new_n1188));
  OAI22_X1  g0988(.A1(new_n779), .A2(new_n1124), .B1(new_n1188), .B2(new_n759), .ZN(new_n1189));
  AND2_X1   g0989(.A1(new_n1189), .A2(KEYINPUT116), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n1189), .A2(KEYINPUT116), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1187), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  OR2_X1    g0992(.A1(new_n1192), .A2(KEYINPUT59), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT117), .ZN(new_n1194));
  OR2_X1    g0994(.A1(new_n1194), .A2(G124), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(G124), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n756), .A2(new_n1195), .A3(new_n1196), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(G33), .A2(G41), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n1197), .B(new_n1198), .C1(new_n790), .C2(new_n765), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1199), .B1(new_n1192), .B2(KEYINPUT59), .ZN(new_n1200));
  AND2_X1   g1000(.A1(new_n1193), .A2(new_n1200), .ZN(new_n1201));
  AOI211_X1 g1001(.A(new_n1184), .B(new_n1201), .C1(KEYINPUT58), .C2(new_n1183), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n1202), .A2(new_n749), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(new_n1203), .B(KEYINPUT118), .ZN(new_n1204));
  AOI211_X1 g1004(.A(new_n744), .B(new_n693), .C1(new_n324), .C2(new_n823), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n1204), .B(new_n1205), .C1(new_n1148), .C2(new_n804), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1207), .B1(new_n1208), .B2(new_n744), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1174), .A2(new_n1209), .ZN(G375));
  NAND2_X1  g1010(.A1(new_n910), .A2(new_n803), .ZN(new_n1211));
  OAI22_X1  g1011(.A1(new_n763), .A2(new_n1124), .B1(new_n835), .B2(new_n771), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1178), .B1(new_n324), .B2(new_n769), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n282), .B1(new_n752), .B2(new_n308), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n759), .A2(new_n839), .B1(new_n755), .B2(new_n1188), .ZN(new_n1215));
  NOR4_X1   g1015(.A1(new_n1212), .A2(new_n1213), .A3(new_n1214), .A4(new_n1215), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1216), .B1(new_n781), .B2(new_n790), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(new_n780), .A2(G97), .B1(G303), .B2(new_n756), .ZN(new_n1218));
  XNOR2_X1  g1018(.A(new_n1218), .B(KEYINPUT122), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n763), .A2(new_n437), .B1(new_n771), .B2(new_n770), .ZN(new_n1220));
  OAI221_X1 g1020(.A(new_n378), .B1(new_n752), .B2(new_n284), .C1(new_n766), .C2(new_n759), .ZN(new_n1221));
  OAI22_X1  g1021(.A1(new_n769), .A2(new_n242), .B1(new_n765), .B2(new_n247), .ZN(new_n1222));
  OR3_X1    g1022(.A1(new_n1220), .A2(new_n1221), .A3(new_n1222), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1217), .B1(new_n1219), .B2(new_n1223), .ZN(new_n1224));
  AND2_X1   g1024(.A1(new_n1224), .A2(new_n748), .ZN(new_n1225));
  AOI211_X1 g1025(.A(new_n802), .B(new_n1225), .C1(new_n328), .C2(new_n823), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n1093), .A2(new_n744), .B1(new_n1211), .B2(new_n1226), .ZN(new_n1227));
  XNOR2_X1  g1027(.A(new_n955), .B(KEYINPUT121), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1096), .A2(new_n1228), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1227), .B1(new_n1229), .B2(new_n1230), .ZN(G381));
  INV_X1    g1031(.A(G396), .ZN(new_n1232));
  OAI211_X1 g1032(.A(new_n1036), .B(new_n1232), .C1(new_n1038), .C2(new_n1039), .ZN(new_n1233));
  NOR4_X1   g1033(.A1(G390), .A2(G384), .A3(G381), .A4(new_n1233), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(G387), .A2(G378), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1234), .A2(new_n1174), .A3(new_n1209), .A4(new_n1235), .ZN(G407));
  INV_X1    g1036(.A(G378), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n668), .A2(new_n664), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  OAI211_X1 g1039(.A(G407), .B(G213), .C1(G375), .C2(new_n1239), .ZN(new_n1240));
  XOR2_X1   g1040(.A(new_n1240), .B(KEYINPUT123), .Z(G409));
  INV_X1    g1041(.A(KEYINPUT126), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(G393), .A2(G396), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1243), .A2(new_n1233), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(G387), .A2(G390), .ZN(new_n1245));
  NAND4_X1  g1045(.A1(new_n971), .A2(new_n1069), .A3(new_n1003), .A4(new_n1071), .ZN(new_n1246));
  AOI211_X1 g1046(.A(KEYINPUT125), .B(new_n1244), .C1(new_n1245), .C2(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT125), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1243), .A2(new_n1248), .A3(new_n1233), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1244), .A2(KEYINPUT125), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1245), .A2(new_n1249), .A3(new_n1246), .A4(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1251), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1242), .B1(new_n1247), .B2(new_n1252), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1245), .A2(new_n1246), .A3(new_n1250), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1249), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1256), .A2(KEYINPUT126), .A3(new_n1251), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1253), .A2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT61), .ZN(new_n1259));
  AND2_X1   g1059(.A1(new_n1096), .A2(KEYINPUT60), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(new_n1230), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(new_n693), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1260), .A2(new_n1230), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1227), .B1(new_n1262), .B2(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(G384), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  OAI211_X1 g1066(.A(G384), .B(new_n1227), .C1(new_n1262), .C2(new_n1263), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1238), .A2(G2897), .ZN(new_n1268));
  AND3_X1   g1068(.A1(new_n1266), .A2(new_n1267), .A3(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1268), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1172), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1207), .B1(new_n1272), .B2(new_n1228), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n744), .B1(new_n1161), .B2(new_n1163), .ZN(new_n1274));
  AOI21_X1  g1074(.A(G378), .B1(new_n1273), .B2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1169), .A2(KEYINPUT57), .ZN(new_n1276));
  OAI21_X1  g1076(.A(KEYINPUT119), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1276), .B1(new_n1162), .B2(new_n1277), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1173), .B1(new_n1278), .B2(new_n1166), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1167), .ZN(new_n1280));
  OAI211_X1 g1080(.A(G378), .B(new_n1209), .C1(new_n1279), .C2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(KEYINPUT124), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT124), .ZN(new_n1283));
  NAND4_X1  g1083(.A1(new_n1174), .A2(new_n1283), .A3(G378), .A4(new_n1209), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1275), .B1(new_n1282), .B2(new_n1284), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1271), .B1(new_n1285), .B2(new_n1238), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1287));
  NOR3_X1   g1087(.A1(new_n1285), .A2(new_n1238), .A3(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT62), .ZN(new_n1289));
  OAI211_X1 g1089(.A(new_n1259), .B(new_n1286), .C1(new_n1288), .C2(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1282), .A2(new_n1284), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1275), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1238), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1287), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1293), .A2(new_n1294), .A3(new_n1295), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n1296), .A2(KEYINPUT62), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1258), .B1(new_n1290), .B2(new_n1297), .ZN(new_n1298));
  AND2_X1   g1098(.A1(new_n1286), .A2(new_n1259), .ZN(new_n1299));
  NOR2_X1   g1099(.A1(new_n1247), .A2(new_n1252), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT63), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1296), .A2(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1288), .A2(KEYINPUT63), .ZN(new_n1303));
  NAND4_X1  g1103(.A1(new_n1299), .A2(new_n1300), .A3(new_n1302), .A4(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1298), .A2(new_n1304), .ZN(G405));
  NAND2_X1  g1105(.A1(G375), .A2(new_n1237), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1291), .A2(new_n1306), .ZN(new_n1307));
  XNOR2_X1  g1107(.A(new_n1307), .B(new_n1295), .ZN(new_n1308));
  XNOR2_X1  g1108(.A(new_n1258), .B(new_n1308), .ZN(G402));
endmodule


