//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 1 1 0 1 0 0 0 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 1 1 1 0 0 1 0 0 1 0 1 1 0 0 1 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n806, new_n807, new_n808, new_n809, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n828,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n847, new_n848, new_n849, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n896, new_n897,
    new_n899, new_n900, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n979,
    new_n980, new_n981, new_n982, new_n984, new_n985, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n996,
    new_n997, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1020, new_n1021, new_n1022, new_n1023, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1030, new_n1031;
  INV_X1    g000(.A(KEYINPUT92), .ZN(new_n202));
  INV_X1    g001(.A(G29gat), .ZN(new_n203));
  INV_X1    g002(.A(G36gat), .ZN(new_n204));
  NAND3_X1  g003(.A1(new_n203), .A2(new_n204), .A3(KEYINPUT91), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT91), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n206), .B1(G29gat), .B2(G36gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n205), .A2(new_n207), .A3(KEYINPUT14), .ZN(new_n208));
  NAND2_X1  g007(.A1(G29gat), .A2(G36gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT14), .ZN(new_n210));
  OAI211_X1 g009(.A(new_n206), .B(new_n210), .C1(G29gat), .C2(G36gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n208), .A2(new_n209), .A3(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G43gat), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n213), .A2(G50gat), .ZN(new_n214));
  INV_X1    g013(.A(G50gat), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n215), .A2(G43gat), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  AND3_X1   g016(.A1(new_n212), .A2(KEYINPUT15), .A3(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT15), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n219), .B1(new_n214), .B2(new_n216), .ZN(new_n220));
  NAND4_X1  g019(.A1(new_n220), .A2(new_n208), .A3(new_n209), .A4(new_n211), .ZN(new_n221));
  NOR3_X1   g020(.A1(new_n214), .A2(new_n216), .A3(new_n219), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n202), .B1(new_n218), .B2(new_n223), .ZN(new_n224));
  AND2_X1   g023(.A1(new_n208), .A2(new_n211), .ZN(new_n225));
  INV_X1    g024(.A(new_n222), .ZN(new_n226));
  NAND4_X1  g025(.A1(new_n225), .A2(new_n226), .A3(new_n220), .A4(new_n209), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n221), .A2(new_n222), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n227), .A2(new_n228), .A3(KEYINPUT92), .ZN(new_n229));
  XNOR2_X1  g028(.A(KEYINPUT93), .B(KEYINPUT17), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n224), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  XNOR2_X1  g030(.A(G15gat), .B(G22gat), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT16), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n232), .B1(new_n233), .B2(G1gat), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n234), .B1(G1gat), .B2(new_n232), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(G8gat), .ZN(new_n236));
  INV_X1    g035(.A(G8gat), .ZN(new_n237));
  OAI211_X1 g036(.A(new_n234), .B(new_n237), .C1(G1gat), .C2(new_n232), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n218), .A2(new_n223), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n239), .B1(new_n240), .B2(KEYINPUT17), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n231), .A2(new_n241), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n224), .A2(new_n229), .A3(new_n239), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT18), .ZN(new_n244));
  AOI22_X1  g043(.A1(new_n244), .A2(KEYINPUT95), .B1(G229gat), .B2(G233gat), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n242), .A2(new_n243), .A3(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT94), .ZN(new_n247));
  AOI21_X1  g046(.A(KEYINPUT95), .B1(new_n247), .B2(new_n244), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n246), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(G229gat), .A2(G233gat), .ZN(new_n251));
  XOR2_X1   g050(.A(new_n251), .B(KEYINPUT13), .Z(new_n252));
  INV_X1    g051(.A(new_n243), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n239), .B1(new_n224), .B2(new_n229), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n252), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NAND4_X1  g054(.A1(new_n242), .A2(new_n243), .A3(new_n248), .A4(new_n245), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n250), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(G113gat), .B(G141gat), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n258), .B(KEYINPUT90), .ZN(new_n259));
  XOR2_X1   g058(.A(KEYINPUT89), .B(KEYINPUT11), .Z(new_n260));
  XNOR2_X1  g059(.A(new_n259), .B(new_n260), .ZN(new_n261));
  XOR2_X1   g060(.A(G169gat), .B(G197gat), .Z(new_n262));
  XNOR2_X1  g061(.A(new_n261), .B(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(new_n263), .B(KEYINPUT12), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n257), .A2(new_n265), .ZN(new_n266));
  NAND4_X1  g065(.A1(new_n264), .A2(new_n255), .A3(new_n256), .A4(new_n250), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n239), .ZN(new_n269));
  XNOR2_X1  g068(.A(G57gat), .B(G64gat), .ZN(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(G71gat), .A2(G78gat), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT9), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  OR2_X1    g073(.A1(G71gat), .A2(G78gat), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(new_n272), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n271), .A2(new_n274), .A3(new_n276), .ZN(new_n277));
  OAI211_X1 g076(.A(new_n272), .B(new_n275), .C1(new_n270), .C2(new_n273), .ZN(new_n278));
  AND2_X1   g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(KEYINPUT21), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n269), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(G183gat), .ZN(new_n282));
  INV_X1    g081(.A(G183gat), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n269), .A2(new_n283), .A3(new_n280), .ZN(new_n284));
  INV_X1    g083(.A(G231gat), .ZN(new_n285));
  INV_X1    g084(.A(G233gat), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n282), .A2(new_n284), .A3(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n288), .B1(new_n282), .B2(new_n284), .ZN(new_n291));
  XNOR2_X1  g090(.A(KEYINPUT96), .B(KEYINPUT21), .ZN(new_n292));
  OAI22_X1  g091(.A1(new_n290), .A2(new_n291), .B1(new_n279), .B2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n291), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n279), .A2(new_n292), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n294), .A2(new_n295), .A3(new_n289), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n293), .A2(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(G127gat), .B(G155gat), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n298), .B(G211gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(new_n299), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n293), .A2(new_n296), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  XNOR2_X1  g102(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n300), .A2(new_n304), .A3(new_n302), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  XOR2_X1   g107(.A(G190gat), .B(G218gat), .Z(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(G232gat), .A2(G233gat), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT41), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n224), .A2(new_n229), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT98), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT7), .ZN(new_n317));
  INV_X1    g116(.A(G85gat), .ZN(new_n318));
  INV_X1    g117(.A(G92gat), .ZN(new_n319));
  OAI221_X1 g118(.A(KEYINPUT99), .B1(new_n316), .B2(new_n317), .C1(new_n318), .C2(new_n319), .ZN(new_n320));
  OR2_X1    g119(.A1(new_n317), .A2(KEYINPUT99), .ZN(new_n321));
  OAI21_X1  g120(.A(KEYINPUT99), .B1(new_n316), .B2(new_n317), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n318), .A2(new_n319), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n321), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(G99gat), .A2(G106gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(KEYINPUT8), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n318), .A2(new_n319), .ZN(new_n327));
  AND3_X1   g126(.A1(new_n326), .A2(KEYINPUT100), .A3(new_n327), .ZN(new_n328));
  AOI21_X1  g127(.A(KEYINPUT100), .B1(new_n326), .B2(new_n327), .ZN(new_n329));
  OAI211_X1 g128(.A(new_n320), .B(new_n324), .C1(new_n328), .C2(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(G99gat), .B(G106gat), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT100), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT8), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n335), .B1(G99gat), .B2(G106gat), .ZN(new_n336));
  NOR2_X1   g135(.A1(G85gat), .A2(G92gat), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n334), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n326), .A2(KEYINPUT100), .A3(new_n327), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND4_X1  g139(.A1(new_n340), .A2(new_n331), .A3(new_n320), .A4(new_n324), .ZN(new_n341));
  AND3_X1   g140(.A1(new_n333), .A2(new_n341), .A3(KEYINPUT101), .ZN(new_n342));
  AOI21_X1  g141(.A(KEYINPUT101), .B1(new_n333), .B2(new_n341), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n313), .B1(new_n315), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n333), .A2(new_n341), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT101), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n333), .A2(new_n341), .A3(KEYINPUT101), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n240), .A2(KEYINPUT17), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n350), .A2(new_n231), .A3(new_n351), .ZN(new_n352));
  AND3_X1   g151(.A1(new_n345), .A2(KEYINPUT102), .A3(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(KEYINPUT102), .B1(new_n345), .B2(new_n352), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n310), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT102), .ZN(new_n356));
  INV_X1    g155(.A(new_n352), .ZN(new_n357));
  OAI22_X1  g156(.A1(new_n350), .A2(new_n314), .B1(new_n312), .B2(new_n311), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n356), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n345), .A2(KEYINPUT102), .A3(new_n352), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n359), .A2(new_n309), .A3(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n355), .A2(KEYINPUT97), .A3(new_n361), .ZN(new_n362));
  XNOR2_X1  g161(.A(G134gat), .B(G162gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n311), .A2(new_n312), .ZN(new_n364));
  XOR2_X1   g163(.A(new_n363), .B(new_n364), .Z(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n362), .A2(new_n366), .ZN(new_n367));
  NAND4_X1  g166(.A1(new_n355), .A2(new_n361), .A3(KEYINPUT97), .A4(new_n365), .ZN(new_n368));
  AND2_X1   g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(G230gat), .A2(G233gat), .ZN(new_n370));
  OR2_X1    g169(.A1(new_n331), .A2(KEYINPUT103), .ZN(new_n371));
  AND3_X1   g170(.A1(new_n277), .A2(new_n278), .A3(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n333), .A2(new_n372), .A3(new_n341), .ZN(new_n373));
  INV_X1    g172(.A(new_n373), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n372), .B1(new_n333), .B2(new_n341), .ZN(new_n375));
  NOR3_X1   g174(.A1(new_n374), .A2(new_n375), .A3(KEYINPUT10), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n279), .A2(KEYINPUT10), .ZN(new_n377));
  NOR3_X1   g176(.A1(new_n342), .A2(new_n343), .A3(new_n377), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n370), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n372), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n346), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n370), .B1(new_n381), .B2(new_n373), .ZN(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  XNOR2_X1  g182(.A(G120gat), .B(G148gat), .ZN(new_n384));
  XNOR2_X1  g183(.A(G176gat), .B(G204gat), .ZN(new_n385));
  XNOR2_X1  g184(.A(new_n384), .B(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n379), .A2(new_n383), .A3(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(new_n370), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT10), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n381), .A2(new_n390), .A3(new_n373), .ZN(new_n391));
  INV_X1    g190(.A(new_n377), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n348), .A2(new_n392), .A3(new_n349), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n389), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n386), .B1(new_n394), .B2(new_n382), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n388), .A2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT104), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n388), .A2(new_n395), .A3(KEYINPUT104), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  NOR3_X1   g200(.A1(new_n308), .A2(new_n369), .A3(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT36), .ZN(new_n403));
  INV_X1    g202(.A(G127gat), .ZN(new_n404));
  INV_X1    g203(.A(G134gat), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(KEYINPUT69), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT69), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(G134gat), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n404), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n405), .A2(G127gat), .ZN(new_n410));
  OAI21_X1  g209(.A(KEYINPUT70), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT70), .ZN(new_n412));
  INV_X1    g211(.A(new_n410), .ZN(new_n413));
  XNOR2_X1  g212(.A(KEYINPUT69), .B(G134gat), .ZN(new_n414));
  OAI211_X1 g213(.A(new_n412), .B(new_n413), .C1(new_n414), .C2(new_n404), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n411), .A2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT1), .ZN(new_n417));
  INV_X1    g216(.A(G113gat), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n418), .A2(G120gat), .ZN(new_n419));
  INV_X1    g218(.A(G120gat), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n420), .A2(G113gat), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n417), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n416), .A2(new_n422), .ZN(new_n423));
  OAI21_X1  g222(.A(KEYINPUT71), .B1(new_n418), .B2(G120gat), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT71), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n425), .A2(new_n420), .A3(G113gat), .ZN(new_n426));
  OAI211_X1 g225(.A(new_n424), .B(new_n426), .C1(G113gat), .C2(new_n420), .ZN(new_n427));
  AND2_X1   g226(.A1(new_n427), .A2(new_n417), .ZN(new_n428));
  XNOR2_X1  g227(.A(G127gat), .B(G134gat), .ZN(new_n429));
  XNOR2_X1  g228(.A(new_n429), .B(KEYINPUT72), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n423), .A2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT25), .ZN(new_n433));
  NAND3_X1  g232(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT66), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND4_X1  g235(.A1(KEYINPUT66), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NOR2_X1   g237(.A1(G183gat), .A2(G190gat), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT24), .ZN(new_n440));
  NAND2_X1  g239(.A1(G183gat), .A2(G190gat), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n439), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  AND3_X1   g241(.A1(new_n438), .A2(KEYINPUT67), .A3(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(KEYINPUT67), .B1(new_n438), .B2(new_n442), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(G169gat), .A2(G176gat), .ZN(new_n446));
  NOR2_X1   g245(.A1(G169gat), .A2(G176gat), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n446), .B1(new_n447), .B2(KEYINPUT23), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT65), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  OAI21_X1  g249(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n448), .B1(new_n452), .B2(KEYINPUT23), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n433), .B1(new_n445), .B2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT64), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n434), .A2(new_n455), .ZN(new_n456));
  NAND4_X1  g255(.A1(KEYINPUT64), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n448), .B1(new_n458), .B2(new_n442), .ZN(new_n459));
  INV_X1    g258(.A(G169gat), .ZN(new_n460));
  INV_X1    g259(.A(G176gat), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n460), .A2(new_n461), .A3(KEYINPUT23), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n459), .A2(new_n433), .A3(new_n462), .ZN(new_n463));
  OAI21_X1  g262(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(new_n446), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT68), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n464), .A2(KEYINPUT68), .A3(new_n446), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(KEYINPUT26), .B1(new_n450), .B2(new_n451), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n441), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  XNOR2_X1  g270(.A(KEYINPUT27), .B(G183gat), .ZN(new_n472));
  INV_X1    g271(.A(G190gat), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(KEYINPUT28), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT28), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n472), .A2(new_n476), .A3(new_n473), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n463), .B1(new_n471), .B2(new_n478), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n432), .B1(new_n454), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n462), .A2(new_n433), .ZN(new_n481));
  AOI211_X1 g280(.A(new_n448), .B(new_n481), .C1(new_n442), .C2(new_n458), .ZN(new_n482));
  AND3_X1   g281(.A1(new_n464), .A2(KEYINPUT68), .A3(new_n446), .ZN(new_n483));
  AOI21_X1  g282(.A(KEYINPUT68), .B1(new_n464), .B2(new_n446), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(new_n470), .ZN(new_n486));
  AOI22_X1  g285(.A1(new_n485), .A2(new_n486), .B1(G183gat), .B2(G190gat), .ZN(new_n487));
  AND2_X1   g286(.A1(new_n475), .A2(new_n477), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n482), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n438), .A2(new_n442), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT67), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n438), .A2(KEYINPUT67), .A3(new_n442), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n492), .A2(new_n453), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(KEYINPUT25), .ZN(new_n495));
  AOI22_X1  g294(.A1(new_n416), .A2(new_n422), .B1(new_n428), .B2(new_n430), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n489), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n480), .A2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(G227gat), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n499), .A2(new_n286), .ZN(new_n500));
  AOI21_X1  g299(.A(KEYINPUT73), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT73), .ZN(new_n502));
  INV_X1    g301(.A(new_n500), .ZN(new_n503));
  AOI211_X1 g302(.A(new_n502), .B(new_n503), .C1(new_n480), .C2(new_n497), .ZN(new_n504));
  OAI21_X1  g303(.A(KEYINPUT32), .B1(new_n501), .B2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT33), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n506), .B1(new_n501), .B2(new_n504), .ZN(new_n507));
  XNOR2_X1  g306(.A(G15gat), .B(G43gat), .ZN(new_n508));
  XNOR2_X1  g307(.A(G71gat), .B(G99gat), .ZN(new_n509));
  XOR2_X1   g308(.A(new_n508), .B(new_n509), .Z(new_n510));
  NAND3_X1  g309(.A1(new_n505), .A2(new_n507), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(KEYINPUT74), .ZN(new_n512));
  AND2_X1   g311(.A1(new_n510), .A2(KEYINPUT33), .ZN(new_n513));
  OR2_X1    g312(.A1(new_n505), .A2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT74), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n505), .A2(new_n507), .A3(new_n515), .A4(new_n510), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n512), .A2(new_n514), .A3(new_n516), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n480), .A2(new_n503), .A3(new_n497), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n518), .B(KEYINPUT34), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(new_n519), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n512), .A2(new_n521), .A3(new_n514), .A4(new_n516), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n403), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT75), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n520), .A2(new_n524), .A3(new_n522), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n517), .A2(KEYINPUT75), .A3(new_n519), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n523), .B1(new_n527), .B2(new_n403), .ZN(new_n528));
  XNOR2_X1  g327(.A(G78gat), .B(G106gat), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n529), .B(new_n215), .ZN(new_n530));
  XNOR2_X1  g329(.A(KEYINPUT82), .B(KEYINPUT31), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n530), .B(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(G22gat), .ZN(new_n533));
  INV_X1    g332(.A(G228gat), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n534), .A2(new_n286), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT80), .ZN(new_n536));
  XOR2_X1   g335(.A(G141gat), .B(G148gat), .Z(new_n537));
  INV_X1    g336(.A(G155gat), .ZN(new_n538));
  INV_X1    g337(.A(G162gat), .ZN(new_n539));
  OAI21_X1  g338(.A(KEYINPUT2), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n537), .A2(new_n540), .ZN(new_n541));
  XNOR2_X1  g340(.A(G155gat), .B(G162gat), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n537), .A2(new_n540), .A3(new_n542), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n536), .B1(new_n546), .B2(KEYINPUT3), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT3), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n544), .A2(KEYINPUT80), .A3(new_n548), .A4(new_n545), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT29), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(G197gat), .B(G204gat), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT22), .ZN(new_n554));
  INV_X1    g353(.A(G211gat), .ZN(new_n555));
  INV_X1    g354(.A(G218gat), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n554), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n553), .A2(new_n557), .ZN(new_n558));
  XOR2_X1   g357(.A(G211gat), .B(G218gat), .Z(new_n559));
  XOR2_X1   g358(.A(new_n558), .B(new_n559), .Z(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(KEYINPUT76), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT76), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n558), .A2(new_n562), .A3(new_n559), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n552), .A2(new_n564), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n548), .B1(new_n560), .B2(KEYINPUT29), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(new_n546), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n535), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n561), .A2(new_n551), .A3(new_n563), .ZN(new_n570));
  AND2_X1   g369(.A1(new_n570), .A2(new_n548), .ZN(new_n571));
  INV_X1    g370(.A(new_n546), .ZN(new_n572));
  OAI211_X1 g371(.A(new_n535), .B(new_n565), .C1(new_n571), .C2(new_n572), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n533), .B1(new_n569), .B2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT83), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n532), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n565), .ZN(new_n577));
  INV_X1    g376(.A(new_n535), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n572), .B1(new_n570), .B2(new_n548), .ZN(new_n579));
  NOR3_X1   g378(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  OAI21_X1  g379(.A(G22gat), .B1(new_n580), .B2(new_n568), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n569), .A2(new_n573), .A3(new_n533), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n581), .A2(KEYINPUT83), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n576), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n581), .A2(new_n532), .A3(new_n582), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT84), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND4_X1  g386(.A1(new_n581), .A2(KEYINPUT84), .A3(new_n532), .A4(new_n582), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n584), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n546), .A2(KEYINPUT3), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n550), .A2(new_n432), .A3(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT4), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n592), .B1(new_n432), .B2(new_n546), .ZN(new_n593));
  NAND2_X1  g392(.A1(G225gat), .A2(G233gat), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n496), .A2(KEYINPUT4), .A3(new_n572), .ZN(new_n595));
  NAND4_X1  g394(.A1(new_n591), .A2(new_n593), .A3(new_n594), .A4(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n596), .A2(KEYINPUT81), .ZN(new_n597));
  INV_X1    g396(.A(new_n594), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n432), .A2(new_n546), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n496), .A2(new_n572), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n598), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(KEYINPUT5), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n597), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n602), .A2(new_n596), .A3(KEYINPUT81), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(G1gat), .B(G29gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(G85gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(KEYINPUT0), .B(G57gat), .ZN(new_n609));
  XOR2_X1   g408(.A(new_n608), .B(new_n609), .Z(new_n610));
  AOI21_X1  g409(.A(KEYINPUT6), .B1(new_n606), .B2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n610), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n604), .A2(new_n605), .A3(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n611), .B(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(G226gat), .A2(G233gat), .ZN(new_n615));
  OAI211_X1 g414(.A(new_n551), .B(new_n615), .C1(new_n454), .C2(new_n479), .ZN(new_n616));
  NAND4_X1  g415(.A1(new_n489), .A2(new_n495), .A3(G226gat), .A4(G233gat), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n564), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n616), .A2(new_n564), .A3(new_n617), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(KEYINPUT78), .B(G92gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(KEYINPUT77), .B(G64gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n624), .B(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(G8gat), .B(G36gat), .ZN(new_n627));
  XOR2_X1   g426(.A(new_n626), .B(new_n627), .Z(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n623), .A2(KEYINPUT79), .A3(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT30), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT79), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n632), .B1(new_n622), .B2(new_n628), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n630), .A2(new_n631), .A3(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n623), .A2(KEYINPUT30), .A3(new_n629), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n622), .A2(new_n628), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n634), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n589), .B1(new_n614), .B2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  AOI21_X1  g439(.A(KEYINPUT85), .B1(new_n528), .B2(new_n640), .ZN(new_n641));
  AOI21_X1  g440(.A(KEYINPUT36), .B1(new_n525), .B2(new_n526), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT85), .ZN(new_n643));
  NOR4_X1   g442(.A1(new_n642), .A2(new_n643), .A3(new_n639), .A4(new_n523), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT38), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n629), .B1(new_n622), .B2(KEYINPUT37), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  OR2_X1    g446(.A1(new_n647), .A2(KEYINPUT88), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n622), .A2(KEYINPUT37), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n649), .B1(new_n647), .B2(KEYINPUT88), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n645), .B1(new_n648), .B2(new_n650), .ZN(new_n651));
  XOR2_X1   g450(.A(new_n610), .B(KEYINPUT86), .Z(new_n652));
  NAND3_X1  g451(.A1(new_n604), .A2(new_n605), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n611), .A2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT6), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n613), .A2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  AND2_X1   g456(.A1(new_n630), .A2(new_n633), .ZN(new_n658));
  OAI211_X1 g457(.A(new_n646), .B(new_n645), .C1(KEYINPUT37), .C2(new_n622), .ZN(new_n659));
  NAND4_X1  g458(.A1(new_n654), .A2(new_n657), .A3(new_n658), .A4(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT87), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n656), .B1(new_n611), .B2(new_n653), .ZN(new_n663));
  NAND4_X1  g462(.A1(new_n663), .A2(KEYINPUT87), .A3(new_n658), .A4(new_n659), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n651), .B1(new_n662), .B2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n589), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n591), .A2(new_n593), .A3(new_n595), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT39), .ZN(new_n668));
  AND2_X1   g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n667), .A2(new_n668), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n598), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n652), .ZN(new_n672));
  OAI211_X1 g471(.A(KEYINPUT39), .B(new_n594), .C1(new_n599), .C2(new_n600), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n671), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT40), .ZN(new_n675));
  OR2_X1    g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n674), .A2(new_n675), .ZN(new_n677));
  NAND4_X1  g476(.A1(new_n676), .A2(new_n637), .A3(new_n653), .A4(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  NOR3_X1   g478(.A1(new_n665), .A2(new_n666), .A3(new_n679), .ZN(new_n680));
  NOR3_X1   g479(.A1(new_n641), .A2(new_n644), .A3(new_n680), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n614), .A2(KEYINPUT35), .A3(new_n638), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n589), .A2(new_n520), .A3(new_n522), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n663), .A2(new_n637), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n527), .A2(new_n589), .A3(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT35), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n684), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  OAI211_X1 g488(.A(new_n268), .B(new_n402), .C1(new_n681), .C2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n690), .A2(KEYINPUT105), .ZN(new_n691));
  AND2_X1   g490(.A1(new_n266), .A2(new_n267), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n527), .A2(new_n403), .ZN(new_n693));
  INV_X1    g492(.A(new_n523), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n693), .A2(new_n640), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(new_n643), .ZN(new_n696));
  AND2_X1   g495(.A1(new_n662), .A2(new_n664), .ZN(new_n697));
  OAI211_X1 g496(.A(new_n678), .B(new_n589), .C1(new_n697), .C2(new_n651), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n528), .A2(KEYINPUT85), .A3(new_n640), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n696), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n692), .B1(new_n700), .B2(new_n688), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT105), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n701), .A2(new_n702), .A3(new_n402), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n691), .A2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n614), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n706), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g506(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n233), .A2(new_n237), .ZN(new_n709));
  NAND4_X1  g508(.A1(new_n704), .A2(new_n637), .A3(new_n708), .A4(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT42), .ZN(new_n711));
  OR2_X1    g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  AND2_X1   g511(.A1(new_n691), .A2(new_n703), .ZN(new_n713));
  OAI21_X1  g512(.A(G8gat), .B1(new_n713), .B2(new_n638), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n710), .A2(new_n711), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n712), .A2(new_n714), .A3(new_n715), .ZN(G1325gat));
  AOI21_X1  g515(.A(G15gat), .B1(new_n704), .B2(new_n527), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT106), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n528), .A2(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(KEYINPUT106), .B1(new_n642), .B2(new_n523), .ZN(new_n720));
  AND2_X1   g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n713), .A2(new_n721), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n717), .B1(new_n722), .B2(G15gat), .ZN(G1326gat));
  XNOR2_X1  g522(.A(KEYINPUT43), .B(G22gat), .ZN(new_n724));
  OAI21_X1  g523(.A(KEYINPUT107), .B1(new_n713), .B2(new_n589), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT107), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n704), .A2(new_n726), .A3(new_n666), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n724), .B1(new_n725), .B2(new_n727), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n726), .B1(new_n704), .B2(new_n666), .ZN(new_n729));
  AOI211_X1 g528(.A(KEYINPUT107), .B(new_n589), .C1(new_n691), .C2(new_n703), .ZN(new_n730));
  INV_X1    g529(.A(new_n724), .ZN(new_n731));
  NOR3_X1   g530(.A1(new_n729), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n728), .A2(new_n732), .ZN(G1327gat));
  NAND4_X1  g532(.A1(new_n719), .A2(new_n698), .A3(new_n640), .A4(new_n720), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT109), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n688), .A2(new_n735), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n666), .B1(new_n525), .B2(new_n526), .ZN(new_n737));
  AOI21_X1  g536(.A(KEYINPUT35), .B1(new_n737), .B2(new_n685), .ZN(new_n738));
  NOR3_X1   g537(.A1(new_n738), .A2(KEYINPUT109), .A3(new_n684), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n734), .B1(new_n736), .B2(new_n739), .ZN(new_n740));
  AOI21_X1  g539(.A(KEYINPUT44), .B1(new_n740), .B2(new_n369), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n367), .A2(new_n368), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n742), .B1(new_n700), .B2(new_n688), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n741), .B1(KEYINPUT44), .B2(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(new_n308), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n746), .A2(new_n401), .ZN(new_n747));
  INV_X1    g546(.A(new_n747), .ZN(new_n748));
  AND3_X1   g547(.A1(new_n266), .A2(KEYINPUT108), .A3(new_n267), .ZN(new_n749));
  AOI21_X1  g548(.A(KEYINPUT108), .B1(new_n266), .B2(new_n267), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n748), .A2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(new_n753), .ZN(new_n754));
  NOR3_X1   g553(.A1(new_n745), .A2(new_n614), .A3(new_n754), .ZN(new_n755));
  OAI211_X1 g554(.A(new_n268), .B(new_n747), .C1(new_n681), .C2(new_n689), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n756), .A2(new_n742), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n757), .A2(new_n203), .A3(new_n705), .ZN(new_n758));
  AND2_X1   g557(.A1(new_n758), .A2(KEYINPUT45), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n758), .A2(KEYINPUT45), .ZN(new_n760));
  OAI22_X1  g559(.A1(new_n755), .A2(new_n203), .B1(new_n759), .B2(new_n760), .ZN(G1328gat));
  NOR4_X1   g560(.A1(new_n756), .A2(G36gat), .A3(new_n638), .A4(new_n742), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT46), .ZN(new_n763));
  OR2_X1    g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n762), .A2(new_n763), .ZN(new_n765));
  NOR3_X1   g564(.A1(new_n745), .A2(new_n638), .A3(new_n754), .ZN(new_n766));
  OAI211_X1 g565(.A(new_n764), .B(new_n765), .C1(new_n766), .C2(new_n204), .ZN(G1329gat));
  INV_X1    g566(.A(KEYINPUT110), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n757), .A2(new_n768), .A3(new_n213), .A4(new_n527), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n701), .A2(new_n213), .A3(new_n369), .A4(new_n747), .ZN(new_n770));
  INV_X1    g569(.A(new_n527), .ZN(new_n771));
  OAI21_X1  g570(.A(KEYINPUT110), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  AND2_X1   g571(.A1(new_n769), .A2(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT44), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n680), .A2(new_n639), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n686), .A2(new_n687), .ZN(new_n776));
  INV_X1    g575(.A(new_n684), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n776), .A2(new_n735), .A3(new_n777), .ZN(new_n778));
  OAI21_X1  g577(.A(KEYINPUT109), .B1(new_n738), .B2(new_n684), .ZN(new_n779));
  AOI22_X1  g578(.A1(new_n721), .A2(new_n775), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n774), .B1(new_n780), .B2(new_n742), .ZN(new_n781));
  INV_X1    g580(.A(new_n721), .ZN(new_n782));
  OAI211_X1 g581(.A(KEYINPUT44), .B(new_n369), .C1(new_n681), .C2(new_n689), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n781), .A2(new_n782), .A3(new_n753), .A4(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(G43gat), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT111), .ZN(new_n786));
  OAI211_X1 g585(.A(new_n773), .B(new_n785), .C1(new_n786), .C2(KEYINPUT47), .ZN(new_n787));
  AOI21_X1  g586(.A(KEYINPUT47), .B1(new_n785), .B2(new_n786), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n785), .A2(new_n772), .A3(new_n769), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n787), .A2(new_n790), .ZN(G1330gat));
  NOR2_X1   g590(.A1(new_n589), .A2(new_n215), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n781), .A2(new_n753), .A3(new_n783), .A4(new_n792), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n701), .A2(new_n666), .A3(new_n369), .A4(new_n747), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(new_n215), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT48), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n793), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT112), .ZN(new_n798));
  AND2_X1   g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n797), .A2(new_n798), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n793), .A2(new_n795), .ZN(new_n801));
  AOI21_X1  g600(.A(KEYINPUT113), .B1(new_n801), .B2(KEYINPUT48), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT113), .ZN(new_n803));
  AOI211_X1 g602(.A(new_n803), .B(new_n796), .C1(new_n793), .C2(new_n795), .ZN(new_n804));
  OAI22_X1  g603(.A1(new_n799), .A2(new_n800), .B1(new_n802), .B2(new_n804), .ZN(G1331gat));
  NOR2_X1   g604(.A1(new_n308), .A2(new_n369), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n751), .A2(new_n400), .ZN(new_n807));
  AND3_X1   g606(.A1(new_n740), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(new_n705), .ZN(new_n809));
  XNOR2_X1  g608(.A(new_n809), .B(G57gat), .ZN(G1332gat));
  INV_X1    g609(.A(new_n808), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n811), .A2(new_n638), .ZN(new_n812));
  NOR2_X1   g611(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n813));
  AND2_X1   g612(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n812), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n815), .B1(new_n812), .B2(new_n813), .ZN(G1333gat));
  INV_X1    g615(.A(KEYINPUT50), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n740), .A2(new_n527), .A3(new_n806), .A4(new_n807), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT114), .ZN(new_n819));
  XNOR2_X1  g618(.A(new_n818), .B(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(G71gat), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n821), .B1(new_n808), .B2(new_n782), .ZN(new_n823));
  INV_X1    g622(.A(new_n823), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n817), .B1(new_n822), .B2(new_n824), .ZN(new_n825));
  AOI211_X1 g624(.A(KEYINPUT50), .B(new_n823), .C1(new_n820), .C2(new_n821), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n825), .A2(new_n826), .ZN(G1334gat));
  NAND2_X1  g626(.A1(new_n808), .A2(new_n666), .ZN(new_n828));
  XNOR2_X1  g627(.A(new_n828), .B(G78gat), .ZN(G1335gat));
  NAND4_X1  g628(.A1(new_n781), .A2(new_n308), .A3(new_n783), .A4(new_n807), .ZN(new_n830));
  NOR3_X1   g629(.A1(new_n830), .A2(new_n318), .A3(new_n614), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n746), .A2(new_n751), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n740), .A2(new_n369), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(KEYINPUT51), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT51), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n740), .A2(new_n835), .A3(new_n369), .A4(new_n832), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n834), .A2(new_n705), .A3(new_n401), .A4(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n831), .B1(new_n318), .B2(new_n837), .ZN(G1336gat));
  OAI21_X1  g637(.A(G92gat), .B1(new_n830), .B2(new_n638), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n638), .A2(G92gat), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n834), .A2(new_n401), .A3(new_n836), .A4(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(KEYINPUT52), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT52), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n839), .A2(new_n844), .A3(new_n841), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n843), .A2(new_n845), .ZN(G1337gat));
  OAI21_X1  g645(.A(G99gat), .B1(new_n830), .B2(new_n721), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n771), .A2(G99gat), .ZN(new_n848));
  NAND4_X1  g647(.A1(new_n834), .A2(new_n401), .A3(new_n836), .A4(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n847), .A2(new_n849), .ZN(G1338gat));
  NAND4_X1  g649(.A1(new_n834), .A2(new_n666), .A3(new_n401), .A4(new_n836), .ZN(new_n851));
  INV_X1    g650(.A(G106gat), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n589), .A2(new_n852), .ZN(new_n854));
  NAND4_X1  g653(.A1(new_n744), .A2(new_n308), .A3(new_n807), .A4(new_n854), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT53), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n853), .A2(new_n855), .A3(KEYINPUT53), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(G1339gat));
  NAND3_X1  g659(.A1(new_n391), .A2(new_n393), .A3(new_n389), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n379), .A2(KEYINPUT54), .A3(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT54), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n387), .B1(new_n394), .B2(new_n863), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n862), .A2(new_n864), .A3(KEYINPUT55), .ZN(new_n865));
  AND2_X1   g664(.A1(new_n865), .A2(new_n388), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n862), .A2(new_n864), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT55), .ZN(new_n868));
  AOI21_X1  g667(.A(KEYINPUT115), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT115), .ZN(new_n870));
  AOI211_X1 g669(.A(new_n870), .B(KEYINPUT55), .C1(new_n862), .C2(new_n864), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n866), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(KEYINPUT116), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT116), .ZN(new_n874));
  OAI211_X1 g673(.A(new_n866), .B(new_n874), .C1(new_n869), .C2(new_n871), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n873), .A2(new_n751), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n251), .B1(new_n242), .B2(new_n243), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n253), .A2(new_n254), .A3(new_n252), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n263), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND4_X1  g678(.A1(new_n398), .A2(new_n879), .A3(new_n267), .A4(new_n399), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n369), .B1(new_n876), .B2(new_n880), .ZN(new_n881));
  AND2_X1   g680(.A1(new_n267), .A2(new_n879), .ZN(new_n882));
  NAND4_X1  g681(.A1(new_n369), .A2(new_n873), .A3(new_n875), .A4(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(new_n883), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n308), .B1(new_n881), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n402), .A2(new_n752), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n614), .A2(new_n637), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n889), .A2(new_n683), .ZN(new_n890));
  AOI21_X1  g689(.A(G113gat), .B1(new_n890), .B2(new_n751), .ZN(new_n891));
  INV_X1    g690(.A(new_n737), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n889), .A2(new_n892), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n692), .A2(new_n418), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n891), .B1(new_n893), .B2(new_n894), .ZN(G1340gat));
  AOI21_X1  g694(.A(G120gat), .B1(new_n890), .B2(new_n401), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n400), .A2(new_n420), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n896), .B1(new_n893), .B2(new_n897), .ZN(G1341gat));
  NAND3_X1  g697(.A1(new_n890), .A2(new_n404), .A3(new_n746), .ZN(new_n899));
  NOR3_X1   g698(.A1(new_n889), .A2(new_n892), .A3(new_n308), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n899), .B1(new_n404), .B2(new_n900), .ZN(G1342gat));
  INV_X1    g700(.A(new_n414), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n890), .A2(new_n902), .A3(new_n369), .ZN(new_n903));
  OR2_X1    g702(.A1(new_n903), .A2(KEYINPUT56), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(KEYINPUT56), .ZN(new_n905));
  NOR3_X1   g704(.A1(new_n889), .A2(new_n892), .A3(new_n742), .ZN(new_n906));
  OAI211_X1 g705(.A(new_n904), .B(new_n905), .C1(new_n405), .C2(new_n906), .ZN(G1343gat));
  INV_X1    g706(.A(KEYINPUT121), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT118), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n861), .A2(KEYINPUT54), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n910), .A2(new_n394), .ZN(new_n911));
  OAI211_X1 g710(.A(new_n863), .B(new_n370), .C1(new_n376), .C2(new_n378), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(new_n386), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n868), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n914), .A2(new_n388), .A3(new_n865), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n880), .B1(new_n692), .B2(new_n915), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT117), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OAI211_X1 g717(.A(new_n880), .B(KEYINPUT117), .C1(new_n692), .C2(new_n915), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n918), .A2(new_n742), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(new_n883), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n909), .B1(new_n921), .B2(new_n308), .ZN(new_n922));
  AOI211_X1 g721(.A(KEYINPUT118), .B(new_n746), .C1(new_n920), .C2(new_n883), .ZN(new_n923));
  INV_X1    g722(.A(new_n886), .ZN(new_n924));
  NOR3_X1   g723(.A1(new_n922), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT57), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n589), .A2(new_n926), .ZN(new_n927));
  INV_X1    g726(.A(new_n927), .ZN(new_n928));
  OAI21_X1  g727(.A(KEYINPUT119), .B1(new_n925), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n887), .A2(new_n666), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n930), .A2(new_n926), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n921), .A2(new_n308), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(KEYINPUT118), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n921), .A2(new_n909), .A3(new_n308), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n933), .A2(new_n886), .A3(new_n934), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT119), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n935), .A2(new_n936), .A3(new_n927), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n929), .A2(new_n931), .A3(new_n937), .ZN(new_n938));
  AND3_X1   g737(.A1(new_n719), .A2(new_n720), .A3(new_n888), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n938), .A2(new_n751), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(G141gat), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n719), .A2(new_n720), .A3(new_n888), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n930), .A2(new_n942), .ZN(new_n943));
  INV_X1    g742(.A(G141gat), .ZN(new_n944));
  NAND4_X1  g743(.A1(new_n943), .A2(KEYINPUT120), .A3(new_n944), .A4(new_n268), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n589), .B1(new_n885), .B2(new_n886), .ZN(new_n946));
  NAND4_X1  g745(.A1(new_n939), .A2(new_n944), .A3(new_n268), .A4(new_n946), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT120), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n945), .A2(new_n949), .ZN(new_n950));
  INV_X1    g749(.A(new_n950), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n941), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n908), .B1(new_n952), .B2(KEYINPUT58), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n950), .B1(new_n940), .B2(G141gat), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT58), .ZN(new_n955));
  NOR3_X1   g754(.A1(new_n954), .A2(KEYINPUT121), .A3(new_n955), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT122), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n938), .A2(new_n268), .A3(new_n939), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n958), .A2(G141gat), .ZN(new_n959));
  AND4_X1   g758(.A1(new_n957), .A2(new_n959), .A3(new_n955), .A4(new_n947), .ZN(new_n960));
  AOI21_X1  g759(.A(KEYINPUT58), .B1(new_n958), .B2(G141gat), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n957), .B1(new_n961), .B2(new_n947), .ZN(new_n962));
  OAI22_X1  g761(.A1(new_n953), .A2(new_n956), .B1(new_n960), .B2(new_n962), .ZN(G1344gat));
  INV_X1    g762(.A(G148gat), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n943), .A2(new_n964), .A3(new_n401), .ZN(new_n965));
  XOR2_X1   g764(.A(new_n965), .B(KEYINPUT123), .Z(new_n966));
  AND2_X1   g765(.A1(new_n938), .A2(new_n939), .ZN(new_n967));
  AOI211_X1 g766(.A(KEYINPUT59), .B(new_n964), .C1(new_n967), .C2(new_n401), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT59), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n369), .A2(new_n882), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n920), .B1(new_n872), .B2(new_n970), .ZN(new_n971));
  AOI22_X1  g770(.A1(new_n971), .A2(new_n308), .B1(new_n692), .B2(new_n402), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n926), .B1(new_n972), .B2(new_n589), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n973), .B1(new_n930), .B2(new_n926), .ZN(new_n974));
  AND2_X1   g773(.A1(new_n974), .A2(new_n401), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n975), .A2(new_n939), .ZN(new_n976));
  AOI21_X1  g775(.A(new_n969), .B1(new_n976), .B2(G148gat), .ZN(new_n977));
  OAI21_X1  g776(.A(new_n966), .B1(new_n968), .B2(new_n977), .ZN(G1345gat));
  NAND3_X1  g777(.A1(new_n938), .A2(new_n746), .A3(new_n939), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n979), .A2(G155gat), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n943), .A2(new_n538), .A3(new_n746), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  XNOR2_X1  g781(.A(new_n982), .B(KEYINPUT124), .ZN(G1346gat));
  AOI21_X1  g782(.A(G162gat), .B1(new_n943), .B2(new_n369), .ZN(new_n984));
  NOR2_X1   g783(.A1(new_n742), .A2(new_n539), .ZN(new_n985));
  AOI21_X1  g784(.A(new_n984), .B1(new_n967), .B2(new_n985), .ZN(G1347gat));
  NOR2_X1   g785(.A1(new_n705), .A2(new_n638), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n887), .A2(new_n987), .ZN(new_n988));
  NOR2_X1   g787(.A1(new_n988), .A2(new_n683), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n989), .A2(new_n460), .A3(new_n751), .ZN(new_n990));
  XNOR2_X1  g789(.A(new_n990), .B(KEYINPUT125), .ZN(new_n991));
  NOR2_X1   g790(.A1(new_n988), .A2(new_n892), .ZN(new_n992));
  XNOR2_X1  g791(.A(new_n992), .B(KEYINPUT126), .ZN(new_n993));
  AND2_X1   g792(.A1(new_n993), .A2(new_n268), .ZN(new_n994));
  OAI21_X1  g793(.A(new_n991), .B1(new_n994), .B2(new_n460), .ZN(G1348gat));
  AOI21_X1  g794(.A(G176gat), .B1(new_n989), .B2(new_n401), .ZN(new_n996));
  NOR2_X1   g795(.A1(new_n400), .A2(new_n461), .ZN(new_n997));
  AOI21_X1  g796(.A(new_n996), .B1(new_n993), .B2(new_n997), .ZN(G1349gat));
  NAND3_X1  g797(.A1(new_n989), .A2(new_n472), .A3(new_n746), .ZN(new_n999));
  AND2_X1   g798(.A1(new_n993), .A2(new_n746), .ZN(new_n1000));
  OAI21_X1  g799(.A(new_n999), .B1(new_n1000), .B2(new_n283), .ZN(new_n1001));
  NAND2_X1  g800(.A1(new_n1001), .A2(KEYINPUT60), .ZN(new_n1002));
  INV_X1    g801(.A(KEYINPUT60), .ZN(new_n1003));
  OAI211_X1 g802(.A(new_n999), .B(new_n1003), .C1(new_n1000), .C2(new_n283), .ZN(new_n1004));
  NAND2_X1  g803(.A1(new_n1002), .A2(new_n1004), .ZN(G1350gat));
  NAND3_X1  g804(.A1(new_n989), .A2(new_n473), .A3(new_n369), .ZN(new_n1006));
  INV_X1    g805(.A(KEYINPUT61), .ZN(new_n1007));
  NAND2_X1  g806(.A1(new_n993), .A2(new_n369), .ZN(new_n1008));
  AOI21_X1  g807(.A(new_n1007), .B1(new_n1008), .B2(G190gat), .ZN(new_n1009));
  AOI211_X1 g808(.A(KEYINPUT61), .B(new_n473), .C1(new_n993), .C2(new_n369), .ZN(new_n1010));
  OAI21_X1  g809(.A(new_n1006), .B1(new_n1009), .B2(new_n1010), .ZN(G1351gat));
  NAND2_X1  g810(.A1(new_n721), .A2(new_n987), .ZN(new_n1012));
  XNOR2_X1  g811(.A(new_n1012), .B(KEYINPUT127), .ZN(new_n1013));
  NAND2_X1  g812(.A1(new_n1013), .A2(new_n974), .ZN(new_n1014));
  OAI21_X1  g813(.A(G197gat), .B1(new_n1014), .B2(new_n692), .ZN(new_n1015));
  NOR2_X1   g814(.A1(new_n1012), .A2(new_n930), .ZN(new_n1016));
  INV_X1    g815(.A(G197gat), .ZN(new_n1017));
  NAND3_X1  g816(.A1(new_n1016), .A2(new_n1017), .A3(new_n751), .ZN(new_n1018));
  NAND2_X1  g817(.A1(new_n1015), .A2(new_n1018), .ZN(G1352gat));
  INV_X1    g818(.A(G204gat), .ZN(new_n1020));
  NAND3_X1  g819(.A1(new_n1016), .A2(new_n1020), .A3(new_n401), .ZN(new_n1021));
  XNOR2_X1  g820(.A(new_n1021), .B(KEYINPUT62), .ZN(new_n1022));
  AOI21_X1  g821(.A(new_n1020), .B1(new_n1013), .B2(new_n975), .ZN(new_n1023));
  OR2_X1    g822(.A1(new_n1022), .A2(new_n1023), .ZN(G1353gat));
  NAND3_X1  g823(.A1(new_n1016), .A2(new_n555), .A3(new_n746), .ZN(new_n1025));
  NAND3_X1  g824(.A1(new_n1013), .A2(new_n974), .A3(new_n746), .ZN(new_n1026));
  AND3_X1   g825(.A1(new_n1026), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1027));
  AOI21_X1  g826(.A(KEYINPUT63), .B1(new_n1026), .B2(G211gat), .ZN(new_n1028));
  OAI21_X1  g827(.A(new_n1025), .B1(new_n1027), .B2(new_n1028), .ZN(G1354gat));
  OAI21_X1  g828(.A(G218gat), .B1(new_n1014), .B2(new_n742), .ZN(new_n1030));
  NAND3_X1  g829(.A1(new_n1016), .A2(new_n556), .A3(new_n369), .ZN(new_n1031));
  NAND2_X1  g830(.A1(new_n1030), .A2(new_n1031), .ZN(G1355gat));
endmodule


