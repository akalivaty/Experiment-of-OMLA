

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X1 U560 ( .A1(n759), .A2(n758), .ZN(n760) );
  INV_X1 U561 ( .A(n742), .ZN(n527) );
  NOR2_X2 U562 ( .A1(n697), .A2(G1384), .ZN(n793) );
  NOR2_X2 U563 ( .A1(n552), .A2(n551), .ZN(n697) );
  OR2_X2 U564 ( .A1(n699), .A2(n698), .ZN(n700) );
  INV_X1 U565 ( .A(KEYINPUT17), .ZN(n546) );
  AND2_X1 U566 ( .A1(n790), .A2(n529), .ZN(n823) );
  NAND2_X1 U567 ( .A1(n583), .A2(n582), .ZN(n701) );
  NOR2_X2 U568 ( .A1(G2104), .A2(G2105), .ZN(n547) );
  INV_X2 U569 ( .A(G2105), .ZN(n548) );
  NOR2_X2 U570 ( .A1(n701), .A2(n700), .ZN(n791) );
  INV_X1 U571 ( .A(KEYINPUT89), .ZN(n542) );
  XNOR2_X1 U572 ( .A(n595), .B(n594), .ZN(n596) );
  NOR2_X1 U573 ( .A1(G543), .A2(n536), .ZN(n531) );
  NOR2_X1 U574 ( .A1(n777), .A2(n776), .ZN(n528) );
  OR2_X1 U575 ( .A1(n789), .A2(n788), .ZN(n529) );
  XOR2_X1 U576 ( .A(n762), .B(KEYINPUT97), .Z(n530) );
  INV_X1 U577 ( .A(KEYINPUT93), .ZN(n715) );
  XNOR2_X1 U578 ( .A(n715), .B(KEYINPUT27), .ZN(n716) );
  XNOR2_X1 U579 ( .A(n717), .B(n716), .ZN(n719) );
  NOR2_X1 U580 ( .A1(n722), .A2(n723), .ZN(n724) );
  INV_X1 U581 ( .A(n988), .ZN(n776) );
  NAND2_X1 U582 ( .A1(n664), .A2(G54), .ZN(n602) );
  XNOR2_X1 U583 ( .A(KEYINPUT14), .B(KEYINPUT71), .ZN(n594) );
  NOR2_X1 U584 ( .A1(n649), .A2(G651), .ZN(n532) );
  INV_X1 U585 ( .A(KEYINPUT103), .ZN(n827) );
  XOR2_X1 U586 ( .A(KEYINPUT0), .B(G543), .Z(n649) );
  NAND2_X1 U587 ( .A1(n624), .A2(G137), .ZN(n585) );
  INV_X1 U588 ( .A(G651), .ZN(n536) );
  XOR2_X2 U589 ( .A(KEYINPUT1), .B(n531), .Z(n661) );
  NAND2_X1 U590 ( .A1(G64), .A2(n661), .ZN(n534) );
  XNOR2_X2 U591 ( .A(KEYINPUT64), .B(n532), .ZN(n664) );
  NAND2_X1 U592 ( .A1(G52), .A2(n664), .ZN(n533) );
  NAND2_X1 U593 ( .A1(n534), .A2(n533), .ZN(n541) );
  NOR2_X1 U594 ( .A1(G543), .A2(G651), .ZN(n660) );
  NAND2_X1 U595 ( .A1(n660), .A2(G90), .ZN(n535) );
  XOR2_X1 U596 ( .A(KEYINPUT67), .B(n535), .Z(n538) );
  NOR2_X2 U597 ( .A1(n649), .A2(n536), .ZN(n657) );
  NAND2_X1 U598 ( .A1(n657), .A2(G77), .ZN(n537) );
  NAND2_X1 U599 ( .A1(n538), .A2(n537), .ZN(n539) );
  XOR2_X1 U600 ( .A(KEYINPUT9), .B(n539), .Z(n540) );
  NOR2_X1 U601 ( .A1(n541), .A2(n540), .ZN(G171) );
  AND2_X1 U602 ( .A1(G452), .A2(G94), .ZN(G173) );
  NOR2_X2 U603 ( .A1(G2104), .A2(n548), .ZN(n895) );
  NAND2_X1 U604 ( .A1(n895), .A2(G126), .ZN(n545) );
  AND2_X4 U605 ( .A1(n548), .A2(G2104), .ZN(n619) );
  NAND2_X1 U606 ( .A1(G102), .A2(n619), .ZN(n543) );
  XNOR2_X1 U607 ( .A(n543), .B(n542), .ZN(n544) );
  NAND2_X1 U608 ( .A1(n545), .A2(n544), .ZN(n552) );
  XNOR2_X2 U609 ( .A(n547), .B(n546), .ZN(n624) );
  NAND2_X1 U610 ( .A1(G138), .A2(n624), .ZN(n550) );
  AND2_X1 U611 ( .A1(G2104), .A2(G2105), .ZN(n894) );
  NAND2_X1 U612 ( .A1(G114), .A2(n894), .ZN(n549) );
  NAND2_X1 U613 ( .A1(n550), .A2(n549), .ZN(n551) );
  BUF_X1 U614 ( .A(n697), .Z(G164) );
  INV_X1 U615 ( .A(G57), .ZN(G237) );
  NAND2_X1 U616 ( .A1(G62), .A2(n661), .ZN(n554) );
  NAND2_X1 U617 ( .A1(G50), .A2(n664), .ZN(n553) );
  NAND2_X1 U618 ( .A1(n554), .A2(n553), .ZN(n559) );
  NAND2_X1 U619 ( .A1(G88), .A2(n660), .ZN(n556) );
  NAND2_X1 U620 ( .A1(G75), .A2(n657), .ZN(n555) );
  NAND2_X1 U621 ( .A1(n556), .A2(n555), .ZN(n557) );
  XOR2_X1 U622 ( .A(KEYINPUT85), .B(n557), .Z(n558) );
  NOR2_X1 U623 ( .A1(n559), .A2(n558), .ZN(G166) );
  NAND2_X1 U624 ( .A1(G91), .A2(n660), .ZN(n561) );
  NAND2_X1 U625 ( .A1(G78), .A2(n657), .ZN(n560) );
  NAND2_X1 U626 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U627 ( .A(KEYINPUT68), .B(n562), .Z(n566) );
  NAND2_X1 U628 ( .A1(n664), .A2(G53), .ZN(n564) );
  NAND2_X1 U629 ( .A1(G65), .A2(n661), .ZN(n563) );
  AND2_X1 U630 ( .A1(n564), .A2(n563), .ZN(n565) );
  NAND2_X1 U631 ( .A1(n566), .A2(n565), .ZN(G299) );
  XNOR2_X1 U632 ( .A(KEYINPUT73), .B(KEYINPUT74), .ZN(n572) );
  NAND2_X1 U633 ( .A1(n660), .A2(G89), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n567), .B(KEYINPUT4), .ZN(n569) );
  NAND2_X1 U635 ( .A1(G76), .A2(n657), .ZN(n568) );
  NAND2_X1 U636 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n570), .B(KEYINPUT5), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(n577) );
  NAND2_X1 U639 ( .A1(G63), .A2(n661), .ZN(n574) );
  NAND2_X1 U640 ( .A1(G51), .A2(n664), .ZN(n573) );
  NAND2_X1 U641 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U642 ( .A(KEYINPUT6), .B(n575), .ZN(n576) );
  NOR2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n579) );
  XNOR2_X1 U644 ( .A(KEYINPUT7), .B(KEYINPUT75), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n579), .B(n578), .ZN(G168) );
  XOR2_X1 U646 ( .A(G168), .B(KEYINPUT8), .Z(n580) );
  XNOR2_X1 U647 ( .A(KEYINPUT76), .B(n580), .ZN(G286) );
  NAND2_X1 U648 ( .A1(n894), .A2(G113), .ZN(n583) );
  NAND2_X1 U649 ( .A1(G101), .A2(n619), .ZN(n581) );
  XOR2_X1 U650 ( .A(KEYINPUT23), .B(n581), .Z(n582) );
  NAND2_X1 U651 ( .A1(G125), .A2(n895), .ZN(n584) );
  NAND2_X1 U652 ( .A1(n585), .A2(n584), .ZN(n699) );
  NOR2_X1 U653 ( .A1(n701), .A2(n699), .ZN(G160) );
  XOR2_X1 U654 ( .A(KEYINPUT69), .B(KEYINPUT10), .Z(n587) );
  NAND2_X1 U655 ( .A1(G7), .A2(G661), .ZN(n586) );
  XNOR2_X1 U656 ( .A(n587), .B(n586), .ZN(G223) );
  XOR2_X1 U657 ( .A(KEYINPUT70), .B(KEYINPUT11), .Z(n589) );
  INV_X1 U658 ( .A(G223), .ZN(n844) );
  NAND2_X1 U659 ( .A1(G567), .A2(n844), .ZN(n588) );
  XNOR2_X1 U660 ( .A(n589), .B(n588), .ZN(G234) );
  NAND2_X1 U661 ( .A1(n660), .A2(G81), .ZN(n590) );
  XNOR2_X1 U662 ( .A(n590), .B(KEYINPUT12), .ZN(n592) );
  NAND2_X1 U663 ( .A1(G68), .A2(n657), .ZN(n591) );
  NAND2_X1 U664 ( .A1(n592), .A2(n591), .ZN(n593) );
  XOR2_X1 U665 ( .A(KEYINPUT13), .B(n593), .Z(n597) );
  NAND2_X1 U666 ( .A1(G56), .A2(n661), .ZN(n595) );
  NOR2_X1 U667 ( .A1(n597), .A2(n596), .ZN(n599) );
  NAND2_X1 U668 ( .A1(G43), .A2(n664), .ZN(n598) );
  NAND2_X1 U669 ( .A1(n599), .A2(n598), .ZN(n992) );
  INV_X1 U670 ( .A(G860), .ZN(n612) );
  OR2_X1 U671 ( .A1(n992), .A2(n612), .ZN(G153) );
  INV_X1 U672 ( .A(G171), .ZN(G301) );
  INV_X1 U673 ( .A(G868), .ZN(n678) );
  NAND2_X1 U674 ( .A1(G92), .A2(n660), .ZN(n601) );
  NAND2_X1 U675 ( .A1(G79), .A2(n657), .ZN(n600) );
  NAND2_X1 U676 ( .A1(n601), .A2(n600), .ZN(n605) );
  NAND2_X1 U677 ( .A1(G66), .A2(n661), .ZN(n603) );
  NAND2_X1 U678 ( .A1(n603), .A2(n602), .ZN(n604) );
  NOR2_X1 U679 ( .A1(n605), .A2(n604), .ZN(n606) );
  XOR2_X2 U680 ( .A(KEYINPUT15), .B(n606), .Z(n991) );
  AND2_X1 U681 ( .A1(n678), .A2(n991), .ZN(n608) );
  NOR2_X1 U682 ( .A1(n678), .A2(G301), .ZN(n607) );
  NOR2_X1 U683 ( .A1(n608), .A2(n607), .ZN(n609) );
  XNOR2_X1 U684 ( .A(KEYINPUT72), .B(n609), .ZN(G284) );
  NAND2_X1 U685 ( .A1(G868), .A2(G286), .ZN(n611) );
  NAND2_X1 U686 ( .A1(G299), .A2(n678), .ZN(n610) );
  NAND2_X1 U687 ( .A1(n611), .A2(n610), .ZN(G297) );
  NAND2_X1 U688 ( .A1(n612), .A2(G559), .ZN(n613) );
  NAND2_X1 U689 ( .A1(n613), .A2(n991), .ZN(n614) );
  XNOR2_X1 U690 ( .A(n614), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U691 ( .A1(G868), .A2(n992), .ZN(n617) );
  NAND2_X1 U692 ( .A1(G868), .A2(n991), .ZN(n615) );
  NOR2_X1 U693 ( .A1(G559), .A2(n615), .ZN(n616) );
  NOR2_X1 U694 ( .A1(n617), .A2(n616), .ZN(n618) );
  XOR2_X1 U695 ( .A(KEYINPUT77), .B(n618), .Z(G282) );
  NAND2_X1 U696 ( .A1(G99), .A2(n619), .ZN(n621) );
  NAND2_X1 U697 ( .A1(G111), .A2(n894), .ZN(n620) );
  NAND2_X1 U698 ( .A1(n621), .A2(n620), .ZN(n622) );
  XNOR2_X1 U699 ( .A(KEYINPUT78), .B(n622), .ZN(n628) );
  NAND2_X1 U700 ( .A1(G123), .A2(n895), .ZN(n623) );
  XNOR2_X1 U701 ( .A(n623), .B(KEYINPUT18), .ZN(n626) );
  NAND2_X1 U702 ( .A1(n624), .A2(G135), .ZN(n625) );
  NAND2_X1 U703 ( .A1(n626), .A2(n625), .ZN(n627) );
  NOR2_X1 U704 ( .A1(n628), .A2(n627), .ZN(n944) );
  XNOR2_X1 U705 ( .A(G2096), .B(n944), .ZN(n630) );
  INV_X1 U706 ( .A(G2100), .ZN(n629) );
  NAND2_X1 U707 ( .A1(n630), .A2(n629), .ZN(G156) );
  NAND2_X1 U708 ( .A1(n664), .A2(G55), .ZN(n631) );
  XNOR2_X1 U709 ( .A(n631), .B(KEYINPUT80), .ZN(n638) );
  NAND2_X1 U710 ( .A1(G80), .A2(n657), .ZN(n633) );
  NAND2_X1 U711 ( .A1(G67), .A2(n661), .ZN(n632) );
  NAND2_X1 U712 ( .A1(n633), .A2(n632), .ZN(n636) );
  NAND2_X1 U713 ( .A1(G93), .A2(n660), .ZN(n634) );
  XNOR2_X1 U714 ( .A(KEYINPUT79), .B(n634), .ZN(n635) );
  NOR2_X1 U715 ( .A1(n636), .A2(n635), .ZN(n637) );
  NAND2_X1 U716 ( .A1(n638), .A2(n637), .ZN(n679) );
  NAND2_X1 U717 ( .A1(n991), .A2(G559), .ZN(n676) );
  XNOR2_X1 U718 ( .A(n992), .B(n676), .ZN(n639) );
  NOR2_X1 U719 ( .A1(G860), .A2(n639), .ZN(n640) );
  XOR2_X1 U720 ( .A(n679), .B(n640), .Z(G145) );
  NAND2_X1 U721 ( .A1(n660), .A2(G85), .ZN(n641) );
  XOR2_X1 U722 ( .A(KEYINPUT65), .B(n641), .Z(n643) );
  NAND2_X1 U723 ( .A1(n657), .A2(G72), .ZN(n642) );
  NAND2_X1 U724 ( .A1(n643), .A2(n642), .ZN(n644) );
  XOR2_X1 U725 ( .A(KEYINPUT66), .B(n644), .Z(n648) );
  NAND2_X1 U726 ( .A1(n664), .A2(G47), .ZN(n646) );
  NAND2_X1 U727 ( .A1(G60), .A2(n661), .ZN(n645) );
  AND2_X1 U728 ( .A1(n646), .A2(n645), .ZN(n647) );
  NAND2_X1 U729 ( .A1(n648), .A2(n647), .ZN(G290) );
  NAND2_X1 U730 ( .A1(G87), .A2(n649), .ZN(n655) );
  NAND2_X1 U731 ( .A1(G651), .A2(G74), .ZN(n651) );
  NAND2_X1 U732 ( .A1(G49), .A2(n664), .ZN(n650) );
  NAND2_X1 U733 ( .A1(n651), .A2(n650), .ZN(n652) );
  NOR2_X1 U734 ( .A1(n661), .A2(n652), .ZN(n653) );
  XOR2_X1 U735 ( .A(KEYINPUT81), .B(n653), .Z(n654) );
  NAND2_X1 U736 ( .A1(n655), .A2(n654), .ZN(n656) );
  XNOR2_X1 U737 ( .A(n656), .B(KEYINPUT82), .ZN(G288) );
  XOR2_X1 U738 ( .A(KEYINPUT2), .B(KEYINPUT83), .Z(n659) );
  NAND2_X1 U739 ( .A1(G73), .A2(n657), .ZN(n658) );
  XNOR2_X1 U740 ( .A(n659), .B(n658), .ZN(n669) );
  NAND2_X1 U741 ( .A1(G86), .A2(n660), .ZN(n663) );
  NAND2_X1 U742 ( .A1(G61), .A2(n661), .ZN(n662) );
  NAND2_X1 U743 ( .A1(n663), .A2(n662), .ZN(n667) );
  NAND2_X1 U744 ( .A1(n664), .A2(G48), .ZN(n665) );
  XOR2_X1 U745 ( .A(KEYINPUT84), .B(n665), .Z(n666) );
  NOR2_X1 U746 ( .A1(n667), .A2(n666), .ZN(n668) );
  NAND2_X1 U747 ( .A1(n669), .A2(n668), .ZN(G305) );
  INV_X1 U748 ( .A(G299), .ZN(n723) );
  XNOR2_X1 U749 ( .A(n723), .B(G290), .ZN(n675) );
  XNOR2_X1 U750 ( .A(n679), .B(KEYINPUT19), .ZN(n671) );
  XNOR2_X1 U751 ( .A(G166), .B(G288), .ZN(n670) );
  XNOR2_X1 U752 ( .A(n671), .B(n670), .ZN(n672) );
  XOR2_X1 U753 ( .A(n672), .B(G305), .Z(n673) );
  XNOR2_X1 U754 ( .A(n992), .B(n673), .ZN(n674) );
  XNOR2_X1 U755 ( .A(n675), .B(n674), .ZN(n913) );
  XNOR2_X1 U756 ( .A(n913), .B(n676), .ZN(n677) );
  NOR2_X1 U757 ( .A1(n678), .A2(n677), .ZN(n681) );
  NOR2_X1 U758 ( .A1(G868), .A2(n679), .ZN(n680) );
  NOR2_X1 U759 ( .A1(n681), .A2(n680), .ZN(G295) );
  NAND2_X1 U760 ( .A1(G2078), .A2(G2084), .ZN(n682) );
  XOR2_X1 U761 ( .A(KEYINPUT20), .B(n682), .Z(n683) );
  NAND2_X1 U762 ( .A1(G2090), .A2(n683), .ZN(n684) );
  XNOR2_X1 U763 ( .A(KEYINPUT21), .B(n684), .ZN(n685) );
  NAND2_X1 U764 ( .A1(n685), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U765 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U766 ( .A1(G69), .A2(G120), .ZN(n686) );
  NOR2_X1 U767 ( .A1(G237), .A2(n686), .ZN(n687) );
  NAND2_X1 U768 ( .A1(G108), .A2(n687), .ZN(n935) );
  NAND2_X1 U769 ( .A1(G567), .A2(n935), .ZN(n694) );
  NAND2_X1 U770 ( .A1(G132), .A2(G82), .ZN(n688) );
  XNOR2_X1 U771 ( .A(n688), .B(KEYINPUT86), .ZN(n689) );
  XNOR2_X1 U772 ( .A(n689), .B(KEYINPUT22), .ZN(n690) );
  NOR2_X1 U773 ( .A1(G218), .A2(n690), .ZN(n691) );
  XOR2_X1 U774 ( .A(KEYINPUT87), .B(n691), .Z(n692) );
  NAND2_X1 U775 ( .A1(G96), .A2(n692), .ZN(n934) );
  NAND2_X1 U776 ( .A1(G2106), .A2(n934), .ZN(n693) );
  NAND2_X1 U777 ( .A1(n694), .A2(n693), .ZN(n870) );
  NAND2_X1 U778 ( .A1(G661), .A2(G483), .ZN(n695) );
  XNOR2_X1 U779 ( .A(KEYINPUT88), .B(n695), .ZN(n696) );
  NOR2_X1 U780 ( .A1(n870), .A2(n696), .ZN(n848) );
  NAND2_X1 U781 ( .A1(n848), .A2(G36), .ZN(G176) );
  INV_X1 U782 ( .A(G166), .ZN(G303) );
  INV_X1 U783 ( .A(G40), .ZN(n698) );
  NAND2_X1 U784 ( .A1(n793), .A2(n791), .ZN(n734) );
  INV_X1 U785 ( .A(n734), .ZN(n702) );
  NAND2_X1 U786 ( .A1(G1996), .A2(n702), .ZN(n703) );
  XNOR2_X1 U787 ( .A(n703), .B(KEYINPUT26), .ZN(n705) );
  BUF_X2 U788 ( .A(n734), .Z(n742) );
  NAND2_X1 U789 ( .A1(G1341), .A2(n742), .ZN(n704) );
  NAND2_X1 U790 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U791 ( .A(n706), .B(KEYINPUT94), .ZN(n707) );
  NOR2_X1 U792 ( .A1(n707), .A2(n992), .ZN(n712) );
  NAND2_X1 U793 ( .A1(n712), .A2(n991), .ZN(n711) );
  NOR2_X1 U794 ( .A1(n527), .A2(G1348), .ZN(n709) );
  NOR2_X1 U795 ( .A1(G2067), .A2(n742), .ZN(n708) );
  NOR2_X1 U796 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U797 ( .A1(n711), .A2(n710), .ZN(n714) );
  OR2_X1 U798 ( .A1(n991), .A2(n712), .ZN(n713) );
  NAND2_X1 U799 ( .A1(n714), .A2(n713), .ZN(n721) );
  NAND2_X1 U800 ( .A1(n527), .A2(G2072), .ZN(n717) );
  AND2_X1 U801 ( .A1(n742), .A2(G1956), .ZN(n718) );
  NOR2_X1 U802 ( .A1(n719), .A2(n718), .ZN(n722) );
  NAND2_X1 U803 ( .A1(n723), .A2(n722), .ZN(n720) );
  NAND2_X1 U804 ( .A1(n721), .A2(n720), .ZN(n726) );
  XOR2_X1 U805 ( .A(n724), .B(KEYINPUT28), .Z(n725) );
  NAND2_X1 U806 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U807 ( .A(n727), .B(KEYINPUT29), .ZN(n731) );
  XNOR2_X1 U808 ( .A(G2078), .B(KEYINPUT25), .ZN(n963) );
  NOR2_X1 U809 ( .A1(n742), .A2(n963), .ZN(n729) );
  INV_X1 U810 ( .A(G1961), .ZN(n1013) );
  NOR2_X1 U811 ( .A1(n527), .A2(n1013), .ZN(n728) );
  NOR2_X1 U812 ( .A1(n729), .A2(n728), .ZN(n733) );
  AND2_X1 U813 ( .A1(G171), .A2(n733), .ZN(n730) );
  NOR2_X2 U814 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U815 ( .A(n732), .B(KEYINPUT95), .ZN(n754) );
  NOR2_X1 U816 ( .A1(G171), .A2(n733), .ZN(n740) );
  NAND2_X1 U817 ( .A1(G8), .A2(n734), .ZN(n789) );
  NOR2_X1 U818 ( .A1(G1966), .A2(n789), .ZN(n756) );
  NOR2_X1 U819 ( .A1(G2084), .A2(n742), .ZN(n755) );
  NOR2_X1 U820 ( .A1(n756), .A2(n755), .ZN(n735) );
  XNOR2_X1 U821 ( .A(KEYINPUT96), .B(n735), .ZN(n736) );
  NAND2_X1 U822 ( .A1(n736), .A2(G8), .ZN(n737) );
  XNOR2_X1 U823 ( .A(KEYINPUT30), .B(n737), .ZN(n738) );
  NOR2_X1 U824 ( .A1(G168), .A2(n738), .ZN(n739) );
  NOR2_X1 U825 ( .A1(n740), .A2(n739), .ZN(n741) );
  XOR2_X1 U826 ( .A(KEYINPUT31), .B(n741), .Z(n753) );
  NOR2_X1 U827 ( .A1(G1971), .A2(n789), .ZN(n744) );
  NOR2_X1 U828 ( .A1(G2090), .A2(n742), .ZN(n743) );
  NOR2_X1 U829 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U830 ( .A1(G303), .A2(n745), .ZN(n747) );
  AND2_X1 U831 ( .A1(n753), .A2(n747), .ZN(n746) );
  NAND2_X1 U832 ( .A1(n754), .A2(n746), .ZN(n751) );
  INV_X1 U833 ( .A(n747), .ZN(n748) );
  OR2_X1 U834 ( .A1(n748), .A2(G286), .ZN(n749) );
  AND2_X1 U835 ( .A1(n749), .A2(G8), .ZN(n750) );
  NAND2_X1 U836 ( .A1(n751), .A2(n750), .ZN(n752) );
  XNOR2_X1 U837 ( .A(n752), .B(KEYINPUT32), .ZN(n761) );
  AND2_X1 U838 ( .A1(n754), .A2(n753), .ZN(n759) );
  AND2_X1 U839 ( .A1(G8), .A2(n755), .ZN(n757) );
  OR2_X1 U840 ( .A1(n757), .A2(n756), .ZN(n758) );
  NAND2_X1 U841 ( .A1(n760), .A2(n761), .ZN(n779) );
  NOR2_X1 U842 ( .A1(G1976), .A2(G288), .ZN(n1003) );
  NOR2_X1 U843 ( .A1(G1971), .A2(G303), .ZN(n762) );
  NOR2_X1 U844 ( .A1(n1003), .A2(n530), .ZN(n763) );
  NAND2_X1 U845 ( .A1(n779), .A2(n763), .ZN(n764) );
  NAND2_X1 U846 ( .A1(G1976), .A2(G288), .ZN(n1004) );
  NAND2_X1 U847 ( .A1(n764), .A2(n1004), .ZN(n765) );
  XNOR2_X1 U848 ( .A(n765), .B(KEYINPUT98), .ZN(n767) );
  OR2_X1 U849 ( .A1(n789), .A2(KEYINPUT99), .ZN(n766) );
  NOR2_X1 U850 ( .A1(n767), .A2(n766), .ZN(n768) );
  INV_X1 U851 ( .A(n768), .ZN(n770) );
  INV_X1 U852 ( .A(KEYINPUT33), .ZN(n769) );
  NAND2_X1 U853 ( .A1(n770), .A2(n769), .ZN(n778) );
  INV_X1 U854 ( .A(KEYINPUT99), .ZN(n772) );
  NAND2_X1 U855 ( .A1(n1003), .A2(KEYINPUT33), .ZN(n771) );
  NAND2_X1 U856 ( .A1(n772), .A2(n771), .ZN(n774) );
  NAND2_X1 U857 ( .A1(n1003), .A2(KEYINPUT99), .ZN(n773) );
  NAND2_X1 U858 ( .A1(n774), .A2(n773), .ZN(n775) );
  NOR2_X1 U859 ( .A1(n789), .A2(n775), .ZN(n777) );
  XOR2_X1 U860 ( .A(G1981), .B(G305), .Z(n988) );
  NAND2_X1 U861 ( .A1(n778), .A2(n528), .ZN(n785) );
  NOR2_X1 U862 ( .A1(G2090), .A2(G303), .ZN(n780) );
  NAND2_X1 U863 ( .A1(G8), .A2(n780), .ZN(n781) );
  NAND2_X1 U864 ( .A1(n779), .A2(n781), .ZN(n782) );
  XNOR2_X1 U865 ( .A(n782), .B(KEYINPUT100), .ZN(n783) );
  NAND2_X1 U866 ( .A1(n783), .A2(n789), .ZN(n784) );
  NAND2_X1 U867 ( .A1(n785), .A2(n784), .ZN(n786) );
  XNOR2_X1 U868 ( .A(n786), .B(KEYINPUT101), .ZN(n790) );
  NOR2_X1 U869 ( .A1(G1981), .A2(G305), .ZN(n787) );
  XOR2_X1 U870 ( .A(n787), .B(KEYINPUT24), .Z(n788) );
  INV_X1 U871 ( .A(n791), .ZN(n792) );
  NOR2_X1 U872 ( .A1(n793), .A2(n792), .ZN(n839) );
  NAND2_X1 U873 ( .A1(G104), .A2(n619), .ZN(n795) );
  NAND2_X1 U874 ( .A1(G140), .A2(n624), .ZN(n794) );
  NAND2_X1 U875 ( .A1(n795), .A2(n794), .ZN(n796) );
  XNOR2_X1 U876 ( .A(KEYINPUT34), .B(n796), .ZN(n801) );
  NAND2_X1 U877 ( .A1(G116), .A2(n894), .ZN(n798) );
  NAND2_X1 U878 ( .A1(G128), .A2(n895), .ZN(n797) );
  NAND2_X1 U879 ( .A1(n798), .A2(n797), .ZN(n799) );
  XOR2_X1 U880 ( .A(KEYINPUT35), .B(n799), .Z(n800) );
  NOR2_X1 U881 ( .A1(n801), .A2(n800), .ZN(n802) );
  XNOR2_X1 U882 ( .A(KEYINPUT36), .B(n802), .ZN(n911) );
  XNOR2_X1 U883 ( .A(KEYINPUT37), .B(G2067), .ZN(n837) );
  NOR2_X1 U884 ( .A1(n911), .A2(n837), .ZN(n942) );
  NAND2_X1 U885 ( .A1(n839), .A2(n942), .ZN(n835) );
  NAND2_X1 U886 ( .A1(G95), .A2(n619), .ZN(n804) );
  NAND2_X1 U887 ( .A1(G107), .A2(n894), .ZN(n803) );
  NAND2_X1 U888 ( .A1(n804), .A2(n803), .ZN(n808) );
  NAND2_X1 U889 ( .A1(G131), .A2(n624), .ZN(n806) );
  NAND2_X1 U890 ( .A1(G119), .A2(n895), .ZN(n805) );
  NAND2_X1 U891 ( .A1(n806), .A2(n805), .ZN(n807) );
  OR2_X1 U892 ( .A1(n808), .A2(n807), .ZN(n880) );
  NAND2_X1 U893 ( .A1(G1991), .A2(n880), .ZN(n819) );
  XOR2_X1 U894 ( .A(KEYINPUT90), .B(KEYINPUT38), .Z(n810) );
  NAND2_X1 U895 ( .A1(G105), .A2(n619), .ZN(n809) );
  XNOR2_X1 U896 ( .A(n810), .B(n809), .ZN(n814) );
  NAND2_X1 U897 ( .A1(G117), .A2(n894), .ZN(n812) );
  NAND2_X1 U898 ( .A1(G129), .A2(n895), .ZN(n811) );
  NAND2_X1 U899 ( .A1(n812), .A2(n811), .ZN(n813) );
  NOR2_X1 U900 ( .A1(n814), .A2(n813), .ZN(n815) );
  XOR2_X1 U901 ( .A(KEYINPUT91), .B(n815), .Z(n817) );
  NAND2_X1 U902 ( .A1(n624), .A2(G141), .ZN(n816) );
  NAND2_X1 U903 ( .A1(n817), .A2(n816), .ZN(n903) );
  NAND2_X1 U904 ( .A1(G1996), .A2(n903), .ZN(n818) );
  NAND2_X1 U905 ( .A1(n819), .A2(n818), .ZN(n820) );
  XOR2_X1 U906 ( .A(KEYINPUT92), .B(n820), .Z(n955) );
  INV_X1 U907 ( .A(n955), .ZN(n821) );
  NAND2_X1 U908 ( .A1(n839), .A2(n821), .ZN(n829) );
  NAND2_X1 U909 ( .A1(n835), .A2(n829), .ZN(n822) );
  NOR2_X1 U910 ( .A1(n823), .A2(n822), .ZN(n824) );
  XNOR2_X1 U911 ( .A(n824), .B(KEYINPUT102), .ZN(n826) );
  XNOR2_X1 U912 ( .A(G1986), .B(G290), .ZN(n999) );
  NAND2_X1 U913 ( .A1(n839), .A2(n999), .ZN(n825) );
  NAND2_X1 U914 ( .A1(n826), .A2(n825), .ZN(n828) );
  XNOR2_X1 U915 ( .A(n828), .B(n827), .ZN(n842) );
  NOR2_X1 U916 ( .A1(G1996), .A2(n903), .ZN(n952) );
  INV_X1 U917 ( .A(n829), .ZN(n832) );
  NOR2_X1 U918 ( .A1(G1986), .A2(G290), .ZN(n830) );
  NOR2_X1 U919 ( .A1(G1991), .A2(n880), .ZN(n948) );
  NOR2_X1 U920 ( .A1(n830), .A2(n948), .ZN(n831) );
  NOR2_X1 U921 ( .A1(n832), .A2(n831), .ZN(n833) );
  NOR2_X1 U922 ( .A1(n952), .A2(n833), .ZN(n834) );
  XNOR2_X1 U923 ( .A(n834), .B(KEYINPUT39), .ZN(n836) );
  NAND2_X1 U924 ( .A1(n836), .A2(n835), .ZN(n838) );
  NAND2_X1 U925 ( .A1(n911), .A2(n837), .ZN(n945) );
  NAND2_X1 U926 ( .A1(n838), .A2(n945), .ZN(n840) );
  NAND2_X1 U927 ( .A1(n840), .A2(n839), .ZN(n841) );
  NAND2_X1 U928 ( .A1(n842), .A2(n841), .ZN(n843) );
  XNOR2_X1 U929 ( .A(n843), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U930 ( .A1(n844), .A2(G2106), .ZN(n845) );
  XOR2_X1 U931 ( .A(KEYINPUT105), .B(n845), .Z(G217) );
  AND2_X1 U932 ( .A1(G15), .A2(G2), .ZN(n846) );
  NAND2_X1 U933 ( .A1(G661), .A2(n846), .ZN(G259) );
  NAND2_X1 U934 ( .A1(G3), .A2(G1), .ZN(n847) );
  NAND2_X1 U935 ( .A1(n848), .A2(n847), .ZN(G188) );
  XOR2_X1 U936 ( .A(G1976), .B(G1971), .Z(n850) );
  XNOR2_X1 U937 ( .A(G1986), .B(G1956), .ZN(n849) );
  XNOR2_X1 U938 ( .A(n850), .B(n849), .ZN(n860) );
  XOR2_X1 U939 ( .A(KEYINPUT41), .B(KEYINPUT108), .Z(n852) );
  XNOR2_X1 U940 ( .A(G1996), .B(KEYINPUT107), .ZN(n851) );
  XNOR2_X1 U941 ( .A(n852), .B(n851), .ZN(n856) );
  XOR2_X1 U942 ( .A(G1961), .B(G1966), .Z(n854) );
  XNOR2_X1 U943 ( .A(G1991), .B(G1981), .ZN(n853) );
  XNOR2_X1 U944 ( .A(n854), .B(n853), .ZN(n855) );
  XOR2_X1 U945 ( .A(n856), .B(n855), .Z(n858) );
  XNOR2_X1 U946 ( .A(G2474), .B(KEYINPUT109), .ZN(n857) );
  XNOR2_X1 U947 ( .A(n858), .B(n857), .ZN(n859) );
  XOR2_X1 U948 ( .A(n860), .B(n859), .Z(G229) );
  XOR2_X1 U949 ( .A(G2096), .B(KEYINPUT43), .Z(n862) );
  XNOR2_X1 U950 ( .A(G2090), .B(G2678), .ZN(n861) );
  XNOR2_X1 U951 ( .A(n862), .B(n861), .ZN(n863) );
  XOR2_X1 U952 ( .A(n863), .B(KEYINPUT106), .Z(n865) );
  XNOR2_X1 U953 ( .A(G2067), .B(G2072), .ZN(n864) );
  XNOR2_X1 U954 ( .A(n865), .B(n864), .ZN(n869) );
  XOR2_X1 U955 ( .A(KEYINPUT42), .B(G2100), .Z(n867) );
  XNOR2_X1 U956 ( .A(G2078), .B(G2084), .ZN(n866) );
  XNOR2_X1 U957 ( .A(n867), .B(n866), .ZN(n868) );
  XNOR2_X1 U958 ( .A(n869), .B(n868), .ZN(G227) );
  INV_X1 U959 ( .A(n870), .ZN(G319) );
  NAND2_X1 U960 ( .A1(n895), .A2(G124), .ZN(n871) );
  XNOR2_X1 U961 ( .A(n871), .B(KEYINPUT44), .ZN(n873) );
  NAND2_X1 U962 ( .A1(G136), .A2(n624), .ZN(n872) );
  NAND2_X1 U963 ( .A1(n873), .A2(n872), .ZN(n874) );
  XNOR2_X1 U964 ( .A(KEYINPUT110), .B(n874), .ZN(n878) );
  NAND2_X1 U965 ( .A1(G100), .A2(n619), .ZN(n876) );
  NAND2_X1 U966 ( .A1(G112), .A2(n894), .ZN(n875) );
  NAND2_X1 U967 ( .A1(n876), .A2(n875), .ZN(n877) );
  NOR2_X1 U968 ( .A1(n878), .A2(n877), .ZN(n879) );
  XOR2_X1 U969 ( .A(KEYINPUT111), .B(n879), .Z(G162) );
  XNOR2_X1 U970 ( .A(KEYINPUT114), .B(KEYINPUT46), .ZN(n882) );
  XNOR2_X1 U971 ( .A(n880), .B(KEYINPUT113), .ZN(n881) );
  XNOR2_X1 U972 ( .A(n882), .B(n881), .ZN(n883) );
  XOR2_X1 U973 ( .A(n883), .B(KEYINPUT48), .Z(n893) );
  NAND2_X1 U974 ( .A1(G103), .A2(n619), .ZN(n885) );
  NAND2_X1 U975 ( .A1(G139), .A2(n624), .ZN(n884) );
  NAND2_X1 U976 ( .A1(n885), .A2(n884), .ZN(n891) );
  NAND2_X1 U977 ( .A1(G115), .A2(n894), .ZN(n887) );
  NAND2_X1 U978 ( .A1(G127), .A2(n895), .ZN(n886) );
  NAND2_X1 U979 ( .A1(n887), .A2(n886), .ZN(n888) );
  XOR2_X1 U980 ( .A(KEYINPUT47), .B(n888), .Z(n889) );
  XNOR2_X1 U981 ( .A(KEYINPUT112), .B(n889), .ZN(n890) );
  NOR2_X1 U982 ( .A1(n891), .A2(n890), .ZN(n937) );
  XNOR2_X1 U983 ( .A(G164), .B(n937), .ZN(n892) );
  XNOR2_X1 U984 ( .A(n893), .B(n892), .ZN(n906) );
  NAND2_X1 U985 ( .A1(G118), .A2(n894), .ZN(n897) );
  NAND2_X1 U986 ( .A1(G130), .A2(n895), .ZN(n896) );
  NAND2_X1 U987 ( .A1(n897), .A2(n896), .ZN(n902) );
  NAND2_X1 U988 ( .A1(G106), .A2(n619), .ZN(n899) );
  NAND2_X1 U989 ( .A1(G142), .A2(n624), .ZN(n898) );
  NAND2_X1 U990 ( .A1(n899), .A2(n898), .ZN(n900) );
  XOR2_X1 U991 ( .A(n900), .B(KEYINPUT45), .Z(n901) );
  NOR2_X1 U992 ( .A1(n902), .A2(n901), .ZN(n904) );
  XNOR2_X1 U993 ( .A(n904), .B(n903), .ZN(n905) );
  XOR2_X1 U994 ( .A(n906), .B(n905), .Z(n908) );
  XNOR2_X1 U995 ( .A(G160), .B(n944), .ZN(n907) );
  XNOR2_X1 U996 ( .A(n908), .B(n907), .ZN(n909) );
  XOR2_X1 U997 ( .A(G162), .B(n909), .Z(n910) );
  XNOR2_X1 U998 ( .A(n911), .B(n910), .ZN(n912) );
  NOR2_X1 U999 ( .A1(G37), .A2(n912), .ZN(G395) );
  XOR2_X1 U1000 ( .A(KEYINPUT115), .B(n913), .Z(n915) );
  XNOR2_X1 U1001 ( .A(G171), .B(n991), .ZN(n914) );
  XNOR2_X1 U1002 ( .A(n915), .B(n914), .ZN(n916) );
  XOR2_X1 U1003 ( .A(n916), .B(G286), .Z(n917) );
  NOR2_X1 U1004 ( .A1(G37), .A2(n917), .ZN(G397) );
  NOR2_X1 U1005 ( .A1(G229), .A2(G227), .ZN(n919) );
  XNOR2_X1 U1006 ( .A(KEYINPUT49), .B(KEYINPUT116), .ZN(n918) );
  XNOR2_X1 U1007 ( .A(n919), .B(n918), .ZN(n931) );
  XOR2_X1 U1008 ( .A(G2443), .B(G2451), .Z(n921) );
  XNOR2_X1 U1009 ( .A(G2446), .B(G2454), .ZN(n920) );
  XNOR2_X1 U1010 ( .A(n921), .B(n920), .ZN(n922) );
  XOR2_X1 U1011 ( .A(n922), .B(G2427), .Z(n924) );
  XNOR2_X1 U1012 ( .A(G1341), .B(G1348), .ZN(n923) );
  XNOR2_X1 U1013 ( .A(n924), .B(n923), .ZN(n928) );
  XOR2_X1 U1014 ( .A(G2435), .B(KEYINPUT104), .Z(n926) );
  XNOR2_X1 U1015 ( .A(G2430), .B(G2438), .ZN(n925) );
  XNOR2_X1 U1016 ( .A(n926), .B(n925), .ZN(n927) );
  XOR2_X1 U1017 ( .A(n928), .B(n927), .Z(n929) );
  NAND2_X1 U1018 ( .A1(G14), .A2(n929), .ZN(n936) );
  NAND2_X1 U1019 ( .A1(G319), .A2(n936), .ZN(n930) );
  NOR2_X1 U1020 ( .A1(n931), .A2(n930), .ZN(n933) );
  NOR2_X1 U1021 ( .A1(G395), .A2(G397), .ZN(n932) );
  NAND2_X1 U1022 ( .A1(n933), .A2(n932), .ZN(G225) );
  XNOR2_X1 U1023 ( .A(KEYINPUT117), .B(G225), .ZN(G308) );
  INV_X1 U1025 ( .A(G132), .ZN(G219) );
  INV_X1 U1026 ( .A(G120), .ZN(G236) );
  INV_X1 U1027 ( .A(G96), .ZN(G221) );
  INV_X1 U1028 ( .A(G82), .ZN(G220) );
  INV_X1 U1029 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1030 ( .A1(n935), .A2(n934), .ZN(G325) );
  INV_X1 U1031 ( .A(G325), .ZN(G261) );
  INV_X1 U1032 ( .A(G108), .ZN(G238) );
  INV_X1 U1033 ( .A(n936), .ZN(G401) );
  XOR2_X1 U1034 ( .A(G2072), .B(n937), .Z(n939) );
  XOR2_X1 U1035 ( .A(G164), .B(G2078), .Z(n938) );
  NOR2_X1 U1036 ( .A1(n939), .A2(n938), .ZN(n940) );
  XOR2_X1 U1037 ( .A(KEYINPUT50), .B(n940), .Z(n941) );
  NOR2_X1 U1038 ( .A1(n942), .A2(n941), .ZN(n950) );
  XOR2_X1 U1039 ( .A(G2084), .B(G160), .Z(n943) );
  NOR2_X1 U1040 ( .A1(n944), .A2(n943), .ZN(n946) );
  NAND2_X1 U1041 ( .A1(n946), .A2(n945), .ZN(n947) );
  NOR2_X1 U1042 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1043 ( .A1(n950), .A2(n949), .ZN(n958) );
  XOR2_X1 U1044 ( .A(G2090), .B(G162), .Z(n951) );
  NOR2_X1 U1045 ( .A1(n952), .A2(n951), .ZN(n953) );
  XOR2_X1 U1046 ( .A(KEYINPUT51), .B(n953), .Z(n954) );
  XNOR2_X1 U1047 ( .A(n954), .B(KEYINPUT118), .ZN(n956) );
  NAND2_X1 U1048 ( .A1(n956), .A2(n955), .ZN(n957) );
  NOR2_X1 U1049 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1050 ( .A(KEYINPUT52), .B(n959), .ZN(n961) );
  INV_X1 U1051 ( .A(KEYINPUT55), .ZN(n960) );
  NAND2_X1 U1052 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1053 ( .A1(n962), .A2(G29), .ZN(n987) );
  XNOR2_X1 U1054 ( .A(G29), .B(KEYINPUT121), .ZN(n983) );
  XNOR2_X1 U1055 ( .A(KEYINPUT120), .B(KEYINPUT53), .ZN(n975) );
  XNOR2_X1 U1056 ( .A(G27), .B(n963), .ZN(n970) );
  XNOR2_X1 U1057 ( .A(G1991), .B(G25), .ZN(n968) );
  XNOR2_X1 U1058 ( .A(G2067), .B(G26), .ZN(n965) );
  XNOR2_X1 U1059 ( .A(G2072), .B(G33), .ZN(n964) );
  NOR2_X1 U1060 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1061 ( .A(KEYINPUT119), .B(n966), .ZN(n967) );
  NOR2_X1 U1062 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1063 ( .A1(n970), .A2(n969), .ZN(n973) );
  XOR2_X1 U1064 ( .A(G1996), .B(G32), .Z(n971) );
  NAND2_X1 U1065 ( .A1(G28), .A2(n971), .ZN(n972) );
  NOR2_X1 U1066 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1067 ( .A(n975), .B(n974), .ZN(n980) );
  XOR2_X1 U1068 ( .A(G2090), .B(G35), .Z(n978) );
  XOR2_X1 U1069 ( .A(G34), .B(KEYINPUT54), .Z(n976) );
  XNOR2_X1 U1070 ( .A(n976), .B(G2084), .ZN(n977) );
  NAND2_X1 U1071 ( .A1(n978), .A2(n977), .ZN(n979) );
  NOR2_X1 U1072 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1073 ( .A(KEYINPUT55), .B(n981), .ZN(n982) );
  NAND2_X1 U1074 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1075 ( .A1(n984), .A2(G11), .ZN(n985) );
  XOR2_X1 U1076 ( .A(KEYINPUT122), .B(n985), .Z(n986) );
  NAND2_X1 U1077 ( .A1(n987), .A2(n986), .ZN(n1042) );
  XNOR2_X1 U1078 ( .A(G16), .B(KEYINPUT56), .ZN(n1012) );
  XNOR2_X1 U1079 ( .A(G1966), .B(G168), .ZN(n989) );
  NAND2_X1 U1080 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1081 ( .A(n990), .B(KEYINPUT57), .ZN(n1010) );
  XNOR2_X1 U1082 ( .A(n991), .B(G1348), .ZN(n996) );
  XNOR2_X1 U1083 ( .A(G301), .B(G1961), .ZN(n994) );
  XNOR2_X1 U1084 ( .A(n992), .B(G1341), .ZN(n993) );
  NOR2_X1 U1085 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1086 ( .A1(n996), .A2(n995), .ZN(n1008) );
  XNOR2_X1 U1087 ( .A(G1971), .B(KEYINPUT123), .ZN(n997) );
  XNOR2_X1 U1088 ( .A(n997), .B(G303), .ZN(n1001) );
  XNOR2_X1 U1089 ( .A(G1956), .B(G299), .ZN(n998) );
  NOR2_X1 U1090 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1091 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NOR2_X1 U1092 ( .A1(n1003), .A2(n1002), .ZN(n1005) );
  NAND2_X1 U1093 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1094 ( .A(KEYINPUT124), .B(n1006), .ZN(n1007) );
  NOR2_X1 U1095 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1096 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1097 ( .A1(n1012), .A2(n1011), .ZN(n1040) );
  INV_X1 U1098 ( .A(G16), .ZN(n1038) );
  XNOR2_X1 U1099 ( .A(G5), .B(n1013), .ZN(n1028) );
  XNOR2_X1 U1100 ( .A(KEYINPUT59), .B(G1348), .ZN(n1014) );
  XNOR2_X1 U1101 ( .A(n1014), .B(G4), .ZN(n1022) );
  XOR2_X1 U1102 ( .A(G1341), .B(G19), .Z(n1015) );
  XNOR2_X1 U1103 ( .A(KEYINPUT125), .B(n1015), .ZN(n1017) );
  XNOR2_X1 U1104 ( .A(G6), .B(G1981), .ZN(n1016) );
  NOR2_X1 U1105 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XOR2_X1 U1106 ( .A(KEYINPUT126), .B(n1018), .Z(n1020) );
  XNOR2_X1 U1107 ( .A(G1956), .B(G20), .ZN(n1019) );
  NOR2_X1 U1108 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1109 ( .A1(n1022), .A2(n1021), .ZN(n1024) );
  XOR2_X1 U1110 ( .A(KEYINPUT60), .B(KEYINPUT127), .Z(n1023) );
  XNOR2_X1 U1111 ( .A(n1024), .B(n1023), .ZN(n1026) );
  XNOR2_X1 U1112 ( .A(G1966), .B(G21), .ZN(n1025) );
  NOR2_X1 U1113 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1114 ( .A1(n1028), .A2(n1027), .ZN(n1035) );
  XNOR2_X1 U1115 ( .A(G1986), .B(G24), .ZN(n1030) );
  XNOR2_X1 U1116 ( .A(G1971), .B(G22), .ZN(n1029) );
  NOR2_X1 U1117 ( .A1(n1030), .A2(n1029), .ZN(n1032) );
  XOR2_X1 U1118 ( .A(G1976), .B(G23), .Z(n1031) );
  NAND2_X1 U1119 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  XNOR2_X1 U1120 ( .A(KEYINPUT58), .B(n1033), .ZN(n1034) );
  NOR2_X1 U1121 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  XNOR2_X1 U1122 ( .A(KEYINPUT61), .B(n1036), .ZN(n1037) );
  NAND2_X1 U1123 ( .A1(n1038), .A2(n1037), .ZN(n1039) );
  NAND2_X1 U1124 ( .A1(n1040), .A2(n1039), .ZN(n1041) );
  NOR2_X1 U1125 ( .A1(n1042), .A2(n1041), .ZN(n1043) );
  XNOR2_X1 U1126 ( .A(KEYINPUT62), .B(n1043), .ZN(G311) );
  INV_X1 U1127 ( .A(G311), .ZN(G150) );
endmodule

