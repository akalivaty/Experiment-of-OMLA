//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 1 1 1 0 1 0 1 1 1 0 1 0 1 1 0 0 1 0 1 1 0 1 1 0 1 1 1 0 1 0 1 0 0 1 0 1 0 1 1 0 1 0 0 0 1 1 1 0 1 0 0 0 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:39 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n600, new_n602,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n611, new_n612, new_n613, new_n614, new_n615, new_n616, new_n617,
    new_n618, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n724, new_n725, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n768, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020;
  NAND2_X1  g000(.A1(G234), .A2(G237), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n187), .A2(G952), .A3(new_n188), .ZN(new_n189));
  XOR2_X1   g003(.A(KEYINPUT21), .B(G898), .Z(new_n190));
  NAND3_X1  g004(.A1(new_n187), .A2(G902), .A3(G953), .ZN(new_n191));
  OAI21_X1  g005(.A(new_n189), .B1(new_n190), .B2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  OAI21_X1  g007(.A(G214), .B1(G237), .B2(G902), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G104), .ZN(new_n196));
  OAI21_X1  g010(.A(KEYINPUT3), .B1(new_n196), .B2(G107), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT3), .ZN(new_n198));
  INV_X1    g012(.A(G107), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n198), .A2(new_n199), .A3(G104), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n196), .A2(G107), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n197), .A2(new_n200), .A3(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(KEYINPUT78), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT78), .ZN(new_n204));
  NAND4_X1  g018(.A1(new_n197), .A2(new_n200), .A3(new_n204), .A4(new_n201), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n203), .A2(G101), .A3(new_n205), .ZN(new_n206));
  XNOR2_X1  g020(.A(KEYINPUT79), .B(G101), .ZN(new_n207));
  OAI21_X1  g021(.A(KEYINPUT4), .B1(new_n202), .B2(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  NAND4_X1  g023(.A1(new_n203), .A2(KEYINPUT4), .A3(G101), .A4(new_n205), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  XNOR2_X1  g025(.A(G116), .B(G119), .ZN(new_n212));
  XNOR2_X1  g026(.A(KEYINPUT2), .B(G113), .ZN(new_n213));
  XNOR2_X1  g027(.A(new_n212), .B(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n211), .A2(new_n215), .ZN(new_n216));
  AND3_X1   g030(.A1(new_n197), .A2(new_n200), .A3(new_n201), .ZN(new_n217));
  XOR2_X1   g031(.A(KEYINPUT79), .B(G101), .Z(new_n218));
  NAND2_X1  g032(.A1(new_n199), .A2(G104), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n201), .A2(new_n219), .ZN(new_n220));
  AOI22_X1  g034(.A1(new_n217), .A2(new_n218), .B1(G101), .B2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(new_n212), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n222), .A2(new_n213), .ZN(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(G119), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(G116), .ZN(new_n226));
  INV_X1    g040(.A(G116), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(G119), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n226), .A2(new_n228), .A3(KEYINPUT5), .ZN(new_n229));
  OR3_X1    g043(.A1(new_n227), .A2(KEYINPUT5), .A3(G119), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n229), .A2(new_n230), .A3(G113), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(KEYINPUT81), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT81), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n229), .A2(new_n230), .A3(new_n234), .A4(G113), .ZN(new_n235));
  INV_X1    g049(.A(new_n235), .ZN(new_n236));
  OAI211_X1 g050(.A(new_n221), .B(new_n224), .C1(new_n233), .C2(new_n236), .ZN(new_n237));
  XNOR2_X1  g051(.A(G110), .B(G122), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n216), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(new_n238), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n214), .B1(new_n209), .B2(new_n210), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n199), .A2(G104), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n196), .A2(G107), .ZN(new_n243));
  OAI21_X1  g057(.A(G101), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n244), .B1(new_n202), .B2(new_n207), .ZN(new_n245));
  AOI211_X1 g059(.A(new_n223), .B(new_n245), .C1(new_n235), .C2(new_n232), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n240), .B1(new_n241), .B2(new_n246), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n239), .A2(KEYINPUT6), .A3(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT6), .ZN(new_n249));
  OAI211_X1 g063(.A(new_n249), .B(new_n240), .C1(new_n241), .C2(new_n246), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(KEYINPUT82), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT82), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n248), .A2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT64), .ZN(new_n255));
  INV_X1    g069(.A(G143), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n255), .B1(new_n256), .B2(G146), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(G146), .ZN(new_n258));
  INV_X1    g072(.A(G146), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n259), .A2(KEYINPUT64), .A3(G143), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n257), .A2(new_n258), .A3(new_n260), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n256), .A2(G146), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT1), .ZN(new_n263));
  OAI21_X1  g077(.A(G128), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n261), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n259), .A2(G143), .ZN(new_n266));
  NAND4_X1  g080(.A1(new_n266), .A2(new_n258), .A3(new_n263), .A4(G128), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  AND2_X1   g082(.A1(KEYINPUT0), .A2(G128), .ZN(new_n269));
  NOR2_X1   g083(.A1(KEYINPUT0), .A2(G128), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n261), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g086(.A(G143), .B(G146), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(new_n269), .ZN(new_n274));
  AND2_X1   g088(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  MUX2_X1   g089(.A(new_n268), .B(new_n275), .S(G125), .Z(new_n276));
  NAND2_X1  g090(.A1(new_n188), .A2(G224), .ZN(new_n277));
  XNOR2_X1  g091(.A(new_n276), .B(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n252), .A2(new_n254), .A3(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n277), .A2(KEYINPUT7), .ZN(new_n280));
  XNOR2_X1  g094(.A(new_n276), .B(new_n280), .ZN(new_n281));
  XNOR2_X1  g095(.A(new_n238), .B(KEYINPUT8), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n224), .A2(new_n231), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(new_n221), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n224), .B1(new_n233), .B2(new_n236), .ZN(new_n285));
  OAI211_X1 g099(.A(new_n282), .B(new_n284), .C1(new_n285), .C2(new_n221), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n281), .A2(new_n239), .A3(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(G902), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n287), .A2(KEYINPUT83), .A3(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n287), .A2(new_n288), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT83), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n279), .A2(new_n289), .A3(new_n292), .ZN(new_n293));
  OAI21_X1  g107(.A(G210), .B1(G237), .B2(G902), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  NAND4_X1  g110(.A1(new_n279), .A2(new_n294), .A3(new_n292), .A4(new_n289), .ZN(new_n297));
  AOI211_X1 g111(.A(new_n193), .B(new_n195), .C1(new_n296), .C2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(G469), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n188), .A2(G227), .ZN(new_n300));
  XNOR2_X1  g114(.A(new_n300), .B(G140), .ZN(new_n301));
  XNOR2_X1  g115(.A(KEYINPUT77), .B(G110), .ZN(new_n302));
  XNOR2_X1  g116(.A(new_n301), .B(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT80), .ZN(new_n304));
  AND3_X1   g118(.A1(new_n266), .A2(new_n258), .A3(G128), .ZN(new_n305));
  AOI22_X1  g119(.A1(new_n263), .A2(new_n305), .B1(new_n261), .B2(new_n264), .ZN(new_n306));
  OAI21_X1  g120(.A(KEYINPUT10), .B1(new_n306), .B2(new_n245), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT10), .ZN(new_n308));
  INV_X1    g122(.A(G128), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n309), .B1(new_n266), .B2(KEYINPUT1), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n267), .B1(new_n310), .B2(new_n273), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n221), .A2(new_n308), .A3(new_n311), .ZN(new_n312));
  AOI22_X1  g126(.A1(new_n211), .A2(new_n275), .B1(new_n307), .B2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(G134), .ZN(new_n314));
  OAI21_X1  g128(.A(KEYINPUT65), .B1(new_n314), .B2(G137), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(KEYINPUT11), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n314), .A2(G137), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT11), .ZN(new_n318));
  OAI211_X1 g132(.A(KEYINPUT65), .B(new_n318), .C1(new_n314), .C2(G137), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n316), .A2(new_n317), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(G131), .ZN(new_n321));
  INV_X1    g135(.A(G131), .ZN(new_n322));
  NAND4_X1  g136(.A1(new_n316), .A2(new_n322), .A3(new_n317), .A4(new_n319), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n304), .B1(new_n313), .B2(new_n325), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n308), .B1(new_n221), .B2(new_n268), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n218), .A2(new_n201), .A3(new_n197), .A4(new_n200), .ZN(new_n328));
  AND4_X1   g142(.A1(new_n308), .A2(new_n328), .A3(new_n311), .A4(new_n244), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n272), .A2(new_n274), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n331), .B1(new_n209), .B2(new_n210), .ZN(new_n332));
  OAI211_X1 g146(.A(KEYINPUT80), .B(new_n324), .C1(new_n330), .C2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n326), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n211), .A2(new_n275), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n307), .A2(new_n312), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n335), .A2(new_n325), .A3(new_n336), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n303), .B1(new_n334), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n303), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n245), .A2(new_n265), .A3(new_n267), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n328), .A2(new_n311), .A3(new_n244), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(new_n324), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT12), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n342), .A2(KEYINPUT12), .A3(new_n324), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n339), .A2(new_n348), .ZN(new_n349));
  OAI211_X1 g163(.A(new_n299), .B(new_n288), .C1(new_n338), .C2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n303), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n351), .B1(new_n313), .B2(new_n325), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n334), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n303), .B1(new_n347), .B2(new_n337), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n353), .A2(G469), .A3(new_n355), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n299), .A2(new_n288), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n350), .A2(new_n356), .A3(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(G221), .ZN(new_n360));
  XOR2_X1   g174(.A(KEYINPUT9), .B(G234), .Z(new_n361));
  AOI21_X1  g175(.A(new_n360), .B1(new_n361), .B2(new_n288), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n359), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT23), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n366), .B1(new_n225), .B2(G128), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n309), .A2(KEYINPUT23), .A3(G119), .ZN(new_n368));
  AND2_X1   g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT72), .ZN(new_n370));
  INV_X1    g184(.A(G110), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n225), .A2(G128), .ZN(new_n372));
  NAND4_X1  g186(.A1(new_n369), .A2(new_n370), .A3(new_n371), .A4(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n309), .A2(G119), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(new_n372), .ZN(new_n375));
  XNOR2_X1  g189(.A(KEYINPUT24), .B(G110), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n367), .A2(new_n372), .A3(new_n368), .ZN(new_n378));
  OAI21_X1  g192(.A(KEYINPUT72), .B1(new_n378), .B2(G110), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n373), .A2(new_n377), .A3(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT70), .ZN(new_n381));
  INV_X1    g195(.A(G140), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(G125), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n381), .B1(new_n383), .B2(KEYINPUT16), .ZN(new_n384));
  INV_X1    g198(.A(G125), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(G140), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n383), .A2(new_n386), .A3(KEYINPUT16), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT16), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n388), .A2(new_n382), .A3(KEYINPUT70), .A4(G125), .ZN(new_n389));
  NAND4_X1  g203(.A1(new_n384), .A2(new_n387), .A3(G146), .A4(new_n389), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n383), .A2(new_n386), .A3(new_n259), .ZN(new_n391));
  XNOR2_X1  g205(.A(new_n391), .B(KEYINPUT73), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n380), .A2(new_n390), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(KEYINPUT74), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n384), .A2(new_n387), .A3(new_n389), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(new_n259), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n396), .A2(KEYINPUT71), .A3(new_n390), .ZN(new_n397));
  OR2_X1    g211(.A1(new_n375), .A2(new_n376), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT71), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n395), .A2(new_n399), .A3(new_n259), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n378), .A2(G110), .ZN(new_n401));
  NAND4_X1  g215(.A1(new_n397), .A2(new_n398), .A3(new_n400), .A4(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT74), .ZN(new_n403));
  NAND4_X1  g217(.A1(new_n380), .A2(new_n403), .A3(new_n390), .A4(new_n392), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n394), .A2(new_n402), .A3(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n406));
  XNOR2_X1  g220(.A(new_n406), .B(G137), .ZN(new_n407));
  XNOR2_X1  g221(.A(KEYINPUT75), .B(KEYINPUT22), .ZN(new_n408));
  XNOR2_X1  g222(.A(new_n407), .B(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n405), .A2(new_n410), .ZN(new_n411));
  NAND4_X1  g225(.A1(new_n394), .A2(new_n402), .A3(new_n404), .A4(new_n409), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n411), .A2(new_n288), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(KEYINPUT76), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT25), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  XNOR2_X1  g230(.A(KEYINPUT68), .B(G217), .ZN(new_n417));
  INV_X1    g231(.A(G234), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n417), .B1(new_n418), .B2(G902), .ZN(new_n419));
  XNOR2_X1  g233(.A(new_n419), .B(KEYINPUT69), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n413), .A2(KEYINPUT76), .A3(KEYINPUT25), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n416), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  AND2_X1   g237(.A1(new_n411), .A2(new_n412), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n421), .A2(G902), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n423), .A2(new_n426), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n331), .B1(new_n321), .B2(new_n323), .ZN(new_n428));
  INV_X1    g242(.A(new_n317), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n314), .A2(G137), .ZN(new_n430));
  OAI21_X1  g244(.A(G131), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n323), .A2(new_n431), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n432), .A2(new_n306), .ZN(new_n433));
  NOR3_X1   g247(.A1(new_n428), .A2(new_n433), .A3(KEYINPUT30), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT30), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n324), .A2(new_n275), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n268), .A2(new_n323), .A3(new_n431), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n435), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n215), .B1(new_n434), .B2(new_n438), .ZN(new_n439));
  NOR3_X1   g253(.A1(new_n428), .A2(new_n433), .A3(new_n215), .ZN(new_n440));
  NOR2_X1   g254(.A1(G237), .A2(G953), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(G210), .ZN(new_n442));
  XNOR2_X1  g256(.A(new_n442), .B(G101), .ZN(new_n443));
  XNOR2_X1  g257(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n444));
  XNOR2_X1  g258(.A(new_n443), .B(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(KEYINPUT66), .B1(new_n440), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n436), .A2(new_n214), .A3(new_n437), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT66), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n448), .A2(new_n449), .A3(new_n445), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n439), .A2(new_n447), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(KEYINPUT31), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT31), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n439), .A2(new_n447), .A3(new_n453), .A4(new_n450), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n214), .B1(new_n436), .B2(new_n437), .ZN(new_n455));
  OAI21_X1  g269(.A(KEYINPUT28), .B1(new_n440), .B2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT28), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n448), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(new_n446), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n452), .A2(new_n454), .A3(new_n460), .ZN(new_n461));
  NOR2_X1   g275(.A1(G472), .A2(G902), .ZN(new_n462));
  AND3_X1   g276(.A1(new_n461), .A2(KEYINPUT32), .A3(new_n462), .ZN(new_n463));
  AOI21_X1  g277(.A(KEYINPUT32), .B1(new_n461), .B2(new_n462), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND4_X1  g279(.A1(new_n456), .A2(KEYINPUT29), .A3(new_n445), .A4(new_n458), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(new_n288), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT67), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n456), .A2(new_n445), .A3(new_n458), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT29), .ZN(new_n471));
  OAI21_X1  g285(.A(KEYINPUT30), .B1(new_n428), .B2(new_n433), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n436), .A2(new_n435), .A3(new_n437), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n214), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n474), .A2(new_n440), .ZN(new_n475));
  OAI211_X1 g289(.A(new_n470), .B(new_n471), .C1(new_n445), .C2(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n466), .A2(KEYINPUT67), .A3(new_n288), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n469), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(G472), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n427), .B1(new_n465), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n383), .A2(new_n386), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(KEYINPUT19), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT19), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n383), .A2(new_n386), .A3(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n482), .A2(new_n259), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(new_n390), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(KEYINPUT85), .ZN(new_n487));
  INV_X1    g301(.A(G237), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n488), .A2(new_n188), .A3(G214), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(new_n256), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n441), .A2(G143), .A3(G214), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n490), .A2(new_n322), .A3(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n322), .B1(new_n490), .B2(new_n491), .ZN(new_n494));
  OAI21_X1  g308(.A(KEYINPUT84), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT85), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n485), .A2(new_n496), .A3(new_n390), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n490), .A2(new_n491), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(G131), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT84), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n499), .A2(new_n500), .A3(new_n492), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n487), .A2(new_n495), .A3(new_n497), .A4(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n481), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n392), .B1(new_n259), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(KEYINPUT18), .A2(G131), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n490), .A2(new_n491), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n494), .A2(KEYINPUT18), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n504), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n502), .A2(new_n508), .ZN(new_n509));
  XNOR2_X1  g323(.A(G113), .B(G122), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n510), .B(new_n196), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n509), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n397), .A2(new_n400), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n494), .A2(KEYINPUT17), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT17), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n499), .A2(new_n516), .A3(new_n492), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(KEYINPUT86), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT86), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n499), .A2(new_n519), .A3(new_n516), .A4(new_n492), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n514), .A2(new_n515), .A3(new_n518), .A4(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n521), .A2(new_n511), .A3(new_n508), .ZN(new_n522));
  AOI21_X1  g336(.A(G475), .B1(new_n513), .B2(new_n522), .ZN(new_n523));
  AND3_X1   g337(.A1(new_n523), .A2(KEYINPUT20), .A3(new_n288), .ZN(new_n524));
  AOI21_X1  g338(.A(KEYINPUT20), .B1(new_n523), .B2(new_n288), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AND3_X1   g340(.A1(new_n521), .A2(new_n511), .A3(new_n508), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n511), .B1(new_n521), .B2(new_n508), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n288), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT87), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  OAI211_X1 g345(.A(KEYINPUT87), .B(new_n288), .C1(new_n527), .C2(new_n528), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n531), .A2(G475), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n526), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n361), .A2(new_n188), .A3(new_n417), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n227), .A2(KEYINPUT14), .A3(G122), .ZN(new_n537));
  XNOR2_X1  g351(.A(G116), .B(G122), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  OAI211_X1 g353(.A(G107), .B(new_n537), .C1(new_n539), .C2(KEYINPUT14), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n309), .A2(G143), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n541), .B(KEYINPUT88), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n309), .A2(G143), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n542), .A2(new_n314), .A3(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n314), .B1(new_n542), .B2(new_n544), .ZN(new_n547));
  OAI221_X1 g361(.A(new_n540), .B1(G107), .B2(new_n539), .C1(new_n546), .C2(new_n547), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n542), .B1(KEYINPUT13), .B2(new_n543), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n543), .A2(KEYINPUT13), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n550), .B(KEYINPUT89), .ZN(new_n551));
  OAI21_X1  g365(.A(G134), .B1(new_n549), .B2(new_n551), .ZN(new_n552));
  XNOR2_X1  g366(.A(new_n538), .B(new_n199), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n552), .A2(new_n545), .A3(new_n553), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n536), .B1(new_n548), .B2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n548), .A2(new_n554), .A3(new_n536), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(G478), .ZN(new_n559));
  OAI211_X1 g373(.A(new_n558), .B(new_n288), .C1(KEYINPUT15), .C2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  AOI211_X1 g375(.A(KEYINPUT15), .B(new_n559), .C1(new_n558), .C2(new_n288), .ZN(new_n562));
  OR2_X1    g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n534), .A2(new_n563), .ZN(new_n564));
  NAND4_X1  g378(.A1(new_n298), .A2(new_n365), .A3(new_n480), .A4(new_n564), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n565), .B(new_n207), .ZN(G3));
  NAND2_X1  g380(.A1(new_n461), .A2(new_n288), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(G472), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n461), .A2(new_n462), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT90), .ZN(new_n572));
  AND2_X1   g386(.A1(new_n423), .A2(new_n426), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n365), .A2(new_n571), .A3(new_n572), .A4(new_n573), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n359), .A2(new_n568), .A3(new_n363), .A4(new_n569), .ZN(new_n575));
  OAI21_X1  g389(.A(KEYINPUT90), .B1(new_n575), .B2(new_n427), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n577), .B(KEYINPUT91), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n195), .B1(new_n296), .B2(new_n297), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(new_n192), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT33), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n556), .A2(new_n581), .A3(new_n557), .ZN(new_n582));
  INV_X1    g396(.A(new_n557), .ZN(new_n583));
  OAI21_X1  g397(.A(KEYINPUT33), .B1(new_n583), .B2(new_n555), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n582), .A2(new_n584), .A3(G478), .ZN(new_n585));
  NAND2_X1  g399(.A1(G478), .A2(G902), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n558), .A2(new_n559), .A3(new_n288), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n588), .B1(new_n526), .B2(new_n533), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  NOR3_X1   g404(.A1(new_n578), .A2(new_n580), .A3(new_n590), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n591), .B(new_n196), .ZN(new_n592));
  XNOR2_X1  g406(.A(KEYINPUT92), .B(KEYINPUT34), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n592), .B(new_n593), .ZN(G6));
  INV_X1    g408(.A(new_n534), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(new_n563), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n298), .A2(new_n597), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n578), .A2(new_n598), .ZN(new_n599));
  XNOR2_X1  g413(.A(KEYINPUT35), .B(G107), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n599), .B(new_n600), .ZN(G9));
  NOR2_X1   g415(.A1(new_n410), .A2(KEYINPUT36), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n405), .B(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(new_n425), .ZN(new_n604));
  AND3_X1   g418(.A1(new_n423), .A2(KEYINPUT93), .A3(new_n604), .ZN(new_n605));
  AOI21_X1  g419(.A(KEYINPUT93), .B1(new_n423), .B2(new_n604), .ZN(new_n606));
  NOR3_X1   g420(.A1(new_n364), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n607), .A2(new_n298), .A3(new_n564), .A4(new_n571), .ZN(new_n608));
  XOR2_X1   g422(.A(KEYINPUT37), .B(G110), .Z(new_n609));
  XNOR2_X1  g423(.A(new_n608), .B(new_n609), .ZN(G12));
  OAI21_X1  g424(.A(new_n189), .B1(new_n191), .B2(G900), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n596), .A2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT32), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n569), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n461), .A2(KEYINPUT32), .A3(new_n462), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n479), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n607), .A2(new_n613), .A3(new_n617), .A4(new_n579), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(G128), .ZN(G30));
  XNOR2_X1  g433(.A(new_n611), .B(KEYINPUT39), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n365), .A2(new_n620), .ZN(new_n621));
  XOR2_X1   g435(.A(new_n621), .B(KEYINPUT40), .Z(new_n622));
  NOR2_X1   g436(.A1(new_n561), .A2(new_n562), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n623), .B1(new_n533), .B2(new_n526), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n296), .A2(new_n297), .ZN(new_n625));
  XNOR2_X1  g439(.A(KEYINPUT94), .B(KEYINPUT38), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT93), .ZN(new_n628));
  AND3_X1   g442(.A1(new_n413), .A2(KEYINPUT76), .A3(KEYINPUT25), .ZN(new_n629));
  AOI21_X1  g443(.A(KEYINPUT25), .B1(new_n413), .B2(KEYINPUT76), .ZN(new_n630));
  NOR3_X1   g444(.A1(new_n629), .A2(new_n630), .A3(new_n420), .ZN(new_n631));
  INV_X1    g445(.A(new_n604), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n628), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n423), .A2(KEYINPUT93), .A3(new_n604), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n446), .B1(new_n440), .B2(new_n455), .ZN(new_n636));
  AND2_X1   g450(.A1(new_n451), .A2(new_n636), .ZN(new_n637));
  OAI21_X1  g451(.A(G472), .B1(new_n637), .B2(G902), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n615), .A2(new_n616), .A3(new_n638), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n635), .A2(new_n194), .A3(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n622), .A2(new_n624), .A3(new_n627), .A4(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(G143), .ZN(G45));
  AND3_X1   g457(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n644));
  AND3_X1   g458(.A1(new_n531), .A2(G475), .A3(new_n532), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n523), .A2(new_n288), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT20), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n523), .A2(KEYINPUT20), .A3(new_n288), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  OAI211_X1 g464(.A(new_n644), .B(new_n611), .C1(new_n645), .C2(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n651), .A2(KEYINPUT95), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT95), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n653), .B1(new_n589), .B2(new_n611), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n655), .A2(new_n607), .A3(new_n617), .A4(new_n579), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(G146), .ZN(G48));
  AND3_X1   g471(.A1(new_n579), .A2(new_n192), .A3(new_n589), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n335), .A2(new_n336), .ZN(new_n659));
  AOI21_X1  g473(.A(KEYINPUT80), .B1(new_n659), .B2(new_n324), .ZN(new_n660));
  INV_X1    g474(.A(new_n333), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n337), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n349), .B1(new_n662), .B2(new_n351), .ZN(new_n663));
  OAI21_X1  g477(.A(G469), .B1(new_n663), .B2(G902), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT96), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n664), .A2(new_n665), .A3(new_n350), .ZN(new_n666));
  OAI211_X1 g480(.A(KEYINPUT96), .B(G469), .C1(new_n663), .C2(G902), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  AOI21_X1  g482(.A(KEYINPUT97), .B1(new_n668), .B2(new_n363), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT97), .ZN(new_n670));
  AOI211_X1 g484(.A(new_n670), .B(new_n362), .C1(new_n666), .C2(new_n667), .ZN(new_n671));
  OAI211_X1 g485(.A(new_n658), .B(new_n480), .C1(new_n669), .C2(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(KEYINPUT41), .B(G113), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G15));
  INV_X1    g488(.A(KEYINPUT98), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n480), .B1(new_n669), .B2(new_n671), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n675), .B1(new_n676), .B2(new_n598), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n350), .A2(new_n665), .ZN(new_n678));
  AOI22_X1  g492(.A1(new_n326), .A2(new_n333), .B1(new_n325), .B2(new_n313), .ZN(new_n679));
  OAI22_X1  g493(.A1(new_n679), .A2(new_n303), .B1(new_n348), .B2(new_n339), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n299), .B1(new_n680), .B2(new_n288), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(new_n667), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n363), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(new_n670), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n362), .B1(new_n666), .B2(new_n667), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(KEYINPUT97), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n580), .A2(new_n596), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n688), .A2(KEYINPUT98), .A3(new_n689), .A4(new_n480), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n677), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G116), .ZN(G18));
  NOR2_X1   g506(.A1(new_n684), .A2(new_n635), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n693), .A2(new_n617), .A3(new_n298), .A4(new_n564), .ZN(new_n694));
  XNOR2_X1  g508(.A(KEYINPUT99), .B(G119), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(G21));
  INV_X1    g510(.A(KEYINPUT100), .ZN(new_n697));
  AND3_X1   g511(.A1(new_n448), .A2(new_n449), .A3(new_n445), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n449), .B1(new_n448), .B2(new_n445), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n453), .B1(new_n700), .B2(new_n439), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n445), .B1(new_n456), .B2(new_n458), .ZN(new_n702));
  OAI21_X1  g516(.A(new_n697), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n452), .A2(KEYINPUT100), .A3(new_n460), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n703), .A2(new_n454), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(new_n462), .ZN(new_n706));
  AOI21_X1  g520(.A(KEYINPUT101), .B1(new_n567), .B2(G472), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT101), .ZN(new_n708));
  INV_X1    g522(.A(G472), .ZN(new_n709));
  AOI211_X1 g523(.A(new_n708), .B(new_n709), .C1(new_n461), .C2(new_n288), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n706), .B1(new_n707), .B2(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT102), .ZN(new_n712));
  NOR3_X1   g526(.A1(new_n711), .A2(new_n712), .A3(new_n427), .ZN(new_n713));
  AOI22_X1  g527(.A1(new_n451), .A2(KEYINPUT31), .B1(new_n459), .B2(new_n446), .ZN(new_n714));
  AOI21_X1  g528(.A(G902), .B1(new_n714), .B2(new_n454), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n708), .B1(new_n715), .B2(new_n709), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n567), .A2(KEYINPUT101), .A3(G472), .ZN(new_n717));
  AOI22_X1  g531(.A1(new_n716), .A2(new_n717), .B1(new_n462), .B2(new_n705), .ZN(new_n718));
  AOI21_X1  g532(.A(KEYINPUT102), .B1(new_n718), .B2(new_n573), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n298), .B1(new_n713), .B2(new_n719), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n624), .B1(new_n669), .B2(new_n671), .ZN(new_n721));
  OR2_X1    g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G122), .ZN(G24));
  AND2_X1   g537(.A1(new_n718), .A2(new_n579), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n693), .A2(new_n724), .A3(new_n655), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G125), .ZN(G27));
  XOR2_X1   g540(.A(KEYINPUT105), .B(KEYINPUT42), .Z(new_n727));
  INV_X1    g541(.A(KEYINPUT104), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n354), .B1(new_n334), .B2(new_n352), .ZN(new_n729));
  AOI21_X1  g543(.A(KEYINPUT103), .B1(new_n729), .B2(G469), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n339), .B1(new_n326), .B2(new_n333), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT103), .ZN(new_n732));
  NOR4_X1   g546(.A1(new_n731), .A2(new_n732), .A3(new_n299), .A4(new_n354), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n730), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n350), .A2(new_n358), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n728), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n356), .A2(new_n732), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n729), .A2(KEYINPUT103), .A3(G469), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n739), .A2(KEYINPUT104), .A3(new_n350), .A4(new_n358), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n736), .A2(new_n363), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n617), .A2(new_n573), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n296), .A2(new_n194), .A3(new_n297), .ZN(new_n743));
  NOR3_X1   g557(.A1(new_n741), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n727), .B1(new_n744), .B2(new_n655), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT106), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n615), .A2(new_n746), .ZN(new_n747));
  OAI211_X1 g561(.A(new_n479), .B(new_n747), .C1(new_n465), .C2(new_n746), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(new_n573), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n736), .A2(new_n740), .A3(KEYINPUT42), .A4(new_n363), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n651), .A2(KEYINPUT95), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n589), .A2(new_n653), .A3(new_n611), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NOR4_X1   g567(.A1(new_n749), .A2(new_n750), .A3(new_n753), .A4(new_n743), .ZN(new_n754));
  OAI21_X1  g568(.A(KEYINPUT107), .B1(new_n745), .B2(new_n754), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n742), .A2(new_n743), .ZN(new_n756));
  AND3_X1   g570(.A1(new_n736), .A2(new_n363), .A3(new_n740), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n756), .A2(new_n757), .A3(new_n655), .ZN(new_n758));
  INV_X1    g572(.A(new_n727), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n753), .A2(new_n743), .ZN(new_n761));
  INV_X1    g575(.A(new_n750), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n761), .A2(new_n762), .A3(new_n573), .A4(new_n748), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT107), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n760), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n755), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G131), .ZN(G33));
  NAND2_X1  g581(.A1(new_n744), .A2(new_n613), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G134), .ZN(G36));
  NAND2_X1  g583(.A1(new_n595), .A2(new_n644), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT43), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n595), .A2(KEYINPUT43), .A3(new_n644), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n605), .A2(new_n606), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n775), .A2(KEYINPUT110), .A3(new_n570), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT110), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n777), .B1(new_n635), .B2(new_n571), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n774), .A2(new_n776), .A3(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT44), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT108), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n353), .A2(new_n355), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT45), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n782), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n729), .A2(KEYINPUT108), .A3(KEYINPUT45), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n783), .A2(new_n784), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n787), .A2(G469), .A3(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n789), .A2(KEYINPUT46), .A3(new_n358), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n790), .A2(new_n350), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(KEYINPUT109), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT46), .ZN(new_n793));
  INV_X1    g607(.A(new_n789), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n793), .B1(new_n794), .B2(new_n357), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT109), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n790), .A2(new_n796), .A3(new_n350), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n792), .A2(new_n795), .A3(new_n797), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n781), .A2(new_n798), .A3(new_n363), .A4(new_n620), .ZN(new_n799));
  INV_X1    g613(.A(new_n743), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n800), .B1(new_n779), .B2(new_n780), .ZN(new_n801));
  OR2_X1    g615(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(G137), .ZN(G39));
  NAND2_X1  g617(.A1(new_n798), .A2(new_n363), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT47), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n798), .A2(KEYINPUT47), .A3(new_n363), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n617), .A2(new_n573), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n808), .A2(new_n761), .A3(new_n809), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(G140), .ZN(G42));
  AOI21_X1  g625(.A(new_n189), .B1(new_n772), .B2(new_n773), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n684), .A2(new_n743), .ZN(new_n813));
  AND4_X1   g627(.A1(new_n573), .A2(new_n812), .A3(new_n813), .A4(new_n748), .ZN(new_n814));
  XOR2_X1   g628(.A(new_n814), .B(KEYINPUT48), .Z(new_n815));
  NAND2_X1  g629(.A1(new_n668), .A2(new_n362), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n806), .A2(new_n807), .A3(new_n816), .ZN(new_n817));
  OR2_X1    g631(.A1(new_n713), .A2(new_n719), .ZN(new_n818));
  AND2_X1   g632(.A1(new_n818), .A2(new_n812), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n817), .A2(new_n800), .A3(new_n819), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n711), .A2(new_n635), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n812), .A2(new_n813), .A3(new_n821), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n427), .A2(new_n189), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n813), .A2(new_n465), .A3(new_n638), .A4(new_n823), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n824), .A2(new_n534), .A3(new_n644), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n627), .A2(new_n194), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n819), .A2(KEYINPUT50), .A3(new_n686), .A4(new_n826), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n818), .A2(new_n826), .A3(new_n686), .A4(new_n812), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT50), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n825), .B1(new_n827), .B2(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n820), .A2(new_n822), .A3(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT51), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n820), .A2(KEYINPUT51), .A3(new_n822), .A4(new_n831), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n819), .A2(new_n686), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(new_n579), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n837), .A2(KEYINPUT116), .ZN(new_n838));
  OR2_X1    g652(.A1(new_n824), .A2(new_n590), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT116), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n836), .A2(new_n840), .A3(new_n579), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n838), .A2(new_n839), .A3(new_n841), .ZN(new_n842));
  AND4_X1   g656(.A1(new_n815), .A2(new_n834), .A3(new_n835), .A4(new_n842), .ZN(new_n843));
  AND2_X1   g657(.A1(new_n677), .A2(new_n690), .ZN(new_n844));
  NOR3_X1   g658(.A1(new_n534), .A2(new_n563), .A3(new_n612), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n775), .A2(new_n365), .A3(new_n617), .A4(new_n845), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n775), .A2(new_n718), .A3(new_n752), .A4(new_n751), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n846), .B1(new_n847), .B2(new_n741), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(new_n800), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n608), .A2(new_n565), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n596), .A2(new_n590), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n574), .A2(new_n576), .A3(new_n298), .A4(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n849), .A2(new_n850), .A3(new_n852), .ZN(new_n853));
  OAI211_X1 g667(.A(new_n672), .B(new_n694), .C1(new_n720), .C2(new_n721), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n844), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(new_n768), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n856), .B1(new_n755), .B2(new_n765), .ZN(new_n857));
  AND3_X1   g671(.A1(new_n625), .A2(new_n194), .A3(new_n624), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n631), .A2(new_n632), .ZN(new_n859));
  AND3_X1   g673(.A1(new_n639), .A2(new_n859), .A3(new_n611), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n757), .A2(new_n858), .A3(new_n860), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n725), .A2(new_n656), .A3(new_n861), .A4(new_n618), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT52), .ZN(new_n863));
  XNOR2_X1  g677(.A(new_n862), .B(new_n863), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n855), .A2(KEYINPUT53), .A3(new_n857), .A4(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT114), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n760), .A2(new_n763), .A3(new_n764), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n764), .B1(new_n760), .B2(new_n763), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n768), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n821), .A2(new_n757), .A3(new_n655), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n743), .B1(new_n871), .B2(new_n846), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n852), .A2(new_n565), .A3(new_n608), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  AND2_X1   g688(.A1(new_n672), .A2(new_n694), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n874), .A2(new_n691), .A3(new_n722), .A4(new_n875), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n870), .A2(new_n876), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n877), .A2(KEYINPUT114), .A3(KEYINPUT53), .A4(new_n864), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT53), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n854), .B1(new_n677), .B2(new_n690), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n857), .A2(new_n880), .A3(new_n874), .ZN(new_n881));
  AND3_X1   g695(.A1(new_n725), .A2(new_n618), .A3(new_n656), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n882), .A2(KEYINPUT113), .A3(KEYINPUT52), .A4(new_n861), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n862), .A2(new_n863), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT113), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n885), .B1(new_n862), .B2(new_n863), .ZN(new_n886));
  AND3_X1   g700(.A1(new_n883), .A2(new_n884), .A3(new_n886), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n879), .B1(new_n881), .B2(new_n887), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n867), .A2(new_n878), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(KEYINPUT54), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n855), .A2(new_n857), .A3(new_n864), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n891), .A2(new_n879), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT54), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n883), .A2(new_n884), .A3(new_n886), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n879), .B1(new_n760), .B2(new_n763), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n894), .A2(new_n855), .A3(new_n768), .A4(new_n895), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n892), .A2(new_n893), .A3(new_n896), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n843), .A2(new_n890), .A3(KEYINPUT115), .A4(new_n897), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n898), .A2(G952), .A3(new_n188), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n627), .A2(new_n639), .ZN(new_n900));
  INV_X1    g714(.A(new_n770), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n668), .B(KEYINPUT49), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n573), .A2(new_n363), .A3(new_n194), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(KEYINPUT111), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n900), .A2(new_n901), .A3(new_n902), .A4(new_n904), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n905), .B(KEYINPUT112), .Z(new_n906));
  INV_X1    g720(.A(KEYINPUT115), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n843), .A2(new_n890), .A3(new_n907), .A4(new_n897), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(G953), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n899), .A2(new_n906), .A3(new_n909), .ZN(G75));
  AOI21_X1  g724(.A(new_n288), .B1(new_n892), .B2(new_n896), .ZN(new_n911));
  AOI21_X1  g725(.A(KEYINPUT56), .B1(new_n911), .B2(G210), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n252), .A2(new_n254), .ZN(new_n913));
  XOR2_X1   g727(.A(new_n913), .B(new_n278), .Z(new_n914));
  XNOR2_X1  g728(.A(new_n914), .B(KEYINPUT55), .ZN(new_n915));
  INV_X1    g729(.A(new_n915), .ZN(new_n916));
  AND2_X1   g730(.A1(new_n912), .A2(new_n916), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n912), .A2(new_n916), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n188), .A2(G952), .ZN(new_n919));
  NOR3_X1   g733(.A1(new_n917), .A2(new_n918), .A3(new_n919), .ZN(G51));
  NAND2_X1  g734(.A1(new_n892), .A2(new_n896), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(new_n893), .ZN(new_n922));
  XOR2_X1   g736(.A(new_n357), .B(KEYINPUT57), .Z(new_n923));
  OAI21_X1  g737(.A(new_n680), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n911), .A2(new_n794), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n919), .B1(new_n924), .B2(new_n925), .ZN(G54));
  NAND3_X1  g740(.A1(new_n911), .A2(KEYINPUT58), .A3(G475), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n513), .A2(new_n522), .ZN(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  AND2_X1   g743(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n927), .A2(new_n929), .ZN(new_n931));
  NOR3_X1   g745(.A1(new_n930), .A2(new_n931), .A3(new_n919), .ZN(G60));
  NAND2_X1  g746(.A1(new_n582), .A2(new_n584), .ZN(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n586), .B(KEYINPUT59), .Z(new_n935));
  OR2_X1    g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  OAI22_X1  g750(.A1(new_n922), .A2(new_n936), .B1(G952), .B2(new_n188), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n935), .B1(new_n890), .B2(new_n897), .ZN(new_n938));
  OAI21_X1  g752(.A(KEYINPUT117), .B1(new_n938), .B2(new_n933), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT117), .ZN(new_n940));
  AND3_X1   g754(.A1(new_n892), .A2(new_n893), .A3(new_n896), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n941), .B1(KEYINPUT54), .B2(new_n889), .ZN(new_n942));
  OAI211_X1 g756(.A(new_n940), .B(new_n934), .C1(new_n942), .C2(new_n935), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n937), .B1(new_n939), .B2(new_n943), .ZN(G63));
  NAND2_X1  g758(.A1(G217), .A2(G902), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n945), .B(KEYINPUT60), .Z(new_n946));
  AOI21_X1  g760(.A(new_n424), .B1(new_n921), .B2(new_n946), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n947), .A2(new_n919), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n921), .A2(new_n603), .A3(new_n946), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(KEYINPUT118), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT118), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n921), .A2(new_n951), .A3(new_n603), .A4(new_n946), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n948), .A2(new_n950), .A3(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT61), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n948), .A2(new_n950), .A3(KEYINPUT61), .A4(new_n952), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n955), .A2(new_n956), .ZN(G66));
  AOI21_X1  g771(.A(new_n188), .B1(new_n190), .B2(G224), .ZN(new_n958));
  NOR3_X1   g772(.A1(new_n844), .A2(new_n873), .A3(new_n854), .ZN(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n958), .B1(new_n960), .B2(new_n188), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n913), .B1(G898), .B2(new_n188), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n961), .B(new_n962), .Z(G69));
  NOR2_X1   g777(.A1(new_n434), .A2(new_n438), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n482), .A2(new_n484), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n965), .B(KEYINPUT119), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n964), .B(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT123), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n967), .B1(new_n968), .B2(G900), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n969), .B1(new_n968), .B2(G900), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n188), .B1(G227), .B2(G900), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(KEYINPUT124), .ZN(new_n973));
  INV_X1    g787(.A(new_n851), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n621), .B1(new_n974), .B2(KEYINPUT121), .ZN(new_n975));
  OAI211_X1 g789(.A(new_n975), .B(new_n756), .C1(KEYINPUT121), .C2(new_n974), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n976), .B1(new_n799), .B2(new_n801), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n977), .A2(KEYINPUT122), .ZN(new_n978));
  INV_X1    g792(.A(KEYINPUT122), .ZN(new_n979));
  OAI211_X1 g793(.A(new_n979), .B(new_n976), .C1(new_n799), .C2(new_n801), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n725), .A2(new_n618), .A3(new_n656), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT120), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND4_X1  g798(.A1(new_n725), .A2(new_n656), .A3(KEYINPUT120), .A4(new_n618), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n642), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  INV_X1    g800(.A(KEYINPUT62), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND4_X1  g802(.A1(new_n642), .A2(new_n984), .A3(KEYINPUT62), .A4(new_n985), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n981), .A2(new_n810), .A3(new_n990), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n991), .A2(new_n188), .A3(new_n967), .ZN(new_n992));
  INV_X1    g806(.A(new_n971), .ZN(new_n993));
  AND2_X1   g807(.A1(new_n810), .A2(new_n857), .ZN(new_n994));
  AND3_X1   g808(.A1(new_n858), .A2(new_n573), .A3(new_n748), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n798), .A2(new_n363), .A3(new_n620), .A4(new_n995), .ZN(new_n996));
  AND4_X1   g810(.A1(new_n802), .A2(new_n984), .A3(new_n985), .A4(new_n996), .ZN(new_n997));
  AND2_X1   g811(.A1(new_n994), .A2(new_n997), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n993), .B1(new_n998), .B2(G953), .ZN(new_n999));
  OAI211_X1 g813(.A(new_n973), .B(new_n992), .C1(new_n999), .C2(new_n967), .ZN(G72));
  NAND4_X1  g814(.A1(new_n981), .A2(new_n990), .A3(new_n810), .A4(new_n959), .ZN(new_n1001));
  XNOR2_X1  g815(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n1002));
  NAND2_X1  g816(.A1(G472), .A2(G902), .ZN(new_n1003));
  XNOR2_X1  g817(.A(new_n1002), .B(new_n1003), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1001), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g819(.A(new_n475), .ZN(new_n1006));
  NAND3_X1  g820(.A1(new_n1005), .A2(new_n445), .A3(new_n1006), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1007), .A2(KEYINPUT126), .ZN(new_n1008));
  INV_X1    g822(.A(KEYINPUT126), .ZN(new_n1009));
  NAND4_X1  g823(.A1(new_n1005), .A2(new_n1009), .A3(new_n445), .A4(new_n1006), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n451), .B1(new_n475), .B2(new_n445), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n889), .A2(new_n1012), .A3(new_n1004), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1013), .A2(KEYINPUT127), .ZN(new_n1014));
  INV_X1    g828(.A(KEYINPUT127), .ZN(new_n1015));
  NAND4_X1  g829(.A1(new_n889), .A2(new_n1015), .A3(new_n1012), .A4(new_n1004), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g831(.A1(new_n994), .A2(new_n959), .A3(new_n997), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n445), .B1(new_n1018), .B2(new_n1004), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n919), .B1(new_n1019), .B2(new_n475), .ZN(new_n1020));
  AND3_X1   g834(.A1(new_n1011), .A2(new_n1017), .A3(new_n1020), .ZN(G57));
endmodule


