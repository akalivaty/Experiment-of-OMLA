//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 1 0 1 0 1 1 1 1 0 1 0 0 0 0 1 0 1 1 1 1 1 0 0 1 1 0 0 1 0 1 1 1 0 1 1 0 1 0 0 1 0 1 0 0 0 0 0 0 0 0 0 0 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n715, new_n716, new_n717, new_n719, new_n720, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n805, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n894, new_n895, new_n896, new_n898,
    new_n899, new_n900, new_n901, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n993, new_n994, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1046, new_n1047, new_n1048;
  INV_X1    g000(.A(KEYINPUT90), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT89), .ZN(new_n203));
  INV_X1    g002(.A(G1gat), .ZN(new_n204));
  INV_X1    g003(.A(G22gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n205), .A2(G15gat), .ZN(new_n206));
  INV_X1    g005(.A(G15gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n207), .A2(G22gat), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n204), .B1(new_n206), .B2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n207), .A2(G22gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n205), .A2(G15gat), .ZN(new_n211));
  OAI21_X1  g010(.A(KEYINPUT16), .B1(KEYINPUT88), .B2(G1gat), .ZN(new_n212));
  AND2_X1   g011(.A1(KEYINPUT88), .A2(G1gat), .ZN(new_n213));
  OAI211_X1 g012(.A(new_n210), .B(new_n211), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(G8gat), .ZN(new_n215));
  AND3_X1   g014(.A1(new_n209), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  AOI21_X1  g015(.A(new_n215), .B1(new_n209), .B2(new_n214), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n203), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n209), .A2(new_n214), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(G8gat), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n209), .A2(new_n214), .A3(new_n215), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n220), .A2(KEYINPUT89), .A3(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n218), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT14), .ZN(new_n224));
  INV_X1    g023(.A(G29gat), .ZN(new_n225));
  INV_X1    g024(.A(G36gat), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  OAI21_X1  g026(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(G50gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(G43gat), .ZN(new_n231));
  INV_X1    g030(.A(G43gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(G50gat), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n231), .A2(new_n233), .A3(KEYINPUT15), .ZN(new_n234));
  NAND2_X1  g033(.A1(G29gat), .A2(G36gat), .ZN(new_n235));
  AND3_X1   g034(.A1(new_n229), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT15), .ZN(new_n237));
  OR2_X1    g036(.A1(KEYINPUT86), .A2(G43gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(KEYINPUT86), .A2(G43gat), .ZN(new_n239));
  AOI21_X1  g038(.A(G50gat), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT87), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n241), .B1(new_n230), .B2(G43gat), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n232), .A2(KEYINPUT87), .A3(G50gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n237), .B1(new_n240), .B2(new_n244), .ZN(new_n245));
  AND2_X1   g044(.A1(new_n236), .A2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT85), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n227), .A2(new_n247), .ZN(new_n248));
  NOR3_X1   g047(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(KEYINPUT85), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n228), .A2(KEYINPUT84), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT84), .ZN(new_n252));
  OAI211_X1 g051(.A(new_n252), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n253));
  NAND4_X1  g052(.A1(new_n248), .A2(new_n250), .A3(new_n251), .A4(new_n253), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n234), .B1(new_n254), .B2(new_n235), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n246), .A2(new_n255), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n202), .B1(new_n223), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n236), .A2(new_n245), .ZN(new_n258));
  INV_X1    g057(.A(new_n235), .ZN(new_n259));
  AND2_X1   g058(.A1(new_n248), .A2(new_n250), .ZN(new_n260));
  AND2_X1   g059(.A1(new_n251), .A2(new_n253), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n259), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n258), .B1(new_n262), .B2(new_n234), .ZN(new_n263));
  NAND4_X1  g062(.A1(new_n263), .A2(KEYINPUT90), .A3(new_n222), .A4(new_n218), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n220), .A2(new_n221), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT17), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n265), .B1(new_n263), .B2(new_n266), .ZN(new_n267));
  OAI211_X1 g066(.A(KEYINPUT17), .B(new_n258), .C1(new_n262), .C2(new_n234), .ZN(new_n268));
  AOI22_X1  g067(.A1(new_n257), .A2(new_n264), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(G229gat), .A2(G233gat), .ZN(new_n270));
  AOI21_X1  g069(.A(KEYINPUT18), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n257), .A2(new_n264), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n267), .A2(new_n268), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT18), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n274), .B1(G229gat), .B2(G233gat), .ZN(new_n275));
  AND3_X1   g074(.A1(new_n272), .A2(new_n273), .A3(new_n275), .ZN(new_n276));
  XOR2_X1   g075(.A(new_n270), .B(KEYINPUT13), .Z(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n223), .A2(new_n256), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n278), .B1(new_n272), .B2(new_n279), .ZN(new_n280));
  NOR3_X1   g079(.A1(new_n271), .A2(new_n276), .A3(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(G113gat), .B(G141gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(G169gat), .B(G197gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n282), .B(new_n283), .ZN(new_n284));
  XOR2_X1   g083(.A(KEYINPUT83), .B(KEYINPUT11), .Z(new_n285));
  XNOR2_X1  g084(.A(new_n284), .B(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n286), .B(KEYINPUT12), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT91), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n288), .B1(new_n271), .B2(new_n289), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n281), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n272), .A2(new_n270), .A3(new_n273), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(new_n274), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n287), .B1(new_n293), .B2(KEYINPUT91), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n272), .A2(new_n279), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(new_n277), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n269), .A2(new_n275), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n293), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n294), .A2(new_n298), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n291), .A2(new_n299), .ZN(new_n300));
  XNOR2_X1  g099(.A(G211gat), .B(G218gat), .ZN(new_n301));
  OR2_X1    g100(.A1(new_n301), .A2(KEYINPUT70), .ZN(new_n302));
  XNOR2_X1  g101(.A(G197gat), .B(G204gat), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT22), .ZN(new_n304));
  INV_X1    g103(.A(G211gat), .ZN(new_n305));
  INV_X1    g104(.A(G218gat), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n304), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n303), .A2(new_n307), .ZN(new_n308));
  XNOR2_X1  g107(.A(new_n302), .B(new_n308), .ZN(new_n309));
  XOR2_X1   g108(.A(KEYINPUT66), .B(G190gat), .Z(new_n310));
  OR2_X1    g109(.A1(KEYINPUT65), .A2(G183gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(KEYINPUT65), .A2(G183gat), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n311), .A2(KEYINPUT27), .A3(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT67), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(KEYINPUT27), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT27), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(KEYINPUT67), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n315), .A2(new_n317), .A3(G183gat), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT28), .ZN(new_n319));
  NAND4_X1  g118(.A1(new_n310), .A2(new_n313), .A3(new_n318), .A4(new_n319), .ZN(new_n320));
  XOR2_X1   g119(.A(KEYINPUT27), .B(G183gat), .Z(new_n321));
  XNOR2_X1  g120(.A(KEYINPUT66), .B(G190gat), .ZN(new_n322));
  OAI21_X1  g121(.A(KEYINPUT28), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NOR2_X1   g122(.A1(G169gat), .A2(G176gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(KEYINPUT26), .ZN(new_n325));
  NAND2_X1  g124(.A1(G183gat), .A2(G190gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(G169gat), .A2(G176gat), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT26), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n330), .A2(new_n324), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n327), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n320), .A2(new_n323), .A3(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT68), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  OAI211_X1 g134(.A(new_n325), .B(new_n326), .C1(new_n330), .C2(new_n324), .ZN(new_n336));
  XNOR2_X1  g135(.A(KEYINPUT27), .B(G183gat), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n310), .A2(new_n337), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n336), .B1(new_n338), .B2(KEYINPUT28), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n339), .A2(KEYINPUT68), .A3(new_n320), .ZN(new_n340));
  NOR2_X1   g139(.A1(G183gat), .A2(G190gat), .ZN(new_n341));
  XNOR2_X1  g140(.A(new_n341), .B(KEYINPUT64), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n326), .A2(KEYINPUT24), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT24), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n344), .A2(G183gat), .A3(G190gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n342), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n324), .A2(KEYINPUT23), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT23), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n349), .B1(G169gat), .B2(G176gat), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n348), .A2(new_n328), .A3(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n347), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT25), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n311), .A2(new_n312), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n346), .B1(new_n356), .B2(new_n322), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n357), .A2(new_n352), .A3(KEYINPUT25), .ZN(new_n358));
  AOI22_X1  g157(.A1(new_n335), .A2(new_n340), .B1(new_n355), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(G226gat), .A2(G233gat), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n351), .B1(new_n342), .B2(new_n346), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n358), .B1(new_n363), .B2(KEYINPUT25), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(new_n333), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT29), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n365), .A2(new_n366), .A3(new_n360), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n309), .B1(new_n362), .B2(new_n367), .ZN(new_n368));
  OAI211_X1 g167(.A(KEYINPUT71), .B(new_n360), .C1(new_n359), .C2(KEYINPUT29), .ZN(new_n369));
  AOI21_X1  g168(.A(KEYINPUT68), .B1(new_n339), .B2(new_n320), .ZN(new_n370));
  AND4_X1   g169(.A1(KEYINPUT68), .A2(new_n320), .A3(new_n323), .A4(new_n332), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n364), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n361), .B1(new_n372), .B2(new_n366), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT71), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n374), .B1(new_n365), .B2(new_n361), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n369), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n368), .B1(new_n376), .B2(new_n309), .ZN(new_n377));
  XNOR2_X1  g176(.A(G8gat), .B(G36gat), .ZN(new_n378));
  XNOR2_X1  g177(.A(G64gat), .B(G92gat), .ZN(new_n379));
  XOR2_X1   g178(.A(new_n378), .B(new_n379), .Z(new_n380));
  NAND2_X1  g179(.A1(new_n377), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(new_n380), .ZN(new_n382));
  INV_X1    g181(.A(new_n309), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n360), .B1(new_n359), .B2(KEYINPUT29), .ZN(new_n384));
  INV_X1    g183(.A(new_n375), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n383), .B1(new_n386), .B2(new_n369), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n382), .B1(new_n387), .B2(new_n368), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n381), .A2(new_n388), .A3(KEYINPUT30), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT30), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n377), .A2(new_n390), .A3(new_n380), .ZN(new_n391));
  AND2_X1   g190(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  XNOR2_X1  g192(.A(G127gat), .B(G134gat), .ZN(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  XNOR2_X1  g194(.A(G113gat), .B(G120gat), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n395), .B1(KEYINPUT1), .B2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(new_n396), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT1), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n398), .A2(new_n399), .A3(new_n394), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n397), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n372), .A2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(G227gat), .ZN(new_n403));
  INV_X1    g202(.A(G233gat), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n401), .ZN(new_n407));
  OAI211_X1 g206(.A(new_n364), .B(new_n407), .C1(new_n370), .C2(new_n371), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n402), .A2(new_n406), .A3(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT69), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  XOR2_X1   g211(.A(G15gat), .B(G43gat), .Z(new_n413));
  XNOR2_X1  g212(.A(G71gat), .B(G99gat), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n413), .B(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n406), .B1(new_n402), .B2(new_n408), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n415), .B1(new_n416), .B2(KEYINPUT33), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT32), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n402), .A2(new_n408), .ZN(new_n421));
  AOI221_X4 g220(.A(new_n418), .B1(KEYINPUT33), .B2(new_n415), .C1(new_n421), .C2(new_n405), .ZN(new_n422));
  AOI21_X1  g221(.A(KEYINPUT34), .B1(new_n409), .B2(new_n410), .ZN(new_n423));
  NOR3_X1   g222(.A1(new_n420), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n423), .ZN(new_n425));
  INV_X1    g224(.A(new_n408), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n335), .A2(new_n340), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n407), .B1(new_n427), .B2(new_n364), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n405), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(KEYINPUT32), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT33), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n430), .A2(new_n432), .A3(new_n415), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n419), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n425), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n412), .B1(new_n424), .B2(new_n435), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n423), .B1(new_n420), .B2(new_n422), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n433), .A2(new_n434), .A3(new_n425), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n437), .A2(new_n411), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n436), .A2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT81), .ZN(new_n441));
  INV_X1    g240(.A(G155gat), .ZN(new_n442));
  INV_X1    g241(.A(G162gat), .ZN(new_n443));
  OAI21_X1  g242(.A(KEYINPUT2), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT74), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  XNOR2_X1  g245(.A(G155gat), .B(G162gat), .ZN(new_n447));
  OAI211_X1 g246(.A(KEYINPUT74), .B(KEYINPUT2), .C1(new_n442), .C2(new_n443), .ZN(new_n448));
  AND3_X1   g247(.A1(new_n446), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(G148gat), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(G141gat), .ZN(new_n451));
  XNOR2_X1  g250(.A(KEYINPUT73), .B(G141gat), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n451), .B1(new_n452), .B2(new_n450), .ZN(new_n453));
  INV_X1    g252(.A(new_n447), .ZN(new_n454));
  XNOR2_X1  g253(.A(KEYINPUT72), .B(KEYINPUT2), .ZN(new_n455));
  INV_X1    g254(.A(new_n451), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n450), .A2(G141gat), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n455), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  AOI22_X1  g257(.A1(new_n449), .A2(new_n453), .B1(new_n454), .B2(new_n458), .ZN(new_n459));
  XOR2_X1   g258(.A(KEYINPUT76), .B(KEYINPUT3), .Z(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(new_n366), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(new_n309), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n458), .A2(new_n454), .ZN(new_n464));
  XOR2_X1   g263(.A(KEYINPUT73), .B(G141gat), .Z(new_n465));
  AOI21_X1  g264(.A(new_n456), .B1(new_n465), .B2(G148gat), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n446), .A2(new_n447), .A3(new_n448), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n464), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT75), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  OAI211_X1 g269(.A(new_n464), .B(KEYINPUT75), .C1(new_n466), .C2(new_n467), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n309), .A2(KEYINPUT29), .ZN(new_n472));
  OAI211_X1 g271(.A(new_n470), .B(new_n471), .C1(new_n472), .C2(KEYINPUT3), .ZN(new_n473));
  AND4_X1   g272(.A1(G228gat), .A2(new_n463), .A3(new_n473), .A4(G233gat), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT80), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n308), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(KEYINPUT80), .B1(new_n303), .B2(new_n307), .ZN(new_n477));
  NOR3_X1   g276(.A1(new_n476), .A2(new_n301), .A3(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n308), .A2(new_n475), .A3(new_n301), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(new_n366), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n460), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(new_n468), .ZN(new_n482));
  AOI22_X1  g281(.A1(new_n463), .A2(new_n482), .B1(G228gat), .B2(G233gat), .ZN(new_n483));
  OR3_X1    g282(.A1(new_n474), .A2(new_n483), .A3(G22gat), .ZN(new_n484));
  OAI21_X1  g283(.A(G22gat), .B1(new_n474), .B2(new_n483), .ZN(new_n485));
  XOR2_X1   g284(.A(KEYINPUT31), .B(G50gat), .Z(new_n486));
  XNOR2_X1  g285(.A(new_n486), .B(KEYINPUT79), .ZN(new_n487));
  XOR2_X1   g286(.A(G78gat), .B(G106gat), .Z(new_n488));
  XNOR2_X1  g287(.A(new_n487), .B(new_n488), .ZN(new_n489));
  AND4_X1   g288(.A1(new_n441), .A2(new_n484), .A3(new_n485), .A4(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n485), .A2(KEYINPUT81), .ZN(new_n491));
  AOI22_X1  g290(.A1(new_n491), .A2(new_n489), .B1(new_n484), .B2(new_n485), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT6), .ZN(new_n494));
  XNOR2_X1  g293(.A(G1gat), .B(G29gat), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n495), .B(KEYINPUT0), .ZN(new_n496));
  XNOR2_X1  g295(.A(G57gat), .B(G85gat), .ZN(new_n497));
  XOR2_X1   g296(.A(new_n496), .B(new_n497), .Z(new_n498));
  NAND3_X1  g297(.A1(new_n470), .A2(KEYINPUT3), .A3(new_n471), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n407), .B1(new_n459), .B2(new_n460), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(G225gat), .A2(G233gat), .ZN(new_n502));
  INV_X1    g301(.A(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT4), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n459), .A2(new_n407), .A3(new_n504), .ZN(new_n505));
  OAI21_X1  g304(.A(KEYINPUT4), .B1(new_n468), .B2(new_n401), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n503), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n501), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n470), .A2(new_n401), .A3(new_n471), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n459), .A2(new_n407), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(new_n503), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n508), .A2(new_n512), .A3(KEYINPUT5), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n503), .A2(KEYINPUT5), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n504), .B1(new_n459), .B2(new_n407), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT77), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n515), .B1(new_n516), .B2(new_n505), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n510), .A2(new_n516), .A3(KEYINPUT4), .ZN(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  OAI211_X1 g318(.A(new_n501), .B(new_n514), .C1(new_n517), .C2(new_n519), .ZN(new_n520));
  AOI211_X1 g319(.A(new_n494), .B(new_n498), .C1(new_n513), .C2(new_n520), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n498), .B1(new_n513), .B2(new_n520), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n522), .A2(KEYINPUT6), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n513), .A2(new_n520), .A3(new_n498), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n521), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  NAND4_X1  g325(.A1(new_n393), .A2(new_n440), .A3(new_n493), .A4(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT35), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n520), .ZN(new_n530));
  INV_X1    g329(.A(new_n498), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n532), .A2(new_n494), .A3(new_n524), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT78), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n523), .A2(KEYINPUT78), .A3(new_n524), .ZN(new_n536));
  INV_X1    g335(.A(new_n521), .ZN(new_n537));
  AND3_X1   g336(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n538), .A2(new_n528), .ZN(new_n539));
  NAND4_X1  g338(.A1(new_n539), .A2(new_n393), .A3(new_n493), .A4(new_n440), .ZN(new_n540));
  AND2_X1   g339(.A1(new_n529), .A2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT36), .ZN(new_n542));
  NOR3_X1   g341(.A1(new_n424), .A2(new_n435), .A3(new_n412), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n411), .B1(new_n437), .B2(new_n438), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n436), .A2(KEYINPUT36), .A3(new_n439), .ZN(new_n546));
  AND2_X1   g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n501), .B1(new_n517), .B2(new_n519), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT82), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n548), .A2(new_n549), .A3(new_n503), .ZN(new_n550));
  NOR3_X1   g349(.A1(new_n468), .A2(KEYINPUT4), .A3(new_n401), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n506), .B1(new_n551), .B2(KEYINPUT77), .ZN(new_n552));
  AOI22_X1  g351(.A1(new_n552), .A2(new_n518), .B1(new_n499), .B2(new_n500), .ZN(new_n553));
  OAI21_X1  g352(.A(KEYINPUT82), .B1(new_n553), .B2(new_n502), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n550), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT39), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n531), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n509), .A2(new_n502), .A3(new_n510), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n550), .A2(new_n554), .A3(KEYINPUT39), .A4(new_n558), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n557), .A2(KEYINPUT40), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n549), .B1(new_n548), .B2(new_n503), .ZN(new_n561));
  NOR3_X1   g360(.A1(new_n553), .A2(KEYINPUT82), .A3(new_n502), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n556), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n563), .A2(new_n498), .A3(new_n559), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT40), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND4_X1  g365(.A1(new_n392), .A2(new_n532), .A3(new_n560), .A4(new_n566), .ZN(new_n567));
  NOR3_X1   g366(.A1(new_n387), .A2(new_n368), .A3(new_n382), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT37), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n380), .B1(new_n377), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n376), .A2(new_n383), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n362), .A2(new_n367), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n569), .B1(new_n572), .B2(new_n309), .ZN(new_n573));
  AOI21_X1  g372(.A(KEYINPUT38), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n568), .B1(new_n570), .B2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT38), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n382), .A2(KEYINPUT37), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n376), .A2(new_n309), .ZN(new_n578));
  INV_X1    g377(.A(new_n368), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  AOI22_X1  g379(.A1(new_n388), .A2(new_n577), .B1(new_n580), .B2(KEYINPUT37), .ZN(new_n581));
  OAI211_X1 g380(.A(new_n575), .B(new_n525), .C1(new_n576), .C2(new_n581), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n567), .A2(new_n493), .A3(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n493), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n584), .B1(new_n538), .B2(new_n392), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n547), .A2(new_n583), .A3(new_n585), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n300), .B1(new_n541), .B2(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(G134gat), .B(G162gat), .ZN(new_n588));
  AOI21_X1  g387(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n589));
  XOR2_X1   g388(.A(new_n588), .B(new_n589), .Z(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n266), .B1(new_n246), .B2(new_n255), .ZN(new_n592));
  AND2_X1   g391(.A1(G99gat), .A2(G106gat), .ZN(new_n593));
  NOR2_X1   g392(.A1(G99gat), .A2(G106gat), .ZN(new_n594));
  OAI21_X1  g393(.A(KEYINPUT95), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  OR2_X1    g394(.A1(G99gat), .A2(G106gat), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT95), .ZN(new_n597));
  NAND2_X1  g396(.A1(G99gat), .A2(G106gat), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(G85gat), .A2(G92gat), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n600), .A2(KEYINPUT7), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT7), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n602), .A2(G85gat), .A3(G92gat), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(G85gat), .ZN(new_n605));
  INV_X1    g404(.A(G92gat), .ZN(new_n606));
  AOI22_X1  g405(.A1(KEYINPUT8), .A2(new_n598), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  AND4_X1   g406(.A1(new_n595), .A2(new_n599), .A3(new_n604), .A4(new_n607), .ZN(new_n608));
  AOI22_X1  g407(.A1(new_n595), .A2(new_n599), .B1(new_n604), .B2(new_n607), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n592), .A2(new_n268), .A3(new_n611), .ZN(new_n612));
  AND3_X1   g411(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n613), .B1(new_n263), .B2(new_n610), .ZN(new_n614));
  XNOR2_X1  g413(.A(G190gat), .B(G218gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(KEYINPUT96), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n612), .A2(new_n614), .A3(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT97), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n612), .A2(new_n614), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n621), .A2(new_n616), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n591), .B1(new_n620), .B2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT98), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n621), .A2(KEYINPUT98), .A3(new_n616), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n625), .A2(new_n591), .A3(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n618), .B(KEYINPUT97), .ZN(new_n628));
  OAI21_X1  g427(.A(KEYINPUT99), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT99), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n590), .B1(new_n622), .B2(new_n624), .ZN(new_n631));
  NAND4_X1  g430(.A1(new_n620), .A2(new_n630), .A3(new_n631), .A4(new_n626), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n623), .B1(new_n629), .B2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT21), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT92), .ZN(new_n635));
  INV_X1    g434(.A(G64gat), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n635), .B1(new_n636), .B2(G57gat), .ZN(new_n637));
  INV_X1    g436(.A(G57gat), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n638), .A2(KEYINPUT92), .A3(G64gat), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n636), .A2(G57gat), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n637), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  NOR2_X1   g440(.A1(G71gat), .A2(G78gat), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(KEYINPUT9), .ZN(new_n643));
  NAND2_X1  g442(.A1(G71gat), .A2(G78gat), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n641), .A2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n644), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n647), .A2(new_n642), .ZN(new_n648));
  XNOR2_X1  g447(.A(G57gat), .B(G64gat), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT9), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n648), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n646), .A2(new_n651), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n223), .B1(new_n634), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n634), .ZN(new_n654));
  XOR2_X1   g453(.A(KEYINPUT94), .B(KEYINPUT19), .Z(new_n655));
  XNOR2_X1  g454(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n653), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(G127gat), .B(G155gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(KEYINPUT20), .ZN(new_n659));
  NAND2_X1  g458(.A1(G231gat), .A2(G233gat), .ZN(new_n660));
  XOR2_X1   g459(.A(new_n660), .B(KEYINPUT93), .Z(new_n661));
  XNOR2_X1  g460(.A(new_n659), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(G183gat), .B(G211gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n657), .B(new_n664), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n652), .B1(new_n608), .B2(new_n609), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n599), .A2(new_n595), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n604), .A2(new_n607), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND4_X1  g468(.A1(new_n595), .A2(new_n599), .A3(new_n604), .A4(new_n607), .ZN(new_n670));
  NAND4_X1  g469(.A1(new_n669), .A2(new_n646), .A3(new_n670), .A4(new_n651), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT10), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n666), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n652), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n610), .A2(KEYINPUT10), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(G230gat), .A2(G233gat), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n677), .B1(new_n666), .B2(new_n671), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  XNOR2_X1  g479(.A(G120gat), .B(G148gat), .ZN(new_n681));
  XNOR2_X1  g480(.A(G176gat), .B(G204gat), .ZN(new_n682));
  XOR2_X1   g481(.A(new_n681), .B(new_n682), .Z(new_n683));
  NAND3_X1  g482(.A1(new_n678), .A2(new_n680), .A3(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n683), .ZN(new_n685));
  INV_X1    g484(.A(new_n677), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n686), .B1(new_n673), .B2(new_n675), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n685), .B1(new_n687), .B2(new_n679), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n684), .A2(KEYINPUT100), .A3(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT100), .ZN(new_n690));
  OAI211_X1 g489(.A(new_n690), .B(new_n685), .C1(new_n687), .C2(new_n679), .ZN(new_n691));
  AND2_X1   g490(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n633), .A2(new_n665), .A3(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(KEYINPUT101), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT101), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n694), .A2(new_n697), .ZN(new_n698));
  AND2_X1   g497(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n587), .A2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT102), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n587), .A2(KEYINPUT102), .A3(new_n699), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(new_n538), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g505(.A1(new_n704), .A2(new_n392), .ZN(new_n707));
  XNOR2_X1  g506(.A(KEYINPUT16), .B(G8gat), .ZN(new_n708));
  OAI21_X1  g507(.A(KEYINPUT103), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(KEYINPUT42), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT42), .ZN(new_n711));
  OAI211_X1 g510(.A(KEYINPUT103), .B(new_n711), .C1(new_n707), .C2(new_n708), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n707), .A2(G8gat), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n710), .A2(new_n712), .A3(new_n713), .ZN(G1325gat));
  INV_X1    g513(.A(new_n704), .ZN(new_n715));
  OAI21_X1  g514(.A(G15gat), .B1(new_n715), .B2(new_n547), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n704), .A2(new_n207), .A3(new_n440), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(G1326gat));
  NAND2_X1  g517(.A1(new_n704), .A2(new_n584), .ZN(new_n719));
  XNOR2_X1  g518(.A(KEYINPUT43), .B(G22gat), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n719), .B(new_n720), .ZN(G1327gat));
  NOR2_X1   g520(.A1(new_n633), .A2(new_n665), .ZN(new_n722));
  AND3_X1   g521(.A1(new_n587), .A2(new_n693), .A3(new_n722), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n723), .A2(new_n225), .A3(new_n538), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n724), .B(KEYINPUT45), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT44), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n529), .A2(new_n540), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n521), .B1(new_n533), .B2(new_n534), .ZN(new_n728));
  AOI22_X1  g527(.A1(new_n728), .A2(new_n536), .B1(new_n391), .B2(new_n389), .ZN(new_n729));
  OAI211_X1 g528(.A(new_n545), .B(new_n546), .C1(new_n493), .C2(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n582), .A2(new_n493), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n389), .A2(new_n532), .A3(new_n391), .ZN(new_n732));
  AND4_X1   g531(.A1(KEYINPUT40), .A2(new_n563), .A3(new_n498), .A4(new_n559), .ZN(new_n733));
  AOI21_X1  g532(.A(KEYINPUT40), .B1(new_n557), .B2(new_n559), .ZN(new_n734));
  NOR3_X1   g533(.A1(new_n732), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n731), .A2(new_n735), .ZN(new_n736));
  OAI21_X1  g535(.A(KEYINPUT105), .B1(new_n730), .B2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT105), .ZN(new_n738));
  NAND4_X1  g537(.A1(new_n547), .A2(new_n738), .A3(new_n583), .A4(new_n585), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n727), .B1(new_n737), .B2(new_n739), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n726), .B1(new_n740), .B2(new_n633), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n541), .A2(new_n586), .ZN(new_n742));
  INV_X1    g541(.A(new_n633), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n742), .A2(KEYINPUT44), .A3(new_n743), .ZN(new_n744));
  AND2_X1   g543(.A1(new_n741), .A2(new_n744), .ZN(new_n745));
  XOR2_X1   g544(.A(new_n692), .B(KEYINPUT104), .Z(new_n746));
  NOR3_X1   g545(.A1(new_n746), .A2(new_n300), .A3(new_n665), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(new_n538), .ZN(new_n749));
  OAI21_X1  g548(.A(KEYINPUT106), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(G29gat), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n748), .A2(KEYINPUT106), .A3(new_n749), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n725), .B1(new_n751), .B2(new_n752), .ZN(G1328gat));
  OAI21_X1  g552(.A(G36gat), .B1(new_n748), .B2(new_n393), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n723), .A2(new_n226), .A3(new_n392), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT46), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n756), .A2(KEYINPUT107), .ZN(new_n757));
  AND2_X1   g556(.A1(new_n756), .A2(KEYINPUT107), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n755), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  OAI211_X1 g558(.A(new_n754), .B(new_n759), .C1(new_n757), .C2(new_n755), .ZN(G1329gat));
  NAND2_X1  g559(.A1(new_n723), .A2(new_n440), .ZN(new_n761));
  AND2_X1   g560(.A1(new_n238), .A2(new_n239), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  OR2_X1    g562(.A1(new_n547), .A2(new_n762), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n763), .B1(new_n748), .B2(new_n764), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g565(.A1(new_n723), .A2(new_n230), .A3(new_n584), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n741), .A2(new_n584), .A3(new_n744), .A4(new_n747), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT108), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(G50gat), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n768), .A2(new_n769), .ZN(new_n772));
  OAI211_X1 g571(.A(KEYINPUT48), .B(new_n767), .C1(new_n771), .C2(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n768), .A2(G50gat), .ZN(new_n774));
  AND2_X1   g573(.A1(new_n774), .A2(new_n767), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n773), .B1(KEYINPUT48), .B2(new_n775), .ZN(G1331gat));
  INV_X1    g575(.A(new_n300), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n737), .A2(new_n739), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n777), .B1(new_n778), .B2(new_n541), .ZN(new_n779));
  INV_X1    g578(.A(new_n779), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n746), .A2(new_n665), .A3(new_n633), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(new_n538), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n783), .B(G57gat), .ZN(G1332gat));
  INV_X1    g583(.A(new_n782), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n785), .A2(new_n393), .ZN(new_n786));
  NOR2_X1   g585(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n787));
  AND2_X1   g586(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n786), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n789), .B1(new_n786), .B2(new_n787), .ZN(G1333gat));
  INV_X1    g589(.A(G71gat), .ZN(new_n791));
  INV_X1    g590(.A(new_n440), .ZN(new_n792));
  OR2_X1    g591(.A1(new_n792), .A2(KEYINPUT109), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(KEYINPUT109), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(new_n795), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n791), .B1(new_n785), .B2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(new_n547), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n782), .A2(G71gat), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(KEYINPUT50), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT50), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n797), .A2(new_n802), .A3(new_n799), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n801), .A2(new_n803), .ZN(G1334gat));
  NAND2_X1  g603(.A1(new_n782), .A2(new_n584), .ZN(new_n805));
  XNOR2_X1  g604(.A(new_n805), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g605(.A1(new_n777), .A2(new_n665), .A3(new_n693), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n745), .A2(new_n538), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(G85gat), .ZN(new_n809));
  AOI21_X1  g608(.A(KEYINPUT51), .B1(new_n779), .B2(new_n722), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT51), .ZN(new_n811));
  INV_X1    g610(.A(new_n722), .ZN(new_n812));
  NOR4_X1   g611(.A1(new_n740), .A2(new_n811), .A3(new_n777), .A4(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT110), .ZN(new_n814));
  OR3_X1    g613(.A1(new_n810), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n814), .B1(new_n810), .B2(new_n813), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n815), .A2(new_n692), .A3(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n538), .A2(new_n605), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n809), .B1(new_n817), .B2(new_n818), .ZN(G1336gat));
  NAND4_X1  g618(.A1(new_n741), .A2(new_n392), .A3(new_n744), .A4(new_n807), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(G92gat), .ZN(new_n821));
  INV_X1    g620(.A(new_n746), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n393), .A2(new_n822), .A3(G92gat), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n823), .B1(new_n810), .B2(new_n813), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n821), .A2(new_n824), .ZN(new_n825));
  XNOR2_X1  g624(.A(new_n825), .B(KEYINPUT52), .ZN(G1337gat));
  NAND3_X1  g625(.A1(new_n745), .A2(new_n798), .A3(new_n807), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(KEYINPUT111), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(G99gat), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n827), .A2(KEYINPUT111), .ZN(new_n830));
  OR2_X1    g629(.A1(new_n792), .A2(G99gat), .ZN(new_n831));
  OAI22_X1  g630(.A1(new_n829), .A2(new_n830), .B1(new_n817), .B2(new_n831), .ZN(G1338gat));
  NOR3_X1   g631(.A1(new_n822), .A2(new_n493), .A3(G106gat), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n833), .B1(new_n810), .B2(new_n813), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(KEYINPUT112), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT112), .ZN(new_n836));
  OAI211_X1 g635(.A(new_n836), .B(new_n833), .C1(new_n810), .C2(new_n813), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n741), .A2(new_n584), .A3(new_n744), .A4(new_n807), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(G106gat), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n835), .A2(new_n837), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(KEYINPUT53), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n834), .A2(KEYINPUT113), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT53), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT113), .ZN(new_n844));
  OAI211_X1 g643(.A(new_n844), .B(new_n833), .C1(new_n810), .C2(new_n813), .ZN(new_n845));
  NAND4_X1  g644(.A1(new_n842), .A2(new_n843), .A3(new_n839), .A4(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n841), .A2(new_n846), .ZN(G1339gat));
  NOR2_X1   g646(.A1(new_n694), .A2(new_n777), .ZN(new_n848));
  NAND4_X1  g647(.A1(new_n293), .A2(new_n296), .A3(new_n297), .A4(new_n287), .ZN(new_n849));
  AND3_X1   g648(.A1(new_n272), .A2(new_n279), .A3(new_n278), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n270), .B1(new_n272), .B2(new_n273), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n286), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n849), .A2(new_n692), .A3(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(KEYINPUT115), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT115), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n849), .A2(new_n692), .A3(new_n855), .A4(new_n852), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n673), .A2(new_n675), .A3(new_n686), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n678), .A2(KEYINPUT54), .A3(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT54), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n683), .B1(new_n687), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT55), .ZN(new_n863));
  OAI21_X1  g662(.A(KEYINPUT114), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NOR3_X1   g663(.A1(new_n687), .A2(new_n679), .A3(new_n685), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n865), .B1(new_n862), .B2(new_n863), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT114), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n859), .A2(new_n861), .A3(new_n867), .A4(KEYINPUT55), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n864), .A2(new_n866), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n281), .A2(new_n290), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n294), .A2(new_n298), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n869), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n633), .B1(new_n857), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n849), .A2(new_n852), .ZN(new_n874));
  OR3_X1    g673(.A1(new_n633), .A2(new_n869), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n665), .B1(new_n876), .B2(KEYINPUT116), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n633), .A2(new_n869), .A3(new_n874), .ZN(new_n878));
  AND3_X1   g677(.A1(new_n864), .A2(new_n866), .A3(new_n868), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n879), .B1(new_n291), .B2(new_n299), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n880), .A2(new_n856), .A3(new_n854), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n878), .B1(new_n881), .B2(new_n633), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT116), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n848), .B1(new_n877), .B2(new_n884), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n885), .A2(new_n584), .ZN(new_n886));
  NAND4_X1  g685(.A1(new_n886), .A2(new_n538), .A3(new_n393), .A4(new_n440), .ZN(new_n887));
  INV_X1    g686(.A(G113gat), .ZN(new_n888));
  NOR3_X1   g687(.A1(new_n887), .A2(new_n888), .A3(new_n300), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n885), .A2(new_n749), .ZN(new_n890));
  AND4_X1   g689(.A1(new_n393), .A2(new_n890), .A3(new_n493), .A4(new_n440), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(new_n777), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n889), .B1(new_n888), .B2(new_n892), .ZN(G1340gat));
  INV_X1    g692(.A(G120gat), .ZN(new_n894));
  NOR3_X1   g693(.A1(new_n887), .A2(new_n894), .A3(new_n822), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n891), .A2(new_n692), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n895), .B1(new_n894), .B2(new_n896), .ZN(G1341gat));
  INV_X1    g696(.A(G127gat), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n891), .A2(new_n898), .A3(new_n665), .ZN(new_n899));
  INV_X1    g698(.A(new_n665), .ZN(new_n900));
  OAI21_X1  g699(.A(G127gat), .B1(new_n887), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n899), .A2(new_n901), .ZN(G1342gat));
  INV_X1    g701(.A(G134gat), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n891), .A2(new_n903), .A3(new_n743), .ZN(new_n904));
  OR2_X1    g703(.A1(new_n904), .A2(KEYINPUT56), .ZN(new_n905));
  OAI21_X1  g704(.A(G134gat), .B1(new_n887), .B2(new_n633), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n904), .A2(KEYINPUT56), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n905), .A2(new_n906), .A3(new_n907), .ZN(G1343gat));
  INV_X1    g707(.A(KEYINPUT58), .ZN(new_n909));
  NOR3_X1   g708(.A1(new_n798), .A2(new_n392), .A3(new_n493), .ZN(new_n910));
  AND2_X1   g709(.A1(new_n890), .A2(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(G141gat), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n911), .A2(new_n912), .A3(new_n777), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n909), .B1(new_n913), .B2(KEYINPUT120), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n393), .A2(new_n538), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n798), .A2(new_n915), .ZN(new_n916));
  INV_X1    g715(.A(new_n916), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT57), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n918), .B1(new_n885), .B2(new_n493), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n880), .A2(KEYINPUT118), .A3(new_n853), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT118), .ZN(new_n921));
  INV_X1    g720(.A(new_n853), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n921), .B1(new_n872), .B2(new_n922), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n743), .B1(new_n920), .B2(new_n923), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT119), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n875), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  AOI211_X1 g725(.A(KEYINPUT119), .B(new_n743), .C1(new_n920), .C2(new_n923), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n900), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  INV_X1    g727(.A(new_n848), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n493), .A2(new_n918), .ZN(new_n931));
  AOI22_X1  g730(.A1(new_n919), .A2(KEYINPUT117), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n900), .B1(new_n882), .B2(new_n883), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n876), .A2(KEYINPUT116), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n929), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  AOI21_X1  g734(.A(KEYINPUT57), .B1(new_n935), .B2(new_n584), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT117), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n917), .B1(new_n932), .B2(new_n938), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n465), .B1(new_n939), .B2(new_n777), .ZN(new_n940));
  AND3_X1   g739(.A1(new_n911), .A2(new_n912), .A3(new_n777), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n914), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n930), .A2(new_n931), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n943), .B1(new_n937), .B2(new_n936), .ZN(new_n944));
  INV_X1    g743(.A(new_n938), .ZN(new_n945));
  OAI211_X1 g744(.A(new_n777), .B(new_n916), .C1(new_n944), .C2(new_n945), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n946), .A2(new_n452), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT120), .ZN(new_n948));
  OAI21_X1  g747(.A(KEYINPUT58), .B1(new_n941), .B2(new_n948), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n947), .A2(new_n949), .A3(new_n913), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n942), .A2(new_n950), .ZN(G1344gat));
  NAND3_X1  g750(.A1(new_n911), .A2(new_n450), .A3(new_n692), .ZN(new_n952));
  AOI211_X1 g751(.A(KEYINPUT59), .B(new_n450), .C1(new_n939), .C2(new_n692), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT59), .ZN(new_n954));
  INV_X1    g753(.A(new_n931), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n885), .A2(new_n955), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n900), .B1(new_n924), .B2(new_n878), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n696), .A2(new_n300), .A3(new_n698), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  AOI21_X1  g758(.A(KEYINPUT57), .B1(new_n959), .B2(new_n584), .ZN(new_n960));
  OAI211_X1 g759(.A(new_n692), .B(new_n916), .C1(new_n956), .C2(new_n960), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n954), .B1(new_n961), .B2(G148gat), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n952), .B1(new_n953), .B2(new_n962), .ZN(G1345gat));
  NAND3_X1  g762(.A1(new_n911), .A2(new_n442), .A3(new_n665), .ZN(new_n964));
  AND2_X1   g763(.A1(new_n939), .A2(new_n665), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n964), .B1(new_n965), .B2(new_n442), .ZN(G1346gat));
  AOI21_X1  g765(.A(new_n443), .B1(new_n939), .B2(new_n743), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n911), .A2(new_n443), .A3(new_n743), .ZN(new_n968));
  INV_X1    g767(.A(new_n968), .ZN(new_n969));
  OAI21_X1  g768(.A(KEYINPUT121), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  OAI211_X1 g769(.A(new_n743), .B(new_n916), .C1(new_n944), .C2(new_n945), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n971), .A2(G162gat), .ZN(new_n972));
  INV_X1    g771(.A(KEYINPUT121), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n972), .A2(new_n973), .A3(new_n968), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n970), .A2(new_n974), .ZN(G1347gat));
  NOR2_X1   g774(.A1(new_n393), .A2(new_n538), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n886), .A2(new_n795), .A3(new_n976), .ZN(new_n977));
  INV_X1    g776(.A(KEYINPUT123), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND4_X1  g778(.A1(new_n886), .A2(KEYINPUT123), .A3(new_n795), .A4(new_n976), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g780(.A(G169gat), .ZN(new_n982));
  NOR3_X1   g781(.A1(new_n981), .A2(new_n982), .A3(new_n300), .ZN(new_n983));
  OAI21_X1  g782(.A(KEYINPUT122), .B1(new_n885), .B2(new_n538), .ZN(new_n984));
  INV_X1    g783(.A(KEYINPUT122), .ZN(new_n985));
  NAND3_X1  g784(.A1(new_n935), .A2(new_n985), .A3(new_n749), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n984), .A2(new_n986), .ZN(new_n987));
  NOR3_X1   g786(.A1(new_n792), .A2(new_n584), .A3(new_n393), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  INV_X1    g788(.A(new_n989), .ZN(new_n990));
  AOI21_X1  g789(.A(G169gat), .B1(new_n990), .B2(new_n777), .ZN(new_n991));
  NOR2_X1   g790(.A1(new_n983), .A2(new_n991), .ZN(G1348gat));
  OAI21_X1  g791(.A(G176gat), .B1(new_n981), .B2(new_n822), .ZN(new_n993));
  OR2_X1    g792(.A1(new_n693), .A2(G176gat), .ZN(new_n994));
  OAI21_X1  g793(.A(new_n993), .B1(new_n989), .B2(new_n994), .ZN(G1349gat));
  NAND3_X1  g794(.A1(new_n979), .A2(new_n665), .A3(new_n980), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n996), .A2(new_n356), .ZN(new_n997));
  NAND3_X1  g796(.A1(new_n990), .A2(new_n337), .A3(new_n665), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n999), .A2(KEYINPUT60), .ZN(new_n1000));
  INV_X1    g799(.A(KEYINPUT60), .ZN(new_n1001));
  NAND3_X1  g800(.A1(new_n997), .A2(new_n1001), .A3(new_n998), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n1000), .A2(new_n1002), .ZN(G1350gat));
  NAND3_X1  g802(.A1(new_n990), .A2(new_n310), .A3(new_n743), .ZN(new_n1004));
  INV_X1    g803(.A(KEYINPUT124), .ZN(new_n1005));
  NAND3_X1  g804(.A1(new_n979), .A2(new_n743), .A3(new_n980), .ZN(new_n1006));
  INV_X1    g805(.A(KEYINPUT61), .ZN(new_n1007));
  AND4_X1   g806(.A1(new_n1005), .A2(new_n1006), .A3(new_n1007), .A4(G190gat), .ZN(new_n1008));
  INV_X1    g807(.A(G190gat), .ZN(new_n1009));
  AOI21_X1  g808(.A(new_n1009), .B1(KEYINPUT124), .B2(KEYINPUT61), .ZN(new_n1010));
  AOI22_X1  g809(.A1(new_n1006), .A2(new_n1010), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1011));
  OAI21_X1  g810(.A(new_n1004), .B1(new_n1008), .B2(new_n1011), .ZN(G1351gat));
  NAND4_X1  g811(.A1(new_n545), .A2(new_n584), .A3(new_n392), .A4(new_n546), .ZN(new_n1013));
  XNOR2_X1  g812(.A(new_n1013), .B(KEYINPUT125), .ZN(new_n1014));
  AOI21_X1  g813(.A(new_n1014), .B1(new_n984), .B2(new_n986), .ZN(new_n1015));
  AOI21_X1  g814(.A(G197gat), .B1(new_n1015), .B2(new_n777), .ZN(new_n1016));
  NOR2_X1   g815(.A1(new_n956), .A2(new_n960), .ZN(new_n1017));
  INV_X1    g816(.A(new_n976), .ZN(new_n1018));
  NOR3_X1   g817(.A1(new_n1017), .A2(new_n798), .A3(new_n1018), .ZN(new_n1019));
  AND2_X1   g818(.A1(new_n777), .A2(G197gat), .ZN(new_n1020));
  AOI21_X1  g819(.A(new_n1016), .B1(new_n1019), .B2(new_n1020), .ZN(G1352gat));
  NOR2_X1   g820(.A1(new_n693), .A2(G204gat), .ZN(new_n1022));
  INV_X1    g821(.A(new_n1022), .ZN(new_n1023));
  AOI211_X1 g822(.A(new_n1014), .B(new_n1023), .C1(new_n984), .C2(new_n986), .ZN(new_n1024));
  INV_X1    g823(.A(KEYINPUT62), .ZN(new_n1025));
  NOR2_X1   g824(.A1(new_n798), .A2(new_n1018), .ZN(new_n1026));
  OAI211_X1 g825(.A(new_n746), .B(new_n1026), .C1(new_n956), .C2(new_n960), .ZN(new_n1027));
  AOI22_X1  g826(.A1(new_n1024), .A2(new_n1025), .B1(G204gat), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g827(.A(new_n1014), .ZN(new_n1029));
  NOR3_X1   g828(.A1(new_n885), .A2(KEYINPUT122), .A3(new_n538), .ZN(new_n1030));
  AOI21_X1  g829(.A(new_n985), .B1(new_n935), .B2(new_n749), .ZN(new_n1031));
  OAI211_X1 g830(.A(new_n1029), .B(new_n1022), .C1(new_n1030), .C2(new_n1031), .ZN(new_n1032));
  INV_X1    g831(.A(KEYINPUT126), .ZN(new_n1033));
  AND3_X1   g832(.A1(new_n1032), .A2(new_n1033), .A3(KEYINPUT62), .ZN(new_n1034));
  AOI21_X1  g833(.A(new_n1033), .B1(new_n1032), .B2(KEYINPUT62), .ZN(new_n1035));
  OAI21_X1  g834(.A(new_n1028), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g835(.A1(new_n1036), .A2(KEYINPUT127), .ZN(new_n1037));
  INV_X1    g836(.A(KEYINPUT127), .ZN(new_n1038));
  OAI211_X1 g837(.A(new_n1028), .B(new_n1038), .C1(new_n1034), .C2(new_n1035), .ZN(new_n1039));
  NAND2_X1  g838(.A1(new_n1037), .A2(new_n1039), .ZN(G1353gat));
  NAND3_X1  g839(.A1(new_n1015), .A2(new_n305), .A3(new_n665), .ZN(new_n1041));
  NAND2_X1  g840(.A1(new_n1019), .A2(new_n665), .ZN(new_n1042));
  AND3_X1   g841(.A1(new_n1042), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1043));
  AOI21_X1  g842(.A(KEYINPUT63), .B1(new_n1042), .B2(G211gat), .ZN(new_n1044));
  OAI21_X1  g843(.A(new_n1041), .B1(new_n1043), .B2(new_n1044), .ZN(G1354gat));
  NAND3_X1  g844(.A1(new_n1015), .A2(new_n306), .A3(new_n743), .ZN(new_n1046));
  NAND2_X1  g845(.A1(new_n1019), .A2(new_n743), .ZN(new_n1047));
  INV_X1    g846(.A(new_n1047), .ZN(new_n1048));
  OAI21_X1  g847(.A(new_n1046), .B1(new_n1048), .B2(new_n306), .ZN(G1355gat));
endmodule


