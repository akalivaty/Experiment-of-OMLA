//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 1 0 0 0 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 0 1 0 1 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 0 1 0 0 0 0 0 1 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:52 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n670, new_n671, new_n672, new_n673, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n682, new_n683, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n718, new_n719, new_n720, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991;
  INV_X1    g000(.A(KEYINPUT79), .ZN(new_n187));
  XNOR2_X1  g001(.A(G104), .B(G107), .ZN(new_n188));
  INV_X1    g002(.A(G101), .ZN(new_n189));
  OAI21_X1  g003(.A(new_n187), .B1(new_n188), .B2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G104), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G107), .ZN(new_n192));
  INV_X1    g006(.A(G107), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G104), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n195), .A2(KEYINPUT79), .A3(G101), .ZN(new_n196));
  OAI21_X1  g010(.A(KEYINPUT3), .B1(new_n191), .B2(G107), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT3), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n198), .A2(new_n193), .A3(G104), .ZN(new_n199));
  AND3_X1   g013(.A1(new_n197), .A2(new_n199), .A3(new_n192), .ZN(new_n200));
  AOI22_X1  g014(.A1(new_n190), .A2(new_n196), .B1(new_n200), .B2(new_n189), .ZN(new_n201));
  INV_X1    g015(.A(G116), .ZN(new_n202));
  NOR3_X1   g016(.A1(new_n202), .A2(KEYINPUT5), .A3(G119), .ZN(new_n203));
  XNOR2_X1  g017(.A(G116), .B(G119), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n203), .B1(new_n204), .B2(KEYINPUT5), .ZN(new_n205));
  XNOR2_X1  g019(.A(KEYINPUT2), .B(G113), .ZN(new_n206));
  INV_X1    g020(.A(new_n206), .ZN(new_n207));
  AOI22_X1  g021(.A1(new_n205), .A2(G113), .B1(new_n204), .B2(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n201), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(KEYINPUT82), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT83), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n211), .B1(new_n201), .B2(new_n208), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n190), .A2(new_n196), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n197), .A2(new_n199), .A3(new_n189), .A4(new_n192), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n205), .A2(G113), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n207), .A2(new_n204), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n215), .A2(new_n218), .A3(KEYINPUT83), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT82), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n201), .A2(new_n220), .A3(new_n208), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n210), .A2(new_n212), .A3(new_n219), .A4(new_n221), .ZN(new_n222));
  XOR2_X1   g036(.A(G110), .B(G122), .Z(new_n223));
  XOR2_X1   g037(.A(new_n223), .B(KEYINPUT8), .Z(new_n224));
  NAND2_X1  g038(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(KEYINPUT0), .A2(G128), .ZN(new_n226));
  XNOR2_X1  g040(.A(G143), .B(G146), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT64), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n226), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(G146), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G143), .ZN(new_n231));
  INV_X1    g045(.A(G143), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(G146), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  XNOR2_X1  g048(.A(KEYINPUT0), .B(G128), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n234), .A2(new_n235), .A3(KEYINPUT64), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n229), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(G125), .ZN(new_n238));
  INV_X1    g052(.A(G128), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n239), .A2(new_n230), .A3(G143), .ZN(new_n240));
  OAI211_X1 g054(.A(new_n232), .B(G146), .C1(new_n239), .C2(KEYINPUT1), .ZN(new_n241));
  OR2_X1    g055(.A1(new_n239), .A2(KEYINPUT1), .ZN(new_n242));
  OAI211_X1 g056(.A(new_n240), .B(new_n241), .C1(new_n234), .C2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(G125), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n238), .A2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(G953), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(G224), .ZN(new_n248));
  XNOR2_X1  g062(.A(new_n248), .B(KEYINPUT81), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n246), .A2(KEYINPUT7), .A3(new_n249), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n197), .A2(new_n199), .A3(new_n192), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G101), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n252), .A2(KEYINPUT4), .A3(new_n214), .ZN(new_n253));
  INV_X1    g067(.A(new_n204), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(new_n206), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(new_n217), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n251), .A2(new_n257), .A3(G101), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n253), .A2(new_n256), .A3(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n223), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n209), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  AND2_X1   g075(.A1(new_n250), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n249), .A2(KEYINPUT7), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n238), .A2(new_n245), .A3(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n225), .A2(new_n262), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n209), .A2(new_n259), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(new_n223), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n267), .A2(KEYINPUT6), .A3(new_n261), .ZN(new_n268));
  XNOR2_X1  g082(.A(new_n246), .B(new_n249), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT6), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n266), .A2(new_n270), .A3(new_n223), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n268), .A2(new_n269), .A3(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(G902), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n265), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  OAI21_X1  g088(.A(G210), .B1(G237), .B2(G902), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n265), .A2(new_n272), .A3(new_n273), .A4(new_n275), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(KEYINPUT84), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT84), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n278), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  OAI21_X1  g097(.A(G214), .B1(G237), .B2(G902), .ZN(new_n284));
  NAND2_X1  g098(.A1(G234), .A2(G237), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n285), .A2(G952), .A3(new_n247), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  XOR2_X1   g101(.A(KEYINPUT21), .B(G898), .Z(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n285), .A2(G902), .A3(G953), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n287), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n283), .A2(new_n284), .A3(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT20), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT19), .ZN(new_n297));
  AND2_X1   g111(.A1(G125), .A2(G140), .ZN(new_n298));
  NOR2_X1   g112(.A1(G125), .A2(G140), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT74), .ZN(new_n300));
  NOR3_X1   g114(.A1(new_n298), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(G140), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n244), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(G125), .A2(G140), .ZN(new_n304));
  AOI21_X1  g118(.A(KEYINPUT74), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n297), .B1(new_n301), .B2(new_n305), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n303), .A2(KEYINPUT19), .A3(new_n304), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n306), .A2(new_n230), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(KEYINPUT87), .ZN(new_n309));
  OAI21_X1  g123(.A(KEYINPUT16), .B1(new_n298), .B2(new_n299), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT16), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n311), .A2(new_n302), .A3(G125), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n310), .A2(G146), .A3(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT73), .ZN(new_n314));
  XNOR2_X1  g128(.A(new_n313), .B(new_n314), .ZN(new_n315));
  XNOR2_X1  g129(.A(KEYINPUT65), .B(G131), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(G237), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n318), .A2(new_n247), .A3(G214), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n319), .A2(new_n232), .ZN(new_n320));
  NOR2_X1   g134(.A1(G237), .A2(G953), .ZN(new_n321));
  AOI21_X1  g135(.A(G143), .B1(new_n321), .B2(G214), .ZN(new_n322));
  OR3_X1    g136(.A1(new_n317), .A2(new_n320), .A3(new_n322), .ZN(new_n323));
  XNOR2_X1  g137(.A(new_n319), .B(new_n232), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(new_n317), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT87), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n306), .A2(new_n327), .A3(new_n230), .A4(new_n307), .ZN(new_n328));
  NAND4_X1  g142(.A1(new_n309), .A2(new_n315), .A3(new_n326), .A4(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(KEYINPUT18), .A2(G131), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n324), .A2(KEYINPUT85), .A3(new_n330), .ZN(new_n331));
  OAI21_X1  g145(.A(KEYINPUT85), .B1(new_n320), .B2(new_n322), .ZN(new_n332));
  INV_X1    g146(.A(new_n330), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n331), .A2(new_n334), .ZN(new_n335));
  OR2_X1    g149(.A1(new_n324), .A2(KEYINPUT85), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT86), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n230), .B1(new_n301), .B2(new_n305), .ZN(new_n338));
  NOR3_X1   g152(.A1(new_n298), .A2(new_n299), .A3(new_n230), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n337), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n300), .B1(new_n298), .B2(new_n299), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n303), .A2(KEYINPUT74), .A3(new_n304), .ZN(new_n343));
  AOI21_X1  g157(.A(G146), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NOR3_X1   g158(.A1(new_n344), .A2(KEYINPUT86), .A3(new_n339), .ZN(new_n345));
  OAI211_X1 g159(.A(new_n335), .B(new_n336), .C1(new_n341), .C2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n329), .A2(new_n346), .ZN(new_n347));
  XNOR2_X1  g161(.A(G113), .B(G122), .ZN(new_n348));
  XNOR2_X1  g162(.A(new_n348), .B(new_n191), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(KEYINPUT88), .B1(new_n347), .B2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT88), .ZN(new_n352));
  AOI211_X1 g166(.A(new_n352), .B(new_n349), .C1(new_n329), .C2(new_n346), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT89), .ZN(new_n354));
  OAI211_X1 g168(.A(new_n317), .B(KEYINPUT17), .C1(new_n320), .C2(new_n322), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n311), .B1(new_n303), .B2(new_n304), .ZN(new_n357));
  INV_X1    g171(.A(new_n312), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n230), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(new_n313), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n354), .B1(new_n356), .B2(new_n360), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n355), .A2(new_n359), .A3(KEYINPUT89), .A4(new_n313), .ZN(new_n362));
  OAI211_X1 g176(.A(new_n361), .B(new_n362), .C1(KEYINPUT17), .C2(new_n326), .ZN(new_n363));
  AND3_X1   g177(.A1(new_n363), .A2(new_n349), .A3(new_n346), .ZN(new_n364));
  NOR3_X1   g178(.A1(new_n351), .A2(new_n353), .A3(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(G475), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(new_n273), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n296), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  NOR2_X1   g182(.A1(G475), .A2(G902), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n347), .A2(new_n350), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(new_n352), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n347), .A2(KEYINPUT88), .A3(new_n350), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  OAI211_X1 g187(.A(KEYINPUT20), .B(new_n369), .C1(new_n373), .C2(new_n364), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n349), .B1(new_n363), .B2(new_n346), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n273), .B1(new_n364), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(G475), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n368), .A2(new_n374), .A3(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(G122), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(KEYINPUT90), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT90), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(G122), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n202), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n379), .A2(G116), .ZN(new_n384));
  OAI21_X1  g198(.A(G107), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n202), .A2(G122), .ZN(new_n386));
  XNOR2_X1  g200(.A(KEYINPUT90), .B(G122), .ZN(new_n387));
  OAI211_X1 g201(.A(new_n193), .B(new_n386), .C1(new_n387), .C2(new_n202), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n385), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n232), .A2(G128), .ZN(new_n390));
  OR2_X1    g204(.A1(new_n390), .A2(KEYINPUT13), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n239), .A2(G143), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n390), .A2(new_n392), .A3(KEYINPUT13), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n391), .A2(G134), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(KEYINPUT91), .ZN(new_n395));
  AND2_X1   g209(.A1(new_n390), .A2(new_n392), .ZN(new_n396));
  INV_X1    g210(.A(G134), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT91), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n391), .A2(new_n399), .A3(new_n393), .A4(G134), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n389), .A2(new_n395), .A3(new_n398), .A4(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT14), .ZN(new_n402));
  OAI22_X1  g216(.A1(new_n387), .A2(new_n202), .B1(new_n402), .B2(new_n384), .ZN(new_n403));
  OAI21_X1  g217(.A(KEYINPUT92), .B1(new_n386), .B2(KEYINPUT14), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT92), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n384), .A2(new_n405), .A3(new_n402), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  OAI21_X1  g221(.A(G107), .B1(new_n403), .B2(new_n407), .ZN(new_n408));
  XNOR2_X1  g222(.A(new_n396), .B(new_n397), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n408), .A2(new_n409), .A3(new_n388), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n401), .A2(new_n410), .ZN(new_n411));
  XNOR2_X1  g225(.A(KEYINPUT9), .B(G234), .ZN(new_n412));
  INV_X1    g226(.A(G217), .ZN(new_n413));
  NOR3_X1   g227(.A1(new_n412), .A2(new_n413), .A3(G953), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n411), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n401), .A2(new_n410), .A3(new_n414), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(new_n273), .ZN(new_n419));
  INV_X1    g233(.A(G478), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n420), .A2(KEYINPUT15), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n419), .B(new_n421), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n378), .A2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(G221), .ZN(new_n424));
  INV_X1    g238(.A(new_n412), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n424), .B1(new_n425), .B2(new_n273), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  XOR2_X1   g241(.A(G110), .B(G140), .Z(new_n428));
  XNOR2_X1  g242(.A(new_n428), .B(KEYINPUT78), .ZN(new_n429));
  INV_X1    g243(.A(G227), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n430), .A2(G953), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n429), .B(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT11), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n433), .B1(new_n397), .B2(G137), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n397), .A2(G137), .ZN(new_n435));
  INV_X1    g249(.A(G137), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n436), .A2(KEYINPUT11), .A3(G134), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n434), .A2(new_n435), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(G131), .ZN(new_n439));
  NAND4_X1  g253(.A1(new_n316), .A2(new_n435), .A3(new_n437), .A4(new_n434), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n253), .A2(new_n237), .A3(new_n258), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT10), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n444), .B1(new_n201), .B2(new_n243), .ZN(new_n445));
  AND4_X1   g259(.A1(new_n444), .A2(new_n213), .A3(new_n243), .A4(new_n214), .ZN(new_n446));
  OAI211_X1 g260(.A(new_n442), .B(new_n443), .C1(new_n445), .C2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n201), .A2(new_n444), .A3(new_n243), .ZN(new_n449));
  AOI21_X1  g263(.A(KEYINPUT79), .B1(new_n195), .B2(G101), .ZN(new_n450));
  AOI211_X1 g264(.A(new_n187), .B(new_n189), .C1(new_n192), .C2(new_n194), .ZN(new_n451));
  OAI211_X1 g265(.A(new_n243), .B(new_n214), .C1(new_n450), .C2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(KEYINPUT10), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n449), .A2(new_n453), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n442), .B1(new_n454), .B2(new_n443), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n432), .B1(new_n448), .B2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT80), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(new_n452), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n243), .B1(new_n213), .B2(new_n214), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n441), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(KEYINPUT12), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT12), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n463), .B(new_n441), .C1(new_n459), .C2(new_n460), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n462), .A2(new_n447), .A3(new_n464), .ZN(new_n465));
  OR2_X1    g279(.A1(new_n465), .A2(new_n432), .ZN(new_n466));
  OAI211_X1 g280(.A(KEYINPUT80), .B(new_n432), .C1(new_n448), .C2(new_n455), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n458), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(G469), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n468), .A2(new_n469), .A3(new_n273), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n469), .A2(new_n273), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  OR3_X1    g286(.A1(new_n448), .A2(new_n455), .A3(new_n432), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n465), .A2(new_n432), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n473), .A2(G469), .A3(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n470), .A2(new_n472), .A3(new_n475), .ZN(new_n476));
  AND3_X1   g290(.A1(new_n423), .A2(new_n427), .A3(new_n476), .ZN(new_n477));
  XOR2_X1   g291(.A(KEYINPUT75), .B(KEYINPUT22), .Z(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(G137), .ZN(new_n479));
  AND3_X1   g293(.A1(new_n247), .A2(G221), .A3(G234), .ZN(new_n480));
  XNOR2_X1  g294(.A(KEYINPUT75), .B(KEYINPUT22), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(new_n436), .ZN(new_n482));
  AND3_X1   g296(.A1(new_n479), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n480), .B1(new_n479), .B2(new_n482), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  XNOR2_X1  g299(.A(KEYINPUT24), .B(G110), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT71), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n486), .B(new_n487), .ZN(new_n488));
  XNOR2_X1  g302(.A(G119), .B(G128), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT23), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n490), .B1(G119), .B2(new_n239), .ZN(new_n491));
  INV_X1    g305(.A(G119), .ZN(new_n492));
  NOR3_X1   g306(.A1(new_n492), .A2(KEYINPUT23), .A3(G128), .ZN(new_n493));
  OAI22_X1  g307(.A1(new_n491), .A2(new_n493), .B1(G119), .B2(new_n239), .ZN(new_n494));
  XNOR2_X1  g308(.A(KEYINPUT72), .B(G110), .ZN(new_n495));
  OAI22_X1  g309(.A1(new_n488), .A2(new_n489), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n315), .A2(new_n496), .A3(new_n338), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n494), .A2(G110), .ZN(new_n498));
  XOR2_X1   g312(.A(KEYINPUT24), .B(G110), .Z(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(new_n487), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n486), .A2(KEYINPUT71), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n500), .A2(new_n489), .A3(new_n501), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n360), .A2(new_n498), .A3(new_n502), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n485), .B1(new_n497), .B2(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n489), .B1(new_n500), .B2(new_n501), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n494), .A2(new_n495), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n338), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  XNOR2_X1  g321(.A(new_n313), .B(KEYINPUT73), .ZN(new_n508));
  OAI211_X1 g322(.A(new_n485), .B(new_n503), .C1(new_n507), .C2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n273), .B1(new_n504), .B2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT76), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n511), .A2(new_n512), .A3(KEYINPUT25), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n503), .B1(new_n507), .B2(new_n508), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n514), .B1(new_n483), .B2(new_n484), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(new_n509), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n512), .A2(KEYINPUT25), .ZN(new_n517));
  OR2_X1    g331(.A1(new_n512), .A2(KEYINPUT25), .ZN(new_n518));
  NAND4_X1  g332(.A1(new_n516), .A2(new_n273), .A3(new_n517), .A4(new_n518), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n413), .B1(G234), .B2(new_n273), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n513), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT77), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n513), .A2(new_n519), .A3(KEYINPUT77), .A4(new_n520), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n520), .A2(G902), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n516), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n523), .A2(new_n524), .A3(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(new_n435), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n397), .A2(G137), .ZN(new_n529));
  OAI21_X1  g343(.A(G131), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n440), .A2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT66), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n440), .A2(KEYINPUT66), .A3(new_n530), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n533), .A2(new_n243), .A3(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n256), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n441), .A2(new_n237), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n243), .A2(new_n440), .A3(new_n530), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n538), .B1(new_n536), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(KEYINPUT28), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT69), .ZN(new_n544));
  INV_X1    g358(.A(new_n538), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n544), .B1(new_n545), .B2(KEYINPUT28), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT28), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n538), .A2(KEYINPUT69), .A3(new_n547), .ZN(new_n548));
  XNOR2_X1  g362(.A(KEYINPUT67), .B(KEYINPUT27), .ZN(new_n549));
  AND3_X1   g363(.A1(new_n318), .A2(new_n247), .A3(G210), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n549), .B(new_n550), .ZN(new_n551));
  XNOR2_X1  g365(.A(KEYINPUT26), .B(G101), .ZN(new_n552));
  XOR2_X1   g366(.A(new_n551), .B(new_n552), .Z(new_n553));
  NAND4_X1  g367(.A1(new_n543), .A2(new_n546), .A3(new_n548), .A4(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT30), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n555), .B1(new_n535), .B2(new_n537), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n540), .A2(KEYINPUT30), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n256), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(new_n538), .ZN(new_n559));
  INV_X1    g373(.A(new_n553), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT29), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n554), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(KEYINPUT70), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n536), .B1(new_n535), .B2(new_n537), .ZN(new_n565));
  OAI21_X1  g379(.A(KEYINPUT28), .B1(new_n545), .B2(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n566), .A2(new_n546), .A3(new_n548), .ZN(new_n567));
  OR3_X1    g381(.A1(new_n567), .A2(new_n562), .A3(new_n560), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT70), .ZN(new_n569));
  NAND4_X1  g383(.A1(new_n554), .A2(new_n561), .A3(new_n569), .A4(new_n562), .ZN(new_n570));
  NAND4_X1  g384(.A1(new_n564), .A2(new_n273), .A3(new_n568), .A4(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(G472), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT68), .ZN(new_n573));
  AND3_X1   g387(.A1(new_n538), .A2(new_n553), .A3(new_n573), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n573), .B1(new_n538), .B2(new_n553), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n576), .A2(KEYINPUT31), .A3(new_n558), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n538), .A2(new_n553), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(KEYINPUT68), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n538), .A2(new_n553), .A3(new_n573), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n579), .A2(new_n558), .A3(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT31), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n543), .A2(new_n546), .A3(new_n548), .ZN(new_n584));
  AOI22_X1  g398(.A1(new_n577), .A2(new_n583), .B1(new_n584), .B2(new_n560), .ZN(new_n585));
  INV_X1    g399(.A(G472), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(new_n273), .ZN(new_n587));
  OAI21_X1  g401(.A(KEYINPUT32), .B1(new_n585), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n584), .A2(new_n560), .ZN(new_n589));
  AOI21_X1  g403(.A(KEYINPUT31), .B1(new_n576), .B2(new_n558), .ZN(new_n590));
  AND4_X1   g404(.A1(KEYINPUT31), .A2(new_n579), .A3(new_n558), .A4(new_n580), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n589), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT32), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n592), .A2(new_n593), .A3(new_n586), .A4(new_n273), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n588), .A2(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n527), .B1(new_n572), .B2(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n295), .A2(new_n477), .A3(new_n596), .ZN(new_n597));
  XNOR2_X1  g411(.A(KEYINPUT93), .B(G101), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n597), .B(new_n598), .ZN(G3));
  NAND2_X1  g413(.A1(new_n476), .A2(new_n427), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n585), .A2(new_n587), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n586), .B1(new_n592), .B2(new_n273), .ZN(new_n602));
  NOR3_X1   g416(.A1(new_n600), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n527), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT33), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n607), .B1(new_n411), .B2(KEYINPUT94), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n608), .A2(new_n417), .A3(new_n416), .ZN(new_n609));
  INV_X1    g423(.A(new_n417), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n414), .B1(new_n401), .B2(new_n410), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT94), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n612), .B1(new_n401), .B2(new_n410), .ZN(new_n613));
  OAI22_X1  g427(.A1(new_n610), .A2(new_n611), .B1(new_n613), .B2(new_n607), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n420), .B1(new_n609), .B2(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n418), .A2(new_n420), .A3(new_n273), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n420), .A2(new_n273), .ZN(new_n618));
  NOR3_X1   g432(.A1(new_n615), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n378), .A2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n284), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n621), .B1(new_n277), .B2(new_n278), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(new_n293), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n620), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(KEYINPUT95), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n606), .A2(new_n625), .ZN(new_n626));
  XOR2_X1   g440(.A(KEYINPUT34), .B(G104), .Z(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(G6));
  AND3_X1   g442(.A1(new_n368), .A2(new_n377), .A3(new_n374), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(new_n422), .ZN(new_n630));
  NOR3_X1   g444(.A1(new_n605), .A2(new_n623), .A3(new_n630), .ZN(new_n631));
  XNOR2_X1  g445(.A(KEYINPUT35), .B(G107), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(G9));
  NOR2_X1   g447(.A1(new_n602), .A2(new_n601), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n485), .A2(KEYINPUT36), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n514), .B(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(new_n525), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n523), .A2(new_n524), .A3(new_n637), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n295), .A2(new_n477), .A3(new_n634), .A4(new_n638), .ZN(new_n639));
  XOR2_X1   g453(.A(new_n639), .B(KEYINPUT37), .Z(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(G110), .ZN(G12));
  INV_X1    g455(.A(new_n638), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n642), .B1(new_n572), .B2(new_n595), .ZN(new_n643));
  INV_X1    g457(.A(G900), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n287), .B1(new_n291), .B2(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n630), .A2(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n622), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n600), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n643), .A2(new_n646), .A3(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(G128), .ZN(G30));
  INV_X1    g464(.A(KEYINPUT96), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n280), .A2(new_n651), .A3(new_n282), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT38), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n651), .B1(new_n280), .B2(new_n282), .ZN(new_n655));
  OR3_X1    g469(.A1(new_n653), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n654), .B1(new_n653), .B2(new_n655), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XOR2_X1   g472(.A(new_n645), .B(KEYINPUT39), .Z(new_n659));
  NAND3_X1  g473(.A1(new_n476), .A2(new_n427), .A3(new_n659), .ZN(new_n660));
  XOR2_X1   g474(.A(new_n660), .B(KEYINPUT40), .Z(new_n661));
  OAI21_X1  g475(.A(new_n560), .B1(new_n545), .B2(new_n565), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(new_n581), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n586), .B1(new_n663), .B2(new_n273), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n664), .B1(new_n588), .B2(new_n594), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n378), .A2(new_n422), .ZN(new_n666));
  NOR3_X1   g480(.A1(new_n665), .A2(new_n638), .A3(new_n666), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n658), .A2(new_n284), .A3(new_n661), .A4(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(G143), .ZN(G45));
  INV_X1    g483(.A(new_n645), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n378), .A2(new_n619), .A3(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n643), .A2(new_n648), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G146), .ZN(G48));
  NAND2_X1  g488(.A1(new_n468), .A2(new_n273), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(G469), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n676), .A2(new_n427), .A3(new_n470), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n625), .A2(new_n596), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(KEYINPUT41), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G113), .ZN(G15));
  NOR3_X1   g495(.A1(new_n630), .A2(new_n677), .A3(new_n623), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n596), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G116), .ZN(G18));
  NOR2_X1   g498(.A1(new_n677), .A2(new_n647), .ZN(new_n685));
  AND2_X1   g499(.A1(new_n685), .A2(new_n423), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT97), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n686), .A2(new_n687), .A3(new_n293), .A4(new_n643), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n685), .A2(new_n293), .A3(new_n423), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n572), .A2(new_n595), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(new_n638), .ZN(new_n691));
  OAI21_X1  g505(.A(KEYINPUT97), .B1(new_n689), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n688), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G119), .ZN(G21));
  XOR2_X1   g508(.A(KEYINPUT98), .B(G472), .Z(new_n695));
  OAI21_X1  g509(.A(new_n695), .B1(new_n585), .B2(G902), .ZN(new_n696));
  AOI22_X1  g510(.A1(new_n577), .A2(new_n583), .B1(new_n560), .B2(new_n567), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n696), .B1(new_n587), .B2(new_n697), .ZN(new_n698));
  NOR3_X1   g512(.A1(new_n698), .A2(new_n677), .A3(new_n527), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n666), .A2(new_n623), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G122), .ZN(G24));
  NOR2_X1   g516(.A1(new_n698), .A2(new_n642), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n703), .A2(new_n672), .A3(new_n685), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G125), .ZN(G27));
  NAND2_X1  g519(.A1(new_n474), .A2(KEYINPUT99), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT99), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n465), .A2(new_n707), .A3(new_n432), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n706), .A2(G469), .A3(new_n473), .A4(new_n708), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n470), .A2(new_n472), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(new_n427), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n280), .A2(new_n284), .A3(new_n282), .ZN(new_n712));
  NOR3_X1   g526(.A1(new_n711), .A2(new_n712), .A3(new_n671), .ZN(new_n713));
  AND3_X1   g527(.A1(new_n713), .A2(KEYINPUT42), .A3(new_n596), .ZN(new_n714));
  AOI21_X1  g528(.A(KEYINPUT42), .B1(new_n713), .B2(new_n596), .ZN(new_n715));
  OR2_X1    g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G131), .ZN(G33));
  INV_X1    g531(.A(new_n711), .ZN(new_n718));
  INV_X1    g532(.A(new_n712), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n596), .A2(new_n646), .A3(new_n718), .A4(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G134), .ZN(G36));
  INV_X1    g535(.A(KEYINPUT101), .ZN(new_n722));
  OAI211_X1 g536(.A(new_n629), .B(new_n619), .C1(new_n722), .C2(KEYINPUT43), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n368), .A2(new_n374), .A3(new_n619), .A4(new_n377), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n368), .A2(new_n374), .A3(new_n722), .A4(new_n377), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT43), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n724), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n723), .A2(new_n727), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n638), .B1(new_n602), .B2(new_n601), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(KEYINPUT102), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT102), .ZN(new_n731));
  OAI211_X1 g545(.A(new_n638), .B(new_n731), .C1(new_n602), .C2(new_n601), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n728), .A2(KEYINPUT44), .A3(new_n730), .A4(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(new_n719), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n706), .A2(KEYINPUT45), .A3(new_n473), .A4(new_n708), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT45), .ZN(new_n736));
  INV_X1    g550(.A(new_n474), .ZN(new_n737));
  NOR3_X1   g551(.A1(new_n448), .A2(new_n455), .A3(new_n432), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n736), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n735), .A2(G469), .A3(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(KEYINPUT100), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT100), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n735), .A2(new_n739), .A3(new_n742), .A4(G469), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n471), .B1(new_n741), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(KEYINPUT46), .ZN(new_n745));
  INV_X1    g559(.A(new_n745), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n470), .B1(new_n744), .B2(KEYINPUT46), .ZN(new_n747));
  OAI211_X1 g561(.A(new_n427), .B(new_n659), .C1(new_n746), .C2(new_n747), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n734), .A2(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT44), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n730), .A2(new_n732), .ZN(new_n751));
  AND3_X1   g565(.A1(new_n724), .A2(new_n725), .A3(new_n726), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n724), .B1(new_n726), .B2(new_n725), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n750), .B1(new_n751), .B2(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT103), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  OAI211_X1 g571(.A(KEYINPUT103), .B(new_n750), .C1(new_n751), .C2(new_n754), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n749), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G137), .ZN(G39));
  NOR2_X1   g574(.A1(new_n712), .A2(new_n671), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n690), .A2(new_n604), .ZN(new_n762));
  INV_X1    g576(.A(new_n470), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n741), .A2(new_n743), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n764), .A2(new_n472), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT46), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n763), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n426), .B1(new_n767), .B2(new_n745), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n768), .A2(KEYINPUT47), .ZN(new_n769));
  OAI211_X1 g583(.A(KEYINPUT47), .B(new_n427), .C1(new_n746), .C2(new_n747), .ZN(new_n770));
  INV_X1    g584(.A(new_n770), .ZN(new_n771));
  OAI211_X1 g585(.A(new_n761), .B(new_n762), .C1(new_n769), .C2(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G140), .ZN(G42));
  NOR4_X1   g587(.A1(new_n658), .A2(new_n621), .A3(new_n426), .A4(new_n724), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n676), .A2(new_n470), .ZN(new_n775));
  XOR2_X1   g589(.A(new_n775), .B(KEYINPUT49), .Z(new_n776));
  NAND4_X1  g590(.A1(new_n774), .A2(new_n604), .A3(new_n665), .A4(new_n776), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n712), .A2(new_n677), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n778), .A2(new_n604), .A3(new_n287), .A4(new_n665), .ZN(new_n779));
  NOR3_X1   g593(.A1(new_n779), .A2(new_n378), .A3(new_n619), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n728), .A2(new_n287), .ZN(new_n781));
  INV_X1    g595(.A(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(new_n699), .ZN(new_n783));
  NOR3_X1   g597(.A1(new_n783), .A2(new_n284), .A3(new_n658), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT111), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n785), .A2(KEYINPUT50), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n784), .B(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n782), .A2(new_n778), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  AOI211_X1 g603(.A(new_n780), .B(new_n787), .C1(new_n703), .C2(new_n789), .ZN(new_n790));
  AOI21_X1  g604(.A(KEYINPUT51), .B1(new_n790), .B2(KEYINPUT110), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n427), .B1(new_n746), .B2(new_n747), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT47), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  OAI211_X1 g608(.A(new_n794), .B(new_n770), .C1(new_n427), .C2(new_n775), .ZN(new_n795));
  NOR3_X1   g609(.A1(new_n781), .A2(new_n527), .A3(new_n698), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n795), .A2(new_n719), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n790), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n791), .A2(new_n798), .ZN(new_n799));
  OAI211_X1 g613(.A(new_n790), .B(new_n797), .C1(KEYINPUT110), .C2(KEYINPUT51), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n423), .A2(new_n476), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n426), .A2(new_n621), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n283), .A2(new_n645), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n802), .A2(new_n690), .A3(new_n803), .A4(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(new_n713), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n805), .B1(new_n806), .B2(new_n698), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(new_n638), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n716), .A2(new_n808), .A3(new_n720), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n630), .A2(new_n620), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n603), .A2(new_n295), .A3(new_n604), .A4(new_n810), .ZN(new_n811));
  AND3_X1   g625(.A1(new_n811), .A2(new_n639), .A3(new_n597), .ZN(new_n812));
  AND2_X1   g626(.A1(new_n683), .A2(new_n701), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n812), .A2(new_n693), .A3(new_n679), .A4(new_n813), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n809), .A2(new_n814), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n523), .A2(new_n524), .A3(new_n637), .A4(new_n670), .ZN(new_n816));
  XOR2_X1   g630(.A(new_n816), .B(KEYINPUT104), .Z(new_n817));
  INV_X1    g631(.A(KEYINPUT105), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n817), .A2(new_n818), .A3(new_n718), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n816), .B(KEYINPUT104), .ZN(new_n820));
  OAI21_X1  g634(.A(KEYINPUT105), .B1(new_n820), .B2(new_n711), .ZN(new_n821));
  INV_X1    g635(.A(new_n665), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n666), .A2(new_n647), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n819), .A2(new_n821), .A3(new_n822), .A4(new_n823), .ZN(new_n824));
  AND3_X1   g638(.A1(new_n649), .A2(new_n673), .A3(new_n704), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT52), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n824), .A2(new_n825), .A3(KEYINPUT52), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n815), .A2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT53), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n815), .A2(new_n830), .A3(KEYINPUT53), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n833), .A2(KEYINPUT106), .A3(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT106), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n831), .A2(new_n836), .A3(new_n832), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n835), .A2(KEYINPUT54), .A3(new_n837), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n693), .A2(KEYINPUT108), .A3(new_n679), .A4(new_n813), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n839), .A2(new_n812), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n693), .A2(new_n679), .A3(new_n813), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT108), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n832), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(new_n809), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n840), .A2(new_n830), .A3(new_n843), .A4(new_n844), .ZN(new_n845));
  XNOR2_X1  g659(.A(KEYINPUT109), .B(KEYINPUT54), .ZN(new_n846));
  INV_X1    g660(.A(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT107), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n848), .B1(new_n831), .B2(new_n832), .ZN(new_n849));
  AOI211_X1 g663(.A(KEYINPUT107), .B(KEYINPUT53), .C1(new_n815), .C2(new_n830), .ZN(new_n850));
  OAI211_X1 g664(.A(new_n845), .B(new_n847), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n789), .A2(KEYINPUT48), .A3(new_n596), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT48), .ZN(new_n853));
  INV_X1    g667(.A(new_n596), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n853), .B1(new_n788), .B2(new_n854), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n838), .A2(new_n851), .A3(new_n852), .A4(new_n855), .ZN(new_n856));
  OAI211_X1 g670(.A(G952), .B(new_n247), .C1(new_n779), .C2(new_n620), .ZN(new_n857));
  INV_X1    g671(.A(new_n783), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n857), .B1(new_n858), .B2(new_n622), .ZN(new_n859));
  XNOR2_X1  g673(.A(new_n859), .B(KEYINPUT112), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n801), .A2(new_n856), .A3(new_n860), .ZN(new_n861));
  NOR2_X1   g675(.A1(G952), .A2(G953), .ZN(new_n862));
  XOR2_X1   g676(.A(new_n862), .B(KEYINPUT113), .Z(new_n863));
  OAI21_X1  g677(.A(new_n777), .B1(new_n861), .B2(new_n863), .ZN(G75));
  OAI21_X1  g678(.A(new_n845), .B1(new_n849), .B2(new_n850), .ZN(new_n865));
  AND2_X1   g679(.A1(new_n865), .A2(G902), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(G210), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT56), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n268), .A2(new_n271), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n869), .B(new_n269), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n870), .B(KEYINPUT55), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n867), .A2(new_n868), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n871), .B1(new_n867), .B2(new_n868), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n247), .A2(G952), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n874), .B(KEYINPUT114), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n872), .A2(new_n873), .A3(new_n875), .ZN(G51));
  NAND2_X1  g690(.A1(new_n865), .A2(new_n846), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT115), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n877), .A2(new_n878), .A3(new_n851), .ZN(new_n879));
  OR3_X1    g693(.A1(new_n865), .A2(new_n878), .A3(new_n846), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n471), .B(KEYINPUT57), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(new_n468), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n866), .A2(new_n743), .A3(new_n741), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n874), .B1(new_n883), .B2(new_n884), .ZN(G54));
  NAND4_X1  g699(.A1(new_n865), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT116), .ZN(new_n887));
  AND3_X1   g701(.A1(new_n886), .A2(new_n887), .A3(new_n365), .ZN(new_n888));
  INV_X1    g702(.A(new_n874), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n889), .B1(new_n886), .B2(new_n365), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n887), .B1(new_n886), .B2(new_n365), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n888), .A2(new_n890), .A3(new_n891), .ZN(G60));
  NAND2_X1  g706(.A1(new_n609), .A2(new_n614), .ZN(new_n893));
  INV_X1    g707(.A(new_n893), .ZN(new_n894));
  XOR2_X1   g708(.A(new_n618), .B(KEYINPUT59), .Z(new_n895));
  AND4_X1   g709(.A1(new_n894), .A2(new_n879), .A3(new_n880), .A4(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n838), .A2(new_n851), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n894), .B1(new_n897), .B2(new_n895), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n896), .A2(new_n875), .A3(new_n898), .ZN(G63));
  NAND2_X1  g713(.A1(G217), .A2(G902), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n900), .B(KEYINPUT117), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(KEYINPUT60), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n516), .B1(new_n865), .B2(new_n902), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n903), .A2(new_n875), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n865), .A2(new_n636), .A3(new_n902), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n905), .A2(KEYINPUT118), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT118), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n865), .A2(new_n907), .A3(new_n636), .A4(new_n902), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n904), .A2(new_n906), .A3(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT61), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n904), .A2(new_n906), .A3(KEYINPUT61), .A4(new_n908), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n911), .A2(new_n912), .ZN(G66));
  NAND2_X1  g727(.A1(new_n814), .A2(new_n247), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n914), .B(KEYINPUT119), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n247), .B1(new_n288), .B2(G224), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n869), .B1(G898), .B2(new_n247), .ZN(new_n918));
  XOR2_X1   g732(.A(new_n917), .B(new_n918), .Z(G69));
  OAI21_X1  g733(.A(G953), .B1(new_n430), .B2(new_n644), .ZN(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT125), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n757), .A2(new_n758), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n768), .A2(new_n659), .A3(new_n719), .A4(new_n733), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n825), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n925), .A2(KEYINPUT123), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT123), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n759), .A2(new_n927), .A3(new_n825), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n720), .B1(new_n714), .B2(new_n715), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(KEYINPUT124), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT124), .ZN(new_n932));
  OAI211_X1 g746(.A(new_n932), .B(new_n720), .C1(new_n714), .C2(new_n715), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n768), .A2(new_n596), .A3(new_n659), .A4(new_n823), .ZN(new_n935));
  AND3_X1   g749(.A1(new_n934), .A2(new_n772), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g750(.A(G953), .B1(new_n929), .B2(new_n936), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n247), .A2(G900), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n922), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n556), .A2(new_n557), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n306), .A2(new_n307), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n940), .B(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(new_n938), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n934), .A2(new_n772), .A3(new_n935), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n944), .B1(new_n926), .B2(new_n928), .ZN(new_n945));
  OAI211_X1 g759(.A(KEYINPUT125), .B(new_n943), .C1(new_n945), .C2(G953), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n939), .A2(new_n942), .A3(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT122), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n668), .A2(new_n825), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT62), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n668), .A2(new_n825), .A3(KEYINPUT62), .ZN(new_n952));
  INV_X1    g766(.A(new_n761), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n953), .B1(new_n794), .B2(new_n770), .ZN(new_n954));
  AOI22_X1  g768(.A1(new_n951), .A2(new_n952), .B1(new_n954), .B2(new_n762), .ZN(new_n955));
  INV_X1    g769(.A(new_n660), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n596), .A2(new_n956), .A3(new_n719), .A4(new_n810), .ZN(new_n957));
  AND3_X1   g771(.A1(new_n759), .A2(KEYINPUT120), .A3(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(KEYINPUT120), .B1(new_n759), .B2(new_n957), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n955), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n960), .A2(KEYINPUT121), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT121), .ZN(new_n962));
  OAI211_X1 g776(.A(new_n955), .B(new_n962), .C1(new_n958), .C2(new_n959), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n942), .A2(G953), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  AND3_X1   g780(.A1(new_n947), .A2(new_n948), .A3(new_n966), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n948), .B1(new_n947), .B2(new_n966), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n921), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n947), .A2(new_n966), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n970), .A2(KEYINPUT122), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n947), .A2(new_n966), .A3(new_n948), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n971), .A2(new_n920), .A3(new_n972), .ZN(new_n973));
  AND2_X1   g787(.A1(new_n969), .A2(new_n973), .ZN(G72));
  NAND2_X1  g788(.A1(G472), .A2(G902), .ZN(new_n975));
  XOR2_X1   g789(.A(new_n975), .B(KEYINPUT63), .Z(new_n976));
  NAND2_X1  g790(.A1(new_n561), .A2(new_n581), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n835), .A2(new_n837), .A3(new_n976), .A4(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n929), .A2(new_n936), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n976), .B1(new_n979), .B2(new_n814), .ZN(new_n980));
  INV_X1    g794(.A(new_n559), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n980), .A2(new_n560), .A3(new_n981), .ZN(new_n982));
  AND3_X1   g796(.A1(new_n982), .A2(KEYINPUT127), .A3(new_n889), .ZN(new_n983));
  AOI21_X1  g797(.A(KEYINPUT127), .B1(new_n982), .B2(new_n889), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n978), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  INV_X1    g799(.A(new_n814), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n961), .A2(new_n986), .A3(new_n963), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n981), .B1(new_n987), .B2(new_n976), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n988), .A2(new_n553), .ZN(new_n989));
  OR2_X1    g803(.A1(new_n989), .A2(KEYINPUT126), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n989), .A2(KEYINPUT126), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n985), .B1(new_n990), .B2(new_n991), .ZN(G57));
endmodule


