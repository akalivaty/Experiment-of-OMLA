//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 0 0 0 0 0 1 1 1 1 1 1 1 1 1 1 0 0 0 0 0 1 1 1 0 0 0 1 0 1 1 1 0 1 1 0 0 1 1 0 1 0 0 1 0 1 0 0 0 1 0 1 1 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n720, new_n721, new_n722, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n730, new_n731, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n741, new_n742,
    new_n743, new_n744, new_n746, new_n747, new_n748, new_n750, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n791, new_n792, new_n793, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n849, new_n850, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n858, new_n859, new_n860, new_n861, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n919, new_n920, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n931, new_n932, new_n933, new_n934,
    new_n936, new_n937, new_n938, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n960,
    new_n961;
  INV_X1    g000(.A(KEYINPUT88), .ZN(new_n202));
  INV_X1    g001(.A(G29gat), .ZN(new_n203));
  INV_X1    g002(.A(G36gat), .ZN(new_n204));
  NAND4_X1  g003(.A1(new_n202), .A2(new_n203), .A3(new_n204), .A4(KEYINPUT14), .ZN(new_n205));
  NAND3_X1  g004(.A1(KEYINPUT89), .A2(G29gat), .A3(G36gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(G29gat), .A2(G36gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT89), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  AND3_X1   g008(.A1(new_n205), .A2(new_n206), .A3(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(G43gat), .B(G50gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(KEYINPUT15), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT15), .ZN(new_n213));
  INV_X1    g012(.A(G50gat), .ZN(new_n214));
  AND2_X1   g013(.A1(new_n214), .A2(G43gat), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n214), .A2(G43gat), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n213), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n202), .A2(KEYINPUT14), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT14), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(KEYINPUT88), .ZN(new_n220));
  OAI211_X1 g019(.A(new_n218), .B(new_n220), .C1(G29gat), .C2(G36gat), .ZN(new_n221));
  NAND4_X1  g020(.A1(new_n210), .A2(new_n212), .A3(new_n217), .A4(new_n221), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n205), .A2(new_n206), .A3(new_n209), .ZN(new_n223));
  OAI22_X1  g022(.A1(new_n219), .A2(KEYINPUT88), .B1(G29gat), .B2(G36gat), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n202), .A2(KEYINPUT14), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI211_X1 g025(.A(KEYINPUT15), .B(new_n211), .C1(new_n223), .C2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n222), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT17), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(G15gat), .B(G22gat), .ZN(new_n231));
  INV_X1    g030(.A(G1gat), .ZN(new_n232));
  AND2_X1   g031(.A1(new_n232), .A2(KEYINPUT16), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n231), .A2(new_n232), .ZN(new_n236));
  OAI211_X1 g035(.A(KEYINPUT90), .B(G8gat), .C1(new_n235), .C2(new_n236), .ZN(new_n237));
  OR2_X1    g036(.A1(new_n231), .A2(new_n232), .ZN(new_n238));
  NAND2_X1  g037(.A1(KEYINPUT90), .A2(G8gat), .ZN(new_n239));
  OR2_X1    g038(.A1(KEYINPUT90), .A2(G8gat), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n238), .A2(new_n234), .A3(new_n239), .A4(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n237), .A2(new_n241), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n222), .A2(KEYINPUT17), .A3(new_n227), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n230), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(G229gat), .A2(G233gat), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n228), .A2(new_n237), .A3(new_n241), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n244), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT18), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n242), .A2(new_n227), .A3(new_n222), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n250), .A2(new_n246), .A3(KEYINPUT91), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n245), .B(KEYINPUT13), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT91), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n242), .A2(new_n254), .A3(new_n227), .A4(new_n222), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n251), .A2(new_n253), .A3(new_n255), .ZN(new_n256));
  NAND4_X1  g055(.A1(new_n244), .A2(KEYINPUT18), .A3(new_n245), .A4(new_n246), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n249), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  XNOR2_X1  g057(.A(KEYINPUT11), .B(G169gat), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n259), .B(G197gat), .ZN(new_n260));
  XNOR2_X1  g059(.A(G113gat), .B(G141gat), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n260), .B(new_n261), .ZN(new_n262));
  XOR2_X1   g061(.A(new_n262), .B(KEYINPUT12), .Z(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n258), .A2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT92), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n258), .A2(KEYINPUT92), .A3(new_n264), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n249), .A2(new_n263), .A3(new_n256), .A4(new_n257), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT93), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n270), .B(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n269), .A2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(KEYINPUT0), .B(G57gat), .ZN(new_n275));
  INV_X1    g074(.A(G85gat), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n275), .B(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(G1gat), .B(G29gat), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n277), .B(new_n278), .ZN(new_n279));
  XOR2_X1   g078(.A(G141gat), .B(G148gat), .Z(new_n280));
  INV_X1    g079(.A(G155gat), .ZN(new_n281));
  INV_X1    g080(.A(G162gat), .ZN(new_n282));
  OAI21_X1  g081(.A(KEYINPUT2), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n280), .A2(new_n283), .ZN(new_n284));
  XNOR2_X1  g083(.A(G155gat), .B(G162gat), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(G113gat), .ZN(new_n288));
  OAI21_X1  g087(.A(KEYINPUT72), .B1(new_n288), .B2(G120gat), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT72), .ZN(new_n290));
  INV_X1    g089(.A(G120gat), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n290), .A2(new_n291), .A3(G113gat), .ZN(new_n292));
  OAI211_X1 g091(.A(new_n289), .B(new_n292), .C1(G113gat), .C2(new_n291), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT1), .ZN(new_n294));
  XNOR2_X1  g093(.A(G127gat), .B(G134gat), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n293), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n280), .A2(new_n285), .A3(new_n283), .ZN(new_n297));
  INV_X1    g096(.A(new_n295), .ZN(new_n298));
  XNOR2_X1  g097(.A(G113gat), .B(G120gat), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n298), .B1(KEYINPUT1), .B2(new_n299), .ZN(new_n300));
  NAND4_X1  g099(.A1(new_n287), .A2(new_n296), .A3(new_n297), .A4(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT78), .ZN(new_n302));
  OR3_X1    g101(.A1(new_n301), .A2(new_n302), .A3(KEYINPUT4), .ZN(new_n303));
  XNOR2_X1  g102(.A(KEYINPUT77), .B(KEYINPUT4), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n302), .B1(new_n301), .B2(KEYINPUT4), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n303), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(G225gat), .A2(G233gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n287), .A2(new_n297), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT3), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n300), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n309), .A2(KEYINPUT3), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n312), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n307), .A2(new_n308), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n309), .A2(new_n313), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n308), .B1(new_n317), .B2(new_n301), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT5), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n320), .A2(KEYINPUT79), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT79), .ZN(new_n322));
  NOR3_X1   g121(.A1(new_n318), .A2(new_n322), .A3(new_n319), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n316), .B1(new_n321), .B2(new_n323), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n315), .A2(KEYINPUT4), .A3(new_n301), .ZN(new_n325));
  OR2_X1    g124(.A1(new_n301), .A2(new_n304), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n327), .A2(new_n319), .A3(new_n308), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n279), .B1(new_n324), .B2(new_n328), .ZN(new_n329));
  XNOR2_X1  g128(.A(KEYINPUT80), .B(KEYINPUT6), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n324), .A2(new_n328), .A3(new_n279), .ZN(new_n332));
  INV_X1    g131(.A(new_n330), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n331), .B1(new_n334), .B2(new_n329), .ZN(new_n335));
  XNOR2_X1  g134(.A(G211gat), .B(G218gat), .ZN(new_n336));
  OR2_X1    g135(.A1(new_n336), .A2(KEYINPUT73), .ZN(new_n337));
  XNOR2_X1  g136(.A(G197gat), .B(G204gat), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT22), .ZN(new_n339));
  INV_X1    g138(.A(G211gat), .ZN(new_n340));
  INV_X1    g139(.A(G218gat), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n339), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n338), .A2(new_n342), .ZN(new_n343));
  XNOR2_X1  g142(.A(new_n337), .B(new_n343), .ZN(new_n344));
  XOR2_X1   g143(.A(KEYINPUT67), .B(G176gat), .Z(new_n345));
  XNOR2_X1  g144(.A(KEYINPUT66), .B(G169gat), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n345), .A2(KEYINPUT23), .A3(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT25), .ZN(new_n348));
  NAND2_X1  g147(.A1(G169gat), .A2(G176gat), .ZN(new_n349));
  AND3_X1   g148(.A1(new_n347), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(G169gat), .ZN(new_n351));
  INV_X1    g150(.A(G176gat), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT23), .ZN(new_n354));
  AND2_X1   g153(.A1(new_n354), .A2(KEYINPUT68), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n354), .A2(KEYINPUT68), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n353), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(G183gat), .A2(G190gat), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT24), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NOR2_X1   g159(.A1(G183gat), .A2(G190gat), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  AOI21_X1  g161(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n363));
  OR2_X1    g162(.A1(new_n363), .A2(KEYINPUT64), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(KEYINPUT64), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n362), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT65), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND4_X1  g167(.A1(new_n362), .A2(new_n364), .A3(KEYINPUT65), .A4(new_n365), .ZN(new_n369));
  NAND4_X1  g168(.A1(new_n350), .A2(new_n357), .A3(new_n368), .A4(new_n369), .ZN(new_n370));
  OR3_X1    g169(.A1(new_n360), .A2(new_n361), .A3(new_n363), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n351), .A2(new_n352), .A3(KEYINPUT23), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n371), .A2(new_n349), .A3(new_n372), .A4(new_n357), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(KEYINPUT25), .ZN(new_n374));
  XNOR2_X1  g173(.A(KEYINPUT27), .B(G183gat), .ZN(new_n375));
  INV_X1    g174(.A(G190gat), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n375), .A2(KEYINPUT28), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(KEYINPUT70), .ZN(new_n378));
  INV_X1    g177(.A(G183gat), .ZN(new_n379));
  OAI21_X1  g178(.A(KEYINPUT27), .B1(new_n379), .B2(KEYINPUT69), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT27), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(G183gat), .ZN(new_n382));
  OAI211_X1 g181(.A(new_n380), .B(new_n376), .C1(KEYINPUT69), .C2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT28), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT70), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n375), .A2(new_n386), .A3(KEYINPUT28), .A4(new_n376), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n378), .A2(new_n385), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n353), .A2(KEYINPUT26), .ZN(new_n389));
  OR3_X1    g188(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n389), .A2(new_n390), .A3(new_n349), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(new_n358), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT71), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n391), .A2(KEYINPUT71), .A3(new_n358), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n388), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n370), .A2(new_n374), .A3(new_n396), .ZN(new_n397));
  AND3_X1   g196(.A1(new_n397), .A2(G226gat), .A3(G233gat), .ZN(new_n398));
  NAND2_X1  g197(.A1(G226gat), .A2(G233gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n399), .B(KEYINPUT74), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT29), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n401), .B1(new_n397), .B2(new_n402), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n344), .B1(new_n398), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n397), .A2(new_n402), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(new_n399), .ZN(new_n406));
  INV_X1    g205(.A(new_n343), .ZN(new_n407));
  XNOR2_X1  g206(.A(new_n407), .B(new_n337), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n397), .A2(new_n401), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n406), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n404), .A2(new_n410), .ZN(new_n411));
  XOR2_X1   g210(.A(G8gat), .B(G36gat), .Z(new_n412));
  XNOR2_X1  g211(.A(new_n412), .B(G64gat), .ZN(new_n413));
  INV_X1    g212(.A(G92gat), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n413), .B(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n411), .A2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n415), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n404), .A2(new_n410), .A3(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT30), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  OAI21_X1  g220(.A(KEYINPUT75), .B1(new_n417), .B2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT76), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n419), .A2(new_n423), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n404), .A2(new_n410), .A3(KEYINPUT76), .A4(new_n418), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n424), .A2(new_n420), .A3(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT75), .ZN(new_n427));
  OAI211_X1 g226(.A(new_n416), .B(new_n427), .C1(new_n420), .C2(new_n419), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n335), .A2(new_n422), .A3(new_n426), .A4(new_n428), .ZN(new_n429));
  XNOR2_X1  g228(.A(G78gat), .B(G106gat), .ZN(new_n430));
  INV_X1    g229(.A(G22gat), .ZN(new_n431));
  XNOR2_X1  g230(.A(new_n430), .B(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n344), .A2(KEYINPUT29), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n311), .B1(new_n434), .B2(KEYINPUT82), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n408), .A2(new_n402), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT82), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n309), .B1(new_n435), .B2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT83), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  OAI211_X1 g240(.A(KEYINPUT83), .B(new_n309), .C1(new_n435), .C2(new_n438), .ZN(new_n442));
  INV_X1    g241(.A(G228gat), .ZN(new_n443));
  INV_X1    g242(.A(G233gat), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n408), .B1(new_n312), .B2(new_n402), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n441), .A2(new_n442), .A3(new_n445), .A4(new_n447), .ZN(new_n448));
  OR2_X1    g247(.A1(new_n343), .A2(new_n336), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n343), .A2(new_n336), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n449), .A2(new_n402), .A3(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n310), .B1(new_n451), .B2(new_n311), .ZN(new_n452));
  OAI22_X1  g251(.A1(new_n446), .A2(new_n452), .B1(new_n443), .B2(new_n444), .ZN(new_n453));
  XNOR2_X1  g252(.A(new_n453), .B(KEYINPUT81), .ZN(new_n454));
  XNOR2_X1  g253(.A(KEYINPUT31), .B(G50gat), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n448), .A2(new_n454), .A3(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n456), .B1(new_n448), .B2(new_n454), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n433), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n448), .A2(new_n454), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(new_n455), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n462), .A2(new_n432), .A3(new_n457), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n460), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n429), .A2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT36), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT34), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n397), .A2(new_n300), .A3(new_n296), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n370), .A2(new_n396), .A3(new_n313), .A4(new_n374), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(G227gat), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n471), .A2(new_n444), .ZN(new_n472));
  INV_X1    g271(.A(new_n472), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n467), .B1(new_n470), .B2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  AOI211_X1 g274(.A(KEYINPUT34), .B(new_n472), .C1(new_n468), .C2(new_n469), .ZN(new_n476));
  INV_X1    g275(.A(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n468), .A2(new_n472), .A3(new_n469), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(KEYINPUT32), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n475), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  OAI211_X1 g279(.A(KEYINPUT32), .B(new_n478), .C1(new_n474), .C2(new_n476), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT33), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n478), .A2(new_n482), .ZN(new_n483));
  XNOR2_X1  g282(.A(G15gat), .B(G43gat), .ZN(new_n484));
  XNOR2_X1  g283(.A(G71gat), .B(G99gat), .ZN(new_n485));
  XOR2_X1   g284(.A(new_n484), .B(new_n485), .Z(new_n486));
  NAND2_X1  g285(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  AND3_X1   g287(.A1(new_n480), .A2(new_n481), .A3(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n488), .B1(new_n480), .B2(new_n481), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n466), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n480), .A2(new_n481), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(new_n487), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n480), .A2(new_n481), .A3(new_n488), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n493), .A2(KEYINPUT36), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n491), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n465), .A2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT84), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  XOR2_X1   g298(.A(new_n279), .B(KEYINPUT85), .Z(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  OR2_X1    g300(.A1(new_n327), .A2(new_n308), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n317), .A2(new_n308), .A3(new_n301), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(KEYINPUT39), .ZN(new_n504));
  XNOR2_X1  g303(.A(new_n504), .B(KEYINPUT86), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n501), .B1(new_n502), .B2(new_n505), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n506), .B1(KEYINPUT39), .B2(new_n502), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT40), .ZN(new_n508));
  OR2_X1    g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n417), .A2(new_n421), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(new_n426), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n324), .A2(new_n328), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(new_n501), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n507), .A2(new_n508), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n509), .A2(new_n511), .A3(new_n513), .A4(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n464), .ZN(new_n516));
  INV_X1    g315(.A(new_n334), .ZN(new_n517));
  AOI22_X1  g316(.A1(new_n517), .A2(new_n513), .B1(new_n329), .B2(new_n330), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT37), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n519), .B1(new_n404), .B2(new_n410), .ZN(new_n520));
  NAND4_X1  g319(.A1(new_n404), .A2(new_n410), .A3(KEYINPUT87), .A4(new_n519), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT87), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n522), .B1(new_n411), .B2(KEYINPUT37), .ZN(new_n523));
  AOI211_X1 g322(.A(new_n418), .B(new_n520), .C1(new_n521), .C2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT38), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n518), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n418), .B1(new_n523), .B2(new_n521), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n408), .B1(new_n398), .B2(new_n403), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n406), .A2(new_n344), .A3(new_n409), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n528), .A2(new_n529), .A3(KEYINPUT37), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n527), .A2(new_n525), .A3(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n531), .A2(new_n424), .A3(new_n425), .ZN(new_n532));
  OAI211_X1 g331(.A(new_n515), .B(new_n516), .C1(new_n526), .C2(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n465), .A2(KEYINPUT84), .A3(new_n496), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n499), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n489), .A2(new_n490), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n536), .A2(new_n463), .A3(new_n460), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  NOR3_X1   g337(.A1(new_n518), .A2(new_n511), .A3(KEYINPUT35), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  OAI21_X1  g339(.A(KEYINPUT35), .B1(new_n537), .B2(new_n429), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n274), .B1(new_n535), .B2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT21), .ZN(new_n544));
  NAND2_X1  g343(.A1(G71gat), .A2(G78gat), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT9), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  OR2_X1    g346(.A1(G57gat), .A2(G64gat), .ZN(new_n548));
  NAND2_X1  g347(.A1(G57gat), .A2(G64gat), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT94), .ZN(new_n551));
  XNOR2_X1  g350(.A(G71gat), .B(G78gat), .ZN(new_n552));
  AND3_X1   g351(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n552), .B1(new_n550), .B2(new_n551), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n242), .B1(new_n544), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(G183gat), .ZN(new_n557));
  OAI211_X1 g356(.A(new_n242), .B(new_n379), .C1(new_n544), .C2(new_n555), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(G57gat), .B(G64gat), .ZN(new_n560));
  AOI21_X1  g359(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n551), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n552), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(KEYINPUT95), .B(KEYINPUT21), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n559), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n566), .A2(new_n567), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n557), .A2(new_n558), .A3(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(G127gat), .B(G155gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n571), .B(G211gat), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  AND3_X1   g372(.A1(new_n568), .A2(new_n570), .A3(new_n573), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n573), .B1(new_n568), .B2(new_n570), .ZN(new_n575));
  XNOR2_X1  g374(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n576));
  NAND2_X1  g375(.A1(G231gat), .A2(G233gat), .ZN(new_n577));
  XOR2_X1   g376(.A(new_n576), .B(new_n577), .Z(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  OR3_X1    g378(.A1(new_n574), .A2(new_n575), .A3(new_n579), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n579), .B1(new_n574), .B2(new_n575), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT101), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT99), .ZN(new_n584));
  XNOR2_X1  g383(.A(G99gat), .B(G106gat), .ZN(new_n585));
  NAND2_X1  g384(.A1(G99gat), .A2(G106gat), .ZN(new_n586));
  AOI22_X1  g385(.A1(KEYINPUT8), .A2(new_n586), .B1(new_n276), .B2(new_n414), .ZN(new_n587));
  NAND3_X1  g386(.A1(KEYINPUT98), .A2(G85gat), .A3(G92gat), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT7), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n588), .A2(KEYINPUT97), .A3(new_n589), .ZN(new_n590));
  AND2_X1   g389(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n588), .A2(KEYINPUT97), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT97), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n593), .A2(G85gat), .A3(G92gat), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n592), .A2(KEYINPUT7), .A3(new_n594), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n585), .B1(new_n591), .B2(new_n595), .ZN(new_n596));
  AND4_X1   g395(.A1(new_n585), .A2(new_n595), .A3(new_n590), .A4(new_n587), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n584), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n595), .A2(new_n590), .A3(new_n587), .ZN(new_n599));
  INV_X1    g398(.A(new_n585), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n591), .A2(new_n585), .A3(new_n595), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n601), .A2(new_n602), .A3(KEYINPUT99), .ZN(new_n603));
  NAND4_X1  g402(.A1(new_n230), .A2(new_n598), .A3(new_n243), .A4(new_n603), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n596), .A2(new_n597), .ZN(new_n605));
  AND2_X1   g404(.A1(G232gat), .A2(G233gat), .ZN(new_n606));
  AOI22_X1  g405(.A1(new_n605), .A2(new_n228), .B1(KEYINPUT41), .B2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT100), .ZN(new_n608));
  AND3_X1   g407(.A1(new_n604), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n608), .B1(new_n604), .B2(new_n607), .ZN(new_n610));
  OAI21_X1  g409(.A(G190gat), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n604), .A2(new_n607), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n612), .A2(KEYINPUT100), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n604), .A2(new_n607), .A3(new_n608), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n613), .A2(new_n376), .A3(new_n614), .ZN(new_n615));
  AND3_X1   g414(.A1(new_n611), .A2(new_n615), .A3(G218gat), .ZN(new_n616));
  AOI21_X1  g415(.A(G218gat), .B1(new_n611), .B2(new_n615), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n583), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NOR3_X1   g417(.A1(new_n609), .A2(new_n610), .A3(G190gat), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n376), .B1(new_n613), .B2(new_n614), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n341), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n611), .A2(new_n615), .A3(G218gat), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n621), .A2(KEYINPUT101), .A3(new_n622), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n606), .A2(KEYINPUT41), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(KEYINPUT96), .ZN(new_n625));
  XNOR2_X1  g424(.A(G134gat), .B(G162gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n618), .A2(new_n623), .A3(new_n628), .ZN(new_n629));
  NAND4_X1  g428(.A1(new_n621), .A2(KEYINPUT101), .A3(new_n622), .A4(new_n627), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n582), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  XOR2_X1   g430(.A(KEYINPUT105), .B(G148gat), .Z(new_n632));
  XNOR2_X1  g431(.A(G176gat), .B(G204gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(KEYINPUT104), .B(G120gat), .ZN(new_n635));
  XOR2_X1   g434(.A(new_n634), .B(new_n635), .Z(new_n636));
  OAI21_X1  g435(.A(new_n555), .B1(new_n597), .B2(new_n596), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n566), .A2(new_n602), .A3(new_n601), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n637), .A2(KEYINPUT102), .A3(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT102), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n605), .A2(new_n640), .A3(new_n566), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT10), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n644), .A2(KEYINPUT103), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n638), .A2(new_n643), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT103), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n642), .A2(new_n648), .A3(new_n643), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n645), .A2(new_n647), .A3(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(G230gat), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n651), .A2(new_n444), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n650), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n642), .A2(new_n653), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n636), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n648), .B1(new_n642), .B2(new_n643), .ZN(new_n658));
  AOI211_X1 g457(.A(KEYINPUT103), .B(KEYINPUT10), .C1(new_n639), .C2(new_n641), .ZN(new_n659));
  NOR3_X1   g458(.A1(new_n658), .A2(new_n659), .A3(new_n646), .ZN(new_n660));
  OAI211_X1 g459(.A(new_n656), .B(new_n636), .C1(new_n660), .C2(new_n652), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n661), .A2(KEYINPUT106), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n655), .B1(new_n650), .B2(new_n653), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT106), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n663), .A2(new_n664), .A3(new_n636), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n657), .B1(new_n662), .B2(new_n665), .ZN(new_n666));
  AND2_X1   g465(.A1(new_n631), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n543), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n668), .A2(new_n335), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(new_n232), .ZN(G1324gat));
  INV_X1    g469(.A(new_n668), .ZN(new_n671));
  NAND2_X1  g470(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n672));
  OR2_X1    g471(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n673));
  NAND4_X1  g472(.A1(new_n671), .A2(new_n511), .A3(new_n672), .A4(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT42), .ZN(new_n675));
  OR2_X1    g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n511), .ZN(new_n677));
  OAI21_X1  g476(.A(G8gat), .B1(new_n668), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n674), .A2(new_n675), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n676), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT107), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n680), .B(new_n681), .ZN(G1325gat));
  AOI21_X1  g481(.A(G15gat), .B1(new_n671), .B2(new_n536), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n683), .B(KEYINPUT108), .ZN(new_n684));
  INV_X1    g483(.A(new_n496), .ZN(new_n685));
  AND2_X1   g484(.A1(new_n685), .A2(G15gat), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n684), .B1(new_n671), .B2(new_n686), .ZN(G1326gat));
  NOR2_X1   g486(.A1(new_n668), .A2(new_n516), .ZN(new_n688));
  XOR2_X1   g487(.A(KEYINPUT43), .B(G22gat), .Z(new_n689));
  XNOR2_X1  g488(.A(new_n688), .B(new_n689), .ZN(G1327gat));
  NAND2_X1  g489(.A1(new_n629), .A2(new_n630), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n691), .B1(new_n535), .B2(new_n542), .ZN(new_n692));
  INV_X1    g491(.A(new_n657), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n661), .A2(KEYINPUT106), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n664), .B1(new_n663), .B2(new_n636), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n693), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n582), .ZN(new_n697));
  NOR3_X1   g496(.A1(new_n696), .A2(new_n697), .A3(new_n274), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n692), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n335), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n700), .A2(new_n203), .A3(new_n701), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(KEYINPUT45), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n535), .A2(new_n542), .ZN(new_n704));
  INV_X1    g503(.A(new_n691), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n704), .A2(KEYINPUT44), .A3(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT44), .ZN(new_n707));
  AND2_X1   g506(.A1(new_n465), .A2(new_n496), .ZN(new_n708));
  AOI22_X1  g507(.A1(new_n533), .A2(new_n708), .B1(new_n540), .B2(new_n541), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n707), .B1(new_n709), .B2(new_n691), .ZN(new_n710));
  AND2_X1   g509(.A1(new_n706), .A2(new_n710), .ZN(new_n711));
  AND3_X1   g510(.A1(new_n269), .A2(new_n272), .A3(KEYINPUT109), .ZN(new_n712));
  AOI21_X1  g511(.A(KEYINPUT109), .B1(new_n269), .B2(new_n272), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n696), .A2(new_n697), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n711), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(G29gat), .B1(new_n717), .B2(new_n335), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n703), .A2(new_n718), .ZN(G1328gat));
  NOR3_X1   g518(.A1(new_n699), .A2(G36gat), .A3(new_n677), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(KEYINPUT46), .ZN(new_n721));
  OAI21_X1  g520(.A(G36gat), .B1(new_n717), .B2(new_n677), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(G1329gat));
  OAI21_X1  g522(.A(G43gat), .B1(new_n717), .B2(new_n496), .ZN(new_n724));
  INV_X1    g523(.A(new_n536), .ZN(new_n725));
  OR3_X1    g524(.A1(new_n699), .A2(G43gat), .A3(new_n725), .ZN(new_n726));
  AOI21_X1  g525(.A(KEYINPUT110), .B1(new_n724), .B2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT47), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n727), .B(new_n728), .ZN(G1330gat));
  OAI21_X1  g528(.A(G50gat), .B1(new_n717), .B2(new_n516), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n700), .A2(new_n214), .A3(new_n464), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  XOR2_X1   g531(.A(KEYINPUT111), .B(KEYINPUT48), .Z(new_n733));
  XNOR2_X1  g532(.A(new_n732), .B(new_n733), .ZN(G1331gat));
  NOR3_X1   g533(.A1(new_n709), .A2(new_n582), .A3(new_n705), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n715), .A2(new_n666), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(new_n701), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g539(.A1(new_n737), .A2(new_n677), .ZN(new_n741));
  NOR2_X1   g540(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n742));
  AND2_X1   g541(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n741), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n744), .B1(new_n741), .B2(new_n742), .ZN(G1333gat));
  NAND3_X1  g544(.A1(new_n738), .A2(G71gat), .A3(new_n685), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n737), .A2(new_n725), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n746), .B1(G71gat), .B2(new_n747), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g548(.A1(new_n738), .A2(new_n464), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g550(.A1(new_n715), .A2(new_n697), .A3(new_n666), .ZN(new_n752));
  AND2_X1   g551(.A1(new_n711), .A2(new_n752), .ZN(new_n753));
  AND2_X1   g552(.A1(new_n753), .A2(new_n701), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n708), .A2(new_n533), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(new_n542), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n715), .A2(new_n697), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n756), .A2(new_n705), .A3(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT51), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT113), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n758), .A2(KEYINPUT113), .A3(new_n759), .ZN(new_n763));
  OAI21_X1  g562(.A(KEYINPUT112), .B1(new_n758), .B2(new_n759), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n709), .A2(new_n691), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT112), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n765), .A2(new_n766), .A3(KEYINPUT51), .A4(new_n757), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n762), .A2(new_n763), .A3(new_n764), .A4(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(new_n768), .ZN(new_n769));
  NOR3_X1   g568(.A1(new_n666), .A2(G85gat), .A3(new_n335), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n770), .B(KEYINPUT114), .ZN(new_n771));
  OAI22_X1  g570(.A1(new_n754), .A2(new_n276), .B1(new_n769), .B2(new_n771), .ZN(G1336gat));
  NOR3_X1   g571(.A1(new_n677), .A2(G92gat), .A3(new_n666), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n768), .A2(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT52), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n706), .A2(new_n511), .A3(new_n710), .A4(new_n752), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(G92gat), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n774), .A2(new_n775), .A3(new_n777), .ZN(new_n778));
  AOI21_X1  g577(.A(KEYINPUT51), .B1(new_n765), .B2(new_n757), .ZN(new_n779));
  AND4_X1   g578(.A1(KEYINPUT51), .A2(new_n756), .A3(new_n705), .A4(new_n757), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n773), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n777), .A2(new_n781), .ZN(new_n782));
  AOI21_X1  g581(.A(KEYINPUT115), .B1(new_n782), .B2(KEYINPUT52), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT115), .ZN(new_n784));
  AOI211_X1 g583(.A(new_n784), .B(new_n775), .C1(new_n777), .C2(new_n781), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n778), .B1(new_n783), .B2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT116), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  OAI211_X1 g587(.A(new_n778), .B(KEYINPUT116), .C1(new_n783), .C2(new_n785), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(G1337gat));
  OR4_X1    g589(.A1(G99gat), .A2(new_n769), .A3(new_n725), .A4(new_n666), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n753), .A2(new_n685), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(G99gat), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n791), .A2(new_n793), .ZN(G1338gat));
  NAND2_X1  g593(.A1(new_n753), .A2(new_n464), .ZN(new_n795));
  INV_X1    g594(.A(G106gat), .ZN(new_n796));
  OR2_X1    g595(.A1(new_n796), .A2(KEYINPUT117), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(KEYINPUT117), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n795), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT53), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n516), .A2(G106gat), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n768), .A2(new_n696), .A3(new_n801), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n799), .A2(new_n800), .A3(new_n802), .ZN(new_n803));
  OAI211_X1 g602(.A(new_n696), .B(new_n801), .C1(new_n779), .C2(new_n780), .ZN(new_n804));
  AND2_X1   g603(.A1(new_n799), .A2(new_n804), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n803), .B1(new_n805), .B2(new_n800), .ZN(G1339gat));
  INV_X1    g605(.A(new_n262), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n253), .B1(new_n251), .B2(new_n255), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n245), .B1(new_n244), .B2(new_n246), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n807), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n272), .A2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(new_n811), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n696), .A2(KEYINPUT119), .A3(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT119), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n814), .B1(new_n666), .B2(new_n811), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT55), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n645), .A2(new_n652), .A3(new_n647), .A4(new_n649), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(KEYINPUT54), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n658), .A2(new_n659), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n652), .B1(new_n820), .B2(new_n647), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT54), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n650), .A2(new_n823), .A3(new_n653), .ZN(new_n824));
  INV_X1    g623(.A(new_n636), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n817), .B1(new_n822), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n662), .A2(new_n665), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n654), .A2(KEYINPUT54), .A3(new_n818), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n829), .A2(KEYINPUT55), .A3(new_n825), .A4(new_n824), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n827), .A2(new_n828), .A3(new_n830), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n714), .A2(new_n831), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n691), .B1(new_n816), .B2(new_n832), .ZN(new_n833));
  OR3_X1    g632(.A1(new_n831), .A2(new_n691), .A3(new_n811), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n697), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n631), .A2(new_n714), .A3(new_n666), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(KEYINPUT118), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT118), .ZN(new_n838));
  NAND4_X1  g637(.A1(new_n631), .A2(new_n714), .A3(new_n838), .A4(new_n666), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  OR2_X1    g639(.A1(new_n835), .A2(new_n840), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n841), .A2(new_n538), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n511), .A2(new_n335), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  XOR2_X1   g643(.A(new_n844), .B(KEYINPUT120), .Z(new_n845));
  NAND3_X1  g644(.A1(new_n845), .A2(new_n288), .A3(new_n715), .ZN(new_n846));
  OAI21_X1  g645(.A(G113gat), .B1(new_n844), .B2(new_n274), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(G1340gat));
  NAND3_X1  g647(.A1(new_n845), .A2(new_n291), .A3(new_n696), .ZN(new_n849));
  OAI21_X1  g648(.A(G120gat), .B1(new_n844), .B2(new_n666), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(G1341gat));
  NAND3_X1  g650(.A1(new_n842), .A2(new_n697), .A3(new_n843), .ZN(new_n852));
  INV_X1    g651(.A(G127gat), .ZN(new_n853));
  OR3_X1    g652(.A1(new_n852), .A2(KEYINPUT121), .A3(new_n853), .ZN(new_n854));
  OAI21_X1  g653(.A(KEYINPUT121), .B1(new_n852), .B2(new_n853), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n856), .B1(new_n853), .B2(new_n852), .ZN(G1342gat));
  NOR2_X1   g656(.A1(new_n844), .A2(new_n691), .ZN(new_n858));
  XNOR2_X1  g657(.A(KEYINPUT56), .B(G134gat), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NOR2_X1   g659(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n860), .B1(new_n858), .B2(new_n861), .ZN(G1343gat));
  INV_X1    g661(.A(KEYINPUT123), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT57), .ZN(new_n864));
  OAI211_X1 g663(.A(new_n864), .B(new_n464), .C1(new_n835), .C2(new_n840), .ZN(new_n865));
  INV_X1    g664(.A(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n496), .A2(new_n843), .ZN(new_n867));
  INV_X1    g666(.A(new_n867), .ZN(new_n868));
  AND2_X1   g667(.A1(new_n837), .A2(new_n839), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n696), .A2(new_n812), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n827), .A2(new_n828), .A3(new_n830), .A4(new_n273), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n705), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NOR3_X1   g671(.A1(new_n831), .A2(new_n691), .A3(new_n811), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n582), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n516), .B1(new_n869), .B2(new_n874), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n868), .B1(new_n875), .B2(new_n864), .ZN(new_n876));
  OAI21_X1  g675(.A(KEYINPUT122), .B1(new_n866), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n870), .A2(new_n871), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(new_n691), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n697), .B1(new_n879), .B2(new_n834), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n464), .B1(new_n880), .B2(new_n840), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n867), .B1(new_n881), .B2(KEYINPUT57), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT122), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n882), .A2(new_n883), .A3(new_n865), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n714), .B1(new_n877), .B2(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(G141gat), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n863), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n841), .A2(new_n464), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(new_n868), .ZN(new_n889));
  INV_X1    g688(.A(new_n889), .ZN(new_n890));
  OAI21_X1  g689(.A(KEYINPUT124), .B1(new_n274), .B2(G141gat), .ZN(new_n891));
  OR3_X1    g690(.A1(new_n274), .A2(KEYINPUT124), .A3(G141gat), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n890), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  AND3_X1   g692(.A1(new_n882), .A2(new_n883), .A3(new_n865), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n883), .B1(new_n882), .B2(new_n865), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n715), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n896), .A2(KEYINPUT123), .A3(G141gat), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n887), .A2(new_n893), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(KEYINPUT58), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT58), .ZN(new_n900));
  NOR3_X1   g699(.A1(new_n866), .A2(new_n876), .A3(new_n274), .ZN(new_n901));
  OAI211_X1 g700(.A(new_n893), .B(new_n900), .C1(new_n886), .C2(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n899), .A2(new_n902), .ZN(G1344gat));
  NOR2_X1   g702(.A1(new_n888), .A2(new_n864), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n667), .A2(new_n274), .ZN(new_n905));
  AOI211_X1 g704(.A(KEYINPUT57), .B(new_n516), .C1(new_n874), .C2(new_n905), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(new_n696), .ZN(new_n908));
  XNOR2_X1  g707(.A(KEYINPUT125), .B(KEYINPUT59), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n868), .A2(new_n909), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n894), .A2(new_n895), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n911), .A2(new_n666), .ZN(new_n912));
  OAI22_X1  g711(.A1(new_n908), .A2(new_n910), .B1(new_n912), .B2(KEYINPUT59), .ZN(new_n913));
  AOI21_X1  g712(.A(G148gat), .B1(new_n890), .B2(new_n696), .ZN(new_n914));
  AOI22_X1  g713(.A1(new_n913), .A2(G148gat), .B1(new_n909), .B2(new_n914), .ZN(G1345gat));
  NOR3_X1   g714(.A1(new_n911), .A2(new_n281), .A3(new_n582), .ZN(new_n916));
  AOI21_X1  g715(.A(G155gat), .B1(new_n890), .B2(new_n697), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n916), .A2(new_n917), .ZN(G1346gat));
  NOR3_X1   g717(.A1(new_n911), .A2(new_n282), .A3(new_n691), .ZN(new_n919));
  AOI21_X1  g718(.A(G162gat), .B1(new_n890), .B2(new_n705), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n919), .A2(new_n920), .ZN(G1347gat));
  NOR2_X1   g720(.A1(new_n677), .A2(new_n701), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n842), .A2(new_n922), .ZN(new_n923));
  OAI21_X1  g722(.A(G169gat), .B1(new_n923), .B2(new_n274), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n715), .A2(new_n346), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n924), .B1(new_n923), .B2(new_n925), .ZN(G1348gat));
  NAND3_X1  g725(.A1(new_n842), .A2(new_n696), .A3(new_n922), .ZN(new_n927));
  AOI21_X1  g726(.A(KEYINPUT126), .B1(new_n927), .B2(new_n352), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n927), .A2(new_n345), .ZN(new_n929));
  MUX2_X1   g728(.A(new_n928), .B(KEYINPUT126), .S(new_n929), .Z(G1349gat));
  OAI21_X1  g729(.A(new_n379), .B1(new_n923), .B2(new_n582), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n842), .A2(new_n697), .A3(new_n922), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n931), .B1(new_n932), .B2(new_n375), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT60), .ZN(new_n934));
  XNOR2_X1  g733(.A(new_n933), .B(new_n934), .ZN(G1350gat));
  XNOR2_X1  g734(.A(KEYINPUT61), .B(G190gat), .ZN(new_n936));
  NAND2_X1  g735(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n923), .A2(new_n691), .ZN(new_n938));
  MUX2_X1   g737(.A(new_n936), .B(new_n937), .S(new_n938), .Z(G1351gat));
  NAND2_X1  g738(.A1(new_n922), .A2(new_n496), .ZN(new_n940));
  INV_X1    g739(.A(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n907), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g741(.A(G197gat), .B1(new_n942), .B2(new_n274), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n888), .A2(new_n941), .ZN(new_n944));
  XNOR2_X1  g743(.A(new_n944), .B(KEYINPUT127), .ZN(new_n945));
  INV_X1    g744(.A(G197gat), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n945), .A2(new_n946), .A3(new_n715), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n943), .A2(new_n947), .ZN(G1352gat));
  NOR3_X1   g747(.A1(new_n944), .A2(G204gat), .A3(new_n666), .ZN(new_n949));
  XNOR2_X1  g748(.A(new_n949), .B(KEYINPUT62), .ZN(new_n950));
  OAI21_X1  g749(.A(G204gat), .B1(new_n908), .B2(new_n940), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n950), .A2(new_n951), .ZN(G1353gat));
  NAND3_X1  g751(.A1(new_n945), .A2(new_n340), .A3(new_n697), .ZN(new_n953));
  INV_X1    g752(.A(new_n904), .ZN(new_n954));
  INV_X1    g753(.A(new_n906), .ZN(new_n955));
  NAND4_X1  g754(.A1(new_n954), .A2(new_n697), .A3(new_n955), .A4(new_n941), .ZN(new_n956));
  AND3_X1   g755(.A1(new_n956), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n957));
  AOI21_X1  g756(.A(KEYINPUT63), .B1(new_n956), .B2(G211gat), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n953), .B1(new_n957), .B2(new_n958), .ZN(G1354gat));
  OAI21_X1  g758(.A(G218gat), .B1(new_n942), .B2(new_n691), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n945), .A2(new_n341), .A3(new_n705), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n960), .A2(new_n961), .ZN(G1355gat));
endmodule


