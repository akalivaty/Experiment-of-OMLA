

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XOR2_X1 U554 ( .A(n694), .B(KEYINPUT28), .Z(n522) );
  AND2_X1 U555 ( .A1(n890), .A2(G126), .ZN(n523) );
  XOR2_X1 U556 ( .A(KEYINPUT13), .B(n578), .Z(n524) );
  OR2_X1 U557 ( .A1(n769), .A2(n768), .ZN(n525) );
  AND2_X1 U558 ( .A1(n752), .A2(n1001), .ZN(n526) );
  OR2_X1 U559 ( .A1(n732), .A2(n690), .ZN(n691) );
  OR2_X1 U560 ( .A1(n702), .A2(n701), .ZN(n705) );
  XNOR2_X1 U561 ( .A(n739), .B(KEYINPUT104), .ZN(n740) );
  AND2_X1 U562 ( .A1(n755), .A2(n753), .ZN(n754) );
  NAND2_X1 U563 ( .A1(n770), .A2(n525), .ZN(n771) );
  XOR2_X1 U564 ( .A(G543), .B(KEYINPUT0), .Z(n650) );
  NOR2_X1 U565 ( .A1(G651), .A2(n650), .ZN(n661) );
  NAND2_X1 U566 ( .A1(n581), .A2(n580), .ZN(n999) );
  NAND2_X1 U567 ( .A1(G2105), .A2(G2104), .ZN(n527) );
  XOR2_X2 U568 ( .A(KEYINPUT64), .B(n527), .Z(n891) );
  NAND2_X1 U569 ( .A1(G114), .A2(n891), .ZN(n534) );
  INV_X1 U570 ( .A(G2105), .ZN(n554) );
  AND2_X1 U571 ( .A1(n554), .A2(G2104), .ZN(n894) );
  NAND2_X1 U572 ( .A1(G102), .A2(n894), .ZN(n531) );
  XNOR2_X1 U573 ( .A(KEYINPUT17), .B(KEYINPUT65), .ZN(n529) );
  NOR2_X1 U574 ( .A1(G2104), .A2(G2105), .ZN(n528) );
  XNOR2_X2 U575 ( .A(n529), .B(n528), .ZN(n895) );
  NAND2_X1 U576 ( .A1(G138), .A2(n895), .ZN(n530) );
  NAND2_X1 U577 ( .A1(n531), .A2(n530), .ZN(n532) );
  NOR2_X1 U578 ( .A1(G2104), .A2(n554), .ZN(n890) );
  NOR2_X1 U579 ( .A1(n532), .A2(n523), .ZN(n533) );
  AND2_X2 U580 ( .A1(n534), .A2(n533), .ZN(G164) );
  NOR2_X1 U581 ( .A1(G651), .A2(G543), .ZN(n654) );
  NAND2_X1 U582 ( .A1(n654), .A2(G89), .ZN(n535) );
  XNOR2_X1 U583 ( .A(n535), .B(KEYINPUT4), .ZN(n538) );
  INV_X1 U584 ( .A(G651), .ZN(n541) );
  OR2_X1 U585 ( .A1(n541), .A2(n650), .ZN(n536) );
  XOR2_X2 U586 ( .A(n536), .B(KEYINPUT66), .Z(n657) );
  NAND2_X1 U587 ( .A1(G76), .A2(n657), .ZN(n537) );
  NAND2_X1 U588 ( .A1(n538), .A2(n537), .ZN(n539) );
  XOR2_X1 U589 ( .A(KEYINPUT5), .B(n539), .Z(n549) );
  NAND2_X1 U590 ( .A1(n661), .A2(G51), .ZN(n540) );
  XOR2_X1 U591 ( .A(KEYINPUT77), .B(n540), .Z(n545) );
  NOR2_X1 U592 ( .A1(G543), .A2(n541), .ZN(n543) );
  XNOR2_X1 U593 ( .A(KEYINPUT1), .B(KEYINPUT67), .ZN(n542) );
  XNOR2_X1 U594 ( .A(n543), .B(n542), .ZN(n653) );
  NAND2_X1 U595 ( .A1(n653), .A2(G63), .ZN(n544) );
  NAND2_X1 U596 ( .A1(n545), .A2(n544), .ZN(n547) );
  XOR2_X1 U597 ( .A(KEYINPUT6), .B(KEYINPUT78), .Z(n546) );
  XOR2_X1 U598 ( .A(n547), .B(n546), .Z(n548) );
  NOR2_X1 U599 ( .A1(n549), .A2(n548), .ZN(n551) );
  XNOR2_X1 U600 ( .A(KEYINPUT7), .B(KEYINPUT79), .ZN(n550) );
  XNOR2_X1 U601 ( .A(n551), .B(n550), .ZN(G168) );
  XOR2_X1 U602 ( .A(G168), .B(KEYINPUT8), .Z(n552) );
  XNOR2_X1 U603 ( .A(KEYINPUT80), .B(n552), .ZN(G286) );
  AND2_X1 U604 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U605 ( .A(G132), .ZN(G219) );
  INV_X1 U606 ( .A(G82), .ZN(G220) );
  INV_X1 U607 ( .A(G57), .ZN(G237) );
  INV_X1 U608 ( .A(G108), .ZN(G238) );
  INV_X1 U609 ( .A(G120), .ZN(G236) );
  NAND2_X1 U610 ( .A1(G113), .A2(n891), .ZN(n557) );
  AND2_X1 U611 ( .A1(G101), .A2(G2104), .ZN(n553) );
  NAND2_X1 U612 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U613 ( .A(KEYINPUT23), .B(n555), .Z(n556) );
  NAND2_X1 U614 ( .A1(n557), .A2(n556), .ZN(n561) );
  NAND2_X1 U615 ( .A1(G137), .A2(n895), .ZN(n559) );
  NAND2_X1 U616 ( .A1(G125), .A2(n890), .ZN(n558) );
  NAND2_X1 U617 ( .A1(n559), .A2(n558), .ZN(n560) );
  NOR2_X1 U618 ( .A1(n561), .A2(n560), .ZN(G160) );
  NAND2_X1 U619 ( .A1(G78), .A2(n657), .ZN(n562) );
  XNOR2_X1 U620 ( .A(n562), .B(KEYINPUT72), .ZN(n564) );
  NAND2_X1 U621 ( .A1(G91), .A2(n654), .ZN(n563) );
  NAND2_X1 U622 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U623 ( .A(KEYINPUT73), .B(n565), .ZN(n569) );
  NAND2_X1 U624 ( .A1(n661), .A2(G53), .ZN(n567) );
  NAND2_X1 U625 ( .A1(G65), .A2(n653), .ZN(n566) );
  AND2_X1 U626 ( .A1(n567), .A2(n566), .ZN(n568) );
  NAND2_X1 U627 ( .A1(n569), .A2(n568), .ZN(G299) );
  NAND2_X1 U628 ( .A1(G7), .A2(G661), .ZN(n570) );
  XNOR2_X1 U629 ( .A(n570), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U630 ( .A(G223), .ZN(n827) );
  NAND2_X1 U631 ( .A1(n827), .A2(G567), .ZN(n571) );
  XOR2_X1 U632 ( .A(KEYINPUT11), .B(n571), .Z(G234) );
  XOR2_X1 U633 ( .A(KEYINPUT74), .B(KEYINPUT14), .Z(n573) );
  NAND2_X1 U634 ( .A1(G56), .A2(n653), .ZN(n572) );
  XNOR2_X1 U635 ( .A(n573), .B(n572), .ZN(n579) );
  NAND2_X1 U636 ( .A1(G81), .A2(n654), .ZN(n574) );
  XOR2_X1 U637 ( .A(KEYINPUT75), .B(n574), .Z(n575) );
  XNOR2_X1 U638 ( .A(n575), .B(KEYINPUT12), .ZN(n577) );
  NAND2_X1 U639 ( .A1(G68), .A2(n657), .ZN(n576) );
  NAND2_X1 U640 ( .A1(n577), .A2(n576), .ZN(n578) );
  NOR2_X1 U641 ( .A1(n579), .A2(n524), .ZN(n581) );
  NAND2_X1 U642 ( .A1(n661), .A2(G43), .ZN(n580) );
  INV_X1 U643 ( .A(G860), .ZN(n603) );
  OR2_X1 U644 ( .A1(n999), .A2(n603), .ZN(G153) );
  NAND2_X1 U645 ( .A1(G90), .A2(n654), .ZN(n583) );
  NAND2_X1 U646 ( .A1(G77), .A2(n657), .ZN(n582) );
  NAND2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U648 ( .A(n584), .B(KEYINPUT9), .ZN(n586) );
  NAND2_X1 U649 ( .A1(G64), .A2(n653), .ZN(n585) );
  NAND2_X1 U650 ( .A1(n586), .A2(n585), .ZN(n589) );
  NAND2_X1 U651 ( .A1(G52), .A2(n661), .ZN(n587) );
  XNOR2_X1 U652 ( .A(KEYINPUT71), .B(n587), .ZN(n588) );
  NOR2_X1 U653 ( .A1(n589), .A2(n588), .ZN(G171) );
  INV_X1 U654 ( .A(G171), .ZN(G301) );
  NAND2_X1 U655 ( .A1(G301), .A2(G868), .ZN(n590) );
  XNOR2_X1 U656 ( .A(n590), .B(KEYINPUT76), .ZN(n599) );
  INV_X1 U657 ( .A(G868), .ZN(n673) );
  NAND2_X1 U658 ( .A1(G54), .A2(n661), .ZN(n592) );
  NAND2_X1 U659 ( .A1(G79), .A2(n657), .ZN(n591) );
  NAND2_X1 U660 ( .A1(n592), .A2(n591), .ZN(n596) );
  NAND2_X1 U661 ( .A1(G66), .A2(n653), .ZN(n594) );
  NAND2_X1 U662 ( .A1(G92), .A2(n654), .ZN(n593) );
  NAND2_X1 U663 ( .A1(n594), .A2(n593), .ZN(n595) );
  NOR2_X1 U664 ( .A1(n596), .A2(n595), .ZN(n597) );
  XNOR2_X1 U665 ( .A(n597), .B(KEYINPUT15), .ZN(n1004) );
  NAND2_X1 U666 ( .A1(n673), .A2(n1004), .ZN(n598) );
  NAND2_X1 U667 ( .A1(n599), .A2(n598), .ZN(G284) );
  XNOR2_X1 U668 ( .A(KEYINPUT81), .B(G868), .ZN(n600) );
  NOR2_X1 U669 ( .A1(G286), .A2(n600), .ZN(n602) );
  NOR2_X1 U670 ( .A1(G868), .A2(G299), .ZN(n601) );
  NOR2_X1 U671 ( .A1(n602), .A2(n601), .ZN(G297) );
  NAND2_X1 U672 ( .A1(n603), .A2(G559), .ZN(n604) );
  INV_X1 U673 ( .A(n1004), .ZN(n911) );
  NAND2_X1 U674 ( .A1(n604), .A2(n911), .ZN(n605) );
  XNOR2_X1 U675 ( .A(n605), .B(KEYINPUT16), .ZN(n606) );
  XNOR2_X1 U676 ( .A(KEYINPUT82), .B(n606), .ZN(G148) );
  NOR2_X1 U677 ( .A1(G868), .A2(n999), .ZN(n607) );
  XOR2_X1 U678 ( .A(KEYINPUT83), .B(n607), .Z(n610) );
  NAND2_X1 U679 ( .A1(G868), .A2(n911), .ZN(n608) );
  NOR2_X1 U680 ( .A1(G559), .A2(n608), .ZN(n609) );
  NOR2_X1 U681 ( .A1(n610), .A2(n609), .ZN(G282) );
  NAND2_X1 U682 ( .A1(G99), .A2(n894), .ZN(n612) );
  NAND2_X1 U683 ( .A1(G111), .A2(n891), .ZN(n611) );
  NAND2_X1 U684 ( .A1(n612), .A2(n611), .ZN(n619) );
  NAND2_X1 U685 ( .A1(G123), .A2(n890), .ZN(n613) );
  XNOR2_X1 U686 ( .A(n613), .B(KEYINPUT18), .ZN(n614) );
  XNOR2_X1 U687 ( .A(n614), .B(KEYINPUT84), .ZN(n616) );
  NAND2_X1 U688 ( .A1(G135), .A2(n895), .ZN(n615) );
  NAND2_X1 U689 ( .A1(n616), .A2(n615), .ZN(n617) );
  XOR2_X1 U690 ( .A(KEYINPUT85), .B(n617), .Z(n618) );
  NOR2_X1 U691 ( .A1(n619), .A2(n618), .ZN(n933) );
  XNOR2_X1 U692 ( .A(n933), .B(G2096), .ZN(n621) );
  INV_X1 U693 ( .A(G2100), .ZN(n620) );
  NAND2_X1 U694 ( .A1(n621), .A2(n620), .ZN(G156) );
  NAND2_X1 U695 ( .A1(G67), .A2(n653), .ZN(n623) );
  NAND2_X1 U696 ( .A1(G93), .A2(n654), .ZN(n622) );
  NAND2_X1 U697 ( .A1(n623), .A2(n622), .ZN(n627) );
  NAND2_X1 U698 ( .A1(G55), .A2(n661), .ZN(n625) );
  NAND2_X1 U699 ( .A1(G80), .A2(n657), .ZN(n624) );
  NAND2_X1 U700 ( .A1(n625), .A2(n624), .ZN(n626) );
  OR2_X1 U701 ( .A1(n627), .A2(n626), .ZN(n672) );
  NAND2_X1 U702 ( .A1(G559), .A2(n911), .ZN(n628) );
  XNOR2_X1 U703 ( .A(n628), .B(n999), .ZN(n669) );
  XNOR2_X1 U704 ( .A(KEYINPUT86), .B(n669), .ZN(n629) );
  NOR2_X1 U705 ( .A1(G860), .A2(n629), .ZN(n630) );
  XOR2_X1 U706 ( .A(n672), .B(n630), .Z(G145) );
  NAND2_X1 U707 ( .A1(G72), .A2(n657), .ZN(n632) );
  NAND2_X1 U708 ( .A1(n654), .A2(G85), .ZN(n631) );
  NAND2_X1 U709 ( .A1(n632), .A2(n631), .ZN(n638) );
  NAND2_X1 U710 ( .A1(n661), .A2(G47), .ZN(n633) );
  XNOR2_X1 U711 ( .A(n633), .B(KEYINPUT68), .ZN(n635) );
  NAND2_X1 U712 ( .A1(G60), .A2(n653), .ZN(n634) );
  NAND2_X1 U713 ( .A1(n635), .A2(n634), .ZN(n636) );
  XOR2_X1 U714 ( .A(KEYINPUT69), .B(n636), .Z(n637) );
  NOR2_X1 U715 ( .A1(n638), .A2(n637), .ZN(n639) );
  XOR2_X1 U716 ( .A(KEYINPUT70), .B(n639), .Z(G290) );
  NAND2_X1 U717 ( .A1(G48), .A2(n661), .ZN(n641) );
  NAND2_X1 U718 ( .A1(G86), .A2(n654), .ZN(n640) );
  NAND2_X1 U719 ( .A1(n641), .A2(n640), .ZN(n644) );
  NAND2_X1 U720 ( .A1(n657), .A2(G73), .ZN(n642) );
  XOR2_X1 U721 ( .A(KEYINPUT2), .B(n642), .Z(n643) );
  NOR2_X1 U722 ( .A1(n644), .A2(n643), .ZN(n646) );
  NAND2_X1 U723 ( .A1(n653), .A2(G61), .ZN(n645) );
  NAND2_X1 U724 ( .A1(n646), .A2(n645), .ZN(G305) );
  NAND2_X1 U725 ( .A1(G49), .A2(n661), .ZN(n648) );
  NAND2_X1 U726 ( .A1(G74), .A2(G651), .ZN(n647) );
  NAND2_X1 U727 ( .A1(n648), .A2(n647), .ZN(n649) );
  NOR2_X1 U728 ( .A1(n653), .A2(n649), .ZN(n652) );
  NAND2_X1 U729 ( .A1(n650), .A2(G87), .ZN(n651) );
  NAND2_X1 U730 ( .A1(n652), .A2(n651), .ZN(G288) );
  NAND2_X1 U731 ( .A1(G62), .A2(n653), .ZN(n656) );
  NAND2_X1 U732 ( .A1(G88), .A2(n654), .ZN(n655) );
  NAND2_X1 U733 ( .A1(n656), .A2(n655), .ZN(n660) );
  NAND2_X1 U734 ( .A1(G75), .A2(n657), .ZN(n658) );
  XNOR2_X1 U735 ( .A(KEYINPUT87), .B(n658), .ZN(n659) );
  NOR2_X1 U736 ( .A1(n660), .A2(n659), .ZN(n663) );
  NAND2_X1 U737 ( .A1(n661), .A2(G50), .ZN(n662) );
  NAND2_X1 U738 ( .A1(n663), .A2(n662), .ZN(G303) );
  INV_X1 U739 ( .A(G303), .ZN(G166) );
  XNOR2_X1 U740 ( .A(n672), .B(KEYINPUT19), .ZN(n664) );
  XNOR2_X1 U741 ( .A(G288), .B(n664), .ZN(n665) );
  XNOR2_X1 U742 ( .A(G305), .B(n665), .ZN(n667) );
  INV_X1 U743 ( .A(G299), .ZN(n707) );
  XNOR2_X1 U744 ( .A(G166), .B(n707), .ZN(n666) );
  XNOR2_X1 U745 ( .A(n667), .B(n666), .ZN(n668) );
  XOR2_X1 U746 ( .A(G290), .B(n668), .Z(n910) );
  XNOR2_X1 U747 ( .A(KEYINPUT88), .B(n669), .ZN(n670) );
  XNOR2_X1 U748 ( .A(n910), .B(n670), .ZN(n671) );
  NAND2_X1 U749 ( .A1(n671), .A2(G868), .ZN(n675) );
  NAND2_X1 U750 ( .A1(n673), .A2(n672), .ZN(n674) );
  NAND2_X1 U751 ( .A1(n675), .A2(n674), .ZN(G295) );
  NAND2_X1 U752 ( .A1(G2078), .A2(G2084), .ZN(n676) );
  XOR2_X1 U753 ( .A(KEYINPUT20), .B(n676), .Z(n677) );
  NAND2_X1 U754 ( .A1(G2090), .A2(n677), .ZN(n678) );
  XNOR2_X1 U755 ( .A(KEYINPUT21), .B(n678), .ZN(n679) );
  NAND2_X1 U756 ( .A1(n679), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U757 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U758 ( .A1(G236), .A2(G238), .ZN(n680) );
  NAND2_X1 U759 ( .A1(G69), .A2(n680), .ZN(n681) );
  NOR2_X1 U760 ( .A1(n681), .A2(G237), .ZN(n682) );
  XNOR2_X1 U761 ( .A(n682), .B(KEYINPUT89), .ZN(n832) );
  NAND2_X1 U762 ( .A1(n832), .A2(G567), .ZN(n687) );
  NOR2_X1 U763 ( .A1(G220), .A2(G219), .ZN(n683) );
  XOR2_X1 U764 ( .A(KEYINPUT22), .B(n683), .Z(n684) );
  NOR2_X1 U765 ( .A1(G218), .A2(n684), .ZN(n685) );
  NAND2_X1 U766 ( .A1(G96), .A2(n685), .ZN(n833) );
  NAND2_X1 U767 ( .A1(n833), .A2(G2106), .ZN(n686) );
  NAND2_X1 U768 ( .A1(n687), .A2(n686), .ZN(n921) );
  NAND2_X1 U769 ( .A1(G483), .A2(G661), .ZN(n688) );
  NOR2_X1 U770 ( .A1(n921), .A2(n688), .ZN(n831) );
  NAND2_X1 U771 ( .A1(n831), .A2(G36), .ZN(G176) );
  XNOR2_X1 U772 ( .A(G1981), .B(G305), .ZN(n997) );
  NOR2_X2 U773 ( .A1(G164), .A2(G1384), .ZN(n785) );
  NAND2_X1 U774 ( .A1(G160), .A2(G40), .ZN(n784) );
  INV_X1 U775 ( .A(n784), .ZN(n689) );
  NAND2_X2 U776 ( .A1(n785), .A2(n689), .ZN(n732) );
  INV_X1 U777 ( .A(G2072), .ZN(n690) );
  XNOR2_X1 U778 ( .A(n691), .B(KEYINPUT27), .ZN(n693) );
  AND2_X1 U779 ( .A1(G1956), .A2(n732), .ZN(n692) );
  NOR2_X1 U780 ( .A1(n693), .A2(n692), .ZN(n706) );
  NOR2_X1 U781 ( .A1(n707), .A2(n706), .ZN(n694) );
  INV_X1 U782 ( .A(G1996), .ZN(n951) );
  NOR2_X1 U783 ( .A1(n732), .A2(n951), .ZN(n695) );
  XOR2_X1 U784 ( .A(n695), .B(KEYINPUT26), .Z(n697) );
  NAND2_X1 U785 ( .A1(n732), .A2(G1341), .ZN(n696) );
  NAND2_X1 U786 ( .A1(n697), .A2(n696), .ZN(n698) );
  NOR2_X1 U787 ( .A1(n999), .A2(n698), .ZN(n702) );
  NAND2_X1 U788 ( .A1(G1348), .A2(n732), .ZN(n700) );
  INV_X1 U789 ( .A(n732), .ZN(n713) );
  NAND2_X1 U790 ( .A1(G2067), .A2(n713), .ZN(n699) );
  NAND2_X1 U791 ( .A1(n700), .A2(n699), .ZN(n703) );
  NOR2_X1 U792 ( .A1(n1004), .A2(n703), .ZN(n701) );
  NAND2_X1 U793 ( .A1(n1004), .A2(n703), .ZN(n704) );
  NAND2_X1 U794 ( .A1(n705), .A2(n704), .ZN(n709) );
  NAND2_X1 U795 ( .A1(n707), .A2(n706), .ZN(n708) );
  NAND2_X1 U796 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U797 ( .A1(n522), .A2(n710), .ZN(n711) );
  XNOR2_X1 U798 ( .A(n711), .B(KEYINPUT29), .ZN(n717) );
  XNOR2_X1 U799 ( .A(G2078), .B(KEYINPUT25), .ZN(n712) );
  XNOR2_X1 U800 ( .A(n712), .B(KEYINPUT99), .ZN(n957) );
  NOR2_X1 U801 ( .A1(n957), .A2(n732), .ZN(n715) );
  NOR2_X1 U802 ( .A1(n713), .A2(G1961), .ZN(n714) );
  NOR2_X1 U803 ( .A1(n715), .A2(n714), .ZN(n724) );
  NOR2_X1 U804 ( .A1(G301), .A2(n724), .ZN(n716) );
  NOR2_X1 U805 ( .A1(n717), .A2(n716), .ZN(n729) );
  NAND2_X1 U806 ( .A1(G8), .A2(n732), .ZN(n769) );
  NOR2_X1 U807 ( .A1(G1966), .A2(n769), .ZN(n743) );
  NOR2_X1 U808 ( .A1(G2084), .A2(n732), .ZN(n719) );
  INV_X1 U809 ( .A(KEYINPUT98), .ZN(n718) );
  XNOR2_X1 U810 ( .A(n719), .B(n718), .ZN(n745) );
  NAND2_X1 U811 ( .A1(G8), .A2(n745), .ZN(n720) );
  NOR2_X1 U812 ( .A1(n743), .A2(n720), .ZN(n722) );
  XOR2_X1 U813 ( .A(KEYINPUT30), .B(KEYINPUT100), .Z(n721) );
  XNOR2_X1 U814 ( .A(n722), .B(n721), .ZN(n723) );
  NOR2_X1 U815 ( .A1(G168), .A2(n723), .ZN(n726) );
  AND2_X1 U816 ( .A1(G301), .A2(n724), .ZN(n725) );
  NOR2_X1 U817 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U818 ( .A(n727), .B(KEYINPUT31), .ZN(n728) );
  NOR2_X1 U819 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U820 ( .A(n730), .B(KEYINPUT101), .ZN(n741) );
  NAND2_X1 U821 ( .A1(n741), .A2(G286), .ZN(n737) );
  NOR2_X1 U822 ( .A1(G1971), .A2(n769), .ZN(n731) );
  XNOR2_X1 U823 ( .A(KEYINPUT103), .B(n731), .ZN(n735) );
  NOR2_X1 U824 ( .A1(G2090), .A2(n732), .ZN(n733) );
  NOR2_X1 U825 ( .A1(G166), .A2(n733), .ZN(n734) );
  NAND2_X1 U826 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U827 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U828 ( .A1(n738), .A2(G8), .ZN(n739) );
  XNOR2_X1 U829 ( .A(n740), .B(KEYINPUT32), .ZN(n750) );
  INV_X1 U830 ( .A(n741), .ZN(n742) );
  NOR2_X1 U831 ( .A1(n743), .A2(n742), .ZN(n744) );
  XNOR2_X1 U832 ( .A(n744), .B(KEYINPUT102), .ZN(n748) );
  INV_X1 U833 ( .A(n745), .ZN(n746) );
  NAND2_X1 U834 ( .A1(G8), .A2(n746), .ZN(n747) );
  NAND2_X1 U835 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U836 ( .A1(n750), .A2(n749), .ZN(n764) );
  NOR2_X1 U837 ( .A1(G1976), .A2(G288), .ZN(n756) );
  NOR2_X1 U838 ( .A1(G1971), .A2(G303), .ZN(n751) );
  NOR2_X1 U839 ( .A1(n756), .A2(n751), .ZN(n1006) );
  NAND2_X1 U840 ( .A1(n764), .A2(n1006), .ZN(n752) );
  NAND2_X1 U841 ( .A1(G1976), .A2(G288), .ZN(n1001) );
  INV_X1 U842 ( .A(n769), .ZN(n755) );
  INV_X1 U843 ( .A(KEYINPUT33), .ZN(n753) );
  NAND2_X1 U844 ( .A1(n526), .A2(n754), .ZN(n759) );
  NAND2_X1 U845 ( .A1(n756), .A2(n755), .ZN(n757) );
  NAND2_X1 U846 ( .A1(n757), .A2(KEYINPUT33), .ZN(n758) );
  NAND2_X1 U847 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U848 ( .A(KEYINPUT105), .B(n760), .ZN(n761) );
  NOR2_X1 U849 ( .A1(n997), .A2(n761), .ZN(n772) );
  NOR2_X1 U850 ( .A1(G2090), .A2(G303), .ZN(n762) );
  XNOR2_X1 U851 ( .A(n762), .B(KEYINPUT106), .ZN(n763) );
  NAND2_X1 U852 ( .A1(n763), .A2(G8), .ZN(n765) );
  NAND2_X1 U853 ( .A1(n765), .A2(n764), .ZN(n766) );
  NAND2_X1 U854 ( .A1(n766), .A2(n769), .ZN(n770) );
  NOR2_X1 U855 ( .A1(G1981), .A2(G305), .ZN(n767) );
  XOR2_X1 U856 ( .A(n767), .B(KEYINPUT24), .Z(n768) );
  NOR2_X1 U857 ( .A1(n772), .A2(n771), .ZN(n808) );
  XNOR2_X1 U858 ( .A(G2067), .B(KEYINPUT37), .ZN(n820) );
  NAND2_X1 U859 ( .A1(G104), .A2(n894), .ZN(n774) );
  NAND2_X1 U860 ( .A1(G140), .A2(n895), .ZN(n773) );
  NAND2_X1 U861 ( .A1(n774), .A2(n773), .ZN(n775) );
  XNOR2_X1 U862 ( .A(KEYINPUT34), .B(n775), .ZN(n781) );
  NAND2_X1 U863 ( .A1(n890), .A2(G128), .ZN(n777) );
  NAND2_X1 U864 ( .A1(G116), .A2(n891), .ZN(n776) );
  NAND2_X1 U865 ( .A1(n777), .A2(n776), .ZN(n778) );
  XNOR2_X1 U866 ( .A(KEYINPUT91), .B(n778), .ZN(n779) );
  XNOR2_X1 U867 ( .A(KEYINPUT35), .B(n779), .ZN(n780) );
  NOR2_X1 U868 ( .A1(n781), .A2(n780), .ZN(n782) );
  XNOR2_X1 U869 ( .A(KEYINPUT36), .B(n782), .ZN(n907) );
  NOR2_X1 U870 ( .A1(n820), .A2(n907), .ZN(n783) );
  XNOR2_X1 U871 ( .A(n783), .B(KEYINPUT92), .ZN(n944) );
  NOR2_X1 U872 ( .A1(n785), .A2(n784), .ZN(n822) );
  NAND2_X1 U873 ( .A1(n944), .A2(n822), .ZN(n786) );
  XOR2_X1 U874 ( .A(KEYINPUT93), .B(n786), .Z(n819) );
  NAND2_X1 U875 ( .A1(G95), .A2(n894), .ZN(n788) );
  NAND2_X1 U876 ( .A1(G107), .A2(n891), .ZN(n787) );
  NAND2_X1 U877 ( .A1(n788), .A2(n787), .ZN(n791) );
  NAND2_X1 U878 ( .A1(n890), .A2(G119), .ZN(n789) );
  XOR2_X1 U879 ( .A(KEYINPUT94), .B(n789), .Z(n790) );
  NOR2_X1 U880 ( .A1(n791), .A2(n790), .ZN(n793) );
  NAND2_X1 U881 ( .A1(n895), .A2(G131), .ZN(n792) );
  NAND2_X1 U882 ( .A1(n793), .A2(n792), .ZN(n904) );
  AND2_X1 U883 ( .A1(n904), .A2(G1991), .ZN(n804) );
  XOR2_X1 U884 ( .A(KEYINPUT96), .B(KEYINPUT38), .Z(n795) );
  NAND2_X1 U885 ( .A1(G105), .A2(n894), .ZN(n794) );
  XNOR2_X1 U886 ( .A(n795), .B(n794), .ZN(n800) );
  NAND2_X1 U887 ( .A1(n890), .A2(G129), .ZN(n797) );
  NAND2_X1 U888 ( .A1(G117), .A2(n891), .ZN(n796) );
  NAND2_X1 U889 ( .A1(n797), .A2(n796), .ZN(n798) );
  XOR2_X1 U890 ( .A(KEYINPUT95), .B(n798), .Z(n799) );
  NOR2_X1 U891 ( .A1(n800), .A2(n799), .ZN(n802) );
  NAND2_X1 U892 ( .A1(n895), .A2(G141), .ZN(n801) );
  NAND2_X1 U893 ( .A1(n802), .A2(n801), .ZN(n885) );
  AND2_X1 U894 ( .A1(n885), .A2(G1996), .ZN(n803) );
  NOR2_X1 U895 ( .A1(n804), .A2(n803), .ZN(n931) );
  INV_X1 U896 ( .A(n822), .ZN(n805) );
  NOR2_X1 U897 ( .A1(n931), .A2(n805), .ZN(n814) );
  XNOR2_X1 U898 ( .A(KEYINPUT97), .B(n814), .ZN(n806) );
  NAND2_X1 U899 ( .A1(n819), .A2(n806), .ZN(n807) );
  NOR2_X1 U900 ( .A1(n808), .A2(n807), .ZN(n811) );
  XNOR2_X1 U901 ( .A(G1986), .B(G290), .ZN(n1012) );
  NAND2_X1 U902 ( .A1(n1012), .A2(n822), .ZN(n809) );
  XNOR2_X1 U903 ( .A(n809), .B(KEYINPUT90), .ZN(n810) );
  NAND2_X1 U904 ( .A1(n811), .A2(n810), .ZN(n825) );
  NOR2_X1 U905 ( .A1(G1996), .A2(n885), .ZN(n937) );
  NOR2_X1 U906 ( .A1(G1991), .A2(n904), .ZN(n929) );
  NOR2_X1 U907 ( .A1(G1986), .A2(G290), .ZN(n812) );
  NOR2_X1 U908 ( .A1(n929), .A2(n812), .ZN(n813) );
  NOR2_X1 U909 ( .A1(n814), .A2(n813), .ZN(n815) );
  NOR2_X1 U910 ( .A1(n937), .A2(n815), .ZN(n816) );
  XOR2_X1 U911 ( .A(n816), .B(KEYINPUT39), .Z(n817) );
  XNOR2_X1 U912 ( .A(KEYINPUT107), .B(n817), .ZN(n818) );
  NAND2_X1 U913 ( .A1(n819), .A2(n818), .ZN(n821) );
  NAND2_X1 U914 ( .A1(n907), .A2(n820), .ZN(n934) );
  NAND2_X1 U915 ( .A1(n821), .A2(n934), .ZN(n823) );
  NAND2_X1 U916 ( .A1(n823), .A2(n822), .ZN(n824) );
  NAND2_X1 U917 ( .A1(n825), .A2(n824), .ZN(n826) );
  XNOR2_X1 U918 ( .A(n826), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U919 ( .A1(G2106), .A2(n827), .ZN(G217) );
  NAND2_X1 U920 ( .A1(G15), .A2(G2), .ZN(n828) );
  XOR2_X1 U921 ( .A(KEYINPUT110), .B(n828), .Z(n829) );
  NAND2_X1 U922 ( .A1(G661), .A2(n829), .ZN(G259) );
  NAND2_X1 U923 ( .A1(G3), .A2(G1), .ZN(n830) );
  NAND2_X1 U924 ( .A1(n831), .A2(n830), .ZN(G188) );
  INV_X1 U926 ( .A(G96), .ZN(G221) );
  NOR2_X1 U927 ( .A1(n833), .A2(n832), .ZN(G325) );
  INV_X1 U928 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U929 ( .A(G2454), .B(G2451), .ZN(n842) );
  XNOR2_X1 U930 ( .A(G2430), .B(G2446), .ZN(n840) );
  XOR2_X1 U931 ( .A(G2435), .B(G2427), .Z(n835) );
  XNOR2_X1 U932 ( .A(KEYINPUT108), .B(G2438), .ZN(n834) );
  XNOR2_X1 U933 ( .A(n835), .B(n834), .ZN(n836) );
  XOR2_X1 U934 ( .A(n836), .B(G2443), .Z(n838) );
  XNOR2_X1 U935 ( .A(G1341), .B(G1348), .ZN(n837) );
  XNOR2_X1 U936 ( .A(n838), .B(n837), .ZN(n839) );
  XNOR2_X1 U937 ( .A(n840), .B(n839), .ZN(n841) );
  XNOR2_X1 U938 ( .A(n842), .B(n841), .ZN(n843) );
  NAND2_X1 U939 ( .A1(n843), .A2(G14), .ZN(n844) );
  XNOR2_X1 U940 ( .A(KEYINPUT109), .B(n844), .ZN(G401) );
  XNOR2_X1 U941 ( .A(G1961), .B(KEYINPUT41), .ZN(n854) );
  XOR2_X1 U942 ( .A(G1976), .B(G1981), .Z(n846) );
  XNOR2_X1 U943 ( .A(G1956), .B(G1966), .ZN(n845) );
  XNOR2_X1 U944 ( .A(n846), .B(n845), .ZN(n850) );
  XOR2_X1 U945 ( .A(G1971), .B(G1986), .Z(n848) );
  XNOR2_X1 U946 ( .A(G1996), .B(G1991), .ZN(n847) );
  XNOR2_X1 U947 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U948 ( .A(n850), .B(n849), .Z(n852) );
  XNOR2_X1 U949 ( .A(KEYINPUT112), .B(G2474), .ZN(n851) );
  XNOR2_X1 U950 ( .A(n852), .B(n851), .ZN(n853) );
  XNOR2_X1 U951 ( .A(n854), .B(n853), .ZN(G229) );
  XOR2_X1 U952 ( .A(KEYINPUT42), .B(G2084), .Z(n856) );
  XNOR2_X1 U953 ( .A(G2090), .B(G2072), .ZN(n855) );
  XNOR2_X1 U954 ( .A(n856), .B(n855), .ZN(n857) );
  XOR2_X1 U955 ( .A(n857), .B(G2100), .Z(n859) );
  XNOR2_X1 U956 ( .A(G2067), .B(G2078), .ZN(n858) );
  XNOR2_X1 U957 ( .A(n859), .B(n858), .ZN(n863) );
  XOR2_X1 U958 ( .A(G2096), .B(KEYINPUT43), .Z(n861) );
  XNOR2_X1 U959 ( .A(G2678), .B(KEYINPUT111), .ZN(n860) );
  XNOR2_X1 U960 ( .A(n861), .B(n860), .ZN(n862) );
  XOR2_X1 U961 ( .A(n863), .B(n862), .Z(G227) );
  NAND2_X1 U962 ( .A1(G100), .A2(n894), .ZN(n865) );
  NAND2_X1 U963 ( .A1(G112), .A2(n891), .ZN(n864) );
  NAND2_X1 U964 ( .A1(n865), .A2(n864), .ZN(n866) );
  XNOR2_X1 U965 ( .A(n866), .B(KEYINPUT113), .ZN(n868) );
  NAND2_X1 U966 ( .A1(G136), .A2(n895), .ZN(n867) );
  NAND2_X1 U967 ( .A1(n868), .A2(n867), .ZN(n871) );
  NAND2_X1 U968 ( .A1(n890), .A2(G124), .ZN(n869) );
  XOR2_X1 U969 ( .A(KEYINPUT44), .B(n869), .Z(n870) );
  NOR2_X1 U970 ( .A1(n871), .A2(n870), .ZN(n872) );
  XNOR2_X1 U971 ( .A(KEYINPUT114), .B(n872), .ZN(G162) );
  NAND2_X1 U972 ( .A1(G103), .A2(n894), .ZN(n874) );
  NAND2_X1 U973 ( .A1(G139), .A2(n895), .ZN(n873) );
  NAND2_X1 U974 ( .A1(n874), .A2(n873), .ZN(n881) );
  XNOR2_X1 U975 ( .A(KEYINPUT47), .B(KEYINPUT118), .ZN(n879) );
  NAND2_X1 U976 ( .A1(n890), .A2(G127), .ZN(n877) );
  NAND2_X1 U977 ( .A1(G115), .A2(n891), .ZN(n875) );
  XOR2_X1 U978 ( .A(KEYINPUT117), .B(n875), .Z(n876) );
  NAND2_X1 U979 ( .A1(n877), .A2(n876), .ZN(n878) );
  XOR2_X1 U980 ( .A(n879), .B(n878), .Z(n880) );
  NOR2_X1 U981 ( .A1(n881), .A2(n880), .ZN(n922) );
  XNOR2_X1 U982 ( .A(n922), .B(n933), .ZN(n889) );
  XOR2_X1 U983 ( .A(KEYINPUT119), .B(KEYINPUT116), .Z(n883) );
  XNOR2_X1 U984 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n882) );
  XNOR2_X1 U985 ( .A(n883), .B(n882), .ZN(n884) );
  XNOR2_X1 U986 ( .A(G162), .B(n884), .ZN(n887) );
  XOR2_X1 U987 ( .A(G164), .B(n885), .Z(n886) );
  XNOR2_X1 U988 ( .A(n887), .B(n886), .ZN(n888) );
  XNOR2_X1 U989 ( .A(n889), .B(n888), .ZN(n903) );
  NAND2_X1 U990 ( .A1(n890), .A2(G130), .ZN(n893) );
  NAND2_X1 U991 ( .A1(G118), .A2(n891), .ZN(n892) );
  NAND2_X1 U992 ( .A1(n893), .A2(n892), .ZN(n901) );
  NAND2_X1 U993 ( .A1(G106), .A2(n894), .ZN(n897) );
  NAND2_X1 U994 ( .A1(G142), .A2(n895), .ZN(n896) );
  NAND2_X1 U995 ( .A1(n897), .A2(n896), .ZN(n898) );
  XNOR2_X1 U996 ( .A(KEYINPUT115), .B(n898), .ZN(n899) );
  XNOR2_X1 U997 ( .A(KEYINPUT45), .B(n899), .ZN(n900) );
  NOR2_X1 U998 ( .A1(n901), .A2(n900), .ZN(n902) );
  XOR2_X1 U999 ( .A(n903), .B(n902), .Z(n906) );
  XOR2_X1 U1000 ( .A(G160), .B(n904), .Z(n905) );
  XNOR2_X1 U1001 ( .A(n906), .B(n905), .ZN(n908) );
  XOR2_X1 U1002 ( .A(n908), .B(n907), .Z(n909) );
  NOR2_X1 U1003 ( .A1(G37), .A2(n909), .ZN(G395) );
  XNOR2_X1 U1004 ( .A(n911), .B(n910), .ZN(n913) );
  XNOR2_X1 U1005 ( .A(G286), .B(G171), .ZN(n912) );
  XNOR2_X1 U1006 ( .A(n913), .B(n912), .ZN(n914) );
  XOR2_X1 U1007 ( .A(n914), .B(n999), .Z(n915) );
  NOR2_X1 U1008 ( .A1(G37), .A2(n915), .ZN(G397) );
  OR2_X1 U1009 ( .A1(n921), .A2(G401), .ZN(n918) );
  NOR2_X1 U1010 ( .A1(G229), .A2(G227), .ZN(n916) );
  XNOR2_X1 U1011 ( .A(KEYINPUT49), .B(n916), .ZN(n917) );
  NOR2_X1 U1012 ( .A1(n918), .A2(n917), .ZN(n920) );
  NOR2_X1 U1013 ( .A1(G395), .A2(G397), .ZN(n919) );
  NAND2_X1 U1014 ( .A1(n920), .A2(n919), .ZN(G225) );
  INV_X1 U1015 ( .A(G225), .ZN(G308) );
  INV_X1 U1016 ( .A(n921), .ZN(G319) );
  INV_X1 U1017 ( .A(G69), .ZN(G235) );
  XNOR2_X1 U1018 ( .A(G164), .B(G2078), .ZN(n925) );
  XNOR2_X1 U1019 ( .A(G2072), .B(n922), .ZN(n923) );
  XNOR2_X1 U1020 ( .A(n923), .B(KEYINPUT120), .ZN(n924) );
  NAND2_X1 U1021 ( .A1(n925), .A2(n924), .ZN(n926) );
  XNOR2_X1 U1022 ( .A(n926), .B(KEYINPUT50), .ZN(n927) );
  XNOR2_X1 U1023 ( .A(KEYINPUT121), .B(n927), .ZN(n942) );
  XOR2_X1 U1024 ( .A(G160), .B(G2084), .Z(n928) );
  NOR2_X1 U1025 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1026 ( .A1(n931), .A2(n930), .ZN(n932) );
  NOR2_X1 U1027 ( .A1(n933), .A2(n932), .ZN(n935) );
  NAND2_X1 U1028 ( .A1(n935), .A2(n934), .ZN(n940) );
  XOR2_X1 U1029 ( .A(G2090), .B(G162), .Z(n936) );
  NOR2_X1 U1030 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1031 ( .A(n938), .B(KEYINPUT51), .ZN(n939) );
  NOR2_X1 U1032 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1033 ( .A1(n942), .A2(n941), .ZN(n943) );
  NOR2_X1 U1034 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1035 ( .A(KEYINPUT52), .B(n945), .ZN(n946) );
  INV_X1 U1036 ( .A(KEYINPUT55), .ZN(n967) );
  NAND2_X1 U1037 ( .A1(n946), .A2(n967), .ZN(n947) );
  NAND2_X1 U1038 ( .A1(n947), .A2(G29), .ZN(n1025) );
  XNOR2_X1 U1039 ( .A(G2090), .B(G35), .ZN(n962) );
  XNOR2_X1 U1040 ( .A(G1991), .B(G25), .ZN(n949) );
  XNOR2_X1 U1041 ( .A(G33), .B(G2072), .ZN(n948) );
  NOR2_X1 U1042 ( .A1(n949), .A2(n948), .ZN(n956) );
  XOR2_X1 U1043 ( .A(G2067), .B(G26), .Z(n950) );
  NAND2_X1 U1044 ( .A1(n950), .A2(G28), .ZN(n954) );
  XOR2_X1 U1045 ( .A(G32), .B(n951), .Z(n952) );
  XNOR2_X1 U1046 ( .A(KEYINPUT122), .B(n952), .ZN(n953) );
  NOR2_X1 U1047 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1048 ( .A1(n956), .A2(n955), .ZN(n959) );
  XNOR2_X1 U1049 ( .A(G27), .B(n957), .ZN(n958) );
  NOR2_X1 U1050 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1051 ( .A(KEYINPUT53), .B(n960), .ZN(n961) );
  NOR2_X1 U1052 ( .A1(n962), .A2(n961), .ZN(n965) );
  XOR2_X1 U1053 ( .A(G2084), .B(G34), .Z(n963) );
  XNOR2_X1 U1054 ( .A(KEYINPUT54), .B(n963), .ZN(n964) );
  NAND2_X1 U1055 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1056 ( .A(n967), .B(n966), .ZN(n969) );
  INV_X1 U1057 ( .A(G29), .ZN(n968) );
  NAND2_X1 U1058 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1059 ( .A1(G11), .A2(n970), .ZN(n1023) );
  XOR2_X1 U1060 ( .A(G1971), .B(G22), .Z(n973) );
  XOR2_X1 U1061 ( .A(G23), .B(KEYINPUT126), .Z(n971) );
  XNOR2_X1 U1062 ( .A(n971), .B(G1976), .ZN(n972) );
  NAND2_X1 U1063 ( .A1(n973), .A2(n972), .ZN(n975) );
  XNOR2_X1 U1064 ( .A(G24), .B(G1986), .ZN(n974) );
  NOR2_X1 U1065 ( .A1(n975), .A2(n974), .ZN(n976) );
  XOR2_X1 U1066 ( .A(KEYINPUT58), .B(n976), .Z(n992) );
  XOR2_X1 U1067 ( .A(G1961), .B(G5), .Z(n987) );
  XNOR2_X1 U1068 ( .A(G1348), .B(KEYINPUT59), .ZN(n977) );
  XNOR2_X1 U1069 ( .A(n977), .B(G4), .ZN(n981) );
  XNOR2_X1 U1070 ( .A(G1341), .B(G19), .ZN(n979) );
  XNOR2_X1 U1071 ( .A(G1956), .B(G20), .ZN(n978) );
  NOR2_X1 U1072 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1073 ( .A1(n981), .A2(n980), .ZN(n984) );
  XNOR2_X1 U1074 ( .A(KEYINPUT124), .B(G1981), .ZN(n982) );
  XNOR2_X1 U1075 ( .A(G6), .B(n982), .ZN(n983) );
  NOR2_X1 U1076 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1077 ( .A(KEYINPUT60), .B(n985), .ZN(n986) );
  NAND2_X1 U1078 ( .A1(n987), .A2(n986), .ZN(n989) );
  XNOR2_X1 U1079 ( .A(G21), .B(G1966), .ZN(n988) );
  NOR2_X1 U1080 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1081 ( .A(KEYINPUT125), .B(n990), .ZN(n991) );
  NOR2_X1 U1082 ( .A1(n992), .A2(n991), .ZN(n993) );
  XOR2_X1 U1083 ( .A(KEYINPUT61), .B(n993), .Z(n994) );
  NOR2_X1 U1084 ( .A1(G16), .A2(n994), .ZN(n995) );
  XNOR2_X1 U1085 ( .A(KEYINPUT127), .B(n995), .ZN(n1021) );
  XNOR2_X1 U1086 ( .A(KEYINPUT56), .B(G16), .ZN(n1019) );
  XOR2_X1 U1087 ( .A(G1966), .B(G168), .Z(n996) );
  NOR2_X1 U1088 ( .A1(n997), .A2(n996), .ZN(n998) );
  XOR2_X1 U1089 ( .A(KEYINPUT57), .B(n998), .Z(n1017) );
  XNOR2_X1 U1090 ( .A(n999), .B(G1341), .ZN(n1015) );
  NAND2_X1 U1091 ( .A1(G1971), .A2(G303), .ZN(n1000) );
  NAND2_X1 U1092 ( .A1(n1001), .A2(n1000), .ZN(n1003) );
  XNOR2_X1 U1093 ( .A(G1961), .B(G301), .ZN(n1002) );
  NOR2_X1 U1094 ( .A1(n1003), .A2(n1002), .ZN(n1010) );
  XOR2_X1 U1095 ( .A(G1348), .B(n1004), .Z(n1005) );
  NAND2_X1 U1096 ( .A1(n1006), .A2(n1005), .ZN(n1008) );
  XNOR2_X1 U1097 ( .A(G1956), .B(G299), .ZN(n1007) );
  NOR2_X1 U1098 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1099 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NOR2_X1 U1100 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1101 ( .A(KEYINPUT123), .B(n1013), .ZN(n1014) );
  NOR2_X1 U1102 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1103 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1104 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1105 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NOR2_X1 U1106 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1107 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XOR2_X1 U1108 ( .A(KEYINPUT62), .B(n1026), .Z(G311) );
  INV_X1 U1109 ( .A(G311), .ZN(G150) );
endmodule

