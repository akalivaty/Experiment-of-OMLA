

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U551 ( .A(n735), .ZN(n722) );
  XOR2_X1 U552 ( .A(KEYINPUT66), .B(n524), .Z(n892) );
  INV_X1 U553 ( .A(KEYINPUT29), .ZN(n719) );
  AND2_X1 U554 ( .A1(n740), .A2(n739), .ZN(n517) );
  NAND2_X1 U555 ( .A1(n924), .A2(n833), .ZN(n518) );
  XNOR2_X1 U556 ( .A(n693), .B(KEYINPUT26), .ZN(n695) );
  INV_X1 U557 ( .A(KEYINPUT30), .ZN(n727) );
  OR2_X1 U558 ( .A1(n734), .A2(n748), .ZN(n740) );
  AND2_X1 U559 ( .A1(n718), .A2(n717), .ZN(n720) );
  XNOR2_X1 U560 ( .A(n720), .B(n719), .ZN(n746) );
  NAND2_X1 U561 ( .A1(n741), .A2(n517), .ZN(n742) );
  NOR2_X1 U562 ( .A1(KEYINPUT33), .A2(n762), .ZN(n763) );
  NAND2_X1 U563 ( .A1(n691), .A2(n690), .ZN(n735) );
  NOR2_X1 U564 ( .A1(n689), .A2(G1384), .ZN(n794) );
  AND2_X1 U565 ( .A1(n523), .A2(G2104), .ZN(n886) );
  AND2_X1 U566 ( .A1(n817), .A2(n518), .ZN(n818) );
  NOR2_X1 U567 ( .A1(G651), .A2(n648), .ZN(n652) );
  XNOR2_X1 U568 ( .A(n520), .B(n519), .ZN(n887) );
  XOR2_X1 U569 ( .A(KEYINPUT1), .B(n541), .Z(n659) );
  BUF_X1 U570 ( .A(n689), .Z(G164) );
  INV_X1 U571 ( .A(G2105), .ZN(n523) );
  NAND2_X1 U572 ( .A1(G102), .A2(n886), .ZN(n522) );
  XNOR2_X1 U573 ( .A(KEYINPUT17), .B(KEYINPUT67), .ZN(n520) );
  NOR2_X1 U574 ( .A1(G2105), .A2(G2104), .ZN(n519) );
  NAND2_X1 U575 ( .A1(G138), .A2(n887), .ZN(n521) );
  NAND2_X1 U576 ( .A1(n522), .A2(n521), .ZN(n528) );
  NOR2_X1 U577 ( .A1(G2104), .A2(n523), .ZN(n891) );
  NAND2_X1 U578 ( .A1(n891), .A2(G126), .ZN(n526) );
  NAND2_X1 U579 ( .A1(G2104), .A2(G2105), .ZN(n524) );
  NAND2_X1 U580 ( .A1(G114), .A2(n892), .ZN(n525) );
  NAND2_X1 U581 ( .A1(n526), .A2(n525), .ZN(n527) );
  NOR2_X1 U582 ( .A1(n528), .A2(n527), .ZN(n689) );
  NAND2_X1 U583 ( .A1(G101), .A2(n886), .ZN(n529) );
  XNOR2_X1 U584 ( .A(n529), .B(KEYINPUT23), .ZN(n530) );
  XNOR2_X1 U585 ( .A(n530), .B(KEYINPUT65), .ZN(n532) );
  NAND2_X1 U586 ( .A1(G113), .A2(n892), .ZN(n531) );
  NAND2_X1 U587 ( .A1(n532), .A2(n531), .ZN(n536) );
  NAND2_X1 U588 ( .A1(G137), .A2(n887), .ZN(n534) );
  NAND2_X1 U589 ( .A1(G125), .A2(n891), .ZN(n533) );
  NAND2_X1 U590 ( .A1(n534), .A2(n533), .ZN(n535) );
  NOR2_X1 U591 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U592 ( .A(n537), .B(KEYINPUT64), .ZN(n690) );
  BUF_X1 U593 ( .A(n690), .Z(G160) );
  NOR2_X1 U594 ( .A1(G543), .A2(G651), .ZN(n651) );
  NAND2_X1 U595 ( .A1(G85), .A2(n651), .ZN(n539) );
  XOR2_X1 U596 ( .A(G543), .B(KEYINPUT0), .Z(n648) );
  INV_X1 U597 ( .A(G651), .ZN(n540) );
  NOR2_X1 U598 ( .A1(n648), .A2(n540), .ZN(n655) );
  NAND2_X1 U599 ( .A1(G72), .A2(n655), .ZN(n538) );
  NAND2_X1 U600 ( .A1(n539), .A2(n538), .ZN(n545) );
  NAND2_X1 U601 ( .A1(G47), .A2(n652), .ZN(n543) );
  NOR2_X1 U602 ( .A1(G543), .A2(n540), .ZN(n541) );
  NAND2_X1 U603 ( .A1(G60), .A2(n659), .ZN(n542) );
  NAND2_X1 U604 ( .A1(n543), .A2(n542), .ZN(n544) );
  OR2_X1 U605 ( .A1(n545), .A2(n544), .ZN(G290) );
  XOR2_X1 U606 ( .A(G2446), .B(G2451), .Z(n547) );
  XNOR2_X1 U607 ( .A(G2454), .B(KEYINPUT105), .ZN(n546) );
  XNOR2_X1 U608 ( .A(n547), .B(n546), .ZN(n554) );
  XOR2_X1 U609 ( .A(G2438), .B(G2430), .Z(n549) );
  XNOR2_X1 U610 ( .A(G2435), .B(G2443), .ZN(n548) );
  XNOR2_X1 U611 ( .A(n549), .B(n548), .ZN(n550) );
  XOR2_X1 U612 ( .A(n550), .B(G2427), .Z(n552) );
  XNOR2_X1 U613 ( .A(G1341), .B(G1348), .ZN(n551) );
  XNOR2_X1 U614 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U615 ( .A(n554), .B(n553), .ZN(n555) );
  AND2_X1 U616 ( .A1(n555), .A2(G14), .ZN(G401) );
  AND2_X1 U617 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U618 ( .A(G57), .ZN(G237) );
  NAND2_X1 U619 ( .A1(G52), .A2(n652), .ZN(n557) );
  NAND2_X1 U620 ( .A1(G64), .A2(n659), .ZN(n556) );
  NAND2_X1 U621 ( .A1(n557), .A2(n556), .ZN(n564) );
  NAND2_X1 U622 ( .A1(n651), .A2(G90), .ZN(n558) );
  XNOR2_X1 U623 ( .A(n558), .B(KEYINPUT68), .ZN(n560) );
  NAND2_X1 U624 ( .A1(G77), .A2(n655), .ZN(n559) );
  NAND2_X1 U625 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U626 ( .A(KEYINPUT9), .B(n561), .ZN(n562) );
  XNOR2_X1 U627 ( .A(KEYINPUT69), .B(n562), .ZN(n563) );
  NOR2_X1 U628 ( .A1(n564), .A2(n563), .ZN(G171) );
  NAND2_X1 U629 ( .A1(G88), .A2(n651), .ZN(n566) );
  NAND2_X1 U630 ( .A1(G75), .A2(n655), .ZN(n565) );
  NAND2_X1 U631 ( .A1(n566), .A2(n565), .ZN(n570) );
  NAND2_X1 U632 ( .A1(G50), .A2(n652), .ZN(n568) );
  NAND2_X1 U633 ( .A1(G62), .A2(n659), .ZN(n567) );
  NAND2_X1 U634 ( .A1(n568), .A2(n567), .ZN(n569) );
  NOR2_X1 U635 ( .A1(n570), .A2(n569), .ZN(G166) );
  NAND2_X1 U636 ( .A1(n651), .A2(G89), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n571), .B(KEYINPUT4), .ZN(n573) );
  NAND2_X1 U638 ( .A1(G76), .A2(n655), .ZN(n572) );
  NAND2_X1 U639 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n574), .B(KEYINPUT5), .ZN(n579) );
  NAND2_X1 U641 ( .A1(G51), .A2(n652), .ZN(n576) );
  NAND2_X1 U642 ( .A1(G63), .A2(n659), .ZN(n575) );
  NAND2_X1 U643 ( .A1(n576), .A2(n575), .ZN(n577) );
  XOR2_X1 U644 ( .A(KEYINPUT6), .B(n577), .Z(n578) );
  NAND2_X1 U645 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n580), .B(KEYINPUT7), .ZN(G168) );
  XNOR2_X1 U647 ( .A(G168), .B(KEYINPUT8), .ZN(n581) );
  XNOR2_X1 U648 ( .A(n581), .B(KEYINPUT73), .ZN(G286) );
  NAND2_X1 U649 ( .A1(G7), .A2(G661), .ZN(n582) );
  XNOR2_X1 U650 ( .A(n582), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U651 ( .A(G223), .ZN(n838) );
  NAND2_X1 U652 ( .A1(n838), .A2(G567), .ZN(n583) );
  XOR2_X1 U653 ( .A(KEYINPUT11), .B(n583), .Z(G234) );
  NAND2_X1 U654 ( .A1(n651), .A2(G81), .ZN(n584) );
  XNOR2_X1 U655 ( .A(n584), .B(KEYINPUT12), .ZN(n586) );
  NAND2_X1 U656 ( .A1(G68), .A2(n655), .ZN(n585) );
  NAND2_X1 U657 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U658 ( .A(n587), .B(KEYINPUT13), .ZN(n589) );
  NAND2_X1 U659 ( .A1(G43), .A2(n652), .ZN(n588) );
  NAND2_X1 U660 ( .A1(n589), .A2(n588), .ZN(n592) );
  NAND2_X1 U661 ( .A1(n659), .A2(G56), .ZN(n590) );
  XOR2_X1 U662 ( .A(KEYINPUT14), .B(n590), .Z(n591) );
  NOR2_X1 U663 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U664 ( .A(KEYINPUT71), .B(n593), .ZN(n936) );
  INV_X1 U665 ( .A(G860), .ZN(n634) );
  NOR2_X1 U666 ( .A1(n936), .A2(n634), .ZN(n594) );
  XOR2_X1 U667 ( .A(KEYINPUT72), .B(n594), .Z(G153) );
  INV_X1 U668 ( .A(G171), .ZN(G301) );
  NAND2_X1 U669 ( .A1(G868), .A2(G301), .ZN(n603) );
  NAND2_X1 U670 ( .A1(G92), .A2(n651), .ZN(n596) );
  NAND2_X1 U671 ( .A1(G79), .A2(n655), .ZN(n595) );
  NAND2_X1 U672 ( .A1(n596), .A2(n595), .ZN(n600) );
  NAND2_X1 U673 ( .A1(G54), .A2(n652), .ZN(n598) );
  NAND2_X1 U674 ( .A1(G66), .A2(n659), .ZN(n597) );
  NAND2_X1 U675 ( .A1(n598), .A2(n597), .ZN(n599) );
  NOR2_X1 U676 ( .A1(n600), .A2(n599), .ZN(n601) );
  XOR2_X1 U677 ( .A(KEYINPUT15), .B(n601), .Z(n921) );
  INV_X1 U678 ( .A(n921), .ZN(n617) );
  INV_X1 U679 ( .A(G868), .ZN(n619) );
  NAND2_X1 U680 ( .A1(n617), .A2(n619), .ZN(n602) );
  NAND2_X1 U681 ( .A1(n603), .A2(n602), .ZN(G284) );
  NAND2_X1 U682 ( .A1(G91), .A2(n651), .ZN(n605) );
  NAND2_X1 U683 ( .A1(G78), .A2(n655), .ZN(n604) );
  NAND2_X1 U684 ( .A1(n605), .A2(n604), .ZN(n608) );
  NAND2_X1 U685 ( .A1(n652), .A2(G53), .ZN(n606) );
  XOR2_X1 U686 ( .A(KEYINPUT70), .B(n606), .Z(n607) );
  NOR2_X1 U687 ( .A1(n608), .A2(n607), .ZN(n610) );
  NAND2_X1 U688 ( .A1(n659), .A2(G65), .ZN(n609) );
  NAND2_X1 U689 ( .A1(n610), .A2(n609), .ZN(G299) );
  XNOR2_X1 U690 ( .A(KEYINPUT74), .B(n619), .ZN(n611) );
  NOR2_X1 U691 ( .A1(G286), .A2(n611), .ZN(n613) );
  NOR2_X1 U692 ( .A1(G868), .A2(G299), .ZN(n612) );
  NOR2_X1 U693 ( .A1(n613), .A2(n612), .ZN(G297) );
  NAND2_X1 U694 ( .A1(n634), .A2(G559), .ZN(n614) );
  NAND2_X1 U695 ( .A1(n614), .A2(n921), .ZN(n615) );
  XNOR2_X1 U696 ( .A(n615), .B(KEYINPUT16), .ZN(n616) );
  XOR2_X1 U697 ( .A(KEYINPUT75), .B(n616), .Z(G148) );
  OR2_X1 U698 ( .A1(G559), .A2(n617), .ZN(n618) );
  NAND2_X1 U699 ( .A1(n618), .A2(G868), .ZN(n621) );
  NAND2_X1 U700 ( .A1(n936), .A2(n619), .ZN(n620) );
  NAND2_X1 U701 ( .A1(n621), .A2(n620), .ZN(G282) );
  NAND2_X1 U702 ( .A1(G99), .A2(n886), .ZN(n623) );
  NAND2_X1 U703 ( .A1(G111), .A2(n892), .ZN(n622) );
  NAND2_X1 U704 ( .A1(n623), .A2(n622), .ZN(n624) );
  XNOR2_X1 U705 ( .A(KEYINPUT76), .B(n624), .ZN(n627) );
  NAND2_X1 U706 ( .A1(n891), .A2(G123), .ZN(n625) );
  XOR2_X1 U707 ( .A(KEYINPUT18), .B(n625), .Z(n626) );
  NOR2_X1 U708 ( .A1(n627), .A2(n626), .ZN(n629) );
  NAND2_X1 U709 ( .A1(n887), .A2(G135), .ZN(n628) );
  NAND2_X1 U710 ( .A1(n629), .A2(n628), .ZN(n630) );
  XNOR2_X1 U711 ( .A(KEYINPUT77), .B(n630), .ZN(n1003) );
  XNOR2_X1 U712 ( .A(G2096), .B(n1003), .ZN(n632) );
  INV_X1 U713 ( .A(G2100), .ZN(n631) );
  NAND2_X1 U714 ( .A1(n632), .A2(n631), .ZN(G156) );
  NAND2_X1 U715 ( .A1(G559), .A2(n921), .ZN(n633) );
  XOR2_X1 U716 ( .A(n936), .B(n633), .Z(n668) );
  NAND2_X1 U717 ( .A1(n634), .A2(n668), .ZN(n644) );
  NAND2_X1 U718 ( .A1(n652), .A2(G55), .ZN(n635) );
  XOR2_X1 U719 ( .A(KEYINPUT79), .B(n635), .Z(n637) );
  NAND2_X1 U720 ( .A1(n659), .A2(G67), .ZN(n636) );
  NAND2_X1 U721 ( .A1(n637), .A2(n636), .ZN(n638) );
  XNOR2_X1 U722 ( .A(KEYINPUT80), .B(n638), .ZN(n643) );
  NAND2_X1 U723 ( .A1(n651), .A2(G93), .ZN(n639) );
  XNOR2_X1 U724 ( .A(n639), .B(KEYINPUT78), .ZN(n641) );
  NAND2_X1 U725 ( .A1(G80), .A2(n655), .ZN(n640) );
  NAND2_X1 U726 ( .A1(n641), .A2(n640), .ZN(n642) );
  NOR2_X1 U727 ( .A1(n643), .A2(n642), .ZN(n670) );
  XOR2_X1 U728 ( .A(n644), .B(n670), .Z(G145) );
  NAND2_X1 U729 ( .A1(G49), .A2(n652), .ZN(n646) );
  NAND2_X1 U730 ( .A1(G74), .A2(G651), .ZN(n645) );
  NAND2_X1 U731 ( .A1(n646), .A2(n645), .ZN(n647) );
  NOR2_X1 U732 ( .A1(n659), .A2(n647), .ZN(n650) );
  NAND2_X1 U733 ( .A1(n648), .A2(G87), .ZN(n649) );
  NAND2_X1 U734 ( .A1(n650), .A2(n649), .ZN(G288) );
  NAND2_X1 U735 ( .A1(G86), .A2(n651), .ZN(n654) );
  NAND2_X1 U736 ( .A1(G48), .A2(n652), .ZN(n653) );
  NAND2_X1 U737 ( .A1(n654), .A2(n653), .ZN(n658) );
  NAND2_X1 U738 ( .A1(n655), .A2(G73), .ZN(n656) );
  XOR2_X1 U739 ( .A(KEYINPUT2), .B(n656), .Z(n657) );
  NOR2_X1 U740 ( .A1(n658), .A2(n657), .ZN(n661) );
  NAND2_X1 U741 ( .A1(n659), .A2(G61), .ZN(n660) );
  NAND2_X1 U742 ( .A1(n661), .A2(n660), .ZN(G305) );
  XNOR2_X1 U743 ( .A(G166), .B(G290), .ZN(n667) );
  INV_X1 U744 ( .A(G299), .ZN(n714) );
  XNOR2_X1 U745 ( .A(KEYINPUT81), .B(KEYINPUT19), .ZN(n663) );
  XNOR2_X1 U746 ( .A(G288), .B(n670), .ZN(n662) );
  XNOR2_X1 U747 ( .A(n663), .B(n662), .ZN(n664) );
  XNOR2_X1 U748 ( .A(n714), .B(n664), .ZN(n665) );
  XNOR2_X1 U749 ( .A(n665), .B(G305), .ZN(n666) );
  XNOR2_X1 U750 ( .A(n667), .B(n666), .ZN(n910) );
  XNOR2_X1 U751 ( .A(n668), .B(n910), .ZN(n669) );
  NAND2_X1 U752 ( .A1(n669), .A2(G868), .ZN(n672) );
  OR2_X1 U753 ( .A1(G868), .A2(n670), .ZN(n671) );
  NAND2_X1 U754 ( .A1(n672), .A2(n671), .ZN(n673) );
  XNOR2_X1 U755 ( .A(KEYINPUT82), .B(n673), .ZN(G295) );
  NAND2_X1 U756 ( .A1(G2078), .A2(G2084), .ZN(n674) );
  XOR2_X1 U757 ( .A(KEYINPUT20), .B(n674), .Z(n675) );
  NAND2_X1 U758 ( .A1(G2090), .A2(n675), .ZN(n676) );
  XNOR2_X1 U759 ( .A(KEYINPUT21), .B(n676), .ZN(n677) );
  NAND2_X1 U760 ( .A1(n677), .A2(G2072), .ZN(G158) );
  XOR2_X1 U761 ( .A(KEYINPUT83), .B(G44), .Z(n678) );
  XNOR2_X1 U762 ( .A(KEYINPUT3), .B(n678), .ZN(G218) );
  NAND2_X1 U763 ( .A1(G132), .A2(G82), .ZN(n679) );
  XNOR2_X1 U764 ( .A(n679), .B(KEYINPUT84), .ZN(n680) );
  XNOR2_X1 U765 ( .A(n680), .B(KEYINPUT22), .ZN(n681) );
  NOR2_X1 U766 ( .A1(G218), .A2(n681), .ZN(n682) );
  NAND2_X1 U767 ( .A1(G96), .A2(n682), .ZN(n843) );
  NAND2_X1 U768 ( .A1(G2106), .A2(n843), .ZN(n683) );
  XOR2_X1 U769 ( .A(KEYINPUT85), .B(n683), .Z(n687) );
  NAND2_X1 U770 ( .A1(G69), .A2(G120), .ZN(n684) );
  NOR2_X1 U771 ( .A1(G237), .A2(n684), .ZN(n685) );
  NAND2_X1 U772 ( .A1(G108), .A2(n685), .ZN(n844) );
  NAND2_X1 U773 ( .A1(G567), .A2(n844), .ZN(n686) );
  NAND2_X1 U774 ( .A1(n687), .A2(n686), .ZN(n845) );
  NAND2_X1 U775 ( .A1(G483), .A2(G661), .ZN(n688) );
  NOR2_X1 U776 ( .A1(n845), .A2(n688), .ZN(n842) );
  NAND2_X1 U777 ( .A1(n842), .A2(G36), .ZN(G176) );
  INV_X1 U778 ( .A(G166), .ZN(G303) );
  AND2_X1 U779 ( .A1(G40), .A2(n794), .ZN(n691) );
  INV_X1 U780 ( .A(n735), .ZN(n692) );
  NAND2_X1 U781 ( .A1(G1996), .A2(n692), .ZN(n693) );
  NAND2_X1 U782 ( .A1(G1341), .A2(n735), .ZN(n694) );
  NAND2_X1 U783 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U784 ( .A(KEYINPUT94), .B(n696), .ZN(n697) );
  NOR2_X1 U785 ( .A1(n697), .A2(n936), .ZN(n704) );
  NAND2_X1 U786 ( .A1(n704), .A2(n921), .ZN(n702) );
  AND2_X1 U787 ( .A1(n722), .A2(G2067), .ZN(n698) );
  XNOR2_X1 U788 ( .A(n698), .B(KEYINPUT95), .ZN(n700) );
  NAND2_X1 U789 ( .A1(n735), .A2(G1348), .ZN(n699) );
  NAND2_X1 U790 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U791 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U792 ( .A(n703), .B(KEYINPUT96), .ZN(n712) );
  OR2_X1 U793 ( .A1(n704), .A2(n921), .ZN(n710) );
  NAND2_X1 U794 ( .A1(n722), .A2(G2072), .ZN(n705) );
  XNOR2_X1 U795 ( .A(n705), .B(KEYINPUT27), .ZN(n707) );
  XNOR2_X1 U796 ( .A(G1956), .B(KEYINPUT93), .ZN(n947) );
  NOR2_X1 U797 ( .A1(n947), .A2(n722), .ZN(n706) );
  NOR2_X1 U798 ( .A1(n707), .A2(n706), .ZN(n713) );
  NOR2_X1 U799 ( .A1(n714), .A2(n713), .ZN(n708) );
  XNOR2_X1 U800 ( .A(n708), .B(KEYINPUT28), .ZN(n716) );
  INV_X1 U801 ( .A(n716), .ZN(n709) );
  AND2_X1 U802 ( .A1(n710), .A2(n709), .ZN(n711) );
  NAND2_X1 U803 ( .A1(n712), .A2(n711), .ZN(n718) );
  NAND2_X1 U804 ( .A1(n714), .A2(n713), .ZN(n715) );
  OR2_X1 U805 ( .A1(n716), .A2(n715), .ZN(n717) );
  NOR2_X1 U806 ( .A1(n722), .A2(G1961), .ZN(n721) );
  XOR2_X1 U807 ( .A(KEYINPUT92), .B(n721), .Z(n724) );
  XNOR2_X1 U808 ( .A(G2078), .B(KEYINPUT25), .ZN(n974) );
  NAND2_X1 U809 ( .A1(n722), .A2(n974), .ZN(n723) );
  NAND2_X1 U810 ( .A1(n724), .A2(n723), .ZN(n730) );
  NAND2_X1 U811 ( .A1(n730), .A2(G171), .ZN(n747) );
  AND2_X1 U812 ( .A1(n747), .A2(G286), .ZN(n725) );
  NAND2_X1 U813 ( .A1(n746), .A2(n725), .ZN(n741) );
  INV_X1 U814 ( .A(G286), .ZN(n734) );
  NAND2_X1 U815 ( .A1(n735), .A2(G8), .ZN(n778) );
  NOR2_X1 U816 ( .A1(G1966), .A2(n778), .ZN(n751) );
  NOR2_X1 U817 ( .A1(G2084), .A2(n735), .ZN(n745) );
  NOR2_X1 U818 ( .A1(n751), .A2(n745), .ZN(n726) );
  AND2_X1 U819 ( .A1(n726), .A2(G8), .ZN(n728) );
  XNOR2_X1 U820 ( .A(n728), .B(n727), .ZN(n729) );
  NOR2_X1 U821 ( .A1(G168), .A2(n729), .ZN(n732) );
  NOR2_X1 U822 ( .A1(G171), .A2(n730), .ZN(n731) );
  NOR2_X1 U823 ( .A1(n732), .A2(n731), .ZN(n733) );
  XOR2_X1 U824 ( .A(KEYINPUT31), .B(n733), .Z(n748) );
  NOR2_X1 U825 ( .A1(G1971), .A2(n778), .ZN(n737) );
  NOR2_X1 U826 ( .A1(G2090), .A2(n735), .ZN(n736) );
  NOR2_X1 U827 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U828 ( .A1(n738), .A2(G303), .ZN(n739) );
  NAND2_X1 U829 ( .A1(n742), .A2(G8), .ZN(n744) );
  XOR2_X1 U830 ( .A(KEYINPUT32), .B(KEYINPUT97), .Z(n743) );
  XNOR2_X1 U831 ( .A(n744), .B(n743), .ZN(n770) );
  NAND2_X1 U832 ( .A1(G8), .A2(n745), .ZN(n753) );
  NAND2_X1 U833 ( .A1(n747), .A2(n746), .ZN(n749) );
  AND2_X1 U834 ( .A1(n749), .A2(n748), .ZN(n750) );
  NOR2_X1 U835 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U836 ( .A1(n753), .A2(n752), .ZN(n771) );
  NAND2_X1 U837 ( .A1(G1976), .A2(G288), .ZN(n929) );
  AND2_X1 U838 ( .A1(n771), .A2(n929), .ZN(n754) );
  NAND2_X1 U839 ( .A1(n770), .A2(n754), .ZN(n761) );
  INV_X1 U840 ( .A(n929), .ZN(n759) );
  NOR2_X1 U841 ( .A1(G288), .A2(G1976), .ZN(n755) );
  XNOR2_X1 U842 ( .A(n755), .B(KEYINPUT98), .ZN(n932) );
  NOR2_X1 U843 ( .A1(G1971), .A2(G303), .ZN(n756) );
  XOR2_X1 U844 ( .A(n756), .B(KEYINPUT99), .Z(n757) );
  NOR2_X1 U845 ( .A1(n932), .A2(n757), .ZN(n758) );
  OR2_X1 U846 ( .A1(n759), .A2(n758), .ZN(n760) );
  AND2_X1 U847 ( .A1(n761), .A2(n760), .ZN(n762) );
  INV_X1 U848 ( .A(n778), .ZN(n764) );
  NAND2_X1 U849 ( .A1(n763), .A2(n764), .ZN(n767) );
  NAND2_X1 U850 ( .A1(n932), .A2(n764), .ZN(n765) );
  NAND2_X1 U851 ( .A1(n765), .A2(KEYINPUT33), .ZN(n766) );
  NAND2_X1 U852 ( .A1(n767), .A2(n766), .ZN(n768) );
  XNOR2_X1 U853 ( .A(n768), .B(KEYINPUT100), .ZN(n769) );
  XOR2_X1 U854 ( .A(G1981), .B(G305), .Z(n939) );
  AND2_X1 U855 ( .A1(n769), .A2(n939), .ZN(n782) );
  NAND2_X1 U856 ( .A1(n771), .A2(n770), .ZN(n774) );
  NOR2_X1 U857 ( .A1(G2090), .A2(G303), .ZN(n772) );
  NAND2_X1 U858 ( .A1(G8), .A2(n772), .ZN(n773) );
  NAND2_X1 U859 ( .A1(n774), .A2(n773), .ZN(n775) );
  NAND2_X1 U860 ( .A1(n775), .A2(n778), .ZN(n780) );
  NOR2_X1 U861 ( .A1(G1981), .A2(G305), .ZN(n776) );
  XOR2_X1 U862 ( .A(n776), .B(KEYINPUT24), .Z(n777) );
  OR2_X1 U863 ( .A1(n778), .A2(n777), .ZN(n779) );
  NAND2_X1 U864 ( .A1(n780), .A2(n779), .ZN(n781) );
  NOR2_X1 U865 ( .A1(n782), .A2(n781), .ZN(n783) );
  INV_X1 U866 ( .A(n783), .ZN(n819) );
  NAND2_X1 U867 ( .A1(n887), .A2(G140), .ZN(n784) );
  XOR2_X1 U868 ( .A(KEYINPUT87), .B(n784), .Z(n786) );
  NAND2_X1 U869 ( .A1(n886), .A2(G104), .ZN(n785) );
  NAND2_X1 U870 ( .A1(n786), .A2(n785), .ZN(n787) );
  XNOR2_X1 U871 ( .A(KEYINPUT34), .B(n787), .ZN(n792) );
  NAND2_X1 U872 ( .A1(n891), .A2(G128), .ZN(n789) );
  NAND2_X1 U873 ( .A1(G116), .A2(n892), .ZN(n788) );
  NAND2_X1 U874 ( .A1(n789), .A2(n788), .ZN(n790) );
  XOR2_X1 U875 ( .A(KEYINPUT35), .B(n790), .Z(n791) );
  NOR2_X1 U876 ( .A1(n792), .A2(n791), .ZN(n793) );
  XNOR2_X1 U877 ( .A(KEYINPUT36), .B(n793), .ZN(n885) );
  XNOR2_X1 U878 ( .A(KEYINPUT37), .B(G2067), .ZN(n831) );
  NOR2_X1 U879 ( .A1(n885), .A2(n831), .ZN(n1017) );
  NAND2_X1 U880 ( .A1(G40), .A2(G160), .ZN(n795) );
  NOR2_X1 U881 ( .A1(n795), .A2(n794), .ZN(n796) );
  XNOR2_X1 U882 ( .A(n796), .B(KEYINPUT86), .ZN(n833) );
  NAND2_X1 U883 ( .A1(n1017), .A2(n833), .ZN(n829) );
  INV_X1 U884 ( .A(n829), .ZN(n815) );
  NAND2_X1 U885 ( .A1(G95), .A2(n886), .ZN(n798) );
  NAND2_X1 U886 ( .A1(G107), .A2(n892), .ZN(n797) );
  NAND2_X1 U887 ( .A1(n798), .A2(n797), .ZN(n802) );
  NAND2_X1 U888 ( .A1(G131), .A2(n887), .ZN(n800) );
  NAND2_X1 U889 ( .A1(G119), .A2(n891), .ZN(n799) );
  NAND2_X1 U890 ( .A1(n800), .A2(n799), .ZN(n801) );
  OR2_X1 U891 ( .A1(n802), .A2(n801), .ZN(n904) );
  NAND2_X1 U892 ( .A1(G1991), .A2(n904), .ZN(n803) );
  XNOR2_X1 U893 ( .A(n803), .B(KEYINPUT88), .ZN(n813) );
  NAND2_X1 U894 ( .A1(n891), .A2(G129), .ZN(n805) );
  NAND2_X1 U895 ( .A1(G117), .A2(n892), .ZN(n804) );
  NAND2_X1 U896 ( .A1(n805), .A2(n804), .ZN(n809) );
  NAND2_X1 U897 ( .A1(G105), .A2(n886), .ZN(n806) );
  XNOR2_X1 U898 ( .A(n806), .B(KEYINPUT89), .ZN(n807) );
  XNOR2_X1 U899 ( .A(n807), .B(KEYINPUT38), .ZN(n808) );
  NOR2_X1 U900 ( .A1(n809), .A2(n808), .ZN(n811) );
  NAND2_X1 U901 ( .A1(n887), .A2(G141), .ZN(n810) );
  NAND2_X1 U902 ( .A1(n811), .A2(n810), .ZN(n898) );
  NAND2_X1 U903 ( .A1(G1996), .A2(n898), .ZN(n812) );
  NAND2_X1 U904 ( .A1(n813), .A2(n812), .ZN(n1006) );
  NAND2_X1 U905 ( .A1(n833), .A2(n1006), .ZN(n823) );
  XOR2_X1 U906 ( .A(KEYINPUT90), .B(n823), .Z(n814) );
  NOR2_X1 U907 ( .A1(n815), .A2(n814), .ZN(n816) );
  XOR2_X1 U908 ( .A(n816), .B(KEYINPUT91), .Z(n817) );
  XNOR2_X1 U909 ( .A(G1986), .B(G290), .ZN(n924) );
  NAND2_X1 U910 ( .A1(n819), .A2(n818), .ZN(n836) );
  NOR2_X1 U911 ( .A1(G1991), .A2(n904), .ZN(n1004) );
  NOR2_X1 U912 ( .A1(G1986), .A2(G290), .ZN(n820) );
  NOR2_X1 U913 ( .A1(n1004), .A2(n820), .ZN(n821) );
  XOR2_X1 U914 ( .A(KEYINPUT102), .B(n821), .Z(n822) );
  NAND2_X1 U915 ( .A1(n823), .A2(n822), .ZN(n825) );
  NOR2_X1 U916 ( .A1(n898), .A2(G1996), .ZN(n824) );
  XNOR2_X1 U917 ( .A(n824), .B(KEYINPUT101), .ZN(n1009) );
  NAND2_X1 U918 ( .A1(n825), .A2(n1009), .ZN(n827) );
  XNOR2_X1 U919 ( .A(KEYINPUT103), .B(KEYINPUT104), .ZN(n826) );
  XNOR2_X1 U920 ( .A(n827), .B(n826), .ZN(n828) );
  XNOR2_X1 U921 ( .A(n828), .B(KEYINPUT39), .ZN(n830) );
  NAND2_X1 U922 ( .A1(n830), .A2(n829), .ZN(n832) );
  NAND2_X1 U923 ( .A1(n885), .A2(n831), .ZN(n1019) );
  NAND2_X1 U924 ( .A1(n832), .A2(n1019), .ZN(n834) );
  NAND2_X1 U925 ( .A1(n834), .A2(n833), .ZN(n835) );
  NAND2_X1 U926 ( .A1(n836), .A2(n835), .ZN(n837) );
  XNOR2_X1 U927 ( .A(KEYINPUT40), .B(n837), .ZN(G329) );
  NAND2_X1 U928 ( .A1(n838), .A2(G2106), .ZN(n839) );
  XNOR2_X1 U929 ( .A(n839), .B(KEYINPUT106), .ZN(G217) );
  AND2_X1 U930 ( .A1(G15), .A2(G2), .ZN(n840) );
  NAND2_X1 U931 ( .A1(G661), .A2(n840), .ZN(G259) );
  NAND2_X1 U932 ( .A1(G3), .A2(G1), .ZN(n841) );
  NAND2_X1 U933 ( .A1(n842), .A2(n841), .ZN(G188) );
  INV_X1 U935 ( .A(G132), .ZN(G219) );
  INV_X1 U936 ( .A(G120), .ZN(G236) );
  INV_X1 U937 ( .A(G82), .ZN(G220) );
  INV_X1 U938 ( .A(G69), .ZN(G235) );
  NOR2_X1 U939 ( .A1(n844), .A2(n843), .ZN(G325) );
  INV_X1 U940 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U941 ( .A(KEYINPUT107), .B(n845), .ZN(G319) );
  XOR2_X1 U942 ( .A(G2096), .B(G2678), .Z(n847) );
  XNOR2_X1 U943 ( .A(G2072), .B(KEYINPUT43), .ZN(n846) );
  XNOR2_X1 U944 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U945 ( .A(n848), .B(KEYINPUT42), .Z(n850) );
  XNOR2_X1 U946 ( .A(G2067), .B(G2090), .ZN(n849) );
  XNOR2_X1 U947 ( .A(n850), .B(n849), .ZN(n854) );
  XOR2_X1 U948 ( .A(KEYINPUT108), .B(G2100), .Z(n852) );
  XNOR2_X1 U949 ( .A(G2078), .B(G2084), .ZN(n851) );
  XNOR2_X1 U950 ( .A(n852), .B(n851), .ZN(n853) );
  XNOR2_X1 U951 ( .A(n854), .B(n853), .ZN(G227) );
  XOR2_X1 U952 ( .A(G1981), .B(G1956), .Z(n856) );
  XNOR2_X1 U953 ( .A(G1986), .B(G1966), .ZN(n855) );
  XNOR2_X1 U954 ( .A(n856), .B(n855), .ZN(n860) );
  XOR2_X1 U955 ( .A(G1976), .B(G1971), .Z(n858) );
  XNOR2_X1 U956 ( .A(G1996), .B(G1991), .ZN(n857) );
  XNOR2_X1 U957 ( .A(n858), .B(n857), .ZN(n859) );
  XOR2_X1 U958 ( .A(n860), .B(n859), .Z(n862) );
  XNOR2_X1 U959 ( .A(KEYINPUT109), .B(KEYINPUT41), .ZN(n861) );
  XNOR2_X1 U960 ( .A(n862), .B(n861), .ZN(n864) );
  XOR2_X1 U961 ( .A(G1961), .B(G2474), .Z(n863) );
  XNOR2_X1 U962 ( .A(n864), .B(n863), .ZN(G229) );
  NAND2_X1 U963 ( .A1(G124), .A2(n891), .ZN(n865) );
  XNOR2_X1 U964 ( .A(n865), .B(KEYINPUT44), .ZN(n868) );
  NAND2_X1 U965 ( .A1(G100), .A2(n886), .ZN(n866) );
  XNOR2_X1 U966 ( .A(n866), .B(KEYINPUT110), .ZN(n867) );
  NAND2_X1 U967 ( .A1(n868), .A2(n867), .ZN(n872) );
  NAND2_X1 U968 ( .A1(G136), .A2(n887), .ZN(n870) );
  NAND2_X1 U969 ( .A1(G112), .A2(n892), .ZN(n869) );
  NAND2_X1 U970 ( .A1(n870), .A2(n869), .ZN(n871) );
  NOR2_X1 U971 ( .A1(n872), .A2(n871), .ZN(G162) );
  NAND2_X1 U972 ( .A1(G103), .A2(n886), .ZN(n874) );
  NAND2_X1 U973 ( .A1(G139), .A2(n887), .ZN(n873) );
  NAND2_X1 U974 ( .A1(n874), .A2(n873), .ZN(n879) );
  NAND2_X1 U975 ( .A1(n891), .A2(G127), .ZN(n876) );
  NAND2_X1 U976 ( .A1(G115), .A2(n892), .ZN(n875) );
  NAND2_X1 U977 ( .A1(n876), .A2(n875), .ZN(n877) );
  XOR2_X1 U978 ( .A(KEYINPUT47), .B(n877), .Z(n878) );
  NOR2_X1 U979 ( .A1(n879), .A2(n878), .ZN(n999) );
  XOR2_X1 U980 ( .A(KEYINPUT112), .B(KEYINPUT114), .Z(n881) );
  XNOR2_X1 U981 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n880) );
  XNOR2_X1 U982 ( .A(n881), .B(n880), .ZN(n882) );
  XOR2_X1 U983 ( .A(n882), .B(KEYINPUT113), .Z(n884) );
  XNOR2_X1 U984 ( .A(n1003), .B(KEYINPUT115), .ZN(n883) );
  XNOR2_X1 U985 ( .A(n884), .B(n883), .ZN(n903) );
  XNOR2_X1 U986 ( .A(G164), .B(n885), .ZN(n901) );
  NAND2_X1 U987 ( .A1(G106), .A2(n886), .ZN(n889) );
  NAND2_X1 U988 ( .A1(G142), .A2(n887), .ZN(n888) );
  NAND2_X1 U989 ( .A1(n889), .A2(n888), .ZN(n890) );
  XNOR2_X1 U990 ( .A(n890), .B(KEYINPUT45), .ZN(n897) );
  NAND2_X1 U991 ( .A1(n891), .A2(G130), .ZN(n894) );
  NAND2_X1 U992 ( .A1(G118), .A2(n892), .ZN(n893) );
  NAND2_X1 U993 ( .A1(n894), .A2(n893), .ZN(n895) );
  XNOR2_X1 U994 ( .A(KEYINPUT111), .B(n895), .ZN(n896) );
  NAND2_X1 U995 ( .A1(n897), .A2(n896), .ZN(n899) );
  XNOR2_X1 U996 ( .A(n899), .B(n898), .ZN(n900) );
  XNOR2_X1 U997 ( .A(n901), .B(n900), .ZN(n902) );
  XNOR2_X1 U998 ( .A(n903), .B(n902), .ZN(n906) );
  XNOR2_X1 U999 ( .A(n904), .B(G162), .ZN(n905) );
  XNOR2_X1 U1000 ( .A(n906), .B(n905), .ZN(n907) );
  XOR2_X1 U1001 ( .A(n999), .B(n907), .Z(n908) );
  XNOR2_X1 U1002 ( .A(G160), .B(n908), .ZN(n909) );
  NOR2_X1 U1003 ( .A1(G37), .A2(n909), .ZN(G395) );
  XOR2_X1 U1004 ( .A(n910), .B(G286), .Z(n912) );
  XNOR2_X1 U1005 ( .A(G171), .B(n921), .ZN(n911) );
  XNOR2_X1 U1006 ( .A(n912), .B(n911), .ZN(n913) );
  XOR2_X1 U1007 ( .A(n913), .B(n936), .Z(n914) );
  NOR2_X1 U1008 ( .A1(G37), .A2(n914), .ZN(G397) );
  NOR2_X1 U1009 ( .A1(G227), .A2(G229), .ZN(n915) );
  XOR2_X1 U1010 ( .A(KEYINPUT49), .B(n915), .Z(n916) );
  NAND2_X1 U1011 ( .A1(G319), .A2(n916), .ZN(n917) );
  NOR2_X1 U1012 ( .A1(G401), .A2(n917), .ZN(n918) );
  XNOR2_X1 U1013 ( .A(KEYINPUT116), .B(n918), .ZN(n920) );
  NOR2_X1 U1014 ( .A1(G395), .A2(G397), .ZN(n919) );
  NAND2_X1 U1015 ( .A1(n920), .A2(n919), .ZN(G225) );
  INV_X1 U1016 ( .A(G225), .ZN(G308) );
  INV_X1 U1017 ( .A(G108), .ZN(G238) );
  INV_X1 U1018 ( .A(G96), .ZN(G221) );
  XNOR2_X1 U1019 ( .A(G16), .B(KEYINPUT56), .ZN(n945) );
  XNOR2_X1 U1020 ( .A(G1348), .B(n921), .ZN(n922) );
  XNOR2_X1 U1021 ( .A(n922), .B(KEYINPUT122), .ZN(n926) );
  XNOR2_X1 U1022 ( .A(G1961), .B(G301), .ZN(n923) );
  NOR2_X1 U1023 ( .A1(n924), .A2(n923), .ZN(n925) );
  NAND2_X1 U1024 ( .A1(n926), .A2(n925), .ZN(n928) );
  XNOR2_X1 U1025 ( .A(G1956), .B(G299), .ZN(n927) );
  NOR2_X1 U1026 ( .A1(n928), .A2(n927), .ZN(n935) );
  XNOR2_X1 U1027 ( .A(G166), .B(G1971), .ZN(n930) );
  NAND2_X1 U1028 ( .A1(n930), .A2(n929), .ZN(n931) );
  NOR2_X1 U1029 ( .A1(n932), .A2(n931), .ZN(n933) );
  XOR2_X1 U1030 ( .A(KEYINPUT123), .B(n933), .Z(n934) );
  NAND2_X1 U1031 ( .A1(n935), .A2(n934), .ZN(n938) );
  XNOR2_X1 U1032 ( .A(G1341), .B(n936), .ZN(n937) );
  NOR2_X1 U1033 ( .A1(n938), .A2(n937), .ZN(n943) );
  XNOR2_X1 U1034 ( .A(G1966), .B(G168), .ZN(n940) );
  NAND2_X1 U1035 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1036 ( .A(n941), .B(KEYINPUT57), .ZN(n942) );
  NAND2_X1 U1037 ( .A1(n943), .A2(n942), .ZN(n944) );
  NAND2_X1 U1038 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1039 ( .A(KEYINPUT124), .B(n946), .ZN(n998) );
  XNOR2_X1 U1040 ( .A(G20), .B(n947), .ZN(n951) );
  XNOR2_X1 U1041 ( .A(G1341), .B(G19), .ZN(n949) );
  XNOR2_X1 U1042 ( .A(G1981), .B(G6), .ZN(n948) );
  NOR2_X1 U1043 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1044 ( .A1(n951), .A2(n950), .ZN(n955) );
  XNOR2_X1 U1045 ( .A(KEYINPUT59), .B(KEYINPUT125), .ZN(n952) );
  XNOR2_X1 U1046 ( .A(n952), .B(G4), .ZN(n953) );
  XNOR2_X1 U1047 ( .A(n953), .B(G1348), .ZN(n954) );
  NOR2_X1 U1048 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1049 ( .A(KEYINPUT60), .B(n956), .ZN(n957) );
  XNOR2_X1 U1050 ( .A(n957), .B(KEYINPUT126), .ZN(n961) );
  XNOR2_X1 U1051 ( .A(G1966), .B(G21), .ZN(n959) );
  XNOR2_X1 U1052 ( .A(G1961), .B(G5), .ZN(n958) );
  NOR2_X1 U1053 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1054 ( .A1(n961), .A2(n960), .ZN(n968) );
  XNOR2_X1 U1055 ( .A(G1971), .B(G22), .ZN(n963) );
  XNOR2_X1 U1056 ( .A(G23), .B(G1976), .ZN(n962) );
  NOR2_X1 U1057 ( .A1(n963), .A2(n962), .ZN(n965) );
  XOR2_X1 U1058 ( .A(G1986), .B(G24), .Z(n964) );
  NAND2_X1 U1059 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1060 ( .A(KEYINPUT58), .B(n966), .ZN(n967) );
  NOR2_X1 U1061 ( .A1(n968), .A2(n967), .ZN(n970) );
  XOR2_X1 U1062 ( .A(KEYINPUT127), .B(KEYINPUT61), .Z(n969) );
  XNOR2_X1 U1063 ( .A(n970), .B(n969), .ZN(n972) );
  INV_X1 U1064 ( .A(G16), .ZN(n971) );
  NAND2_X1 U1065 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1066 ( .A1(n973), .A2(G11), .ZN(n996) );
  XNOR2_X1 U1067 ( .A(G27), .B(n974), .ZN(n985) );
  XOR2_X1 U1068 ( .A(G1991), .B(G25), .Z(n975) );
  NAND2_X1 U1069 ( .A1(G28), .A2(n975), .ZN(n976) );
  XNOR2_X1 U1070 ( .A(n976), .B(KEYINPUT119), .ZN(n980) );
  XNOR2_X1 U1071 ( .A(G2067), .B(G26), .ZN(n978) );
  XNOR2_X1 U1072 ( .A(G2072), .B(G33), .ZN(n977) );
  NOR2_X1 U1073 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1074 ( .A1(n980), .A2(n979), .ZN(n983) );
  XNOR2_X1 U1075 ( .A(G32), .B(G1996), .ZN(n981) );
  XNOR2_X1 U1076 ( .A(KEYINPUT120), .B(n981), .ZN(n982) );
  NOR2_X1 U1077 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1078 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1079 ( .A(n986), .B(KEYINPUT53), .ZN(n989) );
  XOR2_X1 U1080 ( .A(G2084), .B(KEYINPUT54), .Z(n987) );
  XNOR2_X1 U1081 ( .A(G34), .B(n987), .ZN(n988) );
  NAND2_X1 U1082 ( .A1(n989), .A2(n988), .ZN(n991) );
  XNOR2_X1 U1083 ( .A(G35), .B(G2090), .ZN(n990) );
  NOR2_X1 U1084 ( .A1(n991), .A2(n990), .ZN(n992) );
  XOR2_X1 U1085 ( .A(KEYINPUT55), .B(n992), .Z(n993) );
  NOR2_X1 U1086 ( .A1(G29), .A2(n993), .ZN(n994) );
  XOR2_X1 U1087 ( .A(KEYINPUT121), .B(n994), .Z(n995) );
  NOR2_X1 U1088 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1089 ( .A1(n998), .A2(n997), .ZN(n1027) );
  XOR2_X1 U1090 ( .A(G2072), .B(n999), .Z(n1001) );
  XOR2_X1 U1091 ( .A(G164), .B(G2078), .Z(n1000) );
  NOR2_X1 U1092 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1093 ( .A(KEYINPUT50), .B(n1002), .ZN(n1015) );
  NOR2_X1 U1094 ( .A1(n1004), .A2(n1003), .ZN(n1008) );
  XOR2_X1 U1095 ( .A(G2084), .B(G160), .Z(n1005) );
  NOR2_X1 U1096 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1097 ( .A1(n1008), .A2(n1007), .ZN(n1013) );
  XNOR2_X1 U1098 ( .A(G162), .B(G2090), .ZN(n1010) );
  NAND2_X1 U1099 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XOR2_X1 U1100 ( .A(KEYINPUT51), .B(n1011), .Z(n1012) );
  NOR2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1102 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NOR2_X1 U1103 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1104 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1105 ( .A(n1020), .B(KEYINPUT52), .ZN(n1021) );
  XNOR2_X1 U1106 ( .A(KEYINPUT117), .B(n1021), .ZN(n1023) );
  INV_X1 U1107 ( .A(KEYINPUT55), .ZN(n1022) );
  NAND2_X1 U1108 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1109 ( .A1(n1024), .A2(G29), .ZN(n1025) );
  XOR2_X1 U1110 ( .A(KEYINPUT118), .B(n1025), .Z(n1026) );
  NOR2_X1 U1111 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XNOR2_X1 U1112 ( .A(KEYINPUT62), .B(n1028), .ZN(G311) );
  INV_X1 U1113 ( .A(G311), .ZN(G150) );
endmodule

