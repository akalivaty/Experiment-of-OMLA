//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 1 0 1 0 0 1 0 0 1 0 0 0 0 0 0 1 1 0 1 1 0 0 1 1 1 0 0 1 1 0 0 0 1 0 1 0 0 0 1 1 0 1 0 1 1 1 0 0 0 0 1 0 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:11 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1239, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1317,
    new_n1318;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  NOR2_X1   g0001(.A1(G97), .A2(G107), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n203), .A2(G87), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  INV_X1    g0006(.A(G264), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(G87), .ZN(new_n209));
  INV_X1    g0009(.A(G250), .ZN(new_n210));
  INV_X1    g0010(.A(G97), .ZN(new_n211));
  INV_X1    g0011(.A(G257), .ZN(new_n212));
  OAI22_X1  g0012(.A1(new_n209), .A2(new_n210), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  AOI211_X1 g0013(.A(new_n208), .B(new_n213), .C1(G68), .C2(G238), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G50), .A2(G226), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G77), .A2(G244), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G116), .A2(G270), .ZN(new_n217));
  NAND4_X1  g0017(.A1(new_n214), .A2(new_n215), .A3(new_n216), .A4(new_n217), .ZN(new_n218));
  AND2_X1   g0018(.A1(G58), .A2(G232), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n205), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT1), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n205), .A2(G13), .ZN(new_n222));
  OAI211_X1 g0022(.A(new_n222), .B(G250), .C1(G257), .C2(G264), .ZN(new_n223));
  XOR2_X1   g0023(.A(new_n223), .B(KEYINPUT0), .Z(new_n224));
  OAI21_X1  g0024(.A(G50), .B1(G58), .B2(G68), .ZN(new_n225));
  INV_X1    g0025(.A(G20), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  NOR3_X1   g0027(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  NOR3_X1   g0028(.A1(new_n221), .A2(new_n224), .A3(new_n228), .ZN(G361));
  XNOR2_X1  g0029(.A(KEYINPUT2), .B(G226), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XOR2_X1   g0032(.A(new_n231), .B(new_n232), .Z(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT64), .B(G264), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n233), .B(new_n237), .Z(G358));
  XOR2_X1   g0038(.A(G68), .B(G77), .Z(new_n239));
  XNOR2_X1  g0039(.A(G50), .B(G58), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G107), .B(G116), .Z(new_n242));
  XNOR2_X1  g0042(.A(G87), .B(G97), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G351));
  INV_X1    g0045(.A(KEYINPUT3), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(G33), .ZN(new_n247));
  INV_X1    g0047(.A(G33), .ZN(new_n248));
  AND3_X1   g0048(.A1(new_n248), .A2(KEYINPUT78), .A3(KEYINPUT3), .ZN(new_n249));
  AOI21_X1  g0049(.A(KEYINPUT78), .B1(new_n248), .B2(KEYINPUT3), .ZN(new_n250));
  OAI21_X1  g0050(.A(new_n247), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT7), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n251), .A2(new_n252), .A3(new_n226), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n248), .A2(KEYINPUT3), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT78), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n255), .B1(new_n246), .B2(G33), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n248), .A2(KEYINPUT78), .A3(KEYINPUT3), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n254), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  OAI21_X1  g0058(.A(KEYINPUT7), .B1(new_n258), .B2(G20), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n253), .A2(new_n259), .A3(G68), .ZN(new_n260));
  INV_X1    g0060(.A(G58), .ZN(new_n261));
  INV_X1    g0061(.A(G68), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NOR2_X1   g0063(.A1(G58), .A2(G68), .ZN(new_n264));
  OAI21_X1  g0064(.A(G20), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NOR2_X1   g0065(.A1(G20), .A2(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G159), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n260), .A2(KEYINPUT16), .A3(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT16), .ZN(new_n271));
  OAI21_X1  g0071(.A(KEYINPUT79), .B1(new_n248), .B2(KEYINPUT3), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT79), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n273), .A2(new_n246), .A3(G33), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n248), .A2(KEYINPUT3), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n272), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n276), .A2(KEYINPUT7), .A3(new_n226), .ZN(new_n277));
  XNOR2_X1  g0077(.A(KEYINPUT3), .B(G33), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n252), .B1(new_n278), .B2(G20), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n262), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n271), .B1(new_n280), .B2(new_n268), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n227), .B1(new_n205), .B2(new_n248), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n270), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G1), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(G20), .ZN(new_n285));
  INV_X1    g0085(.A(G13), .ZN(new_n286));
  OAI21_X1  g0086(.A(KEYINPUT68), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT68), .ZN(new_n288));
  NAND4_X1  g0088(.A1(new_n288), .A2(new_n284), .A3(G13), .A4(G20), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(new_n282), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n290), .A2(new_n291), .A3(new_n285), .ZN(new_n292));
  XOR2_X1   g0092(.A(KEYINPUT8), .B(G58), .Z(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  AND2_X1   g0094(.A1(new_n287), .A2(new_n289), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n294), .B1(new_n295), .B2(new_n293), .ZN(new_n296));
  AND2_X1   g0096(.A1(new_n283), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G200), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n256), .A2(new_n257), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n299), .A2(G226), .A3(G1698), .A4(new_n247), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(KEYINPUT80), .ZN(new_n301));
  INV_X1    g0101(.A(G1698), .ZN(new_n302));
  AND2_X1   g0102(.A1(new_n302), .A2(G223), .ZN(new_n303));
  AOI22_X1  g0103(.A1(new_n258), .A2(new_n303), .B1(G33), .B2(G87), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT80), .ZN(new_n305));
  NAND4_X1  g0105(.A1(new_n258), .A2(new_n305), .A3(G226), .A4(G1698), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n301), .A2(new_n304), .A3(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n227), .B1(G33), .B2(G41), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(G41), .ZN(new_n310));
  INV_X1    g0110(.A(G45), .ZN(new_n311));
  AOI21_X1  g0111(.A(G1), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n308), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(G232), .ZN(new_n314));
  XOR2_X1   g0114(.A(KEYINPUT65), .B(G45), .Z(new_n315));
  OAI211_X1 g0115(.A(new_n284), .B(G274), .C1(new_n315), .C2(G41), .ZN(new_n316));
  AND2_X1   g0116(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n298), .B1(new_n309), .B2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n309), .A2(G190), .A3(new_n317), .ZN(new_n320));
  NAND4_X1  g0120(.A1(new_n297), .A2(KEYINPUT81), .A3(new_n319), .A4(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT81), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n320), .A2(new_n283), .A3(new_n296), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n322), .B1(new_n323), .B2(new_n318), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n321), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(KEYINPUT17), .ZN(new_n326));
  AND3_X1   g0126(.A1(new_n320), .A2(new_n283), .A3(new_n296), .ZN(new_n327));
  XNOR2_X1  g0127(.A(KEYINPUT82), .B(KEYINPUT17), .ZN(new_n328));
  AND3_X1   g0128(.A1(new_n327), .A2(new_n319), .A3(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n326), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n309), .A2(new_n317), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(G169), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n309), .A2(G179), .A3(new_n317), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n283), .A2(new_n296), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  XOR2_X1   g0137(.A(new_n337), .B(KEYINPUT18), .Z(new_n338));
  NAND2_X1  g0138(.A1(new_n313), .A2(G244), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n278), .A2(G238), .A3(G1698), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n278), .A2(G232), .A3(new_n302), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n247), .A2(new_n275), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(G107), .ZN(new_n343));
  AND3_X1   g0143(.A1(new_n340), .A2(new_n341), .A3(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(new_n227), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n345), .B1(new_n248), .B2(new_n310), .ZN(new_n346));
  OAI211_X1 g0146(.A(new_n339), .B(new_n316), .C1(new_n344), .C2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(G169), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT69), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT67), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n351), .B1(new_n248), .B2(G20), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n226), .A2(KEYINPUT67), .A3(G33), .ZN(new_n353));
  AND2_X1   g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  XNOR2_X1  g0154(.A(KEYINPUT15), .B(G87), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n350), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  AOI22_X1  g0156(.A1(new_n293), .A2(new_n266), .B1(G20), .B2(G77), .ZN(new_n357));
  INV_X1    g0157(.A(new_n355), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n352), .A2(new_n353), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n358), .A2(new_n359), .A3(KEYINPUT69), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n356), .A2(new_n357), .A3(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(new_n282), .ZN(new_n362));
  INV_X1    g0162(.A(G77), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n295), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n290), .A2(new_n291), .A3(G77), .A4(new_n285), .ZN(new_n366));
  XNOR2_X1  g0166(.A(new_n366), .B(KEYINPUT70), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n349), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT73), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  OR2_X1    g0170(.A1(new_n347), .A2(G179), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT70), .ZN(new_n372));
  XNOR2_X1  g0172(.A(new_n366), .B(new_n372), .ZN(new_n373));
  AOI22_X1  g0173(.A1(new_n361), .A2(new_n282), .B1(new_n363), .B2(new_n295), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n375), .A2(KEYINPUT73), .A3(new_n349), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n370), .A2(new_n371), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n375), .A2(KEYINPUT71), .ZN(new_n378));
  INV_X1    g0178(.A(G190), .ZN(new_n379));
  OR2_X1    g0179(.A1(new_n347), .A2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT71), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n373), .A2(new_n374), .A3(new_n381), .ZN(new_n382));
  XOR2_X1   g0182(.A(KEYINPUT72), .B(G200), .Z(new_n383));
  NAND2_X1  g0183(.A1(new_n347), .A2(new_n383), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n378), .A2(new_n380), .A3(new_n382), .A4(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n377), .A2(new_n385), .ZN(new_n386));
  OAI211_X1 g0186(.A(new_n331), .B(new_n338), .C1(KEYINPUT74), .C2(new_n386), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n247), .A2(new_n275), .A3(G222), .A4(new_n302), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT66), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n278), .A2(KEYINPUT66), .A3(G222), .A4(new_n302), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n278), .A2(G223), .A3(G1698), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n342), .A2(G77), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n308), .B1(new_n392), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n313), .A2(G226), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n396), .A2(new_n316), .A3(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(G179), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n290), .A2(new_n291), .A3(G50), .A4(new_n285), .ZN(new_n402));
  INV_X1    g0202(.A(G50), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n295), .A2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(G150), .ZN(new_n405));
  INV_X1    g0205(.A(new_n266), .ZN(new_n406));
  NOR3_X1   g0206(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n407));
  OAI22_X1  g0207(.A1(new_n405), .A2(new_n406), .B1(new_n407), .B2(new_n226), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n408), .B1(new_n293), .B2(new_n359), .ZN(new_n409));
  OAI211_X1 g0209(.A(new_n402), .B(new_n404), .C1(new_n409), .C2(new_n291), .ZN(new_n410));
  OAI211_X1 g0210(.A(new_n401), .B(new_n410), .C1(G169), .C2(new_n399), .ZN(new_n411));
  INV_X1    g0211(.A(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n412), .B1(new_n386), .B2(KEYINPUT74), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT13), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n278), .A2(G232), .A3(G1698), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT77), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(G33), .A2(G97), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n278), .A2(G226), .A3(new_n302), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n278), .A2(KEYINPUT77), .A3(G232), .A4(G1698), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n417), .A2(new_n418), .A3(new_n419), .A4(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(new_n308), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n313), .A2(G238), .ZN(new_n423));
  AND4_X1   g0223(.A1(new_n414), .A2(new_n422), .A3(new_n316), .A4(new_n423), .ZN(new_n424));
  AOI22_X1  g0224(.A1(new_n421), .A2(new_n308), .B1(G238), .B2(new_n313), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n414), .B1(new_n425), .B2(new_n316), .ZN(new_n426));
  OAI21_X1  g0226(.A(G169), .B1(new_n424), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(KEYINPUT14), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n422), .A2(new_n316), .A3(new_n423), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(KEYINPUT13), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n425), .A2(new_n414), .A3(new_n316), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n430), .A2(G179), .A3(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT14), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n433), .B(G169), .C1(new_n424), .C2(new_n426), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n428), .A2(new_n432), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n295), .A2(new_n262), .ZN(new_n436));
  XNOR2_X1  g0236(.A(new_n436), .B(KEYINPUT12), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n354), .A2(new_n363), .ZN(new_n438));
  OAI22_X1  g0238(.A1(new_n406), .A2(new_n403), .B1(new_n226), .B2(G68), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n282), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT11), .ZN(new_n441));
  OR2_X1    g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n440), .A2(new_n441), .ZN(new_n443));
  OR2_X1    g0243(.A1(new_n292), .A2(new_n262), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n437), .A2(new_n442), .A3(new_n443), .A4(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n435), .A2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT9), .ZN(new_n447));
  AOI22_X1  g0247(.A1(new_n398), .A2(new_n383), .B1(new_n447), .B2(new_n410), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT75), .ZN(new_n449));
  OR2_X1    g0249(.A1(new_n410), .A2(new_n447), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n396), .A2(G190), .A3(new_n316), .A4(new_n397), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n448), .A2(new_n449), .A3(new_n450), .A4(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT76), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT10), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n448), .A2(KEYINPUT76), .A3(new_n450), .A4(new_n451), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n452), .A2(new_n453), .A3(KEYINPUT10), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n456), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  OAI21_X1  g0259(.A(G200), .B1(new_n424), .B2(new_n426), .ZN(new_n460));
  INV_X1    g0260(.A(new_n445), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n430), .A2(G190), .A3(new_n431), .ZN(new_n462));
  AND3_X1   g0262(.A1(new_n460), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n413), .A2(new_n446), .A3(new_n459), .A4(new_n464), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n387), .A2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n311), .A2(G1), .ZN(new_n468));
  AND2_X1   g0268(.A1(KEYINPUT5), .A2(G41), .ZN(new_n469));
  NOR2_X1   g0269(.A1(KEYINPUT5), .A2(G41), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n471), .A2(new_n346), .A3(G270), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT84), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n284), .A2(G45), .ZN(new_n474));
  INV_X1    g0274(.A(new_n470), .ZN(new_n475));
  NAND2_X1  g0275(.A1(KEYINPUT5), .A2(G41), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n473), .B1(new_n477), .B2(G274), .ZN(new_n478));
  OAI211_X1 g0278(.A(new_n468), .B(G274), .C1(new_n470), .C2(new_n469), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n479), .A2(KEYINPUT84), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n472), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT88), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  XNOR2_X1  g0283(.A(new_n479), .B(KEYINPUT84), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n484), .A2(KEYINPUT88), .A3(new_n472), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(G33), .A2(G283), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n487), .B(new_n226), .C1(G33), .C2(new_n211), .ZN(new_n488));
  INV_X1    g0288(.A(G116), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(G20), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n488), .A2(new_n282), .A3(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT20), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(KEYINPUT89), .ZN(new_n494));
  OR2_X1    g0294(.A1(new_n491), .A2(new_n492), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT89), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n491), .A2(new_n496), .A3(new_n492), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n494), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n284), .A2(G33), .ZN(new_n499));
  AND3_X1   g0299(.A1(new_n290), .A2(new_n291), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(G116), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n295), .A2(new_n489), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n498), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n258), .B1(G264), .B2(new_n302), .ZN(new_n504));
  NOR2_X1   g0304(.A1(G257), .A2(G1698), .ZN(new_n505));
  INV_X1    g0305(.A(G303), .ZN(new_n506));
  OAI22_X1  g0306(.A1(new_n504), .A2(new_n505), .B1(new_n506), .B2(new_n278), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(new_n308), .ZN(new_n508));
  AND4_X1   g0308(.A1(G179), .A2(new_n486), .A3(new_n503), .A4(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n503), .A2(G169), .ZN(new_n510));
  AOI22_X1  g0310(.A1(new_n483), .A2(new_n485), .B1(new_n308), .B2(new_n507), .ZN(new_n511));
  OAI21_X1  g0311(.A(KEYINPUT21), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n481), .A2(new_n482), .ZN(new_n513));
  AOI21_X1  g0313(.A(KEYINPUT88), .B1(new_n484), .B2(new_n472), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n508), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT21), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n515), .A2(new_n516), .A3(G169), .A4(new_n503), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n509), .B1(new_n512), .B2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT19), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n519), .B1(new_n354), .B2(new_n211), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n226), .B1(new_n418), .B2(new_n519), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n521), .B1(G87), .B2(new_n203), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n258), .A2(new_n226), .A3(G68), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n520), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  AOI22_X1  g0324(.A1(new_n524), .A2(new_n282), .B1(new_n295), .B2(new_n355), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n474), .A2(new_n210), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n346), .B(new_n526), .C1(G274), .C2(new_n474), .ZN(new_n527));
  MUX2_X1   g0327(.A(G238), .B(G244), .S(G1698), .Z(new_n528));
  AOI22_X1  g0328(.A1(new_n258), .A2(new_n528), .B1(G33), .B2(G116), .ZN(new_n529));
  OAI211_X1 g0329(.A(G190), .B(new_n527), .C1(new_n529), .C2(new_n346), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n527), .B1(new_n529), .B2(new_n346), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(new_n383), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n500), .A2(G87), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n525), .A2(new_n530), .A3(new_n532), .A4(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n500), .A2(new_n358), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n531), .A2(G169), .ZN(new_n537));
  OAI211_X1 g0337(.A(G179), .B(new_n527), .C1(new_n529), .C2(new_n346), .ZN(new_n538));
  AOI22_X1  g0338(.A1(new_n525), .A2(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n535), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n511), .A2(G190), .ZN(new_n541));
  INV_X1    g0341(.A(new_n503), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n541), .B(new_n542), .C1(new_n298), .C2(new_n511), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n518), .A2(new_n540), .A3(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT25), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n545), .B1(new_n290), .B2(G107), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n295), .A2(KEYINPUT25), .A3(new_n206), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n546), .A2(new_n547), .B1(new_n500), .B2(G107), .ZN(new_n548));
  INV_X1    g0348(.A(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT24), .ZN(new_n550));
  AND3_X1   g0350(.A1(new_n226), .A2(G33), .A3(G116), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT23), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n552), .B1(new_n226), .B2(G107), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n206), .A2(KEYINPUT23), .A3(G20), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n209), .A2(G20), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n555), .A2(new_n247), .A3(new_n275), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT22), .ZN(new_n557));
  AOI221_X4 g0357(.A(new_n551), .B1(new_n553), .B2(new_n554), .C1(new_n556), .C2(new_n557), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n299), .A2(KEYINPUT22), .A3(new_n247), .A4(new_n555), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n550), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n551), .B1(new_n556), .B2(new_n557), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n553), .A2(new_n554), .ZN(new_n562));
  AND4_X1   g0362(.A1(new_n550), .A2(new_n559), .A3(new_n561), .A4(new_n562), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n282), .B1(new_n560), .B2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT90), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n559), .A2(new_n561), .A3(new_n562), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(KEYINPUT24), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n559), .A2(new_n561), .A3(new_n550), .A4(new_n562), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n570), .A2(KEYINPUT90), .A3(new_n282), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n549), .B1(new_n566), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n210), .A2(new_n302), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n258), .B(new_n573), .C1(G257), .C2(new_n302), .ZN(new_n574));
  NAND2_X1  g0374(.A1(G33), .A2(G294), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n346), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n478), .A2(new_n480), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n471), .A2(new_n346), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n578), .A2(new_n207), .ZN(new_n579));
  NOR3_X1   g0379(.A1(new_n576), .A2(new_n577), .A3(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(G200), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n580), .A2(G190), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n572), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  AOI21_X1  g0384(.A(KEYINPUT90), .B1(new_n570), .B2(new_n282), .ZN(new_n585));
  AOI211_X1 g0385(.A(new_n565), .B(new_n291), .C1(new_n568), .C2(new_n569), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n548), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NOR4_X1   g0387(.A1(new_n576), .A2(new_n577), .A3(new_n579), .A4(G179), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n588), .B1(new_n581), .B2(new_n348), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n584), .A2(new_n590), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n544), .A2(new_n591), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n290), .A2(G97), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n500), .A2(G97), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n406), .A2(new_n363), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT6), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n211), .A2(new_n206), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n597), .B1(new_n598), .B2(new_n202), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n206), .A2(KEYINPUT6), .A3(G97), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n226), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n277), .A2(new_n279), .ZN(new_n602));
  AOI211_X1 g0402(.A(new_n596), .B(new_n601), .C1(new_n602), .C2(G107), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n594), .B(new_n595), .C1(new_n603), .C2(new_n291), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(KEYINPUT86), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n601), .B1(new_n602), .B2(G107), .ZN(new_n606));
  INV_X1    g0406(.A(new_n596), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n282), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT86), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n609), .A2(new_n610), .A3(new_n594), .A4(new_n595), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n302), .A2(G244), .ZN(new_n612));
  OAI21_X1  g0412(.A(KEYINPUT83), .B1(new_n251), .B2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT4), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT83), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n258), .A2(new_n615), .A3(G244), .A4(new_n302), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n613), .A2(new_n614), .A3(new_n616), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n278), .A2(KEYINPUT4), .A3(G244), .A4(new_n302), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n278), .A2(G250), .A3(G1698), .ZN(new_n619));
  AND3_X1   g0419(.A1(new_n618), .A2(new_n487), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n617), .A2(new_n620), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n577), .B1(new_n621), .B2(new_n308), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT85), .ZN(new_n623));
  INV_X1    g0423(.A(new_n578), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n623), .B1(new_n624), .B2(G257), .ZN(new_n625));
  NOR3_X1   g0425(.A1(new_n578), .A2(KEYINPUT85), .A3(new_n212), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n348), .B1(new_n622), .B2(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n346), .B1(new_n617), .B2(new_n620), .ZN(new_n630));
  NOR4_X1   g0430(.A1(new_n630), .A2(new_n627), .A3(new_n400), .A4(new_n577), .ZN(new_n631));
  OAI211_X1 g0431(.A(new_n605), .B(new_n611), .C1(new_n629), .C2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n622), .A2(new_n628), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(G200), .ZN(new_n634));
  NOR3_X1   g0434(.A1(new_n630), .A2(new_n627), .A3(new_n577), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(G190), .ZN(new_n636));
  INV_X1    g0436(.A(new_n604), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n634), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  AOI21_X1  g0438(.A(KEYINPUT87), .B1(new_n632), .B2(new_n638), .ZN(new_n639));
  AND3_X1   g0439(.A1(new_n632), .A2(new_n638), .A3(KEYINPUT87), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n592), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n467), .A2(new_n641), .ZN(G372));
  INV_X1    g0442(.A(KEYINPUT94), .ZN(new_n643));
  INV_X1    g0443(.A(new_n377), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n644), .B1(new_n435), .B2(new_n445), .ZN(new_n645));
  OR2_X1    g0445(.A1(new_n645), .A2(new_n463), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n329), .B1(new_n325), .B2(KEYINPUT17), .ZN(new_n647));
  OAI211_X1 g0447(.A(new_n643), .B(new_n338), .C1(new_n646), .C2(new_n647), .ZN(new_n648));
  NOR3_X1   g0448(.A1(new_n645), .A2(new_n647), .A3(new_n463), .ZN(new_n649));
  XNOR2_X1  g0449(.A(new_n337), .B(KEYINPUT18), .ZN(new_n650));
  OAI21_X1  g0450(.A(KEYINPUT94), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT95), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n459), .A2(new_n652), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n456), .A2(KEYINPUT95), .A3(new_n457), .A4(new_n458), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n648), .A2(new_n651), .A3(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT92), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n580), .A2(new_n400), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n658), .B1(G169), .B2(new_n580), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n657), .B1(new_n572), .B2(new_n659), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n587), .A2(KEYINPUT92), .A3(new_n589), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n660), .A2(new_n518), .A3(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT93), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n537), .A2(new_n538), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(KEYINPUT91), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT91), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n537), .A2(new_n667), .A3(new_n538), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n525), .A2(new_n536), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n535), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  AND4_X1   g0471(.A1(new_n584), .A2(new_n632), .A3(new_n638), .A4(new_n671), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n660), .A2(new_n518), .A3(new_n661), .A4(KEYINPUT93), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n664), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n540), .ZN(new_n675));
  OAI21_X1  g0475(.A(KEYINPUT26), .B1(new_n632), .B2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n668), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n667), .B1(new_n537), .B2(new_n538), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n670), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT26), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n621), .A2(new_n308), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n681), .A2(new_n628), .A3(G179), .A4(new_n484), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n682), .B1(new_n635), .B2(new_n348), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n671), .A2(new_n680), .A3(new_n683), .A4(new_n604), .ZN(new_n684));
  AND3_X1   g0484(.A1(new_n676), .A2(new_n679), .A3(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n674), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n466), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n656), .A2(new_n687), .A3(new_n411), .ZN(G369));
  NOR2_X1   g0488(.A1(new_n286), .A2(G20), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(new_n284), .ZN(new_n690));
  OR2_X1    g0490(.A1(new_n690), .A2(KEYINPUT27), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(KEYINPUT27), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n691), .A2(G213), .A3(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(G343), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n587), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n584), .A2(new_n590), .A3(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT96), .ZN(new_n698));
  OR2_X1    g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n697), .A2(new_n698), .ZN(new_n700));
  INV_X1    g0500(.A(new_n695), .ZN(new_n701));
  OAI211_X1 g0501(.A(new_n699), .B(new_n700), .C1(new_n590), .C2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(G330), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n512), .A2(new_n517), .ZN(new_n704));
  INV_X1    g0504(.A(new_n509), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n706), .A2(new_n503), .A3(new_n695), .ZN(new_n707));
  OAI211_X1 g0507(.A(new_n518), .B(new_n543), .C1(new_n542), .C2(new_n701), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n703), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  AND2_X1   g0509(.A1(new_n702), .A2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n518), .A2(new_n695), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n713), .B1(new_n699), .B2(new_n700), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n695), .B1(new_n660), .B2(new_n661), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n711), .A2(new_n716), .ZN(G399));
  INV_X1    g0517(.A(new_n222), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n718), .A2(G41), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NOR3_X1   g0520(.A1(new_n203), .A2(G87), .A3(G116), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n720), .A2(G1), .A3(new_n721), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n722), .B1(new_n225), .B2(new_n720), .ZN(new_n723));
  XNOR2_X1  g0523(.A(new_n723), .B(KEYINPUT28), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n683), .A2(new_n679), .A3(new_n534), .A4(new_n604), .ZN(new_n725));
  AOI22_X1  g0525(.A1(new_n725), .A2(KEYINPUT26), .B1(KEYINPUT98), .B2(new_n679), .ZN(new_n726));
  OR2_X1    g0526(.A1(new_n679), .A2(KEYINPUT98), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n632), .A2(new_n638), .A3(new_n584), .A4(new_n671), .ZN(new_n728));
  AND2_X1   g0528(.A1(new_n518), .A2(new_n590), .ZN(new_n729));
  OAI211_X1 g0529(.A(new_n726), .B(new_n727), .C1(new_n728), .C2(new_n729), .ZN(new_n730));
  NOR3_X1   g0530(.A1(new_n632), .A2(new_n675), .A3(KEYINPUT26), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n701), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n695), .B1(new_n674), .B2(new_n685), .ZN(new_n733));
  OAI211_X1 g0533(.A(new_n732), .B(KEYINPUT29), .C1(new_n733), .C2(KEYINPUT97), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n576), .A2(new_n579), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n511), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n538), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n737), .A2(KEYINPUT30), .A3(new_n738), .A4(new_n635), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT30), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n635), .A2(new_n738), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n740), .B1(new_n741), .B2(new_n736), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n511), .A2(G179), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n743), .A2(new_n633), .A3(new_n581), .A4(new_n531), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n739), .A2(new_n742), .A3(new_n744), .ZN(new_n745));
  AND3_X1   g0545(.A1(new_n745), .A2(KEYINPUT31), .A3(new_n695), .ZN(new_n746));
  AOI21_X1  g0546(.A(KEYINPUT31), .B1(new_n745), .B2(new_n695), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  OAI211_X1 g0548(.A(new_n592), .B(new_n701), .C1(new_n639), .C2(new_n640), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n703), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT29), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT97), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n752), .B1(new_n733), .B2(new_n753), .ZN(new_n754));
  AND3_X1   g0554(.A1(new_n734), .A2(new_n751), .A3(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n724), .B1(new_n755), .B2(G1), .ZN(G364));
  AOI21_X1  g0556(.A(new_n227), .B1(G20), .B2(new_n348), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n226), .A2(new_n379), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n383), .A2(new_n400), .A3(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(G87), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n226), .A2(new_n400), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n762), .A2(new_n379), .A3(G200), .ZN(new_n763));
  NOR2_X1   g0563(.A1(G179), .A2(G200), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n226), .B1(new_n764), .B2(G190), .ZN(new_n765));
  OAI221_X1 g0565(.A(new_n761), .B1(new_n262), .B2(new_n763), .C1(new_n211), .C2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n400), .A2(G200), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n226), .A2(G190), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(new_n363), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n758), .A2(new_n767), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n342), .B1(new_n772), .B2(G58), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n762), .A2(G190), .A3(G200), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n383), .A2(new_n400), .A3(new_n768), .ZN(new_n775));
  OAI221_X1 g0575(.A(new_n773), .B1(new_n403), .B2(new_n774), .C1(new_n206), .C2(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n768), .A2(new_n764), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(G159), .ZN(new_n779));
  XNOR2_X1  g0579(.A(new_n779), .B(KEYINPUT32), .ZN(new_n780));
  NOR4_X1   g0580(.A1(new_n766), .A2(new_n770), .A3(new_n776), .A4(new_n780), .ZN(new_n781));
  AOI22_X1  g0581(.A1(new_n760), .A2(G303), .B1(G329), .B2(new_n778), .ZN(new_n782));
  INV_X1    g0582(.A(G317), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n763), .B1(KEYINPUT33), .B2(new_n783), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n784), .B1(KEYINPUT33), .B2(new_n783), .ZN(new_n785));
  INV_X1    g0585(.A(new_n774), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n278), .B1(new_n786), .B2(G326), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n782), .A2(new_n785), .A3(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(G322), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n771), .A2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(G283), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n775), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(G311), .ZN(new_n793));
  INV_X1    g0593(.A(G294), .ZN(new_n794));
  OAI22_X1  g0594(.A1(new_n769), .A2(new_n793), .B1(new_n765), .B2(new_n794), .ZN(new_n795));
  NOR4_X1   g0595(.A1(new_n788), .A2(new_n790), .A3(new_n792), .A4(new_n795), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n757), .B1(new_n781), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n689), .A2(G45), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n720), .A2(G1), .A3(new_n798), .ZN(new_n799));
  XNOR2_X1  g0599(.A(new_n799), .B(KEYINPUT99), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n718), .A2(new_n342), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(G355), .ZN(new_n803));
  OAI22_X1  g0603(.A1(new_n241), .A2(new_n311), .B1(new_n225), .B2(new_n315), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n258), .A2(new_n718), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  OAI221_X1 g0606(.A(new_n803), .B1(G116), .B2(new_n222), .C1(new_n804), .C2(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(G13), .A2(G33), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n809), .A2(G20), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n810), .A2(new_n757), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n801), .B1(new_n807), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n707), .A2(new_n708), .ZN(new_n813));
  INV_X1    g0613(.A(new_n810), .ZN(new_n814));
  OAI211_X1 g0614(.A(new_n797), .B(new_n812), .C1(new_n813), .C2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n709), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(new_n801), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n813), .A2(G330), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n815), .B1(new_n817), .B2(new_n818), .ZN(G396));
  INV_X1    g0619(.A(KEYINPUT102), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n377), .A2(new_n820), .A3(new_n385), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n375), .A2(new_n695), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n385), .A2(KEYINPUT102), .ZN(new_n824));
  NAND4_X1  g0624(.A1(new_n824), .A2(new_n375), .A3(new_n377), .A4(new_n695), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n733), .A2(new_n827), .ZN(new_n828));
  AOI211_X1 g0628(.A(new_n695), .B(new_n826), .C1(new_n674), .C2(new_n685), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  XNOR2_X1  g0630(.A(new_n830), .B(new_n751), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n831), .A2(new_n801), .ZN(new_n832));
  INV_X1    g0632(.A(new_n769), .ZN(new_n833));
  AOI22_X1  g0633(.A1(G294), .A2(new_n772), .B1(new_n833), .B2(G116), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n834), .B1(new_n206), .B2(new_n759), .C1(new_n506), .C2(new_n774), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n775), .A2(new_n209), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n342), .B1(new_n765), .B2(new_n211), .C1(new_n763), .C2(new_n791), .ZN(new_n837));
  NOR3_X1   g0637(.A1(new_n835), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n838), .B1(new_n793), .B2(new_n777), .ZN(new_n839));
  INV_X1    g0639(.A(new_n763), .ZN(new_n840));
  AOI22_X1  g0640(.A1(new_n840), .A2(G150), .B1(new_n772), .B2(G143), .ZN(new_n841));
  INV_X1    g0641(.A(G137), .ZN(new_n842));
  INV_X1    g0642(.A(G159), .ZN(new_n843));
  OAI221_X1 g0643(.A(new_n841), .B1(new_n842), .B2(new_n774), .C1(new_n843), .C2(new_n769), .ZN(new_n844));
  XNOR2_X1  g0644(.A(new_n844), .B(KEYINPUT34), .ZN(new_n845));
  INV_X1    g0645(.A(G132), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n258), .B1(new_n846), .B2(new_n777), .ZN(new_n847));
  XOR2_X1   g0647(.A(new_n847), .B(KEYINPUT101), .Z(new_n848));
  OAI211_X1 g0648(.A(new_n845), .B(new_n848), .C1(new_n261), .C2(new_n765), .ZN(new_n849));
  INV_X1    g0649(.A(new_n775), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(G68), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n851), .B1(new_n403), .B2(new_n759), .ZN(new_n852));
  XOR2_X1   g0652(.A(new_n852), .B(KEYINPUT100), .Z(new_n853));
  OAI21_X1  g0653(.A(new_n839), .B1(new_n849), .B2(new_n853), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n801), .B1(new_n854), .B2(new_n757), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n757), .A2(new_n808), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  OAI221_X1 g0657(.A(new_n855), .B1(G77), .B2(new_n857), .C1(new_n827), .C2(new_n809), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n832), .A2(new_n858), .ZN(G384));
  NOR2_X1   g0659(.A1(new_n461), .A2(new_n701), .ZN(new_n860));
  AOI211_X1 g0660(.A(new_n860), .B(new_n463), .C1(new_n435), .C2(new_n445), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n446), .A2(new_n701), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n827), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n863), .B1(new_n749), .B2(new_n748), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT104), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n865), .B1(new_n297), .B2(new_n693), .ZN(new_n866));
  INV_X1    g0666(.A(new_n693), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n336), .A2(KEYINPUT104), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n870), .B1(new_n647), .B2(new_n650), .ZN(new_n871));
  AOI21_X1  g0671(.A(KEYINPUT104), .B1(new_n336), .B2(new_n867), .ZN(new_n872));
  AOI211_X1 g0672(.A(new_n865), .B(new_n693), .C1(new_n283), .C2(new_n296), .ZN(new_n873));
  OAI221_X1 g0673(.A(new_n337), .B1(new_n318), .B2(new_n323), .C1(new_n872), .C2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(KEYINPUT37), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT37), .ZN(new_n876));
  NAND4_X1  g0676(.A1(new_n869), .A2(new_n325), .A3(new_n876), .A4(new_n337), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n871), .A2(new_n878), .ZN(new_n879));
  XNOR2_X1  g0679(.A(KEYINPUT105), .B(KEYINPUT38), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n260), .A2(new_n269), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(new_n271), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n883), .A2(new_n282), .A3(new_n270), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n693), .B1(new_n884), .B2(new_n296), .ZN(new_n885));
  AOI22_X1  g0685(.A1(new_n333), .A2(new_n334), .B1(new_n884), .B2(new_n296), .ZN(new_n886));
  AOI211_X1 g0686(.A(new_n885), .B(new_n886), .C1(new_n324), .C2(new_n321), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n877), .B1(new_n887), .B2(new_n876), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n885), .B1(new_n647), .B2(new_n650), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n888), .A2(new_n889), .A3(KEYINPUT38), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n881), .A2(new_n890), .ZN(new_n891));
  AND3_X1   g0691(.A1(new_n864), .A2(new_n891), .A3(KEYINPUT40), .ZN(new_n892));
  XOR2_X1   g0692(.A(KEYINPUT106), .B(KEYINPUT40), .Z(new_n893));
  INV_X1    g0693(.A(KEYINPUT38), .ZN(new_n894));
  INV_X1    g0694(.A(new_n885), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n895), .B1(new_n331), .B2(new_n338), .ZN(new_n896));
  INV_X1    g0696(.A(new_n886), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n325), .A2(new_n895), .A3(new_n897), .ZN(new_n898));
  OAI211_X1 g0698(.A(new_n337), .B(new_n876), .C1(new_n872), .C2(new_n873), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  AOI22_X1  g0700(.A1(KEYINPUT37), .A2(new_n898), .B1(new_n900), .B2(new_n325), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n894), .B1(new_n896), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(new_n890), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n893), .B1(new_n864), .B2(new_n903), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n892), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n748), .A2(new_n749), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n905), .A2(new_n466), .A3(new_n906), .ZN(new_n907));
  NOR3_X1   g0707(.A1(new_n892), .A2(new_n904), .A3(new_n703), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n751), .A2(new_n467), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n907), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT39), .ZN(new_n911));
  AND3_X1   g0711(.A1(new_n888), .A2(new_n889), .A3(KEYINPUT38), .ZN(new_n912));
  INV_X1    g0712(.A(new_n880), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n913), .B1(new_n871), .B2(new_n878), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n911), .B1(new_n912), .B2(new_n914), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n902), .A2(new_n890), .A3(KEYINPUT39), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n446), .A2(new_n695), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n686), .A2(new_n701), .A3(new_n827), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n377), .A2(new_n695), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n861), .A2(new_n862), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n922), .A2(new_n903), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n650), .A2(new_n693), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n918), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n910), .B(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n467), .B1(new_n734), .B2(new_n754), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n656), .A2(new_n411), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n928), .B(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(new_n284), .B2(new_n689), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n599), .A2(new_n600), .ZN(new_n934));
  OAI211_X1 g0734(.A(G20), .B(new_n345), .C1(new_n934), .C2(KEYINPUT35), .ZN(new_n935));
  AOI211_X1 g0735(.A(new_n489), .B(new_n935), .C1(KEYINPUT35), .C2(new_n934), .ZN(new_n936));
  XOR2_X1   g0736(.A(new_n936), .B(KEYINPUT36), .Z(new_n937));
  INV_X1    g0737(.A(KEYINPUT103), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(new_n262), .B2(G50), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n403), .A2(KEYINPUT103), .A3(G68), .ZN(new_n940));
  OAI21_X1  g0740(.A(G77), .B1(new_n261), .B2(new_n262), .ZN(new_n941));
  OAI211_X1 g0741(.A(new_n939), .B(new_n940), .C1(new_n941), .C2(new_n225), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n942), .A2(G1), .A3(new_n286), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n933), .A2(new_n937), .A3(new_n943), .ZN(G367));
  AND2_X1   g0744(.A1(new_n632), .A2(new_n638), .ZN(new_n945));
  AND3_X1   g0745(.A1(new_n714), .A2(KEYINPUT42), .A3(new_n945), .ZN(new_n946));
  AOI21_X1  g0746(.A(KEYINPUT42), .B1(new_n714), .B2(new_n945), .ZN(new_n947));
  OR2_X1    g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n701), .B1(new_n525), .B2(new_n533), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n671), .A2(new_n950), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n951), .B(KEYINPUT107), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n669), .A2(new_n670), .A3(new_n949), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(KEYINPUT108), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT108), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n952), .A2(new_n956), .A3(new_n953), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n958), .A2(KEYINPUT43), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n945), .B1(new_n637), .B2(new_n701), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n683), .A2(new_n604), .A3(new_n695), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n632), .B1(new_n963), .B2(new_n590), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n964), .A2(new_n701), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n948), .A2(new_n959), .A3(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT109), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND4_X1  g0768(.A1(new_n948), .A2(KEYINPUT109), .A3(new_n959), .A4(new_n965), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n711), .A2(new_n963), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n959), .B1(new_n948), .B2(new_n965), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n958), .A2(KEYINPUT43), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  AND3_X1   g0774(.A1(new_n970), .A2(new_n971), .A3(new_n974), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n971), .B1(new_n970), .B2(new_n974), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n719), .B(KEYINPUT41), .ZN(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n714), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n980), .B1(new_n702), .B2(new_n712), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n710), .B1(new_n981), .B2(new_n816), .ZN(new_n982));
  NAND4_X1  g0782(.A1(new_n982), .A2(new_n751), .A3(new_n754), .A4(new_n734), .ZN(new_n983));
  OR2_X1    g0783(.A1(new_n983), .A2(KEYINPUT110), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(KEYINPUT110), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n963), .B1(new_n714), .B2(new_n715), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT44), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n986), .B(new_n987), .ZN(new_n988));
  AND3_X1   g0788(.A1(new_n716), .A2(KEYINPUT45), .A3(new_n962), .ZN(new_n989));
  AOI21_X1  g0789(.A(KEYINPUT45), .B1(new_n716), .B2(new_n962), .ZN(new_n990));
  OAI211_X1 g0790(.A(new_n988), .B(new_n711), .C1(new_n989), .C2(new_n990), .ZN(new_n991));
  OR2_X1    g0791(.A1(new_n986), .A2(KEYINPUT44), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n986), .A2(KEYINPUT44), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n992), .B(new_n993), .C1(new_n989), .C2(new_n990), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(new_n710), .ZN(new_n995));
  NAND4_X1  g0795(.A1(new_n984), .A2(new_n985), .A3(new_n991), .A4(new_n995), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n979), .B1(new_n996), .B2(new_n755), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n798), .A2(G1), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n977), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n955), .A2(new_n810), .A3(new_n957), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(G50), .A2(new_n833), .B1(new_n778), .B2(G137), .ZN(new_n1001));
  INV_X1    g0801(.A(G143), .ZN(new_n1002));
  OAI221_X1 g0802(.A(new_n1001), .B1(new_n1002), .B2(new_n774), .C1(new_n843), .C2(new_n763), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1003), .B1(G58), .B2(new_n760), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n342), .B1(new_n772), .B2(G150), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n765), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1006), .A2(G68), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n850), .A2(G77), .ZN(new_n1008));
  NAND4_X1  g0808(.A1(new_n1004), .A2(new_n1005), .A3(new_n1007), .A4(new_n1008), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n251), .B1(new_n783), .B2(new_n777), .ZN(new_n1010));
  OAI22_X1  g0810(.A1(new_n775), .A2(new_n211), .B1(new_n793), .B2(new_n774), .ZN(new_n1011));
  AOI211_X1 g0811(.A(new_n1010), .B(new_n1011), .C1(G294), .C2(new_n840), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n759), .A2(new_n489), .ZN(new_n1013));
  OR2_X1    g0813(.A1(new_n1013), .A2(KEYINPUT46), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(new_n1013), .A2(KEYINPUT46), .B1(G303), .B2(new_n772), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n833), .A2(G283), .ZN(new_n1016));
  NAND4_X1  g0816(.A1(new_n1012), .A2(new_n1014), .A3(new_n1015), .A4(new_n1016), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n765), .A2(new_n206), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1009), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT47), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1020), .A2(new_n757), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n811), .B1(new_n222), .B2(new_n355), .C1(new_n237), .C2(new_n806), .ZN(new_n1022));
  NAND4_X1  g0822(.A1(new_n1000), .A2(new_n800), .A3(new_n1021), .A4(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n999), .A2(new_n1023), .ZN(G387));
  NOR2_X1   g0824(.A1(new_n702), .A2(new_n814), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n806), .B1(new_n233), .B2(new_n315), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n721), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1026), .B1(new_n1027), .B2(new_n802), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n293), .A2(new_n403), .ZN(new_n1029));
  XOR2_X1   g0829(.A(new_n1029), .B(KEYINPUT111), .Z(new_n1030));
  OR2_X1    g0830(.A1(new_n1030), .A2(KEYINPUT50), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(G68), .A2(G77), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1027), .B1(new_n1030), .B2(KEYINPUT50), .ZN(new_n1033));
  AND4_X1   g0833(.A1(new_n311), .A2(new_n1031), .A3(new_n1032), .A4(new_n1033), .ZN(new_n1034));
  OAI22_X1  g0834(.A1(new_n1028), .A2(new_n1034), .B1(G107), .B2(new_n222), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1035), .A2(new_n811), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1036), .A2(new_n800), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n765), .A2(new_n355), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n775), .A2(new_n211), .B1(new_n843), .B2(new_n774), .ZN(new_n1039));
  AOI211_X1 g0839(.A(new_n1038), .B(new_n1039), .C1(G50), .C2(new_n772), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n760), .A2(G77), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(G68), .A2(new_n833), .B1(new_n778), .B2(G150), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n251), .B1(new_n840), .B2(new_n293), .ZN(new_n1043));
  NAND4_X1  g0843(.A1(new_n1040), .A2(new_n1041), .A3(new_n1042), .A4(new_n1043), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n763), .A2(new_n793), .B1(new_n774), .B2(new_n789), .ZN(new_n1045));
  XOR2_X1   g0845(.A(new_n1045), .B(KEYINPUT112), .Z(new_n1046));
  OAI221_X1 g0846(.A(new_n1046), .B1(new_n506), .B2(new_n769), .C1(new_n783), .C2(new_n771), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT48), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n1048), .B1(new_n791), .B2(new_n765), .C1(new_n794), .C2(new_n759), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT49), .ZN(new_n1050));
  OR2_X1    g0850(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n850), .A2(G116), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n778), .A2(G326), .ZN(new_n1053));
  NAND4_X1  g0853(.A1(new_n1051), .A2(new_n251), .A3(new_n1052), .A4(new_n1053), .ZN(new_n1054));
  AND2_X1   g0854(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1044), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  AOI211_X1 g0856(.A(new_n1025), .B(new_n1037), .C1(new_n1056), .C2(new_n757), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1057), .B1(new_n998), .B2(new_n982), .ZN(new_n1058));
  AND2_X1   g0858(.A1(new_n983), .A2(KEYINPUT110), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n983), .A2(KEYINPUT110), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n1059), .A2(new_n1060), .B1(new_n755), .B2(new_n982), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1058), .B1(new_n1061), .B2(new_n720), .ZN(G393));
  NAND2_X1  g0862(.A1(new_n995), .A2(new_n991), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1063), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1064), .A2(new_n996), .A3(new_n719), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n774), .A2(new_n405), .B1(new_n771), .B2(new_n843), .ZN(new_n1066));
  XOR2_X1   g0866(.A(new_n1066), .B(KEYINPUT51), .Z(new_n1067));
  OAI22_X1  g0867(.A1(new_n759), .A2(new_n262), .B1(new_n1002), .B2(new_n777), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n836), .B1(new_n1068), .B2(KEYINPUT114), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n1069), .B(new_n258), .C1(KEYINPUT114), .C2(new_n1068), .ZN(new_n1070));
  XOR2_X1   g0870(.A(new_n1070), .B(KEYINPUT115), .Z(new_n1071));
  AOI211_X1 g0871(.A(new_n1067), .B(new_n1071), .C1(new_n293), .C2(new_n833), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1006), .A2(G77), .ZN(new_n1073));
  OAI211_X1 g0873(.A(new_n1072), .B(new_n1073), .C1(new_n403), .C2(new_n763), .ZN(new_n1074));
  XOR2_X1   g0874(.A(new_n1074), .B(KEYINPUT116), .Z(new_n1075));
  OAI22_X1  g0875(.A1(new_n774), .A2(new_n783), .B1(new_n771), .B2(new_n793), .ZN(new_n1076));
  XOR2_X1   g0876(.A(new_n1076), .B(KEYINPUT52), .Z(new_n1077));
  OAI22_X1  g0877(.A1(new_n759), .A2(new_n791), .B1(new_n789), .B2(new_n777), .ZN(new_n1078));
  NOR3_X1   g0878(.A1(new_n1077), .A2(new_n278), .A3(new_n1078), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n840), .A2(G303), .B1(new_n1006), .B2(G116), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n1080), .A2(KEYINPUT117), .B1(new_n206), .B2(new_n775), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1081), .B1(KEYINPUT117), .B2(new_n1080), .ZN(new_n1082));
  OAI211_X1 g0882(.A(new_n1079), .B(new_n1082), .C1(new_n794), .C2(new_n769), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1075), .A2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n801), .B1(new_n1084), .B2(new_n757), .ZN(new_n1085));
  OAI221_X1 g0885(.A(new_n811), .B1(new_n211), .B2(new_n222), .C1(new_n244), .C2(new_n806), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n1085), .B(new_n1086), .C1(new_n814), .C2(new_n962), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1063), .A2(KEYINPUT113), .ZN(new_n1088));
  INV_X1    g0888(.A(KEYINPUT113), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n995), .A2(new_n991), .A3(new_n1089), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1088), .A2(new_n998), .A3(new_n1090), .ZN(new_n1091));
  AND3_X1   g0891(.A1(new_n1065), .A2(new_n1087), .A3(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1092), .ZN(G390));
  NOR3_X1   g0893(.A1(new_n929), .A2(new_n930), .A3(new_n909), .ZN(new_n1094));
  AND3_X1   g0894(.A1(new_n750), .A2(new_n827), .A3(new_n924), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n924), .B1(new_n750), .B2(new_n827), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n922), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n750), .A2(new_n827), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(new_n923), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n701), .B(new_n827), .C1(new_n730), .C2(new_n731), .ZN(new_n1100));
  AND2_X1   g0900(.A1(new_n1100), .A2(new_n921), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n750), .A2(new_n827), .A3(new_n924), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1099), .A2(new_n1101), .A3(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1097), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1094), .A2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n924), .B1(new_n829), .B2(new_n920), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n917), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n1106), .A2(new_n1107), .B1(new_n915), .B2(new_n916), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n891), .A2(new_n1107), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n923), .B1(new_n1100), .B2(new_n921), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NOR3_X1   g0911(.A1(new_n1108), .A2(new_n1111), .A3(new_n1095), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n920), .B1(new_n733), .B2(new_n827), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1107), .B1(new_n1113), .B2(new_n923), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n915), .A2(new_n916), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n917), .B1(new_n881), .B2(new_n890), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1117), .B1(new_n1101), .B2(new_n923), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1102), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1105), .B1(new_n1112), .B2(new_n1119), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1095), .B1(new_n1108), .B2(new_n1111), .ZN(new_n1121));
  AND2_X1   g0921(.A1(new_n915), .A2(new_n916), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n917), .B1(new_n922), .B2(new_n924), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n1118), .B(new_n1102), .C1(new_n1122), .C2(new_n1123), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n1121), .A2(new_n1124), .A3(new_n1094), .A4(new_n1104), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1120), .A2(new_n719), .A3(new_n1125), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1121), .A2(new_n998), .A3(new_n1124), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n786), .A2(G283), .ZN(new_n1128));
  NAND4_X1  g0928(.A1(new_n761), .A2(new_n851), .A3(new_n1073), .A4(new_n1128), .ZN(new_n1129));
  OAI221_X1 g0929(.A(new_n342), .B1(new_n769), .B2(new_n211), .C1(new_n763), .C2(new_n206), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  OAI221_X1 g0931(.A(new_n1131), .B1(new_n489), .B2(new_n771), .C1(new_n794), .C2(new_n777), .ZN(new_n1132));
  INV_X1    g0932(.A(G128), .ZN(new_n1133));
  OAI22_X1  g0933(.A1(new_n774), .A2(new_n1133), .B1(new_n771), .B2(new_n846), .ZN(new_n1134));
  XOR2_X1   g0934(.A(new_n1134), .B(KEYINPUT118), .Z(new_n1135));
  XOR2_X1   g0935(.A(KEYINPUT54), .B(G143), .Z(new_n1136));
  AOI21_X1  g0936(.A(new_n1135), .B1(new_n833), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1006), .A2(G159), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n759), .A2(new_n405), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(new_n1139), .B(KEYINPUT53), .ZN(new_n1140));
  OAI221_X1 g0940(.A(new_n278), .B1(new_n842), .B2(new_n763), .C1(new_n775), .C2(new_n403), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n1137), .A2(new_n1138), .A3(new_n1140), .A4(new_n1142), .ZN(new_n1143));
  AND2_X1   g0943(.A1(new_n778), .A2(G125), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1132), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n801), .B1(new_n1145), .B2(new_n757), .ZN(new_n1146));
  OAI221_X1 g0946(.A(new_n1146), .B1(new_n293), .B2(new_n857), .C1(new_n1122), .C2(new_n809), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1127), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1126), .A2(new_n1149), .ZN(G378));
  NAND2_X1  g0950(.A1(new_n905), .A2(G330), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n655), .A2(new_n411), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n410), .A2(new_n867), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(KEYINPUT120), .B(KEYINPUT55), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(new_n1153), .B(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1152), .A2(new_n1155), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(KEYINPUT121), .B(KEYINPUT56), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1155), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n655), .A2(new_n411), .A3(new_n1158), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1156), .A2(new_n1157), .A3(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1157), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1158), .B1(new_n655), .B2(new_n411), .ZN(new_n1162));
  AOI211_X1 g0962(.A(new_n412), .B(new_n1155), .C1(new_n653), .C2(new_n654), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1161), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1160), .A2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n923), .B1(new_n919), .B2(new_n921), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n1166), .A2(new_n903), .B1(new_n650), .B2(new_n693), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1165), .B1(new_n1167), .B2(new_n918), .ZN(new_n1168));
  AND4_X1   g0968(.A1(new_n918), .A2(new_n925), .A3(new_n1165), .A4(new_n926), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1151), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1165), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n927), .A2(new_n1171), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1167), .A2(new_n918), .A3(new_n1165), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1172), .A2(new_n908), .A3(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1170), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1125), .A2(new_n1094), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT57), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1175), .A2(new_n1176), .A3(KEYINPUT57), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1179), .A2(new_n719), .A3(new_n1180), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(new_n760), .A2(new_n1136), .B1(G137), .B2(new_n833), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(new_n840), .A2(G132), .B1(new_n1006), .B2(G150), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1182), .B(new_n1183), .C1(new_n1133), .C2(new_n771), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1184), .B1(G125), .B2(new_n786), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT59), .ZN(new_n1186));
  OR2_X1    g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n850), .A2(G159), .ZN(new_n1188));
  AOI21_X1  g0988(.A(G33), .B1(new_n778), .B2(G124), .ZN(new_n1189));
  NAND4_X1  g0989(.A1(new_n1187), .A2(new_n310), .A3(new_n1188), .A4(new_n1189), .ZN(new_n1190));
  AND2_X1   g0990(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1191));
  AOI21_X1  g0991(.A(G41), .B1(new_n258), .B2(G33), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n1190), .A2(new_n1191), .B1(G50), .B2(new_n1192), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n763), .A2(new_n211), .B1(new_n774), .B2(new_n489), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(G58), .B2(new_n850), .ZN(new_n1195));
  OAI211_X1 g0995(.A(new_n1195), .B(new_n1041), .C1(new_n791), .C2(new_n777), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n258), .B1(new_n833), .B2(new_n358), .ZN(new_n1197));
  OAI211_X1 g0997(.A(new_n1197), .B(new_n1007), .C1(new_n206), .C2(new_n771), .ZN(new_n1198));
  NOR3_X1   g0998(.A1(new_n1196), .A2(G41), .A3(new_n1198), .ZN(new_n1199));
  XNOR2_X1  g0999(.A(new_n1199), .B(KEYINPUT58), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n757), .B1(new_n1193), .B2(new_n1200), .ZN(new_n1201));
  XOR2_X1   g1001(.A(new_n1201), .B(KEYINPUT119), .Z(new_n1202));
  AOI211_X1 g1002(.A(new_n801), .B(new_n1202), .C1(new_n403), .C2(new_n856), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1171), .A2(new_n808), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1206), .B1(new_n1175), .B2(new_n998), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1181), .A2(new_n1207), .ZN(G375));
  OR3_X1    g1008(.A1(new_n929), .A2(new_n930), .A3(new_n909), .ZN(new_n1209));
  AND2_X1   g1009(.A1(new_n1097), .A2(new_n1103), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1211), .A2(new_n978), .A3(new_n1105), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n850), .A2(G58), .B1(G137), .B2(new_n772), .ZN(new_n1213));
  OAI221_X1 g1013(.A(new_n1213), .B1(new_n1133), .B2(new_n777), .C1(new_n843), .C2(new_n759), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n765), .A2(new_n403), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n774), .A2(new_n846), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1136), .ZN(new_n1217));
  OAI221_X1 g1017(.A(new_n258), .B1(new_n405), .B2(new_n769), .C1(new_n1217), .C2(new_n763), .ZN(new_n1218));
  NOR4_X1   g1018(.A1(new_n1214), .A2(new_n1215), .A3(new_n1216), .A4(new_n1218), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n850), .A2(G77), .B1(G303), .B2(new_n778), .ZN(new_n1220));
  OAI221_X1 g1020(.A(new_n1220), .B1(new_n211), .B2(new_n759), .C1(new_n794), .C2(new_n774), .ZN(new_n1221));
  OAI22_X1  g1021(.A1(new_n763), .A2(new_n489), .B1(new_n769), .B2(new_n206), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n1222), .A2(KEYINPUT122), .B1(G283), .B2(new_n772), .ZN(new_n1223));
  OAI221_X1 g1023(.A(new_n1223), .B1(KEYINPUT122), .B2(new_n1222), .C1(new_n355), .C2(new_n765), .ZN(new_n1224));
  NOR3_X1   g1024(.A1(new_n1221), .A2(new_n1224), .A3(new_n278), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n757), .B1(new_n1219), .B2(new_n1225), .ZN(new_n1226));
  OAI211_X1 g1026(.A(new_n1226), .B(new_n800), .C1(G68), .C2(new_n857), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1227), .B1(new_n923), .B2(new_n808), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1228), .B1(new_n1104), .B2(new_n998), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1212), .A2(new_n1229), .ZN(G381));
  NAND3_X1  g1030(.A1(new_n1092), .A2(new_n999), .A3(new_n1023), .ZN(new_n1231));
  NOR3_X1   g1031(.A1(new_n1231), .A2(G396), .A3(G393), .ZN(new_n1232));
  INV_X1    g1032(.A(G384), .ZN(new_n1233));
  NAND4_X1  g1033(.A1(new_n1232), .A2(new_n1233), .A3(new_n1229), .A4(new_n1212), .ZN(new_n1234));
  XNOR2_X1  g1034(.A(new_n1234), .B(KEYINPUT123), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(G375), .A2(G378), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1236), .ZN(new_n1237));
  OR2_X1    g1037(.A1(new_n1235), .A2(new_n1237), .ZN(G407));
  NAND2_X1  g1038(.A1(new_n1236), .A2(new_n694), .ZN(new_n1239));
  OAI211_X1 g1039(.A(new_n1239), .B(G213), .C1(new_n1235), .C2(new_n1237), .ZN(G409));
  XOR2_X1   g1040(.A(G393), .B(G396), .Z(new_n1241));
  AND3_X1   g1041(.A1(new_n1092), .A2(new_n999), .A3(new_n1023), .ZN(new_n1242));
  AND2_X1   g1042(.A1(new_n1091), .A2(new_n1087), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(new_n999), .A2(new_n1023), .B1(new_n1243), .B2(new_n1065), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1241), .B1(new_n1242), .B2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(G387), .A2(G390), .ZN(new_n1246));
  XNOR2_X1  g1046(.A(G393), .B(G396), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1246), .A2(new_n1231), .A3(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1245), .A2(new_n1248), .ZN(new_n1249));
  XNOR2_X1  g1049(.A(new_n1249), .B(KEYINPUT127), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n1112), .A2(new_n1119), .ZN(new_n1251));
  AND2_X1   g1051(.A1(new_n1094), .A2(new_n1104), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n720), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1148), .B1(new_n1253), .B2(new_n1120), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1254), .B1(new_n1181), .B2(new_n1207), .ZN(new_n1255));
  INV_X1    g1055(.A(G213), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1256), .A2(G343), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  AND3_X1   g1058(.A1(new_n1172), .A2(new_n908), .A3(new_n1173), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n908), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1260));
  OAI21_X1  g1060(.A(KEYINPUT124), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT124), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1170), .A2(new_n1262), .A3(new_n1174), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1261), .A2(new_n998), .A3(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1264), .A2(new_n1254), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1205), .B1(new_n1177), .B2(new_n979), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1258), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n1255), .A2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT60), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1211), .A2(new_n1269), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1209), .A2(new_n1210), .A3(KEYINPUT60), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(new_n1270), .A2(new_n719), .A3(new_n1105), .A4(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(new_n1229), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1273), .A2(new_n1233), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1272), .A2(G384), .A3(new_n1229), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1268), .A2(new_n1277), .ZN(new_n1278));
  XNOR2_X1  g1078(.A(new_n1278), .B(KEYINPUT62), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1257), .A2(G2897), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1276), .A2(new_n1280), .ZN(new_n1281));
  NAND4_X1  g1081(.A1(new_n1274), .A2(G2897), .A3(new_n1275), .A4(new_n1257), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1283), .B1(new_n1255), .B2(new_n1267), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT61), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1250), .B1(new_n1279), .B2(new_n1286), .ZN(new_n1287));
  AND3_X1   g1087(.A1(new_n1175), .A2(new_n1176), .A3(KEYINPUT57), .ZN(new_n1288));
  AOI21_X1  g1088(.A(KEYINPUT57), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1289));
  NOR3_X1   g1089(.A1(new_n1288), .A2(new_n1289), .A3(new_n720), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1207), .ZN(new_n1291));
  OAI21_X1  g1091(.A(G378), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1292));
  AND3_X1   g1092(.A1(new_n1170), .A2(new_n1262), .A3(new_n1174), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1262), .B1(new_n1170), .B2(new_n1174), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1295));
  AOI21_X1  g1095(.A(G378), .B1(new_n1295), .B2(new_n998), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1266), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1257), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT125), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1292), .A2(new_n1298), .A3(new_n1299), .ZN(new_n1300));
  OAI21_X1  g1100(.A(KEYINPUT125), .B1(new_n1255), .B2(new_n1267), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1300), .A2(new_n1301), .A3(new_n1283), .ZN(new_n1302));
  NOR3_X1   g1102(.A1(new_n1242), .A2(new_n1244), .A3(new_n1241), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1247), .B1(new_n1246), .B2(new_n1231), .ZN(new_n1304));
  NOR2_X1   g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  AND3_X1   g1105(.A1(new_n1302), .A2(new_n1285), .A3(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT63), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1307), .B1(new_n1268), .B2(new_n1277), .ZN(new_n1308));
  NOR4_X1   g1108(.A1(new_n1255), .A2(new_n1267), .A3(new_n1276), .A4(KEYINPUT63), .ZN(new_n1309));
  OR2_X1    g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  AOI21_X1  g1110(.A(KEYINPUT126), .B1(new_n1306), .B2(new_n1310), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1302), .A2(new_n1305), .A3(new_n1285), .ZN(new_n1312));
  NOR2_X1   g1112(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT126), .ZN(new_n1314));
  NOR3_X1   g1114(.A1(new_n1312), .A2(new_n1313), .A3(new_n1314), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1287), .B1(new_n1311), .B2(new_n1315), .ZN(G405));
  NOR2_X1   g1116(.A1(new_n1236), .A2(new_n1255), .ZN(new_n1317));
  XNOR2_X1  g1117(.A(new_n1249), .B(new_n1317), .ZN(new_n1318));
  XNOR2_X1  g1118(.A(new_n1318), .B(new_n1277), .ZN(G402));
endmodule


