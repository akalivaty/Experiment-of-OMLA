

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766;

  INV_X1 U370 ( .A(n728), .ZN(n347) );
  AND2_X1 U371 ( .A1(n372), .A2(n370), .ZN(n353) );
  NOR2_X1 U372 ( .A1(n706), .A2(n705), .ZN(n711) );
  XNOR2_X1 U373 ( .A(n636), .B(n418), .ZN(n705) );
  XNOR2_X1 U374 ( .A(n450), .B(n358), .ZN(n599) );
  XNOR2_X1 U375 ( .A(G143), .B(G128), .ZN(n501) );
  AND2_X2 U376 ( .A1(n744), .A2(n754), .ZN(n687) );
  XNOR2_X1 U377 ( .A(n346), .B(n472), .ZN(n654) );
  XNOR2_X1 U378 ( .A(n470), .B(G113), .ZN(n346) );
  OR2_X1 U379 ( .A1(n621), .A2(KEYINPUT48), .ZN(n431) );
  XNOR2_X2 U380 ( .A(n740), .B(n530), .ZN(n453) );
  XNOR2_X2 U381 ( .A(n512), .B(KEYINPUT3), .ZN(n514) );
  XNOR2_X1 U382 ( .A(KEYINPUT68), .B(G131), .ZN(n366) );
  INV_X2 U383 ( .A(KEYINPUT70), .ZN(n512) );
  XNOR2_X2 U384 ( .A(n486), .B(n487), .ZN(n573) );
  OR2_X1 U385 ( .A1(n619), .A2(KEYINPUT47), .ZN(n402) );
  NOR2_X1 U386 ( .A1(n764), .A2(n652), .ZN(n611) );
  XNOR2_X1 U387 ( .A(G116), .B(G107), .ZN(n479) );
  AND2_X1 U388 ( .A1(n411), .A2(n410), .ZN(n409) );
  AND2_X2 U389 ( .A1(n352), .A2(n353), .ZN(n754) );
  AND2_X1 U390 ( .A1(n620), .A2(n401), .ZN(n458) );
  NOR2_X1 U391 ( .A1(n371), .A2(n649), .ZN(n370) );
  XNOR2_X1 U392 ( .A(n555), .B(KEYINPUT35), .ZN(n763) );
  NAND2_X2 U393 ( .A1(n392), .A2(n388), .ZN(n696) );
  XNOR2_X1 U394 ( .A(n479), .B(G122), .ZN(n527) );
  INV_X1 U395 ( .A(KEYINPUT16), .ZN(n526) );
  XNOR2_X2 U396 ( .A(G110), .B(G104), .ZN(n506) );
  NAND2_X2 U397 ( .A1(n348), .A2(n356), .ZN(n441) );
  XNOR2_X2 U398 ( .A(n349), .B(n564), .ZN(n348) );
  NAND2_X1 U399 ( .A1(n350), .A2(n763), .ZN(n349) );
  NAND2_X1 U400 ( .A1(n384), .A2(n382), .ZN(n350) );
  NAND2_X1 U401 ( .A1(n351), .A2(n455), .ZN(n454) );
  INV_X1 U402 ( .A(n453), .ZN(n351) );
  XNOR2_X2 U403 ( .A(n529), .B(n528), .ZN(n740) );
  OR2_X1 U404 ( .A1(n375), .A2(n374), .ZN(n352) );
  BUF_X1 U405 ( .A(n576), .Z(n354) );
  XNOR2_X2 U406 ( .A(n589), .B(KEYINPUT19), .ZN(n612) );
  XNOR2_X2 U407 ( .A(n543), .B(n542), .ZN(n591) );
  NAND2_X1 U408 ( .A1(n449), .A2(n448), .ZN(n533) );
  NAND2_X1 U409 ( .A1(n460), .A2(G125), .ZN(n449) );
  NAND2_X1 U410 ( .A1(n459), .A2(G146), .ZN(n448) );
  XNOR2_X1 U411 ( .A(n501), .B(KEYINPUT4), .ZN(n539) );
  INV_X1 U412 ( .A(G214), .ZN(n467) );
  XNOR2_X1 U413 ( .A(n533), .B(n447), .ZN(n753) );
  XNOR2_X1 U414 ( .A(KEYINPUT10), .B(G140), .ZN(n447) );
  XNOR2_X1 U415 ( .A(n539), .B(n396), .ZN(n752) );
  XNOR2_X1 U416 ( .A(n366), .B(n397), .ZN(n396) );
  XNOR2_X1 U417 ( .A(n502), .B(G134), .ZN(n397) );
  INV_X1 U418 ( .A(G137), .ZN(n502) );
  OR2_X1 U419 ( .A1(n735), .A2(G902), .ZN(n450) );
  XNOR2_X1 U420 ( .A(KEYINPUT88), .B(KEYINPUT18), .ZN(n531) );
  XOR2_X1 U421 ( .A(KEYINPUT75), .B(KEYINPUT17), .Z(n532) );
  NAND2_X1 U422 ( .A1(n696), .A2(n629), .ZN(n395) );
  AND2_X1 U423 ( .A1(n621), .A2(n425), .ZN(n424) );
  INV_X1 U424 ( .A(G472), .ZN(n391) );
  NAND2_X1 U425 ( .A1(G902), .A2(G472), .ZN(n393) );
  XOR2_X1 U426 ( .A(KEYINPUT91), .B(G110), .Z(n494) );
  XNOR2_X1 U427 ( .A(G137), .B(G128), .ZN(n493) );
  XNOR2_X1 U428 ( .A(G119), .B(KEYINPUT23), .ZN(n490) );
  XOR2_X1 U429 ( .A(KEYINPUT24), .B(KEYINPUT92), .Z(n491) );
  XNOR2_X1 U430 ( .A(n483), .B(n482), .ZN(n489) );
  XOR2_X1 U431 ( .A(KEYINPUT74), .B(G140), .Z(n505) );
  XNOR2_X1 U432 ( .A(n752), .B(n504), .ZN(n522) );
  XNOR2_X1 U433 ( .A(KEYINPUT64), .B(G953), .ZN(n646) );
  XNOR2_X1 U434 ( .A(n367), .B(KEYINPUT33), .ZN(n715) );
  AND2_X1 U435 ( .A1(n632), .A2(n587), .ZN(n368) );
  INV_X1 U436 ( .A(KEYINPUT108), .ZN(n377) );
  NOR2_X1 U437 ( .A1(n588), .A2(n423), .ZN(n422) );
  AND2_X1 U438 ( .A1(n715), .A2(n552), .ZN(n553) );
  INV_X1 U439 ( .A(KEYINPUT22), .ZN(n451) );
  AND2_X1 U440 ( .A1(n708), .A2(n446), .ZN(n558) );
  XNOR2_X1 U441 ( .A(n595), .B(n406), .ZN(n405) );
  INV_X1 U442 ( .A(KEYINPUT28), .ZN(n406) );
  NAND2_X1 U443 ( .A1(n662), .A2(n657), .ZN(n410) );
  NAND2_X1 U444 ( .A1(n347), .A2(n408), .ZN(n407) );
  NAND2_X1 U445 ( .A1(n379), .A2(n442), .ZN(n385) );
  NOR2_X1 U446 ( .A1(n443), .A2(n599), .ZN(n442) );
  NOR2_X1 U447 ( .A1(n562), .A2(KEYINPUT65), .ZN(n443) );
  XNOR2_X1 U448 ( .A(n398), .B(KEYINPUT77), .ZN(n425) );
  INV_X1 U449 ( .A(G143), .ZN(n376) );
  XNOR2_X1 U450 ( .A(n540), .B(n536), .ZN(n455) );
  XNOR2_X1 U451 ( .A(KEYINPUT15), .B(G902), .ZN(n579) );
  NOR2_X1 U452 ( .A1(n637), .A2(n374), .ZN(n371) );
  NOR2_X1 U453 ( .A1(n686), .A2(KEYINPUT82), .ZN(n373) );
  XNOR2_X1 U454 ( .A(G104), .B(G122), .ZN(n461) );
  XOR2_X1 U455 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n462) );
  INV_X1 U456 ( .A(KEYINPUT66), .ZN(n503) );
  INV_X1 U457 ( .A(KEYINPUT38), .ZN(n418) );
  XNOR2_X1 U458 ( .A(n395), .B(n602), .ZN(n603) );
  XNOR2_X1 U459 ( .A(n476), .B(n475), .ZN(n572) );
  XNOR2_X1 U460 ( .A(n474), .B(n473), .ZN(n475) );
  NOR2_X1 U461 ( .A1(G902), .A2(n654), .ZN(n476) );
  NOR2_X1 U462 ( .A1(n694), .A2(n693), .ZN(n445) );
  XNOR2_X1 U463 ( .A(KEYINPUT93), .B(KEYINPUT94), .ZN(n515) );
  XNOR2_X1 U464 ( .A(KEYINPUT5), .B(G116), .ZN(n516) );
  NOR2_X1 U465 ( .A1(G953), .A2(G237), .ZN(n466) );
  XOR2_X1 U466 ( .A(KEYINPUT9), .B(KEYINPUT100), .Z(n478) );
  XNOR2_X1 U467 ( .A(G134), .B(KEYINPUT7), .ZN(n477) );
  INV_X1 U468 ( .A(KEYINPUT99), .ZN(n421) );
  BUF_X1 U469 ( .A(n658), .Z(n661) );
  INV_X1 U470 ( .A(G953), .ZN(n743) );
  NOR2_X1 U471 ( .A1(n622), .A2(n636), .ZN(n435) );
  XNOR2_X1 U472 ( .A(n571), .B(n570), .ZN(n607) );
  INV_X1 U473 ( .A(KEYINPUT102), .ZN(n570) );
  NOR2_X1 U474 ( .A1(n572), .A2(n573), .ZN(n571) );
  AND2_X1 U475 ( .A1(n394), .A2(n393), .ZN(n392) );
  NAND2_X1 U476 ( .A1(n391), .A2(n390), .ZN(n389) );
  XNOR2_X1 U477 ( .A(n400), .B(n399), .ZN(n735) );
  NAND2_X1 U478 ( .A1(n489), .A2(G221), .ZN(n399) );
  XNOR2_X1 U479 ( .A(n496), .B(n495), .ZN(n400) );
  XNOR2_X1 U480 ( .A(n522), .B(n510), .ZN(n369) );
  NOR2_X1 U481 ( .A1(n590), .A2(n561), .ZN(n684) );
  XNOR2_X1 U482 ( .A(n419), .B(KEYINPUT36), .ZN(n590) );
  AND2_X1 U483 ( .A1(n632), .A2(n694), .ZN(n416) );
  XNOR2_X1 U484 ( .A(n624), .B(KEYINPUT111), .ZN(n650) );
  AND2_X1 U485 ( .A1(n434), .A2(n433), .ZN(n624) );
  INV_X1 U486 ( .A(n623), .ZN(n433) );
  XNOR2_X1 U487 ( .A(n435), .B(KEYINPUT110), .ZN(n434) );
  XNOR2_X1 U488 ( .A(n404), .B(KEYINPUT76), .ZN(n676) );
  NOR2_X1 U489 ( .A1(n614), .A2(n613), .ZN(n404) );
  XNOR2_X1 U490 ( .A(n607), .B(KEYINPUT107), .ZN(n679) );
  INV_X1 U491 ( .A(KEYINPUT60), .ZN(n436) );
  INV_X1 U492 ( .A(KEYINPUT56), .ZN(n412) );
  NAND2_X1 U493 ( .A1(n409), .A2(n407), .ZN(n414) );
  NAND2_X1 U494 ( .A1(n381), .A2(n380), .ZN(n672) );
  AND2_X1 U495 ( .A1(n458), .A2(KEYINPUT48), .ZN(n355) );
  AND2_X1 U496 ( .A1(n578), .A2(n664), .ZN(n356) );
  INV_X1 U497 ( .A(n693), .ZN(n446) );
  AND2_X1 U498 ( .A1(n551), .A2(n550), .ZN(n357) );
  XOR2_X1 U499 ( .A(n498), .B(KEYINPUT25), .Z(n358) );
  AND2_X1 U500 ( .A1(n445), .A2(n632), .ZN(n359) );
  AND2_X1 U501 ( .A1(n562), .A2(KEYINPUT65), .ZN(n360) );
  XOR2_X1 U502 ( .A(KEYINPUT85), .B(KEYINPUT0), .Z(n361) );
  INV_X1 U503 ( .A(G902), .ZN(n390) );
  INV_X1 U504 ( .A(KEYINPUT82), .ZN(n374) );
  XOR2_X1 U505 ( .A(n426), .B(n643), .Z(n362) );
  XNOR2_X1 U506 ( .A(KEYINPUT59), .B(n654), .ZN(n363) );
  XNOR2_X1 U507 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n364) );
  AND2_X1 U508 ( .A1(n646), .A2(n645), .ZN(n739) );
  INV_X1 U509 ( .A(n739), .ZN(n438) );
  NAND2_X2 U510 ( .A1(n365), .A2(n561), .ZN(n576) );
  AND2_X1 U511 ( .A1(n365), .A2(n588), .ZN(n563) );
  XNOR2_X2 U512 ( .A(n560), .B(n451), .ZN(n365) );
  XNOR2_X1 U513 ( .A(n366), .B(n376), .ZN(n468) );
  NAND2_X1 U514 ( .A1(n368), .A2(n445), .ZN(n367) );
  NAND2_X1 U515 ( .A1(n369), .A2(n390), .ZN(n511) );
  XNOR2_X1 U516 ( .A(n369), .B(n364), .ZN(n729) );
  NAND2_X1 U517 ( .A1(n375), .A2(n373), .ZN(n372) );
  NAND2_X1 U518 ( .A1(n428), .A2(n427), .ZN(n375) );
  NAND2_X1 U519 ( .A1(n630), .A2(n589), .ZN(n419) );
  XNOR2_X2 U520 ( .A(n378), .B(n377), .ZN(n630) );
  NAND2_X1 U521 ( .A1(n422), .A2(n679), .ZN(n378) );
  NOR2_X2 U522 ( .A1(n444), .A2(KEYINPUT65), .ZN(n383) );
  NAND2_X1 U523 ( .A1(n385), .A2(n386), .ZN(n384) );
  NAND2_X1 U524 ( .A1(n444), .A2(n360), .ZN(n379) );
  INV_X1 U525 ( .A(n386), .ZN(n766) );
  NAND2_X1 U526 ( .A1(n386), .A2(n383), .ZN(n382) );
  XNOR2_X2 U527 ( .A(n387), .B(KEYINPUT32), .ZN(n386) );
  NAND2_X1 U528 ( .A1(n563), .A2(n416), .ZN(n387) );
  INV_X1 U529 ( .A(n385), .ZN(n380) );
  INV_X1 U530 ( .A(n383), .ZN(n381) );
  NAND2_X1 U531 ( .A1(n414), .A2(n438), .ZN(n413) );
  NAND2_X1 U532 ( .A1(n653), .A2(G475), .ZN(n440) );
  XNOR2_X1 U533 ( .A(n440), .B(n363), .ZN(n439) );
  XNOR2_X1 U534 ( .A(n413), .B(n412), .ZN(G51) );
  OR2_X1 U535 ( .A1(n426), .A2(n389), .ZN(n388) );
  NAND2_X1 U536 ( .A1(n426), .A2(G472), .ZN(n394) );
  NAND2_X1 U537 ( .A1(n627), .A2(n626), .ZN(n398) );
  NAND2_X1 U538 ( .A1(n403), .A2(n402), .ZN(n401) );
  OR2_X1 U539 ( .A1(n616), .A2(n615), .ZN(n403) );
  NAND2_X1 U540 ( .A1(n405), .A2(n596), .ZN(n613) );
  AND2_X1 U541 ( .A1(n415), .A2(G210), .ZN(n408) );
  NAND2_X1 U542 ( .A1(n728), .A2(n662), .ZN(n411) );
  INV_X1 U543 ( .A(n662), .ZN(n415) );
  NAND2_X1 U544 ( .A1(n417), .A2(n454), .ZN(n658) );
  NAND2_X1 U545 ( .A1(n453), .A2(n456), .ZN(n417) );
  XNOR2_X1 U546 ( .A(n535), .B(n540), .ZN(n456) );
  NAND2_X1 U547 ( .A1(n655), .A2(n656), .ZN(n728) );
  NAND2_X1 U548 ( .A1(n642), .A2(n641), .ZN(n655) );
  XNOR2_X1 U549 ( .A(n527), .B(n420), .ZN(n480) );
  XNOR2_X1 U550 ( .A(n501), .B(n421), .ZN(n420) );
  INV_X1 U551 ( .A(n594), .ZN(n423) );
  NAND2_X1 U552 ( .A1(n439), .A2(n438), .ZN(n437) );
  NAND2_X1 U553 ( .A1(n424), .A2(n355), .ZN(n427) );
  XNOR2_X1 U554 ( .A(n522), .B(n521), .ZN(n426) );
  AND2_X1 U555 ( .A1(n431), .A2(n429), .ZN(n428) );
  NAND2_X1 U556 ( .A1(n430), .A2(n628), .ZN(n429) );
  NAND2_X1 U557 ( .A1(n458), .A2(n425), .ZN(n430) );
  NAND2_X1 U558 ( .A1(n603), .A2(n604), .ZN(n622) );
  XNOR2_X1 U559 ( .A(n437), .B(n436), .ZN(G60) );
  XNOR2_X2 U560 ( .A(n441), .B(KEYINPUT45), .ZN(n744) );
  XNOR2_X2 U561 ( .A(n576), .B(KEYINPUT105), .ZN(n444) );
  XNOR2_X2 U562 ( .A(G119), .B(G113), .ZN(n513) );
  INV_X1 U563 ( .A(n445), .ZN(n691) );
  XNOR2_X1 U564 ( .A(n452), .B(n361), .ZN(n559) );
  NOR2_X2 U565 ( .A1(n612), .A2(n357), .ZN(n452) );
  XNOR2_X2 U566 ( .A(n506), .B(KEYINPUT87), .ZN(n524) );
  XNOR2_X1 U567 ( .A(KEYINPUT71), .B(KEYINPUT34), .ZN(n457) );
  INV_X1 U568 ( .A(KEYINPUT48), .ZN(n628) );
  INV_X1 U569 ( .A(KEYINPUT44), .ZN(n564) );
  XNOR2_X1 U570 ( .A(n505), .B(G107), .ZN(n507) );
  INV_X1 U571 ( .A(G475), .ZN(n473) );
  INV_X1 U572 ( .A(G125), .ZN(n459) );
  INV_X1 U573 ( .A(G146), .ZN(n460) );
  XNOR2_X1 U574 ( .A(n462), .B(n461), .ZN(n464) );
  XOR2_X1 U575 ( .A(KEYINPUT96), .B(KEYINPUT97), .Z(n463) );
  XNOR2_X1 U576 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U577 ( .A(n753), .B(n465), .ZN(n472) );
  XNOR2_X1 U578 ( .A(n466), .B(KEYINPUT73), .ZN(n518) );
  NOR2_X1 U579 ( .A1(n518), .A2(n467), .ZN(n469) );
  XOR2_X1 U580 ( .A(n469), .B(n468), .Z(n470) );
  XNOR2_X1 U581 ( .A(KEYINPUT98), .B(KEYINPUT13), .ZN(n474) );
  INV_X1 U582 ( .A(n572), .ZN(n556) );
  XNOR2_X1 U583 ( .A(KEYINPUT101), .B(G478), .ZN(n487) );
  XNOR2_X1 U584 ( .A(n478), .B(n477), .ZN(n481) );
  XOR2_X1 U585 ( .A(n481), .B(n480), .Z(n485) );
  INV_X1 U586 ( .A(n646), .ZN(n755) );
  NAND2_X1 U587 ( .A1(n755), .A2(G234), .ZN(n483) );
  XNOR2_X1 U588 ( .A(KEYINPUT67), .B(KEYINPUT8), .ZN(n482) );
  NAND2_X1 U589 ( .A1(G217), .A2(n489), .ZN(n484) );
  XNOR2_X1 U590 ( .A(n485), .B(n484), .ZN(n732) );
  NOR2_X1 U591 ( .A1(G902), .A2(n732), .ZN(n486) );
  NAND2_X1 U592 ( .A1(n556), .A2(n573), .ZN(n488) );
  XNOR2_X1 U593 ( .A(n488), .B(KEYINPUT106), .ZN(n623) );
  XNOR2_X1 U594 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U595 ( .A(n753), .B(n492), .ZN(n496) );
  XNOR2_X1 U596 ( .A(n494), .B(n493), .ZN(n495) );
  NAND2_X1 U597 ( .A1(n579), .A2(G234), .ZN(n497) );
  XNOR2_X1 U598 ( .A(n497), .B(KEYINPUT20), .ZN(n499) );
  NAND2_X1 U599 ( .A1(G217), .A2(n499), .ZN(n498) );
  INV_X1 U600 ( .A(n599), .ZN(n694) );
  NAND2_X1 U601 ( .A1(G221), .A2(n499), .ZN(n500) );
  XNOR2_X1 U602 ( .A(n500), .B(KEYINPUT21), .ZN(n693) );
  XNOR2_X1 U603 ( .A(n503), .B(G101), .ZN(n530) );
  XNOR2_X1 U604 ( .A(n530), .B(G146), .ZN(n504) );
  NAND2_X1 U605 ( .A1(G227), .A2(n755), .ZN(n509) );
  XNOR2_X1 U606 ( .A(n507), .B(n524), .ZN(n508) );
  XNOR2_X1 U607 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U608 ( .A(n511), .B(G469), .ZN(n596) );
  XNOR2_X1 U609 ( .A(n596), .B(KEYINPUT1), .ZN(n632) );
  XNOR2_X2 U610 ( .A(n514), .B(n513), .ZN(n525) );
  XNOR2_X1 U611 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U612 ( .A(n525), .B(n517), .ZN(n520) );
  INV_X1 U613 ( .A(G210), .ZN(n657) );
  OR2_X1 U614 ( .A1(n518), .A2(n657), .ZN(n519) );
  XNOR2_X1 U615 ( .A(n520), .B(n519), .ZN(n521) );
  INV_X1 U616 ( .A(KEYINPUT6), .ZN(n523) );
  XNOR2_X1 U617 ( .A(n696), .B(n523), .ZN(n587) );
  XNOR2_X2 U618 ( .A(n525), .B(n524), .ZN(n529) );
  XNOR2_X1 U619 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U620 ( .A(n532), .B(n531), .ZN(n534) );
  XOR2_X1 U621 ( .A(n534), .B(n533), .Z(n535) );
  INV_X1 U622 ( .A(n535), .ZN(n536) );
  INV_X1 U623 ( .A(G224), .ZN(n537) );
  NOR2_X1 U624 ( .A1(n646), .A2(n537), .ZN(n538) );
  XNOR2_X1 U625 ( .A(n539), .B(n538), .ZN(n540) );
  NAND2_X1 U626 ( .A1(n658), .A2(n579), .ZN(n543) );
  NOR2_X1 U627 ( .A1(G237), .A2(G902), .ZN(n541) );
  XOR2_X1 U628 ( .A(KEYINPUT72), .B(n541), .Z(n544) );
  NAND2_X1 U629 ( .A1(n544), .A2(G210), .ZN(n542) );
  NAND2_X1 U630 ( .A1(n544), .A2(G214), .ZN(n546) );
  INV_X1 U631 ( .A(KEYINPUT89), .ZN(n545) );
  XNOR2_X1 U632 ( .A(n546), .B(n545), .ZN(n629) );
  INV_X1 U633 ( .A(n629), .ZN(n706) );
  NOR2_X2 U634 ( .A1(n591), .A2(n706), .ZN(n589) );
  NAND2_X1 U635 ( .A1(G234), .A2(G237), .ZN(n547) );
  XNOR2_X1 U636 ( .A(KEYINPUT14), .B(n547), .ZN(n549) );
  NAND2_X1 U637 ( .A1(n549), .A2(G952), .ZN(n548) );
  XNOR2_X1 U638 ( .A(n548), .B(KEYINPUT90), .ZN(n720) );
  NOR2_X1 U639 ( .A1(G953), .A2(n720), .ZN(n584) );
  INV_X1 U640 ( .A(n584), .ZN(n551) );
  AND2_X1 U641 ( .A1(G902), .A2(n549), .ZN(n581) );
  NOR2_X1 U642 ( .A1(G898), .A2(n743), .ZN(n742) );
  NAND2_X1 U643 ( .A1(n581), .A2(n742), .ZN(n550) );
  BUF_X1 U644 ( .A(n559), .Z(n552) );
  XNOR2_X1 U645 ( .A(n553), .B(n457), .ZN(n554) );
  NOR2_X1 U646 ( .A1(n623), .A2(n554), .ZN(n555) );
  NOR2_X1 U647 ( .A1(n556), .A2(n573), .ZN(n557) );
  XNOR2_X1 U648 ( .A(n557), .B(KEYINPUT104), .ZN(n708) );
  NAND2_X1 U649 ( .A1(n559), .A2(n558), .ZN(n560) );
  INV_X1 U650 ( .A(n632), .ZN(n561) );
  INV_X1 U651 ( .A(n696), .ZN(n562) );
  AND2_X1 U652 ( .A1(n359), .A2(n696), .ZN(n700) );
  NAND2_X1 U653 ( .A1(n552), .A2(n700), .ZN(n565) );
  XNOR2_X1 U654 ( .A(KEYINPUT31), .B(n565), .ZN(n682) );
  INV_X1 U655 ( .A(n552), .ZN(n566) );
  NOR2_X1 U656 ( .A1(n566), .A2(n691), .ZN(n568) );
  INV_X1 U657 ( .A(n596), .ZN(n600) );
  NOR2_X1 U658 ( .A1(n600), .A2(n696), .ZN(n567) );
  AND2_X1 U659 ( .A1(n568), .A2(n567), .ZN(n667) );
  NOR2_X1 U660 ( .A1(n682), .A2(n667), .ZN(n569) );
  XNOR2_X1 U661 ( .A(n569), .B(KEYINPUT95), .ZN(n575) );
  NAND2_X1 U662 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U663 ( .A(n574), .B(KEYINPUT103), .Z(n666) );
  NAND2_X1 U664 ( .A1(n607), .A2(n666), .ZN(n710) );
  NAND2_X1 U665 ( .A1(n575), .A2(n710), .ZN(n578) );
  NOR2_X1 U666 ( .A1(n587), .A2(n354), .ZN(n577) );
  NAND2_X1 U667 ( .A1(n577), .A2(n599), .ZN(n664) );
  INV_X1 U668 ( .A(n579), .ZN(n640) );
  NAND2_X1 U669 ( .A1(n744), .A2(n640), .ZN(n580) );
  XNOR2_X1 U670 ( .A(n580), .B(KEYINPUT81), .ZN(n639) );
  NAND2_X1 U671 ( .A1(n581), .A2(n646), .ZN(n582) );
  NOR2_X1 U672 ( .A1(n582), .A2(G900), .ZN(n583) );
  NOR2_X1 U673 ( .A1(n584), .A2(n583), .ZN(n585) );
  NOR2_X1 U674 ( .A1(n585), .A2(n693), .ZN(n598) );
  XNOR2_X1 U675 ( .A(n598), .B(KEYINPUT69), .ZN(n586) );
  NOR2_X1 U676 ( .A1(n599), .A2(n586), .ZN(n594) );
  INV_X1 U677 ( .A(n587), .ZN(n588) );
  XNOR2_X1 U678 ( .A(n684), .B(KEYINPUT83), .ZN(n621) );
  XOR2_X1 U679 ( .A(KEYINPUT114), .B(KEYINPUT41), .Z(n593) );
  BUF_X2 U680 ( .A(n591), .Z(n636) );
  NAND2_X1 U681 ( .A1(n711), .A2(n708), .ZN(n592) );
  XNOR2_X1 U682 ( .A(n593), .B(n592), .ZN(n688) );
  NAND2_X1 U683 ( .A1(n594), .A2(n696), .ZN(n595) );
  NOR2_X1 U684 ( .A1(n688), .A2(n613), .ZN(n597) );
  XNOR2_X1 U685 ( .A(n597), .B(KEYINPUT42), .ZN(n764) );
  NAND2_X1 U686 ( .A1(n599), .A2(n598), .ZN(n601) );
  NOR2_X1 U687 ( .A1(n601), .A2(n600), .ZN(n604) );
  XNOR2_X1 U688 ( .A(KEYINPUT109), .B(KEYINPUT30), .ZN(n602) );
  NOR2_X1 U689 ( .A1(n705), .A2(n622), .ZN(n606) );
  XNOR2_X1 U690 ( .A(KEYINPUT84), .B(KEYINPUT39), .ZN(n605) );
  XNOR2_X1 U691 ( .A(n606), .B(n605), .ZN(n638) );
  NOR2_X1 U692 ( .A1(n607), .A2(n638), .ZN(n610) );
  XOR2_X1 U693 ( .A(KEYINPUT113), .B(KEYINPUT40), .Z(n608) );
  XNOR2_X1 U694 ( .A(n608), .B(KEYINPUT112), .ZN(n609) );
  XNOR2_X1 U695 ( .A(n610), .B(n609), .ZN(n652) );
  XNOR2_X1 U696 ( .A(n611), .B(KEYINPUT46), .ZN(n620) );
  BUF_X1 U697 ( .A(n612), .Z(n614) );
  XNOR2_X1 U698 ( .A(n676), .B(KEYINPUT79), .ZN(n616) );
  INV_X1 U699 ( .A(KEYINPUT47), .ZN(n615) );
  INV_X1 U700 ( .A(KEYINPUT79), .ZN(n618) );
  NAND2_X1 U701 ( .A1(n676), .A2(n710), .ZN(n617) );
  NAND2_X1 U702 ( .A1(n618), .A2(n617), .ZN(n619) );
  XNOR2_X1 U703 ( .A(n650), .B(KEYINPUT80), .ZN(n627) );
  INV_X1 U704 ( .A(n710), .ZN(n625) );
  NAND2_X1 U705 ( .A1(n625), .A2(KEYINPUT47), .ZN(n626) );
  NAND2_X1 U706 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U707 ( .A1(n632), .A2(n631), .ZN(n634) );
  INV_X1 U708 ( .A(KEYINPUT43), .ZN(n633) );
  XNOR2_X1 U709 ( .A(n634), .B(n633), .ZN(n635) );
  AND2_X1 U710 ( .A1(n636), .A2(n635), .ZN(n686) );
  INV_X1 U711 ( .A(n686), .ZN(n637) );
  NOR2_X1 U712 ( .A1(n638), .A2(n666), .ZN(n649) );
  NAND2_X1 U713 ( .A1(n639), .A2(n754), .ZN(n642) );
  NAND2_X1 U714 ( .A1(n640), .A2(KEYINPUT2), .ZN(n641) );
  NAND2_X1 U715 ( .A1(n687), .A2(KEYINPUT2), .ZN(n656) );
  AND2_X2 U716 ( .A1(n655), .A2(n656), .ZN(n653) );
  NAND2_X1 U717 ( .A1(n653), .A2(G472), .ZN(n644) );
  XNOR2_X1 U718 ( .A(KEYINPUT86), .B(KEYINPUT62), .ZN(n643) );
  XNOR2_X1 U719 ( .A(n644), .B(n362), .ZN(n647) );
  INV_X1 U720 ( .A(G952), .ZN(n645) );
  NAND2_X1 U721 ( .A1(n647), .A2(n438), .ZN(n648) );
  XNOR2_X1 U722 ( .A(n648), .B(KEYINPUT63), .ZN(G57) );
  XOR2_X1 U723 ( .A(G134), .B(n649), .Z(G36) );
  XNOR2_X1 U724 ( .A(n650), .B(G143), .ZN(G45) );
  XNOR2_X1 U725 ( .A(G131), .B(KEYINPUT127), .ZN(n651) );
  XNOR2_X1 U726 ( .A(n652), .B(n651), .ZN(G33) );
  XNOR2_X1 U727 ( .A(KEYINPUT78), .B(KEYINPUT54), .ZN(n659) );
  XOR2_X1 U728 ( .A(n659), .B(KEYINPUT55), .Z(n660) );
  XNOR2_X1 U729 ( .A(n661), .B(n660), .ZN(n662) );
  XOR2_X1 U730 ( .A(G101), .B(KEYINPUT115), .Z(n663) );
  XNOR2_X1 U731 ( .A(n664), .B(n663), .ZN(G3) );
  NAND2_X1 U732 ( .A1(n679), .A2(n667), .ZN(n665) );
  XNOR2_X1 U733 ( .A(n665), .B(G104), .ZN(G6) );
  XNOR2_X1 U734 ( .A(G107), .B(KEYINPUT27), .ZN(n671) );
  XOR2_X1 U735 ( .A(KEYINPUT26), .B(KEYINPUT116), .Z(n669) );
  INV_X1 U736 ( .A(n666), .ZN(n681) );
  NAND2_X1 U737 ( .A1(n667), .A2(n681), .ZN(n668) );
  XNOR2_X1 U738 ( .A(n669), .B(n668), .ZN(n670) );
  XNOR2_X1 U739 ( .A(n671), .B(n670), .ZN(G9) );
  XNOR2_X1 U740 ( .A(n672), .B(G110), .ZN(G12) );
  XOR2_X1 U741 ( .A(KEYINPUT29), .B(KEYINPUT117), .Z(n674) );
  NAND2_X1 U742 ( .A1(n681), .A2(n676), .ZN(n673) );
  XNOR2_X1 U743 ( .A(n674), .B(n673), .ZN(n675) );
  XOR2_X1 U744 ( .A(G128), .B(n675), .Z(G30) );
  NAND2_X1 U745 ( .A1(n676), .A2(n679), .ZN(n677) );
  XNOR2_X1 U746 ( .A(n677), .B(KEYINPUT118), .ZN(n678) );
  XNOR2_X1 U747 ( .A(G146), .B(n678), .ZN(G48) );
  NAND2_X1 U748 ( .A1(n679), .A2(n682), .ZN(n680) );
  XNOR2_X1 U749 ( .A(n680), .B(G113), .ZN(G15) );
  NAND2_X1 U750 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U751 ( .A(n683), .B(G116), .ZN(G18) );
  XNOR2_X1 U752 ( .A(G125), .B(n684), .ZN(n685) );
  XNOR2_X1 U753 ( .A(n685), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U754 ( .A(G140), .B(n686), .Z(G42) );
  XNOR2_X1 U755 ( .A(n687), .B(KEYINPUT2), .ZN(n725) );
  INV_X1 U756 ( .A(n688), .ZN(n703) );
  AND2_X1 U757 ( .A1(n703), .A2(n715), .ZN(n689) );
  XNOR2_X1 U758 ( .A(n689), .B(KEYINPUT121), .ZN(n690) );
  NAND2_X1 U759 ( .A1(n743), .A2(n690), .ZN(n723) );
  NAND2_X1 U760 ( .A1(n561), .A2(n691), .ZN(n692) );
  XNOR2_X1 U761 ( .A(n692), .B(KEYINPUT50), .ZN(n699) );
  NAND2_X1 U762 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U763 ( .A(KEYINPUT49), .B(n695), .ZN(n697) );
  NOR2_X1 U764 ( .A1(n697), .A2(n696), .ZN(n698) );
  AND2_X1 U765 ( .A1(n699), .A2(n698), .ZN(n701) );
  NOR2_X1 U766 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U767 ( .A(KEYINPUT51), .B(n702), .ZN(n704) );
  NAND2_X1 U768 ( .A1(n704), .A2(n703), .ZN(n717) );
  NAND2_X1 U769 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U770 ( .A1(n708), .A2(n707), .ZN(n709) );
  XOR2_X1 U771 ( .A(KEYINPUT119), .B(n709), .Z(n713) );
  NAND2_X1 U772 ( .A1(n711), .A2(n710), .ZN(n712) );
  NAND2_X1 U773 ( .A1(n713), .A2(n712), .ZN(n714) );
  NAND2_X1 U774 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U775 ( .A1(n717), .A2(n716), .ZN(n718) );
  XOR2_X1 U776 ( .A(KEYINPUT52), .B(n718), .Z(n719) );
  NOR2_X1 U777 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U778 ( .A(n721), .B(KEYINPUT120), .ZN(n722) );
  NOR2_X1 U779 ( .A1(n723), .A2(n722), .ZN(n724) );
  NAND2_X1 U780 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U781 ( .A(n726), .B(KEYINPUT122), .ZN(n727) );
  XOR2_X1 U782 ( .A(KEYINPUT53), .B(n727), .Z(G75) );
  NAND2_X1 U783 ( .A1(n347), .A2(G469), .ZN(n730) );
  XNOR2_X1 U784 ( .A(n730), .B(n729), .ZN(n731) );
  NOR2_X1 U785 ( .A1(n739), .A2(n731), .ZN(G54) );
  NAND2_X1 U786 ( .A1(n347), .A2(G478), .ZN(n733) );
  XNOR2_X1 U787 ( .A(n733), .B(n732), .ZN(n734) );
  NOR2_X1 U788 ( .A1(n739), .A2(n734), .ZN(G63) );
  NAND2_X1 U789 ( .A1(n347), .A2(G217), .ZN(n737) );
  XOR2_X1 U790 ( .A(n735), .B(KEYINPUT123), .Z(n736) );
  XNOR2_X1 U791 ( .A(n737), .B(n736), .ZN(n738) );
  NOR2_X1 U792 ( .A1(n739), .A2(n738), .ZN(G66) );
  XOR2_X1 U793 ( .A(n740), .B(G101), .Z(n741) );
  NOR2_X1 U794 ( .A1(n742), .A2(n741), .ZN(n751) );
  NAND2_X1 U795 ( .A1(n744), .A2(n743), .ZN(n745) );
  XNOR2_X1 U796 ( .A(n745), .B(KEYINPUT124), .ZN(n749) );
  NAND2_X1 U797 ( .A1(G953), .A2(G224), .ZN(n746) );
  XNOR2_X1 U798 ( .A(KEYINPUT61), .B(n746), .ZN(n747) );
  NAND2_X1 U799 ( .A1(n747), .A2(G898), .ZN(n748) );
  NAND2_X1 U800 ( .A1(n749), .A2(n748), .ZN(n750) );
  XNOR2_X1 U801 ( .A(n751), .B(n750), .ZN(G69) );
  XNOR2_X1 U802 ( .A(n753), .B(n752), .ZN(n757) );
  XNOR2_X1 U803 ( .A(n754), .B(n757), .ZN(n756) );
  NAND2_X1 U804 ( .A1(n756), .A2(n755), .ZN(n761) );
  XOR2_X1 U805 ( .A(G227), .B(n757), .Z(n758) );
  NAND2_X1 U806 ( .A1(n758), .A2(G900), .ZN(n759) );
  NAND2_X1 U807 ( .A1(G953), .A2(n759), .ZN(n760) );
  NAND2_X1 U808 ( .A1(n761), .A2(n760), .ZN(G72) );
  XOR2_X1 U809 ( .A(G122), .B(KEYINPUT125), .Z(n762) );
  XNOR2_X1 U810 ( .A(n763), .B(n762), .ZN(G24) );
  XOR2_X1 U811 ( .A(G137), .B(KEYINPUT126), .Z(n765) );
  XNOR2_X1 U812 ( .A(n764), .B(n765), .ZN(G39) );
  XOR2_X1 U813 ( .A(G119), .B(n766), .Z(G21) );
endmodule

