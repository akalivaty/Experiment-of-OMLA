

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585;

  XNOR2_X1 U323 ( .A(n549), .B(KEYINPUT65), .ZN(n569) );
  XNOR2_X1 U324 ( .A(n412), .B(n411), .ZN(n544) );
  XOR2_X1 U325 ( .A(n318), .B(KEYINPUT76), .Z(n291) );
  XOR2_X1 U326 ( .A(n397), .B(KEYINPUT17), .Z(n292) );
  XOR2_X1 U327 ( .A(KEYINPUT37), .B(n449), .Z(n293) );
  XOR2_X1 U328 ( .A(G71GAT), .B(G57GAT), .Z(n294) );
  XNOR2_X1 U329 ( .A(n497), .B(KEYINPUT46), .ZN(n498) );
  XNOR2_X1 U330 ( .A(KEYINPUT88), .B(KEYINPUT19), .ZN(n396) );
  NOR2_X1 U331 ( .A1(n419), .A2(n418), .ZN(n420) );
  XNOR2_X1 U332 ( .A(n404), .B(G190GAT), .ZN(n405) );
  XNOR2_X1 U333 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U334 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U335 ( .A(n329), .B(n328), .ZN(n573) );
  NOR2_X1 U336 ( .A1(n492), .A2(n480), .ZN(n451) );
  XNOR2_X1 U337 ( .A(n451), .B(KEYINPUT108), .ZN(n452) );
  INV_X1 U338 ( .A(G92GAT), .ZN(n453) );
  XOR2_X1 U339 ( .A(KEYINPUT30), .B(KEYINPUT70), .Z(n296) );
  XNOR2_X1 U340 ( .A(G141GAT), .B(G8GAT), .ZN(n295) );
  XNOR2_X1 U341 ( .A(n296), .B(n295), .ZN(n313) );
  XOR2_X1 U342 ( .A(G197GAT), .B(G113GAT), .Z(n298) );
  XNOR2_X1 U343 ( .A(G169GAT), .B(G43GAT), .ZN(n297) );
  XNOR2_X1 U344 ( .A(n298), .B(n297), .ZN(n300) );
  XOR2_X1 U345 ( .A(G36GAT), .B(G50GAT), .Z(n299) );
  XNOR2_X1 U346 ( .A(n300), .B(n299), .ZN(n309) );
  XNOR2_X1 U347 ( .A(KEYINPUT69), .B(KEYINPUT71), .ZN(n301) );
  XNOR2_X1 U348 ( .A(n301), .B(KEYINPUT29), .ZN(n302) );
  XOR2_X1 U349 ( .A(n302), .B(KEYINPUT72), .Z(n307) );
  XNOR2_X1 U350 ( .A(G29GAT), .B(KEYINPUT8), .ZN(n303) );
  XNOR2_X1 U351 ( .A(n303), .B(KEYINPUT7), .ZN(n334) );
  XOR2_X1 U352 ( .A(KEYINPUT73), .B(G1GAT), .Z(n305) );
  XNOR2_X1 U353 ( .A(G15GAT), .B(G22GAT), .ZN(n304) );
  XNOR2_X1 U354 ( .A(n305), .B(n304), .ZN(n358) );
  XNOR2_X1 U355 ( .A(n334), .B(n358), .ZN(n306) );
  XNOR2_X1 U356 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U357 ( .A(n309), .B(n308), .ZN(n311) );
  NAND2_X1 U358 ( .A1(G229GAT), .A2(G233GAT), .ZN(n310) );
  XNOR2_X1 U359 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U360 ( .A(n313), .B(n312), .ZN(n570) );
  INV_X1 U361 ( .A(n570), .ZN(n530) );
  XOR2_X1 U362 ( .A(G64GAT), .B(KEYINPUT77), .Z(n315) );
  XNOR2_X1 U363 ( .A(G204GAT), .B(G92GAT), .ZN(n314) );
  XNOR2_X1 U364 ( .A(n315), .B(n314), .ZN(n402) );
  XOR2_X1 U365 ( .A(G148GAT), .B(G78GAT), .Z(n366) );
  XOR2_X1 U366 ( .A(n402), .B(n366), .Z(n317) );
  XNOR2_X1 U367 ( .A(G120GAT), .B(G176GAT), .ZN(n316) );
  XNOR2_X1 U368 ( .A(n317), .B(n316), .ZN(n321) );
  XNOR2_X1 U369 ( .A(KEYINPUT13), .B(n294), .ZN(n359) );
  INV_X1 U370 ( .A(n359), .ZN(n318) );
  NAND2_X1 U371 ( .A1(G230GAT), .A2(G233GAT), .ZN(n319) );
  XNOR2_X1 U372 ( .A(n291), .B(n319), .ZN(n320) );
  XOR2_X1 U373 ( .A(n321), .B(n320), .Z(n329) );
  XOR2_X1 U374 ( .A(KEYINPUT74), .B(KEYINPUT75), .Z(n323) );
  XNOR2_X1 U375 ( .A(G106GAT), .B(G85GAT), .ZN(n322) );
  XNOR2_X1 U376 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U377 ( .A(G99GAT), .B(n324), .Z(n339) );
  XOR2_X1 U378 ( .A(KEYINPUT33), .B(KEYINPUT31), .Z(n326) );
  XNOR2_X1 U379 ( .A(KEYINPUT78), .B(KEYINPUT32), .ZN(n325) );
  XNOR2_X1 U380 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U381 ( .A(n339), .B(n327), .ZN(n328) );
  XOR2_X1 U382 ( .A(n573), .B(KEYINPUT41), .Z(n533) );
  INV_X1 U383 ( .A(n533), .ZN(n555) );
  NOR2_X1 U384 ( .A1(n530), .A2(n555), .ZN(n477) );
  XOR2_X1 U385 ( .A(KEYINPUT11), .B(KEYINPUT67), .Z(n331) );
  XNOR2_X1 U386 ( .A(G134GAT), .B(KEYINPUT9), .ZN(n330) );
  XNOR2_X1 U387 ( .A(n331), .B(n330), .ZN(n343) );
  XOR2_X1 U388 ( .A(G36GAT), .B(G218GAT), .Z(n408) );
  XOR2_X1 U389 ( .A(KEYINPUT10), .B(n408), .Z(n333) );
  XOR2_X1 U390 ( .A(G50GAT), .B(G162GAT), .Z(n376) );
  XNOR2_X1 U391 ( .A(n376), .B(G92GAT), .ZN(n332) );
  XNOR2_X1 U392 ( .A(n333), .B(n332), .ZN(n338) );
  XOR2_X1 U393 ( .A(n334), .B(KEYINPUT66), .Z(n336) );
  NAND2_X1 U394 ( .A1(G232GAT), .A2(G233GAT), .ZN(n335) );
  XNOR2_X1 U395 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U396 ( .A(n338), .B(n337), .Z(n341) );
  XOR2_X1 U397 ( .A(G43GAT), .B(G190GAT), .Z(n384) );
  XNOR2_X1 U398 ( .A(n384), .B(n339), .ZN(n340) );
  XNOR2_X1 U399 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U400 ( .A(n343), .B(n342), .Z(n539) );
  INV_X1 U401 ( .A(n539), .ZN(n561) );
  XNOR2_X1 U402 ( .A(KEYINPUT36), .B(n561), .ZN(n583) );
  XOR2_X1 U403 ( .A(G78GAT), .B(G127GAT), .Z(n345) );
  NAND2_X1 U404 ( .A1(G231GAT), .A2(G233GAT), .ZN(n344) );
  XNOR2_X1 U405 ( .A(n345), .B(n344), .ZN(n348) );
  XOR2_X1 U406 ( .A(KEYINPUT79), .B(G211GAT), .Z(n347) );
  XNOR2_X1 U407 ( .A(G8GAT), .B(G183GAT), .ZN(n346) );
  XNOR2_X1 U408 ( .A(n347), .B(n346), .ZN(n401) );
  XOR2_X1 U409 ( .A(n348), .B(n401), .Z(n356) );
  XOR2_X1 U410 ( .A(KEYINPUT14), .B(KEYINPUT80), .Z(n350) );
  XNOR2_X1 U411 ( .A(G155GAT), .B(G64GAT), .ZN(n349) );
  XNOR2_X1 U412 ( .A(n350), .B(n349), .ZN(n354) );
  XOR2_X1 U413 ( .A(KEYINPUT81), .B(KEYINPUT12), .Z(n352) );
  XNOR2_X1 U414 ( .A(KEYINPUT15), .B(KEYINPUT82), .ZN(n351) );
  XNOR2_X1 U415 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U416 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U417 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U418 ( .A(n358), .B(n357), .ZN(n360) );
  XOR2_X1 U419 ( .A(n360), .B(n359), .Z(n537) );
  INV_X1 U420 ( .A(n537), .ZN(n578) );
  INV_X1 U421 ( .A(KEYINPUT100), .ZN(n421) );
  XOR2_X1 U422 ( .A(KEYINPUT91), .B(G204GAT), .Z(n362) );
  XNOR2_X1 U423 ( .A(G22GAT), .B(KEYINPUT22), .ZN(n361) );
  XNOR2_X1 U424 ( .A(n362), .B(n361), .ZN(n380) );
  XOR2_X1 U425 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n364) );
  XNOR2_X1 U426 ( .A(G211GAT), .B(KEYINPUT94), .ZN(n363) );
  XNOR2_X1 U427 ( .A(n364), .B(n363), .ZN(n365) );
  XOR2_X1 U428 ( .A(n365), .B(G106GAT), .Z(n368) );
  XNOR2_X1 U429 ( .A(n366), .B(G218GAT), .ZN(n367) );
  XNOR2_X1 U430 ( .A(n368), .B(n367), .ZN(n372) );
  XOR2_X1 U431 ( .A(G197GAT), .B(KEYINPUT21), .Z(n403) );
  XOR2_X1 U432 ( .A(n403), .B(KEYINPUT93), .Z(n370) );
  NAND2_X1 U433 ( .A1(G228GAT), .A2(G233GAT), .ZN(n369) );
  XNOR2_X1 U434 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U435 ( .A(n372), .B(n371), .Z(n378) );
  XOR2_X1 U436 ( .A(KEYINPUT2), .B(KEYINPUT92), .Z(n374) );
  XNOR2_X1 U437 ( .A(KEYINPUT3), .B(G155GAT), .ZN(n373) );
  XNOR2_X1 U438 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U439 ( .A(G141GAT), .B(n375), .Z(n434) );
  XNOR2_X1 U440 ( .A(n434), .B(n376), .ZN(n377) );
  XNOR2_X1 U441 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U442 ( .A(n380), .B(n379), .Z(n550) );
  XOR2_X1 U443 ( .A(KEYINPUT20), .B(KEYINPUT86), .Z(n382) );
  XNOR2_X1 U444 ( .A(G99GAT), .B(KEYINPUT87), .ZN(n381) );
  XNOR2_X1 U445 ( .A(n382), .B(n381), .ZN(n383) );
  XOR2_X1 U446 ( .A(n384), .B(n383), .Z(n386) );
  NAND2_X1 U447 ( .A1(G227GAT), .A2(G233GAT), .ZN(n385) );
  XNOR2_X1 U448 ( .A(n386), .B(n385), .ZN(n390) );
  XOR2_X1 U449 ( .A(G183GAT), .B(G71GAT), .Z(n388) );
  XNOR2_X1 U450 ( .A(G15GAT), .B(KEYINPUT89), .ZN(n387) );
  XNOR2_X1 U451 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U452 ( .A(n390), .B(n389), .Z(n400) );
  XOR2_X1 U453 ( .A(KEYINPUT84), .B(KEYINPUT0), .Z(n392) );
  XNOR2_X1 U454 ( .A(G134GAT), .B(KEYINPUT85), .ZN(n391) );
  XNOR2_X1 U455 ( .A(n392), .B(n391), .ZN(n393) );
  XOR2_X1 U456 ( .A(n393), .B(G127GAT), .Z(n395) );
  XNOR2_X1 U457 ( .A(G113GAT), .B(G120GAT), .ZN(n394) );
  XNOR2_X1 U458 ( .A(n395), .B(n394), .ZN(n438) );
  XNOR2_X1 U459 ( .A(n396), .B(KEYINPUT18), .ZN(n397) );
  XNOR2_X1 U460 ( .A(G169GAT), .B(G176GAT), .ZN(n398) );
  XNOR2_X1 U461 ( .A(n292), .B(n398), .ZN(n406) );
  XNOR2_X1 U462 ( .A(n438), .B(n406), .ZN(n399) );
  XNOR2_X1 U463 ( .A(n400), .B(n399), .ZN(n552) );
  XNOR2_X1 U464 ( .A(n402), .B(n401), .ZN(n412) );
  XOR2_X1 U465 ( .A(KEYINPUT99), .B(n403), .Z(n404) );
  XOR2_X1 U466 ( .A(n408), .B(n407), .Z(n410) );
  NAND2_X1 U467 ( .A1(G226GAT), .A2(G233GAT), .ZN(n409) );
  XNOR2_X1 U468 ( .A(n410), .B(n409), .ZN(n411) );
  NAND2_X1 U469 ( .A1(n552), .A2(n544), .ZN(n413) );
  NAND2_X1 U470 ( .A1(n550), .A2(n413), .ZN(n414) );
  XNOR2_X1 U471 ( .A(n414), .B(KEYINPUT25), .ZN(n419) );
  INV_X1 U472 ( .A(KEYINPUT27), .ZN(n415) );
  XNOR2_X1 U473 ( .A(n544), .B(n415), .ZN(n443) );
  NOR2_X1 U474 ( .A1(n550), .A2(n552), .ZN(n416) );
  XNOR2_X1 U475 ( .A(n416), .B(KEYINPUT26), .ZN(n568) );
  INV_X1 U476 ( .A(n568), .ZN(n417) );
  NOR2_X1 U477 ( .A1(n443), .A2(n417), .ZN(n418) );
  XNOR2_X1 U478 ( .A(n421), .B(n420), .ZN(n439) );
  XOR2_X1 U479 ( .A(KEYINPUT95), .B(KEYINPUT5), .Z(n423) );
  XNOR2_X1 U480 ( .A(G1GAT), .B(KEYINPUT96), .ZN(n422) );
  XNOR2_X1 U481 ( .A(n423), .B(n422), .ZN(n427) );
  XOR2_X1 U482 ( .A(KEYINPUT6), .B(KEYINPUT4), .Z(n425) );
  XNOR2_X1 U483 ( .A(G57GAT), .B(KEYINPUT1), .ZN(n424) );
  XNOR2_X1 U484 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U485 ( .A(n427), .B(n426), .Z(n436) );
  XOR2_X1 U486 ( .A(G85GAT), .B(G148GAT), .Z(n429) );
  XNOR2_X1 U487 ( .A(G29GAT), .B(G162GAT), .ZN(n428) );
  XNOR2_X1 U488 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U489 ( .A(KEYINPUT97), .B(n430), .Z(n432) );
  NAND2_X1 U490 ( .A1(G225GAT), .A2(G233GAT), .ZN(n431) );
  XNOR2_X1 U491 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U492 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U493 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U494 ( .A(n438), .B(n437), .Z(n442) );
  NAND2_X1 U495 ( .A1(n439), .A2(n442), .ZN(n446) );
  XOR2_X1 U496 ( .A(n550), .B(KEYINPUT68), .Z(n440) );
  XNOR2_X1 U497 ( .A(KEYINPUT28), .B(n440), .ZN(n512) );
  XNOR2_X1 U498 ( .A(KEYINPUT90), .B(n552), .ZN(n441) );
  NOR2_X1 U499 ( .A1(n512), .A2(n441), .ZN(n444) );
  XNOR2_X1 U500 ( .A(KEYINPUT98), .B(n442), .ZN(n548) );
  NOR2_X1 U501 ( .A1(n443), .A2(n548), .ZN(n508) );
  NAND2_X1 U502 ( .A1(n444), .A2(n508), .ZN(n445) );
  NAND2_X1 U503 ( .A1(n446), .A2(n445), .ZN(n447) );
  XOR2_X1 U504 ( .A(KEYINPUT101), .B(n447), .Z(n457) );
  NAND2_X1 U505 ( .A1(n578), .A2(n457), .ZN(n448) );
  NOR2_X1 U506 ( .A1(n583), .A2(n448), .ZN(n449) );
  NAND2_X1 U507 ( .A1(n477), .A2(n293), .ZN(n450) );
  XOR2_X1 U508 ( .A(KEYINPUT107), .B(n450), .Z(n492) );
  INV_X1 U509 ( .A(n544), .ZN(n480) );
  XNOR2_X1 U510 ( .A(n453), .B(n452), .ZN(G1337GAT) );
  NOR2_X1 U511 ( .A1(n573), .A2(n570), .ZN(n466) );
  NOR2_X1 U512 ( .A1(n578), .A2(n539), .ZN(n454) );
  XNOR2_X1 U513 ( .A(n454), .B(KEYINPUT16), .ZN(n455) );
  XOR2_X1 U514 ( .A(KEYINPUT83), .B(n455), .Z(n456) );
  AND2_X1 U515 ( .A1(n457), .A2(n456), .ZN(n476) );
  NAND2_X1 U516 ( .A1(n466), .A2(n476), .ZN(n464) );
  NOR2_X1 U517 ( .A1(n548), .A2(n464), .ZN(n458) );
  XOR2_X1 U518 ( .A(G1GAT), .B(n458), .Z(n459) );
  XNOR2_X1 U519 ( .A(KEYINPUT34), .B(n459), .ZN(G1324GAT) );
  NOR2_X1 U520 ( .A1(n480), .A2(n464), .ZN(n460) );
  XOR2_X1 U521 ( .A(G8GAT), .B(n460), .Z(G1325GAT) );
  INV_X1 U522 ( .A(n552), .ZN(n490) );
  NOR2_X1 U523 ( .A1(n490), .A2(n464), .ZN(n462) );
  XNOR2_X1 U524 ( .A(KEYINPUT102), .B(KEYINPUT35), .ZN(n461) );
  XNOR2_X1 U525 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U526 ( .A(G15GAT), .B(n463), .ZN(G1326GAT) );
  INV_X1 U527 ( .A(n512), .ZN(n493) );
  NOR2_X1 U528 ( .A1(n493), .A2(n464), .ZN(n465) );
  XOR2_X1 U529 ( .A(G22GAT), .B(n465), .Z(G1327GAT) );
  NAND2_X1 U530 ( .A1(n466), .A2(n293), .ZN(n467) );
  XNOR2_X1 U531 ( .A(n467), .B(KEYINPUT38), .ZN(n474) );
  NOR2_X1 U532 ( .A1(n474), .A2(n548), .ZN(n468) );
  XNOR2_X1 U533 ( .A(n468), .B(KEYINPUT39), .ZN(n469) );
  XNOR2_X1 U534 ( .A(G29GAT), .B(n469), .ZN(G1328GAT) );
  NOR2_X1 U535 ( .A1(n474), .A2(n480), .ZN(n471) );
  XNOR2_X1 U536 ( .A(G36GAT), .B(KEYINPUT103), .ZN(n470) );
  XNOR2_X1 U537 ( .A(n471), .B(n470), .ZN(G1329GAT) );
  NOR2_X1 U538 ( .A1(n474), .A2(n490), .ZN(n472) );
  XOR2_X1 U539 ( .A(n472), .B(KEYINPUT40), .Z(n473) );
  XNOR2_X1 U540 ( .A(G43GAT), .B(n473), .ZN(G1330GAT) );
  NOR2_X1 U541 ( .A1(n493), .A2(n474), .ZN(n475) );
  XOR2_X1 U542 ( .A(G50GAT), .B(n475), .Z(G1331GAT) );
  NAND2_X1 U543 ( .A1(n477), .A2(n476), .ZN(n485) );
  NOR2_X1 U544 ( .A1(n548), .A2(n485), .ZN(n478) );
  XOR2_X1 U545 ( .A(G57GAT), .B(n478), .Z(n479) );
  XNOR2_X1 U546 ( .A(KEYINPUT42), .B(n479), .ZN(G1332GAT) );
  NOR2_X1 U547 ( .A1(n480), .A2(n485), .ZN(n481) );
  XOR2_X1 U548 ( .A(G64GAT), .B(n481), .Z(G1333GAT) );
  NOR2_X1 U549 ( .A1(n490), .A2(n485), .ZN(n483) );
  XNOR2_X1 U550 ( .A(KEYINPUT104), .B(KEYINPUT105), .ZN(n482) );
  XNOR2_X1 U551 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U552 ( .A(G71GAT), .B(n484), .ZN(G1334GAT) );
  NOR2_X1 U553 ( .A1(n493), .A2(n485), .ZN(n487) );
  XNOR2_X1 U554 ( .A(KEYINPUT43), .B(KEYINPUT106), .ZN(n486) );
  XNOR2_X1 U555 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U556 ( .A(G78GAT), .B(n488), .ZN(G1335GAT) );
  NOR2_X1 U557 ( .A1(n548), .A2(n492), .ZN(n489) );
  XOR2_X1 U558 ( .A(G85GAT), .B(n489), .Z(G1336GAT) );
  NOR2_X1 U559 ( .A1(n490), .A2(n492), .ZN(n491) );
  XOR2_X1 U560 ( .A(G99GAT), .B(n491), .Z(G1338GAT) );
  NOR2_X1 U561 ( .A1(n493), .A2(n492), .ZN(n495) );
  XNOR2_X1 U562 ( .A(KEYINPUT44), .B(KEYINPUT109), .ZN(n494) );
  XNOR2_X1 U563 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U564 ( .A(G106GAT), .B(n496), .ZN(G1339GAT) );
  XOR2_X1 U565 ( .A(KEYINPUT113), .B(KEYINPUT114), .Z(n514) );
  XNOR2_X1 U566 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n507) );
  NAND2_X1 U567 ( .A1(n530), .A2(n533), .ZN(n497) );
  XNOR2_X1 U568 ( .A(KEYINPUT110), .B(n578), .ZN(n559) );
  NAND2_X1 U569 ( .A1(n498), .A2(n559), .ZN(n499) );
  NOR2_X1 U570 ( .A1(n539), .A2(n499), .ZN(n500) );
  XNOR2_X1 U571 ( .A(n500), .B(KEYINPUT47), .ZN(n505) );
  NOR2_X1 U572 ( .A1(n583), .A2(n578), .ZN(n501) );
  XOR2_X1 U573 ( .A(KEYINPUT45), .B(n501), .Z(n502) );
  NOR2_X1 U574 ( .A1(n573), .A2(n502), .ZN(n503) );
  NAND2_X1 U575 ( .A1(n503), .A2(n570), .ZN(n504) );
  NAND2_X1 U576 ( .A1(n505), .A2(n504), .ZN(n506) );
  XNOR2_X1 U577 ( .A(n507), .B(n506), .ZN(n543) );
  NAND2_X1 U578 ( .A1(n543), .A2(n508), .ZN(n509) );
  XNOR2_X1 U579 ( .A(n509), .B(KEYINPUT111), .ZN(n528) );
  NAND2_X1 U580 ( .A1(n552), .A2(n528), .ZN(n510) );
  XNOR2_X1 U581 ( .A(KEYINPUT112), .B(n510), .ZN(n511) );
  NOR2_X1 U582 ( .A1(n512), .A2(n511), .ZN(n519) );
  NAND2_X1 U583 ( .A1(n519), .A2(n530), .ZN(n513) );
  XNOR2_X1 U584 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U585 ( .A(G113GAT), .B(n515), .ZN(G1340GAT) );
  XOR2_X1 U586 ( .A(KEYINPUT115), .B(KEYINPUT49), .Z(n517) );
  NAND2_X1 U587 ( .A1(n519), .A2(n533), .ZN(n516) );
  XNOR2_X1 U588 ( .A(n517), .B(n516), .ZN(n518) );
  XOR2_X1 U589 ( .A(G120GAT), .B(n518), .Z(G1341GAT) );
  INV_X1 U590 ( .A(n519), .ZN(n523) );
  NOR2_X1 U591 ( .A1(n559), .A2(n523), .ZN(n521) );
  XNOR2_X1 U592 ( .A(KEYINPUT50), .B(KEYINPUT116), .ZN(n520) );
  XNOR2_X1 U593 ( .A(n521), .B(n520), .ZN(n522) );
  XOR2_X1 U594 ( .A(G127GAT), .B(n522), .Z(G1342GAT) );
  NOR2_X1 U595 ( .A1(n523), .A2(n561), .ZN(n527) );
  XOR2_X1 U596 ( .A(KEYINPUT118), .B(KEYINPUT51), .Z(n525) );
  XNOR2_X1 U597 ( .A(G134GAT), .B(KEYINPUT117), .ZN(n524) );
  XNOR2_X1 U598 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U599 ( .A(n527), .B(n526), .ZN(G1343GAT) );
  XNOR2_X1 U600 ( .A(G141GAT), .B(KEYINPUT120), .ZN(n532) );
  NAND2_X1 U601 ( .A1(n568), .A2(n528), .ZN(n529) );
  XNOR2_X1 U602 ( .A(n529), .B(KEYINPUT119), .ZN(n540) );
  NAND2_X1 U603 ( .A1(n530), .A2(n540), .ZN(n531) );
  XNOR2_X1 U604 ( .A(n532), .B(n531), .ZN(G1344GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n535) );
  NAND2_X1 U606 ( .A1(n540), .A2(n533), .ZN(n534) );
  XNOR2_X1 U607 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U608 ( .A(G148GAT), .B(n536), .ZN(G1345GAT) );
  NAND2_X1 U609 ( .A1(n537), .A2(n540), .ZN(n538) );
  XNOR2_X1 U610 ( .A(G155GAT), .B(n538), .ZN(G1346GAT) );
  XOR2_X1 U611 ( .A(G162GAT), .B(KEYINPUT121), .Z(n542) );
  NAND2_X1 U612 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U613 ( .A(n542), .B(n541), .ZN(G1347GAT) );
  NAND2_X1 U614 ( .A1(n544), .A2(n543), .ZN(n546) );
  XOR2_X1 U615 ( .A(KEYINPUT122), .B(KEYINPUT54), .Z(n545) );
  NAND2_X1 U616 ( .A1(n548), .A2(n547), .ZN(n549) );
  NAND2_X1 U617 ( .A1(n550), .A2(n569), .ZN(n551) );
  XNOR2_X1 U618 ( .A(KEYINPUT55), .B(n551), .ZN(n553) );
  NAND2_X1 U619 ( .A1(n553), .A2(n552), .ZN(n562) );
  NOR2_X1 U620 ( .A1(n570), .A2(n562), .ZN(n554) );
  XOR2_X1 U621 ( .A(G169GAT), .B(n554), .Z(G1348GAT) );
  NOR2_X1 U622 ( .A1(n555), .A2(n562), .ZN(n557) );
  XNOR2_X1 U623 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U625 ( .A(G176GAT), .B(n558), .ZN(G1349GAT) );
  NOR2_X1 U626 ( .A1(n559), .A2(n562), .ZN(n560) );
  XOR2_X1 U627 ( .A(G183GAT), .B(n560), .Z(G1350GAT) );
  NOR2_X1 U628 ( .A1(n562), .A2(n561), .ZN(n564) );
  XNOR2_X1 U629 ( .A(KEYINPUT123), .B(KEYINPUT58), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n564), .B(n563), .ZN(n565) );
  XNOR2_X1 U631 ( .A(G190GAT), .B(n565), .ZN(G1351GAT) );
  XOR2_X1 U632 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n567) );
  XNOR2_X1 U633 ( .A(G197GAT), .B(KEYINPUT124), .ZN(n566) );
  XNOR2_X1 U634 ( .A(n567), .B(n566), .ZN(n572) );
  NAND2_X1 U635 ( .A1(n569), .A2(n568), .ZN(n582) );
  NOR2_X1 U636 ( .A1(n570), .A2(n582), .ZN(n571) );
  XOR2_X1 U637 ( .A(n572), .B(n571), .Z(G1352GAT) );
  XOR2_X1 U638 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n576) );
  INV_X1 U639 ( .A(n582), .ZN(n574) );
  NAND2_X1 U640 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(n577) );
  XOR2_X1 U642 ( .A(G204GAT), .B(n577), .Z(G1353GAT) );
  NOR2_X1 U643 ( .A1(n578), .A2(n582), .ZN(n579) );
  XOR2_X1 U644 ( .A(G211GAT), .B(n579), .Z(G1354GAT) );
  XOR2_X1 U645 ( .A(KEYINPUT126), .B(KEYINPUT62), .Z(n581) );
  XNOR2_X1 U646 ( .A(G218GAT), .B(KEYINPUT127), .ZN(n580) );
  XNOR2_X1 U647 ( .A(n581), .B(n580), .ZN(n585) );
  NOR2_X1 U648 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U649 ( .A(n585), .B(n584), .Z(G1355GAT) );
endmodule

