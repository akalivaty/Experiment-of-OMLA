//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 0 0 0 0 0 1 0 0 0 0 1 1 1 1 0 0 1 1 1 1 0 1 1 0 1 1 1 1 1 0 1 1 0 0 1 1 0 0 0 0 1 0 0 0 1 0 0 0 0 0 0 1 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:43 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n666, new_n667, new_n668,
    new_n669, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n681, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n721, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  XNOR2_X1  g001(.A(new_n187), .B(KEYINPUT72), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT30), .ZN(new_n190));
  XNOR2_X1  g004(.A(G143), .B(G146), .ZN(new_n191));
  NAND2_X1  g005(.A1(KEYINPUT0), .A2(G128), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  XOR2_X1   g007(.A(KEYINPUT0), .B(G128), .Z(new_n194));
  OAI21_X1  g008(.A(new_n193), .B1(new_n191), .B2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G137), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n196), .A2(G134), .ZN(new_n197));
  INV_X1    g011(.A(G134), .ZN(new_n198));
  OAI21_X1  g012(.A(KEYINPUT11), .B1(new_n198), .B2(G137), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT11), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n200), .A2(new_n196), .A3(G134), .ZN(new_n201));
  AOI211_X1 g015(.A(G131), .B(new_n197), .C1(new_n199), .C2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G131), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n199), .A2(new_n201), .ZN(new_n204));
  INV_X1    g018(.A(new_n197), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n203), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n195), .B1(new_n202), .B2(new_n206), .ZN(new_n207));
  OAI21_X1  g021(.A(KEYINPUT64), .B1(new_n196), .B2(G134), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT64), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n209), .A2(new_n198), .A3(G137), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n196), .A2(G134), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n208), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G131), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n200), .B1(G134), .B2(new_n196), .ZN(new_n214));
  NOR3_X1   g028(.A1(new_n198), .A2(KEYINPUT11), .A3(G137), .ZN(new_n215));
  OAI211_X1 g029(.A(new_n203), .B(new_n205), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n213), .A2(new_n216), .A3(KEYINPUT65), .ZN(new_n217));
  INV_X1    g031(.A(G146), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G143), .ZN(new_n219));
  INV_X1    g033(.A(G143), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G146), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT1), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n219), .A2(new_n221), .A3(new_n222), .A4(G128), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n218), .A2(G143), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(KEYINPUT1), .ZN(new_n225));
  OAI211_X1 g039(.A(new_n223), .B(new_n225), .C1(G128), .C2(new_n191), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n217), .A2(new_n226), .ZN(new_n227));
  AOI21_X1  g041(.A(KEYINPUT65), .B1(new_n213), .B2(new_n216), .ZN(new_n228));
  OAI211_X1 g042(.A(new_n190), .B(new_n207), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n226), .A2(new_n216), .A3(new_n213), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n207), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(KEYINPUT30), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n229), .A2(new_n232), .ZN(new_n233));
  XNOR2_X1  g047(.A(G116), .B(G119), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  OR2_X1    g049(.A1(KEYINPUT2), .A2(G113), .ZN(new_n236));
  AND3_X1   g050(.A1(KEYINPUT66), .A2(KEYINPUT2), .A3(G113), .ZN(new_n237));
  AOI21_X1  g051(.A(KEYINPUT66), .B1(KEYINPUT2), .B2(G113), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n236), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n235), .A2(new_n239), .ZN(new_n240));
  OAI211_X1 g054(.A(new_n234), .B(new_n236), .C1(new_n238), .C2(new_n237), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n233), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(G237), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(KEYINPUT67), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT67), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G237), .ZN(new_n247));
  OR2_X1    g061(.A1(KEYINPUT68), .A2(G953), .ZN(new_n248));
  NAND2_X1  g062(.A1(KEYINPUT68), .A2(G953), .ZN(new_n249));
  AOI22_X1  g063(.A1(new_n245), .A2(new_n247), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(G210), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G101), .ZN(new_n252));
  INV_X1    g066(.A(G101), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n250), .A2(new_n253), .A3(G210), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  XNOR2_X1  g069(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(new_n242), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n207), .A2(new_n259), .A3(new_n230), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n252), .A2(new_n254), .A3(new_n256), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n258), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n243), .A2(KEYINPUT69), .A3(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT69), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n259), .B1(new_n229), .B2(new_n232), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n265), .B1(new_n266), .B2(new_n262), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n264), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT31), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n243), .A2(new_n269), .A3(new_n263), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT70), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND4_X1  g086(.A1(new_n243), .A2(KEYINPUT70), .A3(new_n269), .A4(new_n263), .ZN(new_n273));
  AOI22_X1  g087(.A1(KEYINPUT31), .A2(new_n268), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n260), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(KEYINPUT28), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT28), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n260), .A2(new_n277), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n207), .B1(new_n227), .B2(new_n228), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(new_n242), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n276), .A2(new_n278), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n258), .A2(new_n261), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  AOI21_X1  g097(.A(KEYINPUT71), .B1(new_n274), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n272), .A2(new_n273), .ZN(new_n285));
  AOI21_X1  g099(.A(KEYINPUT69), .B1(new_n243), .B2(new_n263), .ZN(new_n286));
  NOR3_X1   g100(.A1(new_n266), .A2(new_n265), .A3(new_n262), .ZN(new_n287));
  OAI21_X1  g101(.A(KEYINPUT31), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NAND4_X1  g102(.A1(new_n285), .A2(new_n288), .A3(KEYINPUT71), .A4(new_n283), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n189), .B1(new_n284), .B2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT32), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n266), .A2(new_n275), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(new_n282), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT29), .ZN(new_n297));
  OAI211_X1 g111(.A(new_n296), .B(new_n297), .C1(new_n282), .C2(new_n281), .ZN(new_n298));
  OR2_X1    g112(.A1(new_n298), .A2(KEYINPUT73), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(KEYINPUT73), .ZN(new_n300));
  XNOR2_X1  g114(.A(new_n231), .B(new_n259), .ZN(new_n301));
  OAI211_X1 g115(.A(KEYINPUT74), .B(new_n278), .C1(new_n301), .C2(new_n277), .ZN(new_n302));
  OR2_X1    g116(.A1(new_n278), .A2(KEYINPUT74), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n297), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(new_n282), .ZN(new_n305));
  AOI21_X1  g119(.A(G902), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n299), .A2(new_n300), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(G472), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n285), .A2(new_n283), .A3(new_n288), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT71), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n188), .B1(new_n311), .B2(new_n289), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(KEYINPUT32), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n293), .A2(new_n308), .A3(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(G217), .ZN(new_n315));
  INV_X1    g129(.A(G902), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n315), .B1(G234), .B2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT16), .ZN(new_n318));
  INV_X1    g132(.A(G140), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n318), .A2(new_n319), .A3(G125), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(G125), .ZN(new_n321));
  INV_X1    g135(.A(G125), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(G140), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n320), .B1(new_n324), .B2(new_n318), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(new_n218), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT76), .ZN(new_n327));
  OAI211_X1 g141(.A(G146), .B(new_n320), .C1(new_n324), .C2(new_n318), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n326), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(G119), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n330), .A2(G128), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(KEYINPUT23), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT23), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n333), .B1(new_n330), .B2(G128), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n332), .B1(new_n331), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(KEYINPUT75), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT75), .ZN(new_n337));
  OAI211_X1 g151(.A(new_n332), .B(new_n337), .C1(new_n331), .C2(new_n334), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n336), .A2(G110), .A3(new_n338), .ZN(new_n339));
  XOR2_X1   g153(.A(KEYINPUT24), .B(G110), .Z(new_n340));
  XNOR2_X1  g154(.A(G119), .B(G128), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n325), .A2(KEYINPUT76), .A3(new_n218), .ZN(new_n343));
  NAND4_X1  g157(.A1(new_n329), .A2(new_n339), .A3(new_n342), .A4(new_n343), .ZN(new_n344));
  OAI22_X1  g158(.A1(new_n335), .A2(G110), .B1(new_n341), .B2(new_n340), .ZN(new_n345));
  OAI211_X1 g159(.A(new_n345), .B(new_n328), .C1(G146), .C2(new_n324), .ZN(new_n346));
  XNOR2_X1  g160(.A(KEYINPUT68), .B(G953), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n347), .A2(G221), .A3(G234), .ZN(new_n348));
  XNOR2_X1  g162(.A(KEYINPUT22), .B(G137), .ZN(new_n349));
  XNOR2_X1  g163(.A(new_n348), .B(new_n349), .ZN(new_n350));
  AND3_X1   g164(.A1(new_n344), .A2(new_n346), .A3(new_n350), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n350), .B1(new_n344), .B2(new_n346), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(KEYINPUT25), .B1(new_n353), .B2(new_n316), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT25), .ZN(new_n355));
  NOR4_X1   g169(.A1(new_n351), .A2(new_n352), .A3(new_n355), .A4(G902), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n317), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(new_n353), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n317), .A2(G902), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n357), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT81), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n363), .B1(new_n226), .B2(G125), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n219), .A2(new_n221), .ZN(new_n365));
  INV_X1    g179(.A(G128), .ZN(new_n366));
  AOI22_X1  g180(.A1(new_n365), .A2(new_n366), .B1(KEYINPUT1), .B2(new_n224), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n367), .A2(KEYINPUT81), .A3(new_n322), .A4(new_n223), .ZN(new_n368));
  OAI211_X1 g182(.A(new_n193), .B(G125), .C1(new_n191), .C2(new_n194), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n364), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(G953), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(G224), .ZN(new_n372));
  XOR2_X1   g186(.A(new_n372), .B(KEYINPUT82), .Z(new_n373));
  XNOR2_X1  g187(.A(new_n370), .B(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(G104), .ZN(new_n375));
  OAI21_X1  g189(.A(KEYINPUT3), .B1(new_n375), .B2(G107), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT3), .ZN(new_n377));
  INV_X1    g191(.A(G107), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n377), .A2(new_n378), .A3(G104), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n375), .A2(G107), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n376), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(G101), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n376), .A2(new_n379), .A3(new_n253), .A4(new_n380), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n382), .A2(KEYINPUT4), .A3(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT4), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n381), .A2(new_n385), .A3(G101), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n384), .A2(new_n242), .A3(new_n386), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n375), .A2(G107), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n378), .A2(G104), .ZN(new_n389));
  OAI21_X1  g203(.A(G101), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  AND2_X1   g204(.A1(new_n383), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n234), .A2(KEYINPUT5), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT5), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n393), .A2(new_n330), .A3(G116), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT80), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n393), .A2(new_n330), .A3(KEYINPUT80), .A4(G116), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n392), .A2(G113), .A3(new_n396), .A4(new_n397), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n391), .A2(new_n398), .A3(new_n241), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n387), .A2(new_n399), .ZN(new_n400));
  XOR2_X1   g214(.A(G110), .B(G122), .Z(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(new_n401), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n387), .A2(new_n403), .A3(new_n399), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n402), .A2(KEYINPUT6), .A3(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT6), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n400), .A2(new_n406), .A3(new_n401), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n374), .A2(new_n405), .A3(new_n407), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n391), .A2(new_n398), .A3(KEYINPUT83), .A4(new_n241), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n401), .A2(KEYINPUT8), .ZN(new_n410));
  AND2_X1   g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  OR2_X1    g225(.A1(new_n401), .A2(KEYINPUT8), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n391), .B1(new_n241), .B2(new_n398), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT83), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n399), .A2(new_n414), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n411), .B(new_n412), .C1(new_n413), .C2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n372), .A2(KEYINPUT7), .ZN(new_n417));
  OR2_X1    g231(.A1(new_n370), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n370), .A2(new_n417), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n416), .A2(new_n418), .A3(new_n404), .A4(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n408), .A2(new_n420), .A3(new_n316), .ZN(new_n421));
  OAI21_X1  g235(.A(G210), .B1(G237), .B2(G902), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT84), .ZN(new_n425));
  NAND4_X1  g239(.A1(new_n408), .A2(new_n420), .A3(new_n316), .A4(new_n422), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n424), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(G234), .A2(G237), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n428), .A2(G952), .A3(new_n371), .ZN(new_n429));
  XNOR2_X1  g243(.A(new_n429), .B(KEYINPUT90), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(new_n347), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n432), .A2(G902), .A3(new_n428), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  XNOR2_X1  g248(.A(KEYINPUT21), .B(G898), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n435), .B(KEYINPUT91), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n431), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  OAI21_X1  g251(.A(G214), .B1(G237), .B2(G902), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n421), .A2(KEYINPUT84), .A3(new_n423), .ZN(new_n441));
  AND3_X1   g255(.A1(new_n427), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(G221), .ZN(new_n443));
  XOR2_X1   g257(.A(KEYINPUT9), .B(G234), .Z(new_n444));
  AOI21_X1  g258(.A(new_n443), .B1(new_n444), .B2(new_n316), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n347), .A2(G227), .ZN(new_n446));
  XNOR2_X1  g260(.A(G110), .B(G140), .ZN(new_n447));
  XNOR2_X1  g261(.A(new_n446), .B(new_n447), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n202), .A2(new_n206), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n384), .A2(new_n195), .A3(new_n386), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n391), .A2(KEYINPUT10), .A3(new_n226), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n223), .A2(KEYINPUT77), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT77), .ZN(new_n455));
  NAND4_X1  g269(.A1(new_n191), .A2(new_n455), .A3(new_n222), .A4(G128), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n367), .A2(new_n454), .A3(new_n456), .ZN(new_n457));
  AOI21_X1  g271(.A(KEYINPUT10), .B1(new_n457), .B2(new_n391), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n450), .B1(new_n453), .B2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(new_n458), .ZN(new_n460));
  NAND4_X1  g274(.A1(new_n460), .A2(new_n449), .A3(new_n451), .A4(new_n452), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n448), .B1(new_n459), .B2(new_n461), .ZN(new_n462));
  OR2_X1    g276(.A1(new_n462), .A2(KEYINPUT79), .ZN(new_n463));
  AND2_X1   g277(.A1(new_n461), .A2(new_n448), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n457), .A2(new_n391), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n465), .B1(new_n226), .B2(new_n391), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT12), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT78), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n467), .B1(new_n449), .B2(new_n468), .ZN(new_n469));
  AND3_X1   g283(.A1(new_n466), .A2(new_n450), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n469), .B1(new_n466), .B2(new_n450), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n464), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n462), .A2(KEYINPUT79), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n463), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(G469), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n474), .A2(new_n475), .A3(new_n316), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n461), .B1(new_n470), .B2(new_n471), .ZN(new_n477));
  INV_X1    g291(.A(new_n448), .ZN(new_n478));
  AOI22_X1  g292(.A1(new_n477), .A2(new_n478), .B1(new_n464), .B2(new_n459), .ZN(new_n479));
  OAI21_X1  g293(.A(G469), .B1(new_n479), .B2(G902), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n445), .B1(new_n476), .B2(new_n480), .ZN(new_n481));
  NOR2_X1   g295(.A1(G475), .A2(G902), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT85), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n483), .A2(G143), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n245), .A2(new_n247), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n485), .A2(new_n347), .A3(G214), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n220), .A2(KEYINPUT85), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n484), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(new_n484), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n490), .B1(new_n250), .B2(G214), .ZN(new_n491));
  OAI211_X1 g305(.A(KEYINPUT18), .B(G131), .C1(new_n489), .C2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(KEYINPUT86), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n486), .A2(new_n484), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n487), .B1(new_n250), .B2(G214), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n494), .B1(new_n495), .B2(new_n484), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT86), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n496), .A2(new_n497), .A3(KEYINPUT18), .A4(G131), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n493), .A2(new_n498), .ZN(new_n499));
  XNOR2_X1  g313(.A(new_n324), .B(new_n218), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  OAI211_X1 g315(.A(new_n494), .B(new_n203), .C1(new_n495), .C2(new_n484), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT18), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n494), .B(new_n503), .C1(new_n495), .C2(new_n484), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n499), .A2(new_n501), .A3(new_n506), .ZN(new_n507));
  XNOR2_X1  g321(.A(G113), .B(G122), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n508), .B(new_n375), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT87), .ZN(new_n510));
  OAI21_X1  g324(.A(G131), .B1(new_n489), .B2(new_n491), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT17), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n511), .A2(new_n502), .A3(new_n512), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n329), .A2(new_n343), .ZN(new_n515));
  NAND4_X1  g329(.A1(new_n496), .A2(KEYINPUT87), .A3(KEYINPUT17), .A4(G131), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n513), .A2(new_n514), .A3(new_n515), .A4(new_n516), .ZN(new_n517));
  AND3_X1   g331(.A1(new_n507), .A2(new_n509), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n511), .A2(new_n502), .ZN(new_n519));
  XOR2_X1   g333(.A(new_n324), .B(KEYINPUT19), .Z(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(new_n218), .ZN(new_n521));
  AND3_X1   g335(.A1(new_n519), .A2(new_n328), .A3(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n509), .B1(new_n523), .B2(new_n507), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n482), .B1(new_n518), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(KEYINPUT20), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n507), .A2(new_n509), .A3(new_n517), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n505), .B1(new_n493), .B2(new_n498), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n522), .B1(new_n528), .B2(new_n501), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n527), .B1(new_n529), .B2(new_n509), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT20), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n530), .A2(new_n531), .A3(new_n482), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n509), .B1(new_n507), .B2(new_n517), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n316), .B1(new_n518), .B2(new_n533), .ZN(new_n534));
  AOI22_X1  g348(.A1(new_n526), .A2(new_n532), .B1(G475), .B2(new_n534), .ZN(new_n535));
  XNOR2_X1  g349(.A(G128), .B(G143), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(KEYINPUT13), .ZN(new_n537));
  NOR3_X1   g351(.A1(new_n366), .A2(KEYINPUT13), .A3(G143), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n538), .A2(new_n198), .ZN(new_n539));
  AOI22_X1  g353(.A1(new_n537), .A2(new_n539), .B1(new_n198), .B2(new_n536), .ZN(new_n540));
  INV_X1    g354(.A(G122), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(G116), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n542), .B(KEYINPUT88), .ZN(new_n543));
  OR2_X1    g357(.A1(new_n541), .A2(G116), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n545), .A2(G107), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n378), .B1(new_n543), .B2(new_n544), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n540), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n543), .A2(KEYINPUT14), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n545), .A2(new_n549), .A3(G107), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n536), .B(new_n198), .ZN(new_n551));
  OAI211_X1 g365(.A(new_n543), .B(new_n544), .C1(KEYINPUT14), .C2(new_n378), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n548), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n444), .A2(G217), .A3(new_n371), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(new_n555), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n548), .A2(new_n553), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT89), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n559), .A2(new_n560), .A3(new_n316), .ZN(new_n561));
  INV_X1    g375(.A(G478), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n562), .A2(KEYINPUT15), .ZN(new_n563));
  XOR2_X1   g377(.A(new_n561), .B(new_n563), .Z(new_n564));
  NAND4_X1  g378(.A1(new_n442), .A2(new_n481), .A3(new_n535), .A4(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT92), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n534), .A2(G475), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n531), .B1(new_n530), .B2(new_n482), .ZN(new_n569));
  INV_X1    g383(.A(new_n482), .ZN(new_n570));
  INV_X1    g384(.A(new_n509), .ZN(new_n571));
  AOI211_X1 g385(.A(new_n500), .B(new_n505), .C1(new_n493), .C2(new_n498), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n571), .B1(new_n572), .B2(new_n522), .ZN(new_n573));
  AOI211_X1 g387(.A(KEYINPUT20), .B(new_n570), .C1(new_n573), .C2(new_n527), .ZN(new_n574));
  OAI211_X1 g388(.A(new_n564), .B(new_n568), .C1(new_n569), .C2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  NAND4_X1  g390(.A1(new_n576), .A2(KEYINPUT92), .A3(new_n481), .A4(new_n442), .ZN(new_n577));
  NAND4_X1  g391(.A1(new_n314), .A2(new_n362), .A3(new_n567), .A4(new_n577), .ZN(new_n578));
  XNOR2_X1  g392(.A(KEYINPUT93), .B(G101), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n578), .B(new_n579), .ZN(G3));
  AOI21_X1  g394(.A(G902), .B1(new_n311), .B2(new_n289), .ZN(new_n581));
  INV_X1    g395(.A(G472), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n291), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n481), .ZN(new_n584));
  NOR3_X1   g398(.A1(new_n583), .A2(new_n361), .A3(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n426), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT94), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n439), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n424), .A2(KEYINPUT94), .A3(new_n426), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  OAI21_X1  g405(.A(KEYINPUT33), .B1(new_n557), .B2(KEYINPUT95), .ZN(new_n592));
  AND3_X1   g406(.A1(new_n548), .A2(new_n553), .A3(new_n557), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n557), .B1(new_n548), .B2(new_n553), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n592), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n592), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n556), .A2(new_n558), .A3(new_n596), .ZN(new_n597));
  AND2_X1   g411(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n598), .A2(KEYINPUT96), .A3(G478), .A4(new_n316), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n559), .A2(new_n316), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(new_n562), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n595), .A2(new_n597), .A3(G478), .A4(new_n316), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT96), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n599), .A2(new_n601), .A3(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  OAI21_X1  g420(.A(KEYINPUT97), .B1(new_n535), .B2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n437), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n568), .B1(new_n574), .B2(new_n569), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT97), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n609), .A2(new_n610), .A3(new_n605), .ZN(new_n611));
  AND3_X1   g425(.A1(new_n607), .A2(new_n608), .A3(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n585), .A2(new_n591), .A3(new_n612), .ZN(new_n613));
  XOR2_X1   g427(.A(KEYINPUT34), .B(G104), .Z(new_n614));
  XNOR2_X1  g428(.A(new_n613), .B(new_n614), .ZN(G6));
  XNOR2_X1  g429(.A(new_n561), .B(new_n563), .ZN(new_n616));
  OAI211_X1 g430(.A(new_n616), .B(new_n568), .C1(new_n574), .C2(new_n569), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n617), .A2(new_n437), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n585), .A2(new_n591), .A3(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(KEYINPUT35), .B(G107), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n620), .B(KEYINPUT98), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n619), .B(new_n621), .ZN(G9));
  NAND2_X1  g436(.A1(new_n311), .A2(new_n289), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(new_n316), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n312), .B1(new_n624), .B2(G472), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n344), .A2(new_n346), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT36), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n350), .A2(new_n627), .ZN(new_n628));
  XOR2_X1   g442(.A(new_n626), .B(new_n628), .Z(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(new_n359), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n357), .A2(new_n630), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n567), .A2(new_n625), .A3(new_n577), .A4(new_n631), .ZN(new_n632));
  XOR2_X1   g446(.A(KEYINPUT37), .B(G110), .Z(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G12));
  AOI21_X1  g448(.A(KEYINPUT32), .B1(new_n623), .B2(new_n189), .ZN(new_n635));
  AOI211_X1 g449(.A(new_n292), .B(new_n188), .C1(new_n311), .C2(new_n289), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n584), .B1(new_n637), .B2(new_n308), .ZN(new_n638));
  AND3_X1   g452(.A1(new_n588), .A2(new_n589), .A3(new_n631), .ZN(new_n639));
  INV_X1    g453(.A(G900), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n431), .B1(new_n434), .B2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n639), .A2(new_n616), .A3(new_n535), .A4(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n638), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(KEYINPUT99), .B(G128), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G30));
  NOR2_X1   g461(.A1(new_n535), .A2(new_n564), .ZN(new_n648));
  XOR2_X1   g462(.A(new_n641), .B(KEYINPUT39), .Z(new_n649));
  NAND2_X1  g463(.A1(new_n481), .A2(new_n649), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n648), .B1(new_n650), .B2(KEYINPUT40), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n427), .A2(new_n441), .ZN(new_n652));
  XOR2_X1   g466(.A(KEYINPUT100), .B(KEYINPUT101), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(KEYINPUT38), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n652), .B(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n651), .A2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n631), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n268), .B1(new_n305), .B2(new_n301), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n582), .B1(new_n658), .B2(new_n316), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(KEYINPUT102), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n293), .A2(new_n313), .A3(new_n660), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n439), .B1(new_n650), .B2(KEYINPUT40), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n656), .A2(new_n657), .A3(new_n661), .A4(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(KEYINPUT103), .B(G143), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G45));
  NAND4_X1  g479(.A1(new_n639), .A2(new_n609), .A3(new_n605), .A4(new_n642), .ZN(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n638), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(KEYINPUT104), .B(G146), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n668), .B(new_n669), .ZN(G48));
  NAND2_X1  g484(.A1(new_n474), .A2(new_n316), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT105), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n671), .A2(new_n672), .A3(G469), .ZN(new_n673));
  INV_X1    g487(.A(new_n445), .ZN(new_n674));
  OAI211_X1 g488(.A(new_n474), .B(new_n316), .C1(KEYINPUT105), .C2(new_n475), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n673), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n676), .A2(new_n590), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n314), .A2(new_n612), .A3(new_n362), .A4(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(KEYINPUT41), .B(G113), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n678), .B(new_n679), .ZN(G15));
  NAND4_X1  g494(.A1(new_n314), .A2(new_n362), .A3(new_n618), .A4(new_n677), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G116), .ZN(G18));
  NOR2_X1   g496(.A1(new_n676), .A2(new_n437), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n314), .A2(new_n576), .A3(new_n639), .A4(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G119), .ZN(G21));
  INV_X1    g499(.A(KEYINPUT106), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n624), .A2(new_n686), .A3(G472), .ZN(new_n687));
  OAI21_X1  g501(.A(KEYINPUT106), .B1(new_n581), .B2(new_n582), .ZN(new_n688));
  INV_X1    g502(.A(new_n274), .ZN(new_n689));
  AND3_X1   g503(.A1(new_n302), .A2(new_n282), .A3(new_n303), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n189), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n687), .A2(new_n688), .A3(new_n362), .A4(new_n691), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n683), .A2(new_n591), .A3(new_n648), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(new_n541), .ZN(G24));
  NAND4_X1  g509(.A1(new_n687), .A2(new_n688), .A3(new_n631), .A4(new_n691), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n609), .A2(new_n605), .A3(new_n642), .ZN(new_n697));
  NOR3_X1   g511(.A1(new_n697), .A2(new_n676), .A3(new_n590), .ZN(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(new_n322), .ZN(G27));
  INV_X1    g515(.A(KEYINPUT42), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT108), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n623), .A2(new_n703), .A3(KEYINPUT32), .A4(new_n189), .ZN(new_n704));
  AND2_X1   g518(.A1(new_n308), .A2(new_n704), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n313), .B1(new_n635), .B2(KEYINPUT108), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n361), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n652), .A2(new_n438), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT107), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n652), .A2(KEYINPUT107), .A3(new_n438), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NOR3_X1   g526(.A1(new_n712), .A2(new_n584), .A3(new_n697), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n702), .B1(new_n707), .B2(new_n713), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n314), .A2(new_n702), .A3(new_n362), .A4(new_n481), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n712), .A2(new_n697), .ZN(new_n716));
  INV_X1    g530(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n714), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G131), .ZN(G33));
  NOR2_X1   g534(.A1(new_n617), .A2(new_n641), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n314), .A2(new_n362), .A3(new_n481), .A4(new_n721), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n722), .A2(new_n712), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(new_n198), .ZN(G36));
  OR2_X1    g538(.A1(new_n479), .A2(KEYINPUT45), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n479), .A2(KEYINPUT45), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n725), .A2(G469), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(G469), .A2(G902), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n727), .A2(KEYINPUT46), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(new_n476), .ZN(new_n730));
  AOI21_X1  g544(.A(KEYINPUT46), .B1(new_n727), .B2(new_n728), .ZN(new_n731));
  OAI211_X1 g545(.A(new_n674), .B(new_n649), .C1(new_n730), .C2(new_n731), .ZN(new_n732));
  XOR2_X1   g546(.A(new_n732), .B(KEYINPUT109), .Z(new_n733));
  OAI211_X1 g547(.A(new_n605), .B(new_n568), .C1(new_n569), .C2(new_n574), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(KEYINPUT43), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT43), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n535), .A2(new_n736), .A3(new_n605), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n583), .A2(new_n631), .A3(new_n735), .A4(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT44), .ZN(new_n739));
  OR3_X1    g553(.A1(new_n738), .A2(KEYINPUT110), .A3(new_n739), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n712), .B1(new_n738), .B2(new_n739), .ZN(new_n741));
  OAI21_X1  g555(.A(KEYINPUT110), .B1(new_n738), .B2(new_n739), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n733), .A2(new_n740), .A3(new_n741), .A4(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G137), .ZN(G39));
  OAI21_X1  g558(.A(new_n674), .B1(new_n730), .B2(new_n731), .ZN(new_n745));
  OR2_X1    g559(.A1(new_n745), .A2(KEYINPUT47), .ZN(new_n746));
  INV_X1    g560(.A(new_n746), .ZN(new_n747));
  AND2_X1   g561(.A1(new_n745), .A2(KEYINPUT47), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n314), .A2(new_n362), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n749), .A2(new_n716), .A3(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G140), .ZN(G42));
  NAND2_X1  g566(.A1(new_n673), .A2(new_n675), .ZN(new_n753));
  OR2_X1    g567(.A1(new_n753), .A2(KEYINPUT49), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(KEYINPUT49), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n754), .A2(new_n655), .A3(new_n362), .A4(new_n755), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n535), .A2(new_n674), .A3(new_n438), .A4(new_n605), .ZN(new_n757));
  OR3_X1    g571(.A1(new_n756), .A2(new_n661), .A3(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n609), .A2(new_n605), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n427), .A2(new_n440), .A3(new_n441), .ZN(new_n760));
  OAI21_X1  g574(.A(KEYINPUT111), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT111), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n442), .A2(new_n762), .A3(new_n609), .A4(new_n605), .ZN(new_n763));
  OAI21_X1  g577(.A(KEYINPUT112), .B1(new_n617), .B2(new_n760), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT112), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n442), .A2(new_n765), .A3(new_n535), .A4(new_n616), .ZN(new_n766));
  AND4_X1   g580(.A1(new_n761), .A2(new_n763), .A3(new_n764), .A4(new_n766), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n625), .A2(new_n362), .A3(new_n481), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n632), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n769), .A2(new_n694), .ZN(new_n770));
  AND3_X1   g584(.A1(new_n678), .A2(new_n578), .A3(new_n681), .ZN(new_n771));
  OR2_X1    g585(.A1(new_n722), .A2(new_n712), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n770), .A2(new_n771), .A3(new_n684), .A4(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n707), .A2(new_n713), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(KEYINPUT42), .ZN(new_n775));
  AOI21_X1  g589(.A(KEYINPUT107), .B1(new_n652), .B2(new_n438), .ZN(new_n776));
  AOI211_X1 g590(.A(new_n709), .B(new_n439), .C1(new_n427), .C2(new_n441), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n575), .A2(new_n641), .ZN(new_n779));
  AND4_X1   g593(.A1(new_n314), .A2(new_n778), .A3(new_n481), .A4(new_n779), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n687), .A2(new_n691), .A3(new_n688), .ZN(new_n781));
  INV_X1    g595(.A(new_n697), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n778), .A2(new_n481), .A3(new_n782), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n631), .B1(new_n780), .B2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(new_n718), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n775), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n773), .A2(new_n787), .ZN(new_n788));
  AOI221_X4 g602(.A(new_n584), .B1(new_n643), .B2(new_n666), .C1(new_n637), .C2(new_n308), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n789), .A2(new_n700), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n648), .A2(new_n591), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n791), .A2(new_n584), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n792), .A2(new_n661), .A3(new_n657), .A4(new_n642), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n790), .A2(KEYINPUT113), .A3(KEYINPUT52), .A4(new_n793), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n686), .B1(new_n624), .B2(G472), .ZN(new_n795));
  NOR3_X1   g609(.A1(new_n581), .A2(KEYINPUT106), .A3(new_n582), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n797), .A2(new_n631), .A3(new_n691), .A4(new_n698), .ZN(new_n798));
  OAI211_X1 g612(.A(new_n314), .B(new_n481), .C1(new_n644), .C2(new_n667), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n798), .A2(KEYINPUT52), .A3(new_n799), .A4(new_n793), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT113), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n798), .A2(new_n799), .A3(new_n793), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT52), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n794), .A2(new_n802), .A3(new_n805), .ZN(new_n806));
  AOI21_X1  g620(.A(KEYINPUT53), .B1(new_n788), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n805), .A2(new_n800), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n535), .A2(new_n590), .A3(new_n564), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n683), .A2(new_n809), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n797), .A2(new_n362), .A3(new_n810), .A4(new_n691), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n761), .A2(new_n763), .A3(new_n764), .A4(new_n766), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n585), .A2(new_n812), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n811), .A2(new_n632), .A3(new_n684), .A4(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n678), .A2(new_n578), .A3(new_n681), .ZN(new_n815));
  NOR3_X1   g629(.A1(new_n814), .A2(new_n723), .A3(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n713), .A2(new_n797), .A3(new_n691), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n314), .A2(new_n778), .A3(new_n481), .A4(new_n779), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n657), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n819), .A2(new_n714), .A3(new_n718), .ZN(new_n820));
  AND4_X1   g634(.A1(KEYINPUT53), .A2(new_n808), .A3(new_n816), .A4(new_n820), .ZN(new_n821));
  OAI21_X1  g635(.A(KEYINPUT54), .B1(new_n807), .B2(new_n821), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n712), .A2(new_n676), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n823), .A2(new_n362), .A3(new_n431), .ZN(new_n824));
  NOR4_X1   g638(.A1(new_n824), .A2(new_n609), .A3(new_n605), .A4(new_n661), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n735), .A2(new_n431), .A3(new_n737), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(KEYINPUT115), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT115), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n735), .A2(new_n828), .A3(new_n737), .A4(new_n431), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(new_n692), .ZN(new_n831));
  INV_X1    g645(.A(new_n676), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n655), .A2(new_n439), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n830), .A2(new_n831), .A3(new_n832), .A4(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT50), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n692), .B1(new_n829), .B2(new_n827), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n837), .A2(KEYINPUT50), .A3(new_n832), .A4(new_n833), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n825), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  OAI21_X1  g653(.A(KEYINPUT116), .B1(new_n753), .B2(new_n674), .ZN(new_n840));
  OR3_X1    g654(.A1(new_n753), .A2(KEYINPUT116), .A3(new_n674), .ZN(new_n841));
  OAI211_X1 g655(.A(new_n840), .B(new_n841), .C1(new_n747), .C2(new_n748), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n842), .A2(new_n778), .A3(new_n837), .ZN(new_n843));
  INV_X1    g657(.A(new_n696), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT117), .ZN(new_n845));
  AND3_X1   g659(.A1(new_n830), .A2(new_n845), .A3(new_n823), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n845), .B1(new_n830), .B2(new_n823), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n844), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n839), .A2(new_n843), .A3(new_n848), .ZN(new_n849));
  XNOR2_X1  g663(.A(KEYINPUT114), .B(KEYINPUT51), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n837), .A2(new_n677), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n753), .A2(new_n674), .ZN(new_n853));
  OAI211_X1 g667(.A(new_n778), .B(new_n837), .C1(new_n749), .C2(new_n853), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n839), .A2(KEYINPUT51), .A3(new_n848), .A4(new_n854), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n707), .B1(new_n846), .B2(new_n847), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(KEYINPUT48), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT48), .ZN(new_n858));
  OAI211_X1 g672(.A(new_n858), .B(new_n707), .C1(new_n846), .C2(new_n847), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n607), .A2(new_n611), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n824), .A2(new_n661), .ZN(new_n861));
  AOI22_X1  g675(.A1(new_n857), .A2(new_n859), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  AND4_X1   g676(.A1(new_n851), .A2(new_n852), .A3(new_n855), .A4(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n808), .A2(new_n816), .A3(new_n820), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT53), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n788), .A2(new_n806), .A3(KEYINPUT53), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT54), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n866), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n371), .A2(G952), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n870), .B(KEYINPUT118), .ZN(new_n871));
  AND4_X1   g685(.A1(new_n822), .A2(new_n863), .A3(new_n869), .A4(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(G952), .A2(G953), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n758), .B1(new_n872), .B2(new_n873), .ZN(G75));
  NAND2_X1  g688(.A1(new_n866), .A2(new_n867), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n875), .A2(G210), .A3(G902), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT56), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n405), .A2(new_n407), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n878), .B(new_n374), .ZN(new_n879));
  XOR2_X1   g693(.A(KEYINPUT119), .B(KEYINPUT55), .Z(new_n880));
  XNOR2_X1  g694(.A(new_n879), .B(new_n880), .ZN(new_n881));
  AND3_X1   g695(.A1(new_n876), .A2(new_n877), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n881), .B1(new_n876), .B2(new_n877), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n347), .A2(G952), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(G51));
  XOR2_X1   g699(.A(new_n728), .B(KEYINPUT57), .Z(new_n886));
  AND3_X1   g700(.A1(new_n866), .A2(new_n867), .A3(new_n868), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n868), .B1(new_n866), .B2(new_n867), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n886), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n474), .B(KEYINPUT120), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n316), .B1(new_n866), .B2(new_n867), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n892), .A2(G469), .A3(new_n725), .A4(new_n726), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n884), .B1(new_n891), .B2(new_n893), .ZN(G54));
  AND2_X1   g708(.A1(KEYINPUT58), .A2(G475), .ZN(new_n895));
  OR2_X1    g709(.A1(new_n895), .A2(KEYINPUT121), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n895), .A2(KEYINPUT121), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n892), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(new_n530), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(new_n884), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n892), .A2(new_n530), .A3(new_n896), .A4(new_n897), .ZN(new_n902));
  AND3_X1   g716(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(G60));
  NAND2_X1  g717(.A1(G478), .A2(G902), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n904), .B(KEYINPUT59), .Z(new_n905));
  AOI21_X1  g719(.A(new_n905), .B1(new_n822), .B2(new_n869), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n901), .B1(new_n906), .B2(new_n598), .ZN(new_n907));
  INV_X1    g721(.A(new_n905), .ZN(new_n908));
  OAI211_X1 g722(.A(new_n598), .B(new_n908), .C1(new_n887), .C2(new_n888), .ZN(new_n909));
  INV_X1    g723(.A(new_n909), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n907), .A2(new_n910), .ZN(G63));
  INV_X1    g725(.A(KEYINPUT61), .ZN(new_n912));
  NAND2_X1  g726(.A1(G217), .A2(G902), .ZN(new_n913));
  XOR2_X1   g727(.A(new_n913), .B(KEYINPUT60), .Z(new_n914));
  XOR2_X1   g728(.A(new_n629), .B(KEYINPUT122), .Z(new_n915));
  NAND3_X1  g729(.A1(new_n875), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n916), .A2(new_n901), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n353), .B1(new_n875), .B2(new_n914), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n912), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n875), .A2(new_n914), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(new_n358), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n921), .A2(KEYINPUT61), .A3(new_n901), .A4(new_n916), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n919), .A2(new_n922), .ZN(G66));
  INV_X1    g737(.A(G224), .ZN(new_n924));
  OAI21_X1  g738(.A(G953), .B1(new_n436), .B2(new_n924), .ZN(new_n925));
  OR2_X1    g739(.A1(new_n925), .A2(KEYINPUT123), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n814), .A2(new_n815), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n926), .B1(new_n927), .B2(new_n432), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n928), .B1(KEYINPUT123), .B2(new_n925), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n878), .B1(G898), .B2(new_n347), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n929), .B(new_n930), .Z(G69));
  XNOR2_X1  g745(.A(new_n233), .B(new_n520), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n790), .A2(new_n663), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT62), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n933), .B(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT124), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n361), .B1(new_n637), .B2(new_n308), .ZN(new_n937));
  INV_X1    g751(.A(new_n650), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n759), .A2(new_n617), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n937), .A2(new_n938), .A3(new_n778), .A4(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n936), .B1(new_n743), .B2(new_n940), .ZN(new_n941));
  AND3_X1   g755(.A1(new_n743), .A2(new_n936), .A3(new_n940), .ZN(new_n942));
  OAI211_X1 g756(.A(new_n935), .B(new_n751), .C1(new_n941), .C2(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n932), .B1(new_n943), .B2(new_n347), .ZN(new_n944));
  AND3_X1   g758(.A1(new_n751), .A2(new_n772), .A3(new_n790), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n740), .A2(new_n741), .A3(new_n742), .ZN(new_n946));
  INV_X1    g760(.A(new_n707), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n946), .B1(new_n791), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n948), .A2(new_n733), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n945), .A2(new_n949), .A3(new_n347), .A4(new_n719), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n432), .A2(G900), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n950), .A2(new_n932), .A3(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(G227), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n432), .B1(new_n954), .B2(new_n640), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n955), .B(KEYINPUT125), .Z(new_n956));
  INV_X1    g770(.A(new_n956), .ZN(new_n957));
  OR3_X1    g771(.A1(new_n944), .A2(new_n953), .A3(new_n957), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n957), .B1(new_n944), .B2(new_n953), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n958), .A2(new_n959), .ZN(G72));
  NAND2_X1  g774(.A1(G472), .A2(G902), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n961), .B(KEYINPUT63), .Z(new_n962));
  INV_X1    g776(.A(new_n927), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n962), .B1(new_n943), .B2(new_n963), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n964), .A2(new_n305), .A3(new_n295), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n945), .A2(new_n949), .A3(new_n719), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n962), .B1(new_n966), .B2(new_n963), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n294), .A2(new_n282), .ZN(new_n968));
  XOR2_X1   g782(.A(new_n968), .B(KEYINPUT126), .Z(new_n969));
  AOI21_X1  g783(.A(new_n884), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(new_n296), .ZN(new_n971));
  AOI22_X1  g785(.A1(new_n971), .A2(KEYINPUT127), .B1(new_n267), .B2(new_n264), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n972), .B1(KEYINPUT127), .B2(new_n971), .ZN(new_n973));
  OAI211_X1 g787(.A(new_n962), .B(new_n973), .C1(new_n807), .C2(new_n821), .ZN(new_n974));
  AND3_X1   g788(.A1(new_n965), .A2(new_n970), .A3(new_n974), .ZN(G57));
endmodule


