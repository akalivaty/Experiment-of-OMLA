//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 1 1 0 0 1 0 1 0 0 0 1 0 0 1 0 0 0 1 0 0 1 0 0 1 0 0 1 1 0 1 1 1 0 0 1 1 1 0 0 0 0 0 1 1 1 0 0 1 0 0 1 1 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:54 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n257, new_n258, new_n259, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1225,
    new_n1226, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1283, new_n1284, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291, new_n1292;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n201), .A2(G77), .A3(new_n203), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G250), .ZN(new_n206));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(G257), .ZN(new_n210));
  INV_X1    g0010(.A(G264), .ZN(new_n211));
  AOI211_X1 g0011(.A(new_n206), .B(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  OR2_X1    g0012(.A1(new_n212), .A2(KEYINPUT0), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n212), .A2(KEYINPUT0), .ZN(new_n214));
  AND2_X1   g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(G20), .ZN(new_n216));
  OR2_X1    g0016(.A1(new_n202), .A2(KEYINPUT65), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n202), .A2(KEYINPUT65), .ZN(new_n218));
  NAND3_X1  g0018(.A1(new_n217), .A2(G50), .A3(new_n218), .ZN(new_n219));
  OAI211_X1 g0019(.A(new_n213), .B(new_n214), .C1(new_n216), .C2(new_n219), .ZN(new_n220));
  XOR2_X1   g0020(.A(new_n220), .B(KEYINPUT66), .Z(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n222));
  XOR2_X1   g0022(.A(new_n222), .B(KEYINPUT67), .Z(new_n223));
  NAND2_X1  g0023(.A1(G77), .A2(G244), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G68), .A2(G238), .ZN(new_n225));
  NAND3_X1  g0025(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  OR2_X1    g0026(.A1(new_n226), .A2(KEYINPUT68), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G97), .A2(G257), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n226), .A2(KEYINPUT68), .ZN(new_n229));
  INV_X1    g0029(.A(G58), .ZN(new_n230));
  INV_X1    g0030(.A(G232), .ZN(new_n231));
  INV_X1    g0031(.A(G87), .ZN(new_n232));
  OAI22_X1  g0032(.A1(new_n230), .A2(new_n231), .B1(new_n232), .B2(new_n206), .ZN(new_n233));
  AOI21_X1  g0033(.A(new_n233), .B1(G107), .B2(G264), .ZN(new_n234));
  NAND4_X1  g0034(.A1(new_n227), .A2(new_n228), .A3(new_n229), .A4(new_n234), .ZN(new_n235));
  AND2_X1   g0035(.A1(new_n235), .A2(new_n207), .ZN(new_n236));
  INV_X1    g0036(.A(KEYINPUT1), .ZN(new_n237));
  NAND2_X1  g0037(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NOR2_X1   g0038(.A1(new_n236), .A2(new_n237), .ZN(new_n239));
  OAI21_X1  g0039(.A(new_n238), .B1(new_n239), .B2(KEYINPUT69), .ZN(new_n240));
  AOI211_X1 g0040(.A(new_n221), .B(new_n240), .C1(KEYINPUT69), .C2(new_n239), .ZN(G361));
  XNOR2_X1  g0041(.A(G238), .B(G244), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(new_n231), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(KEYINPUT2), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(G226), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G250), .B(G257), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(G264), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(G270), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G358));
  XNOR2_X1  g0049(.A(G87), .B(G97), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n250), .B(KEYINPUT70), .ZN(new_n251));
  INV_X1    g0051(.A(G107), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G116), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n253), .B(new_n254), .ZN(new_n255));
  XNOR2_X1  g0055(.A(G68), .B(G77), .ZN(new_n256));
  INV_X1    g0056(.A(G50), .ZN(new_n257));
  XNOR2_X1  g0057(.A(new_n256), .B(new_n257), .ZN(new_n258));
  XNOR2_X1  g0058(.A(new_n258), .B(new_n230), .ZN(new_n259));
  XNOR2_X1  g0059(.A(new_n255), .B(new_n259), .ZN(G351));
  XNOR2_X1  g0060(.A(KEYINPUT3), .B(G33), .ZN(new_n261));
  INV_X1    g0061(.A(G1698), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n261), .A2(G226), .A3(new_n262), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n261), .A2(G232), .A3(G1698), .ZN(new_n264));
  INV_X1    g0064(.A(G33), .ZN(new_n265));
  INV_X1    g0065(.A(G97), .ZN(new_n266));
  OAI211_X1 g0066(.A(new_n263), .B(new_n264), .C1(new_n265), .C2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(G33), .A2(G41), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n215), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n267), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G274), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n272), .B1(new_n215), .B2(new_n268), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT71), .ZN(new_n274));
  NOR2_X1   g0074(.A1(G41), .A2(G45), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n274), .B1(new_n275), .B2(G1), .ZN(new_n276));
  INV_X1    g0076(.A(G1), .ZN(new_n277));
  OAI211_X1 g0077(.A(new_n277), .B(KEYINPUT71), .C1(G41), .C2(G45), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n273), .A2(new_n276), .A3(new_n278), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n277), .B1(G41), .B2(G45), .ZN(new_n280));
  AND2_X1   g0080(.A1(new_n269), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(G238), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n271), .A2(new_n279), .A3(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT13), .ZN(new_n284));
  OR2_X1    g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n283), .A2(new_n284), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n285), .A2(G169), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(KEYINPUT14), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n284), .A2(KEYINPUT76), .ZN(new_n289));
  OR2_X1    g0089(.A1(new_n283), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n283), .A2(new_n289), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n290), .A2(G179), .A3(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT14), .ZN(new_n293));
  NAND4_X1  g0093(.A1(new_n285), .A2(new_n293), .A3(G169), .A4(new_n286), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n288), .A2(new_n292), .A3(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G20), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(G33), .ZN(new_n297));
  INV_X1    g0097(.A(G77), .ZN(new_n298));
  OAI22_X1  g0098(.A1(new_n297), .A2(new_n298), .B1(new_n296), .B2(G68), .ZN(new_n299));
  XNOR2_X1  g0099(.A(new_n299), .B(KEYINPUT77), .ZN(new_n300));
  NOR2_X1   g0100(.A1(G20), .A2(G33), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n300), .B1(new_n257), .B2(new_n302), .ZN(new_n303));
  NAND3_X1  g0103(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n304));
  NAND2_X1  g0104(.A1(G1), .A2(G13), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n303), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT11), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n277), .A2(G13), .A3(G20), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(G68), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  XNOR2_X1  g0113(.A(new_n313), .B(KEYINPUT12), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n303), .A2(KEYINPUT11), .A3(new_n306), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n306), .B1(new_n277), .B2(G20), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(G68), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n309), .A2(new_n314), .A3(new_n315), .A4(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n295), .A2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n318), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n285), .A2(G200), .A3(new_n286), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n290), .A2(G190), .A3(new_n291), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT9), .ZN(new_n324));
  OAI21_X1  g0124(.A(G20), .B1(new_n201), .B2(new_n203), .ZN(new_n325));
  INV_X1    g0125(.A(G150), .ZN(new_n326));
  XNOR2_X1  g0126(.A(KEYINPUT8), .B(G58), .ZN(new_n327));
  OAI221_X1 g0127(.A(new_n325), .B1(new_n326), .B2(new_n302), .C1(new_n297), .C2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(new_n306), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n311), .A2(new_n257), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n316), .A2(G50), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n329), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n261), .A2(G223), .A3(G1698), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n261), .A2(new_n262), .ZN(new_n334));
  INV_X1    g0134(.A(G222), .ZN(new_n335));
  OAI221_X1 g0135(.A(new_n333), .B1(new_n298), .B2(new_n261), .C1(new_n334), .C2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(new_n270), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n281), .A2(G226), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n337), .A2(new_n279), .A3(new_n338), .ZN(new_n339));
  AOI22_X1  g0139(.A1(new_n324), .A2(new_n332), .B1(new_n339), .B2(G200), .ZN(new_n340));
  INV_X1    g0140(.A(new_n332), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(KEYINPUT9), .ZN(new_n342));
  INV_X1    g0142(.A(G190), .ZN(new_n343));
  OAI211_X1 g0143(.A(new_n340), .B(new_n342), .C1(new_n343), .C2(new_n339), .ZN(new_n344));
  XNOR2_X1  g0144(.A(new_n344), .B(KEYINPUT10), .ZN(new_n345));
  INV_X1    g0145(.A(G169), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n339), .A2(new_n346), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n339), .A2(G179), .ZN(new_n348));
  AND2_X1   g0148(.A1(new_n348), .A2(KEYINPUT72), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n348), .A2(KEYINPUT72), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n332), .B(new_n347), .C1(new_n349), .C2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(G20), .A2(G77), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n352), .B1(new_n327), .B2(new_n302), .ZN(new_n353));
  OR2_X1    g0153(.A1(KEYINPUT15), .A2(G87), .ZN(new_n354));
  NAND2_X1  g0154(.A1(KEYINPUT15), .A2(G87), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n356), .A2(new_n297), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n306), .B1(new_n353), .B2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT74), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  OAI211_X1 g0160(.A(KEYINPUT74), .B(new_n306), .C1(new_n353), .C2(new_n357), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n310), .A2(G77), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n316), .A2(G77), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n362), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n261), .A2(G238), .A3(G1698), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n261), .A2(G232), .A3(new_n262), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n265), .A2(KEYINPUT3), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT3), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(G33), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(G107), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n367), .A2(new_n368), .A3(new_n373), .ZN(new_n374));
  AND2_X1   g0174(.A1(new_n276), .A2(new_n278), .ZN(new_n375));
  AOI22_X1  g0175(.A1(new_n374), .A2(new_n270), .B1(new_n273), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n281), .A2(G244), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(new_n346), .ZN(new_n379));
  INV_X1    g0179(.A(G179), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n376), .A2(new_n380), .A3(new_n377), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n366), .A2(new_n379), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n374), .A2(new_n270), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n383), .A2(G190), .A3(new_n279), .A4(new_n377), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(KEYINPUT73), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT73), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n376), .A2(new_n386), .A3(G190), .A4(new_n377), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n366), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n378), .A2(G200), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n388), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n345), .A2(new_n351), .A3(new_n382), .A4(new_n391), .ZN(new_n392));
  OAI211_X1 g0192(.A(new_n319), .B(new_n323), .C1(new_n392), .C2(KEYINPUT75), .ZN(new_n393));
  AND2_X1   g0193(.A1(new_n392), .A2(KEYINPUT75), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n269), .A2(G232), .A3(new_n280), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n279), .A2(new_n395), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n369), .A2(new_n371), .A3(G223), .A4(new_n262), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT79), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n261), .A2(KEYINPUT79), .A3(G223), .A4(new_n262), .ZN(new_n400));
  NAND2_X1  g0200(.A1(G33), .A2(G87), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n261), .A2(G226), .A3(G1698), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n399), .A2(new_n400), .A3(new_n401), .A4(new_n402), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n396), .B1(new_n403), .B2(new_n270), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT80), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n404), .A2(new_n405), .A3(new_n380), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT81), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n404), .A2(new_n408), .ZN(new_n409));
  AOI211_X1 g0209(.A(KEYINPUT81), .B(new_n396), .C1(new_n403), .C2(new_n270), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n407), .B1(new_n411), .B2(new_n346), .ZN(new_n412));
  AOI21_X1  g0212(.A(KEYINPUT7), .B1(new_n372), .B2(new_n296), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT7), .ZN(new_n414));
  AOI211_X1 g0214(.A(new_n414), .B(G20), .C1(new_n369), .C2(new_n371), .ZN(new_n415));
  OAI21_X1  g0215(.A(G68), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n230), .A2(new_n312), .ZN(new_n417));
  OAI21_X1  g0217(.A(G20), .B1(new_n417), .B2(new_n202), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n301), .A2(G159), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n416), .A2(KEYINPUT16), .A3(new_n421), .ZN(new_n422));
  OAI21_X1  g0222(.A(KEYINPUT78), .B1(new_n265), .B2(KEYINPUT3), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT78), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n424), .A2(new_n370), .A3(G33), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n423), .A2(new_n425), .A3(new_n369), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n426), .A2(KEYINPUT7), .A3(new_n296), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n414), .B1(new_n261), .B2(G20), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n420), .B1(new_n429), .B2(G68), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n306), .B(new_n422), .C1(new_n430), .C2(KEYINPUT16), .ZN(new_n431));
  INV_X1    g0231(.A(new_n327), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n432), .A2(new_n310), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n433), .B1(new_n316), .B2(new_n432), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n431), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n399), .A2(new_n400), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n402), .A2(new_n401), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n270), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n396), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  OAI21_X1  g0240(.A(KEYINPUT80), .B1(new_n440), .B2(G179), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n412), .A2(KEYINPUT18), .A3(new_n435), .A4(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n440), .A2(KEYINPUT81), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n404), .A2(new_n408), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n443), .A2(new_n346), .A3(new_n444), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n445), .A2(new_n435), .A3(new_n441), .A4(new_n406), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT18), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n442), .A2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n435), .ZN(new_n450));
  XOR2_X1   g0250(.A(KEYINPUT83), .B(KEYINPUT17), .Z(new_n451));
  INV_X1    g0251(.A(G200), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n443), .A2(new_n452), .A3(new_n444), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT82), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n440), .A2(G190), .ZN(new_n455));
  INV_X1    g0255(.A(new_n455), .ZN(new_n456));
  AND3_X1   g0256(.A1(new_n453), .A2(new_n454), .A3(new_n456), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n454), .B1(new_n453), .B2(new_n456), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n450), .B(new_n451), .C1(new_n457), .C2(new_n458), .ZN(new_n459));
  OR2_X1    g0259(.A1(KEYINPUT83), .A2(KEYINPUT17), .ZN(new_n460));
  NOR3_X1   g0260(.A1(new_n409), .A2(new_n410), .A3(G200), .ZN(new_n461));
  OAI21_X1  g0261(.A(KEYINPUT82), .B1(new_n461), .B2(new_n455), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n453), .A2(new_n454), .A3(new_n456), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n435), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n449), .B(new_n459), .C1(new_n460), .C2(new_n464), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n369), .A2(new_n371), .A3(G244), .A4(new_n262), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT4), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n261), .A2(KEYINPUT4), .A3(G244), .A4(new_n262), .ZN(new_n469));
  NAND2_X1  g0269(.A1(G33), .A2(G283), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n261), .A2(G250), .A3(G1698), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n468), .A2(new_n469), .A3(new_n470), .A4(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(new_n270), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT86), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(G45), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n476), .A2(G1), .ZN(new_n477));
  AND2_X1   g0277(.A1(KEYINPUT5), .A2(G41), .ZN(new_n478));
  NOR2_X1   g0278(.A1(KEYINPUT5), .A2(G41), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n480), .A2(G257), .A3(new_n269), .ZN(new_n481));
  XNOR2_X1  g0281(.A(KEYINPUT5), .B(G41), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n273), .A2(new_n477), .A3(new_n482), .ZN(new_n483));
  AND3_X1   g0283(.A1(new_n481), .A2(new_n483), .A3(KEYINPUT87), .ZN(new_n484));
  AOI21_X1  g0284(.A(KEYINPUT87), .B1(new_n481), .B2(new_n483), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n472), .A2(KEYINPUT86), .A3(new_n270), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n475), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(G200), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n311), .A2(new_n266), .ZN(new_n490));
  INV_X1    g0290(.A(new_n306), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n277), .A2(G33), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n491), .A2(new_n310), .A3(new_n492), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n490), .B1(new_n493), .B2(new_n266), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n266), .A2(new_n252), .A3(KEYINPUT6), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT85), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT6), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(G97), .ZN(new_n498));
  AND3_X1   g0298(.A1(new_n495), .A2(new_n496), .A3(new_n498), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n496), .B1(new_n495), .B2(new_n498), .ZN(new_n500));
  NOR3_X1   g0300(.A1(new_n499), .A2(new_n500), .A3(new_n252), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n495), .A2(new_n498), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(KEYINPUT85), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n495), .A2(new_n496), .A3(new_n498), .ZN(new_n504));
  AOI21_X1  g0304(.A(G107), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  OAI21_X1  g0305(.A(G20), .B1(new_n501), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n429), .A2(G107), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n301), .A2(G77), .ZN(new_n508));
  XOR2_X1   g0308(.A(new_n508), .B(KEYINPUT84), .Z(new_n509));
  NAND3_X1  g0309(.A1(new_n506), .A2(new_n507), .A3(new_n509), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n494), .B1(new_n510), .B2(new_n306), .ZN(new_n511));
  INV_X1    g0311(.A(new_n485), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n481), .A2(new_n483), .A3(KEYINPUT87), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n473), .A2(new_n512), .A3(G190), .A4(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT88), .ZN(new_n515));
  AND2_X1   g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n514), .A2(new_n515), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n489), .B(new_n511), .C1(new_n516), .C2(new_n517), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n493), .A2(new_n252), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n369), .A2(new_n371), .A3(new_n296), .A4(G87), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(KEYINPUT22), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT22), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n261), .A2(new_n522), .A3(new_n296), .A4(G87), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n296), .A2(G33), .A3(G116), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n296), .A2(G107), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT23), .ZN(new_n527));
  OAI21_X1  g0327(.A(KEYINPUT92), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT92), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n529), .B(KEYINPUT23), .C1(new_n296), .C2(G107), .ZN(new_n530));
  AOI22_X1  g0330(.A1(new_n528), .A2(new_n530), .B1(new_n527), .B2(new_n526), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n524), .A2(new_n525), .A3(new_n531), .ZN(new_n532));
  XNOR2_X1  g0332(.A(KEYINPUT91), .B(KEYINPUT24), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n524), .A2(new_n533), .A3(new_n531), .A4(new_n525), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n519), .B1(new_n537), .B2(new_n306), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n310), .A2(G107), .ZN(new_n539));
  XNOR2_X1  g0339(.A(new_n539), .B(KEYINPUT25), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n369), .A2(new_n371), .A3(G257), .A4(G1698), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(KEYINPUT93), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT93), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n261), .A2(new_n543), .A3(G257), .A4(G1698), .ZN(new_n544));
  NAND2_X1  g0344(.A1(G33), .A2(G294), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n261), .A2(G250), .A3(new_n262), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n542), .A2(new_n544), .A3(new_n545), .A4(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n480), .A2(new_n269), .ZN(new_n548));
  INV_X1    g0348(.A(new_n548), .ZN(new_n549));
  AOI22_X1  g0349(.A1(new_n547), .A2(new_n270), .B1(G264), .B2(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n550), .A2(G190), .A3(new_n483), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n483), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(G200), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n538), .A2(new_n540), .A3(new_n551), .A4(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n277), .A2(G45), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n269), .A2(G250), .A3(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(new_n556), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n369), .A2(new_n371), .A3(G244), .A4(G1698), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n369), .A2(new_n371), .A3(G238), .A4(new_n262), .ZN(new_n559));
  NAND2_X1  g0359(.A1(G33), .A2(G116), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n557), .B1(new_n561), .B2(new_n270), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n477), .A2(G274), .ZN(new_n563));
  AOI21_X1  g0363(.A(G169), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n296), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n232), .A2(new_n266), .A3(new_n252), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n369), .A2(new_n371), .A3(new_n296), .A4(G68), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n296), .A2(G33), .A3(G97), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT19), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n568), .A2(new_n569), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(new_n306), .ZN(new_n574));
  INV_X1    g0374(.A(new_n356), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n575), .A2(new_n310), .ZN(new_n576));
  INV_X1    g0376(.A(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n574), .A2(new_n577), .A3(KEYINPUT89), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT89), .ZN(new_n579));
  AOI22_X1  g0379(.A1(new_n566), .A2(new_n567), .B1(new_n570), .B2(new_n571), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n491), .B1(new_n580), .B2(new_n569), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n579), .B1(new_n581), .B2(new_n576), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n578), .A2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(new_n493), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n575), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n564), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n562), .A2(new_n380), .A3(new_n563), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n561), .A2(new_n270), .ZN(new_n588));
  AND4_X1   g0388(.A1(G190), .A2(new_n588), .A3(new_n563), .A4(new_n556), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n452), .B1(new_n562), .B2(new_n563), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  AOI22_X1  g0391(.A1(new_n578), .A2(new_n582), .B1(G87), .B2(new_n584), .ZN(new_n592));
  AOI22_X1  g0392(.A1(new_n586), .A2(new_n587), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n486), .A2(new_n473), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n346), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n475), .A2(new_n380), .A3(new_n486), .A4(new_n487), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n252), .B1(new_n499), .B2(new_n500), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n503), .A2(new_n504), .A3(G107), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  AOI22_X1  g0399(.A1(new_n599), .A2(G20), .B1(G107), .B2(new_n429), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n491), .B1(new_n600), .B2(new_n509), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n595), .B(new_n596), .C1(new_n601), .C2(new_n494), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n518), .A2(new_n554), .A3(new_n593), .A4(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT21), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n261), .A2(G264), .A3(G1698), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n372), .A2(G303), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n606), .B(new_n607), .C1(new_n334), .C2(new_n210), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n270), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n549), .A2(G270), .ZN(new_n610));
  AND3_X1   g0410(.A1(new_n609), .A2(new_n610), .A3(new_n483), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n311), .A2(new_n254), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n304), .A2(new_n305), .B1(G20), .B2(new_n254), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n470), .B(new_n296), .C1(G33), .C2(new_n266), .ZN(new_n614));
  AND3_X1   g0414(.A1(new_n613), .A2(KEYINPUT20), .A3(new_n614), .ZN(new_n615));
  AOI21_X1  g0415(.A(KEYINPUT20), .B1(new_n613), .B2(new_n614), .ZN(new_n616));
  OAI221_X1 g0416(.A(new_n612), .B1(new_n493), .B2(new_n254), .C1(new_n615), .C2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(G169), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n605), .B1(new_n611), .B2(new_n618), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n611), .A2(G179), .A3(new_n617), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n609), .A2(new_n610), .A3(new_n483), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n621), .A2(KEYINPUT21), .A3(G169), .A4(new_n617), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n619), .A2(new_n620), .A3(new_n622), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n552), .A2(G179), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n624), .B1(new_n538), .B2(new_n540), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n552), .A2(new_n346), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n623), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n617), .B1(new_n621), .B2(G200), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n628), .B1(new_n343), .B2(new_n621), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT90), .ZN(new_n630));
  XNOR2_X1  g0430(.A(new_n629), .B(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n604), .A2(new_n627), .A3(new_n631), .ZN(new_n632));
  NOR4_X1   g0432(.A1(new_n393), .A2(new_n394), .A3(new_n465), .A4(new_n632), .ZN(G372));
  NOR3_X1   g0433(.A1(new_n393), .A2(new_n394), .A3(new_n465), .ZN(new_n634));
  INV_X1    g0434(.A(new_n596), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n635), .A2(new_n511), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n636), .A2(new_n593), .A3(KEYINPUT26), .A4(new_n595), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT26), .ZN(new_n638));
  AOI21_X1  g0438(.A(KEYINPUT89), .B1(new_n574), .B2(new_n577), .ZN(new_n639));
  NOR3_X1   g0439(.A1(new_n581), .A2(new_n579), .A3(new_n576), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n585), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n564), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n641), .A2(new_n642), .A3(new_n587), .ZN(new_n643));
  INV_X1    g0443(.A(new_n590), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n562), .A2(G190), .A3(new_n563), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n592), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n643), .A2(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n638), .B1(new_n602), .B2(new_n647), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n637), .A2(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n643), .B1(new_n603), .B2(new_n627), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n634), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n319), .A2(new_n382), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(new_n323), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n459), .B1(new_n464), .B2(new_n460), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AND3_X1   g0455(.A1(new_n442), .A2(new_n448), .A3(KEYINPUT94), .ZN(new_n656));
  AOI21_X1  g0456(.A(KEYINPUT94), .B1(new_n442), .B2(new_n448), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n345), .B1(new_n655), .B2(new_n658), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n659), .A2(new_n351), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n651), .A2(new_n660), .ZN(G369));
  INV_X1    g0461(.A(G330), .ZN(new_n662));
  INV_X1    g0462(.A(new_n623), .ZN(new_n663));
  INV_X1    g0463(.A(G13), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n664), .A2(G20), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(new_n277), .ZN(new_n666));
  OR2_X1    g0466(.A1(new_n666), .A2(KEYINPUT27), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(KEYINPUT27), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n667), .A2(G213), .A3(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(G343), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n617), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n663), .B1(new_n631), .B2(new_n673), .ZN(new_n674));
  XNOR2_X1  g0474(.A(new_n674), .B(KEYINPUT96), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n672), .A2(KEYINPUT95), .ZN(new_n676));
  OR2_X1    g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n675), .A2(new_n676), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n662), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n625), .A2(new_n626), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n680), .A2(new_n671), .ZN(new_n681));
  AND2_X1   g0481(.A1(new_n538), .A2(new_n540), .ZN(new_n682));
  INV_X1    g0482(.A(new_n671), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n554), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n681), .B1(new_n680), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n679), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n684), .A2(new_n680), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n663), .A2(new_n671), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n681), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n686), .A2(new_n689), .ZN(G399));
  NOR2_X1   g0490(.A1(new_n209), .A2(G41), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n567), .A2(G116), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n692), .A2(G1), .A3(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n694), .B1(new_n219), .B2(new_n692), .ZN(new_n695));
  XNOR2_X1  g0495(.A(new_n695), .B(KEYINPUT28), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT30), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n611), .A2(G179), .ZN(new_n698));
  INV_X1    g0498(.A(new_n550), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n562), .A2(new_n563), .ZN(new_n700));
  OR3_X1    g0500(.A1(new_n698), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n697), .B1(new_n701), .B2(new_n594), .ZN(new_n702));
  NOR4_X1   g0502(.A1(new_n698), .A2(new_n699), .A3(new_n594), .A4(new_n700), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(KEYINPUT30), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n611), .A2(G179), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n705), .A2(new_n552), .A3(new_n700), .A4(new_n488), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n702), .A2(new_n704), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(new_n671), .ZN(new_n708));
  OAI211_X1 g0508(.A(new_n708), .B(KEYINPUT31), .C1(new_n632), .C2(new_n671), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT31), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n707), .A2(new_n710), .A3(new_n671), .ZN(new_n711));
  AND2_X1   g0511(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(G330), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT97), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n637), .A2(new_n648), .A3(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n602), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n716), .A2(KEYINPUT97), .A3(KEYINPUT26), .A4(new_n593), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n683), .B1(new_n718), .B2(new_n650), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(KEYINPUT29), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n683), .B1(new_n650), .B2(new_n649), .ZN(new_n721));
  OR2_X1    g0521(.A1(new_n721), .A2(KEYINPUT29), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n713), .A2(new_n720), .A3(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n696), .B1(new_n724), .B2(G1), .ZN(G364));
  NAND2_X1  g0525(.A1(new_n665), .A2(G45), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n692), .A2(G1), .A3(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n679), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n677), .A2(new_n678), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n729), .B1(G330), .B2(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n305), .B1(G20), .B2(new_n346), .ZN(new_n732));
  XNOR2_X1  g0532(.A(new_n732), .B(KEYINPUT101), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n296), .A2(G190), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n452), .A2(G179), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(new_n252), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n296), .A2(new_n343), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n380), .A2(G200), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n738), .A2(new_n735), .ZN(new_n741));
  OAI22_X1  g0541(.A1(new_n230), .A2(new_n740), .B1(new_n741), .B2(new_n232), .ZN(new_n742));
  NOR2_X1   g0542(.A1(G179), .A2(G200), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n296), .B1(new_n743), .B2(G190), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  AOI211_X1 g0545(.A(new_n737), .B(new_n742), .C1(G97), .C2(new_n745), .ZN(new_n746));
  NAND3_X1  g0546(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(G190), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(G68), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n734), .A2(new_n743), .ZN(new_n750));
  INV_X1    g0550(.A(G159), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT32), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n747), .A2(new_n343), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  OAI22_X1  g0555(.A1(new_n752), .A2(new_n753), .B1(new_n257), .B2(new_n755), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n756), .B1(new_n753), .B2(new_n752), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n734), .A2(new_n739), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n372), .B1(new_n759), .B2(G77), .ZN(new_n760));
  NAND4_X1  g0560(.A1(new_n746), .A2(new_n749), .A3(new_n757), .A4(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(G303), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n741), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(G311), .ZN(new_n764));
  INV_X1    g0564(.A(G329), .ZN(new_n765));
  OAI22_X1  g0565(.A1(new_n758), .A2(new_n764), .B1(new_n750), .B2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n736), .ZN(new_n767));
  AOI211_X1 g0567(.A(new_n763), .B(new_n766), .C1(G283), .C2(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n754), .A2(G326), .ZN(new_n769));
  INV_X1    g0569(.A(G294), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n372), .B1(new_n744), .B2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n740), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n771), .B1(G322), .B2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(G317), .ZN(new_n774));
  OR2_X1    g0574(.A1(new_n774), .A2(KEYINPUT33), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n774), .A2(KEYINPUT33), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n748), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  NAND4_X1  g0577(.A1(new_n768), .A2(new_n769), .A3(new_n773), .A4(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n733), .B1(new_n761), .B2(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n372), .A2(new_n208), .ZN(new_n780));
  XOR2_X1   g0580(.A(new_n780), .B(KEYINPUT99), .Z(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n259), .A2(G45), .ZN(new_n783));
  INV_X1    g0583(.A(KEYINPUT98), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n782), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  OAI221_X1 g0585(.A(new_n785), .B1(new_n784), .B2(new_n783), .C1(G45), .C2(new_n219), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n209), .A2(new_n372), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(G355), .ZN(new_n788));
  OAI211_X1 g0588(.A(new_n786), .B(new_n788), .C1(G116), .C2(new_n208), .ZN(new_n789));
  NOR2_X1   g0589(.A1(G13), .A2(G33), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(new_n296), .ZN(new_n791));
  XNOR2_X1  g0591(.A(new_n791), .B(KEYINPUT100), .ZN(new_n792));
  AND2_X1   g0592(.A1(new_n733), .A2(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n779), .B1(new_n789), .B2(new_n793), .ZN(new_n794));
  OAI211_X1 g0594(.A(new_n728), .B(new_n794), .C1(new_n730), .C2(new_n792), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n731), .A2(new_n795), .ZN(G396));
  AND3_X1   g0596(.A1(new_n366), .A2(new_n379), .A3(new_n381), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n366), .A2(new_n671), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n797), .B1(new_n391), .B2(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n382), .A2(new_n671), .ZN(new_n800));
  OAI21_X1  g0600(.A(KEYINPUT105), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(KEYINPUT105), .ZN(new_n802));
  INV_X1    g0602(.A(new_n800), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n366), .B1(new_n385), .B2(new_n387), .ZN(new_n804));
  AOI22_X1  g0604(.A1(new_n804), .A2(new_n390), .B1(new_n366), .B2(new_n671), .ZN(new_n805));
  OAI211_X1 g0605(.A(new_n802), .B(new_n803), .C1(new_n805), .C2(new_n797), .ZN(new_n806));
  AND2_X1   g0606(.A1(new_n801), .A2(new_n806), .ZN(new_n807));
  OAI211_X1 g0607(.A(new_n807), .B(new_n683), .C1(new_n649), .C2(new_n650), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n801), .A2(new_n806), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n721), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n713), .A2(new_n811), .ZN(new_n812));
  OR2_X1    g0612(.A1(new_n812), .A2(KEYINPUT106), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n812), .A2(KEYINPUT106), .ZN(new_n814));
  OR2_X1    g0614(.A1(new_n713), .A2(new_n811), .ZN(new_n815));
  NAND4_X1  g0615(.A1(new_n813), .A2(new_n727), .A3(new_n814), .A4(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n741), .ZN(new_n817));
  AOI22_X1  g0617(.A1(G50), .A2(new_n817), .B1(new_n767), .B2(G68), .ZN(new_n818));
  INV_X1    g0618(.A(KEYINPUT103), .ZN(new_n819));
  AND2_X1   g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  OAI221_X1 g0620(.A(new_n261), .B1(new_n230), .B2(new_n744), .C1(new_n818), .C2(new_n819), .ZN(new_n821));
  AOI22_X1  g0621(.A1(new_n759), .A2(G159), .B1(G137), .B2(new_n754), .ZN(new_n822));
  INV_X1    g0622(.A(G143), .ZN(new_n823));
  INV_X1    g0623(.A(new_n748), .ZN(new_n824));
  OAI221_X1 g0624(.A(new_n822), .B1(new_n823), .B2(new_n740), .C1(new_n326), .C2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT34), .ZN(new_n826));
  AOI211_X1 g0626(.A(new_n820), .B(new_n821), .C1(new_n825), .C2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n750), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(G132), .ZN(new_n829));
  OAI211_X1 g0629(.A(new_n827), .B(new_n829), .C1(new_n826), .C2(new_n825), .ZN(new_n830));
  INV_X1    g0630(.A(G283), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n824), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n767), .A2(G87), .ZN(new_n833));
  OAI221_X1 g0633(.A(new_n833), .B1(new_n770), .B2(new_n740), .C1(new_n764), .C2(new_n750), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n834), .B1(G116), .B2(new_n759), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n372), .B1(new_n741), .B2(new_n252), .ZN(new_n836));
  XNOR2_X1  g0636(.A(new_n836), .B(KEYINPUT102), .ZN(new_n837));
  AOI22_X1  g0637(.A1(new_n745), .A2(G97), .B1(G303), .B2(new_n754), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n835), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n830), .B1(new_n832), .B2(new_n839), .ZN(new_n840));
  XNOR2_X1  g0640(.A(new_n840), .B(KEYINPUT104), .ZN(new_n841));
  INV_X1    g0641(.A(new_n733), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n727), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n842), .A2(new_n790), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n790), .ZN(new_n846));
  OAI221_X1 g0646(.A(new_n843), .B1(G77), .B2(new_n845), .C1(new_n846), .C2(new_n807), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n816), .A2(new_n847), .ZN(G384));
  OAI21_X1  g0648(.A(new_n803), .B1(new_n721), .B2(new_n809), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n318), .A2(new_n671), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n319), .A2(new_n323), .A3(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n323), .ZN(new_n852));
  OAI211_X1 g0652(.A(new_n318), .B(new_n671), .C1(new_n852), .C2(new_n295), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n849), .A2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n434), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n416), .A2(new_n421), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT16), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n491), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n372), .A2(KEYINPUT7), .A3(new_n296), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n428), .A2(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n420), .B1(new_n861), .B2(G68), .ZN(new_n862));
  AOI22_X1  g0662(.A1(new_n859), .A2(KEYINPUT107), .B1(KEYINPUT16), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n306), .B1(new_n862), .B2(KEYINPUT16), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT107), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n856), .B1(new_n863), .B2(new_n866), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n867), .A2(new_n669), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT37), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n450), .B1(new_n457), .B2(new_n458), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n450), .A2(new_n669), .ZN(new_n871));
  INV_X1    g0671(.A(new_n871), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n870), .A2(new_n446), .A3(new_n872), .ZN(new_n873));
  AOI22_X1  g0673(.A1(new_n465), .A2(new_n868), .B1(new_n869), .B2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT108), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n445), .A2(new_n441), .A3(new_n406), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n867), .A2(new_n876), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n875), .B1(new_n464), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n859), .A2(KEYINPUT107), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n879), .A2(new_n422), .A3(new_n866), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(new_n434), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n881), .A2(new_n441), .A3(new_n412), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n870), .A2(KEYINPUT108), .A3(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n868), .ZN(new_n884));
  NAND4_X1  g0684(.A1(new_n878), .A2(new_n883), .A3(KEYINPUT37), .A4(new_n884), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n874), .A2(KEYINPUT38), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n465), .A2(new_n868), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n873), .A2(new_n869), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n887), .A2(new_n885), .A3(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT38), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n855), .B1(new_n886), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n658), .A2(new_n669), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(KEYINPUT109), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n854), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n896), .B1(new_n808), .B2(new_n803), .ZN(new_n897));
  AND3_X1   g0697(.A1(new_n874), .A2(KEYINPUT38), .A3(new_n885), .ZN(new_n898));
  AOI21_X1  g0698(.A(KEYINPUT38), .B1(new_n874), .B2(new_n885), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n897), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT109), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n900), .A2(new_n901), .A3(new_n893), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n895), .A2(new_n902), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n871), .B1(new_n658), .B2(new_n654), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n870), .A2(new_n872), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT94), .ZN(new_n906));
  OAI21_X1  g0706(.A(KEYINPUT37), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n462), .A2(new_n463), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n871), .B1(new_n908), .B2(new_n450), .ZN(new_n909));
  AOI21_X1  g0709(.A(KEYINPUT110), .B1(new_n909), .B2(new_n446), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT110), .ZN(new_n911));
  INV_X1    g0711(.A(new_n446), .ZN(new_n912));
  NOR4_X1   g0712(.A1(new_n464), .A2(new_n911), .A3(new_n912), .A4(new_n871), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n907), .B1(new_n910), .B2(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n869), .B1(new_n909), .B2(KEYINPUT94), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n873), .A2(new_n911), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n909), .A2(KEYINPUT110), .A3(new_n446), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n904), .A2(new_n914), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(new_n890), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT39), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n920), .A2(new_n921), .A3(new_n886), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n891), .A2(new_n886), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(KEYINPUT39), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n319), .A2(new_n671), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  AND3_X1   g0727(.A1(new_n903), .A2(new_n927), .A3(KEYINPUT111), .ZN(new_n928));
  AOI21_X1  g0728(.A(KEYINPUT111), .B1(new_n903), .B2(new_n927), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n930), .B(KEYINPUT112), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT40), .ZN(new_n932));
  AND4_X1   g0732(.A1(new_n709), .A2(new_n711), .A3(new_n807), .A4(new_n854), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n923), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  NAND4_X1  g0734(.A1(new_n709), .A2(new_n711), .A3(new_n807), .A4(new_n854), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n935), .B1(new_n920), .B2(new_n886), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n934), .B1(new_n936), .B2(new_n932), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n634), .A2(new_n712), .ZN(new_n938));
  XOR2_X1   g0738(.A(new_n937), .B(new_n938), .Z(new_n939));
  NOR2_X1   g0739(.A1(new_n939), .A2(new_n662), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n931), .B(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n722), .A2(new_n720), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n634), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(new_n660), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n941), .B(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n945), .B1(new_n277), .B2(new_n665), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n254), .B1(new_n599), .B2(KEYINPUT35), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n305), .A2(new_n296), .ZN(new_n948));
  OAI211_X1 g0748(.A(new_n947), .B(new_n948), .C1(KEYINPUT35), .C2(new_n599), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n949), .B(KEYINPUT36), .ZN(new_n950));
  NOR3_X1   g0750(.A1(new_n219), .A2(new_n298), .A3(new_n417), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n201), .A2(new_n312), .ZN(new_n952));
  OAI211_X1 g0752(.A(G1), .B(new_n664), .C1(new_n951), .C2(new_n952), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n946), .A2(new_n950), .A3(new_n953), .ZN(G367));
  OAI211_X1 g0754(.A(new_n518), .B(new_n602), .C1(new_n511), .C2(new_n683), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n716), .A2(new_n671), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n679), .A2(new_n685), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n685), .A2(new_n688), .ZN(new_n959));
  INV_X1    g0759(.A(new_n957), .ZN(new_n960));
  OR3_X1    g0760(.A1(new_n959), .A2(KEYINPUT42), .A3(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n602), .B1(new_n955), .B2(new_n680), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(new_n683), .ZN(new_n963));
  OAI21_X1  g0763(.A(KEYINPUT42), .B1(new_n959), .B2(new_n960), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n961), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n592), .A2(new_n683), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n966), .A2(new_n586), .A3(new_n587), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n967), .B1(new_n647), .B2(new_n966), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n968), .A2(KEYINPUT43), .ZN(new_n969));
  AND2_X1   g0769(.A1(new_n965), .A2(new_n969), .ZN(new_n970));
  OR2_X1    g0770(.A1(new_n958), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n958), .A2(new_n969), .A3(new_n965), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n968), .A2(KEYINPUT43), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n973), .B(new_n974), .ZN(new_n975));
  XOR2_X1   g0775(.A(KEYINPUT113), .B(KEYINPUT41), .Z(new_n976));
  XOR2_X1   g0776(.A(new_n691), .B(new_n976), .Z(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n685), .B(new_n688), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n679), .B(new_n979), .ZN(new_n980));
  AND2_X1   g0780(.A1(new_n980), .A2(new_n724), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n689), .A2(new_n957), .ZN(new_n982));
  XOR2_X1   g0782(.A(new_n982), .B(KEYINPUT44), .Z(new_n983));
  NAND2_X1  g0783(.A1(new_n689), .A2(new_n957), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(KEYINPUT45), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(KEYINPUT114), .B1(new_n686), .B2(new_n986), .ZN(new_n987));
  AND2_X1   g0787(.A1(new_n686), .A2(new_n986), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n686), .A2(new_n986), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  OAI211_X1 g0790(.A(new_n981), .B(new_n987), .C1(KEYINPUT114), .C2(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n978), .B1(new_n991), .B2(new_n724), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n726), .A2(G1), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n975), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n248), .A2(new_n781), .B1(new_n209), .B2(new_n575), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n727), .B1(new_n995), .B2(new_n793), .ZN(new_n996));
  XOR2_X1   g0796(.A(new_n996), .B(KEYINPUT115), .Z(new_n997));
  OAI22_X1  g0797(.A1(new_n758), .A2(new_n831), .B1(new_n744), .B2(new_n252), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n998), .B(KEYINPUT116), .Z(new_n999));
  NOR2_X1   g0799(.A1(new_n736), .A2(new_n266), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n372), .B1(new_n740), .B2(new_n762), .ZN(new_n1001));
  AOI211_X1 g0801(.A(new_n1000), .B(new_n1001), .C1(G317), .C2(new_n828), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(new_n748), .A2(G294), .B1(new_n754), .B2(G311), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n817), .A2(G116), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT46), .ZN(new_n1005));
  NAND4_X1  g0805(.A1(new_n999), .A2(new_n1002), .A3(new_n1003), .A4(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n745), .A2(G68), .ZN(new_n1007));
  OAI221_X1 g0807(.A(new_n1007), .B1(new_n326), .B2(new_n740), .C1(new_n755), .C2(new_n823), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT117), .ZN(new_n1009));
  INV_X1    g0809(.A(G137), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n261), .B1(new_n750), .B2(new_n1010), .C1(new_n230), .C2(new_n741), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n201), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n1012), .A2(new_n758), .B1(new_n824), .B2(new_n751), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT118), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1011), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  OAI211_X1 g0815(.A(new_n1009), .B(new_n1015), .C1(new_n1014), .C2(new_n1013), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n736), .A2(new_n298), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1006), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  XOR2_X1   g0818(.A(new_n1018), .B(KEYINPUT47), .Z(new_n1019));
  OAI221_X1 g0819(.A(new_n997), .B1(new_n792), .B2(new_n968), .C1(new_n1019), .C2(new_n733), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n994), .A2(new_n1020), .ZN(G387));
  NOR2_X1   g0821(.A1(new_n980), .A2(new_n724), .ZN(new_n1022));
  OR3_X1    g0822(.A1(new_n981), .A2(new_n1022), .A3(new_n692), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n980), .A2(new_n993), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n782), .B1(new_n245), .B2(G45), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n693), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1025), .B1(new_n1026), .B2(new_n787), .ZN(new_n1027));
  OR3_X1    g0827(.A1(new_n327), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1028));
  OAI21_X1  g0828(.A(KEYINPUT50), .B1(new_n327), .B2(G50), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n1028), .A2(new_n1029), .A3(new_n476), .A4(new_n693), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1030), .B1(G68), .B2(G77), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n1027), .A2(new_n1031), .B1(G107), .B2(new_n208), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n727), .B1(new_n1032), .B2(new_n793), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT119), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n759), .A2(G303), .B1(G322), .B2(new_n754), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n1035), .B1(new_n764), .B2(new_n824), .C1(new_n774), .C2(new_n740), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT48), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n1037), .B1(new_n831), .B2(new_n744), .C1(new_n770), .C2(new_n741), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT49), .ZN(new_n1039));
  OR2_X1    g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n828), .A2(G326), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n261), .B1(new_n767), .B2(G116), .ZN(new_n1043));
  NAND4_X1  g0843(.A1(new_n1040), .A2(new_n1041), .A3(new_n1042), .A4(new_n1043), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n741), .A2(new_n298), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n744), .A2(new_n356), .ZN(new_n1046));
  AOI211_X1 g0846(.A(new_n1000), .B(new_n1046), .C1(G159), .C2(new_n754), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n758), .A2(new_n312), .B1(new_n750), .B2(new_n326), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1048), .B1(G50), .B2(new_n772), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n372), .B1(new_n432), .B2(new_n748), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1047), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1044), .B1(new_n1045), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1052), .A2(new_n842), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n1034), .B(new_n1053), .C1(new_n685), .C2(new_n792), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1023), .A2(new_n1024), .A3(new_n1054), .ZN(G393));
  OAI211_X1 g0855(.A(new_n991), .B(new_n691), .C1(new_n981), .C2(new_n990), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n255), .A2(new_n781), .B1(G97), .B2(new_n209), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1057), .A2(new_n793), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n957), .A2(new_n792), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n833), .B1(new_n298), .B2(new_n744), .C1(new_n824), .C2(new_n1012), .ZN(new_n1060));
  AOI211_X1 g0860(.A(new_n372), .B(new_n1060), .C1(new_n432), .C2(new_n759), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n755), .A2(new_n326), .B1(new_n740), .B2(new_n751), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1062), .B(KEYINPUT51), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n741), .A2(new_n312), .B1(new_n750), .B2(new_n823), .ZN(new_n1064));
  XOR2_X1   g0864(.A(new_n1064), .B(KEYINPUT120), .Z(new_n1065));
  NAND3_X1  g0865(.A1(new_n1061), .A2(new_n1063), .A3(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n737), .B1(G303), .B2(new_n748), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(G283), .A2(new_n817), .B1(new_n828), .B2(G322), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n261), .B1(new_n745), .B2(G116), .ZN(new_n1069));
  AND3_X1   g0869(.A1(new_n1067), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n755), .A2(new_n774), .B1(new_n740), .B2(new_n764), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT52), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n1070), .B(new_n1072), .C1(new_n770), .C2(new_n758), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n733), .B1(new_n1066), .B2(new_n1073), .ZN(new_n1074));
  NOR3_X1   g0874(.A1(new_n1059), .A2(new_n727), .A3(new_n1074), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n990), .A2(new_n993), .B1(new_n1058), .B2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1056), .A2(new_n1076), .ZN(G390));
  NOR2_X1   g0877(.A1(new_n938), .A2(new_n662), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n1078), .A2(new_n944), .ZN(new_n1079));
  INV_X1    g0879(.A(KEYINPUT122), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n933), .A2(new_n1080), .A3(G330), .ZN(new_n1081));
  OAI21_X1  g0881(.A(KEYINPUT122), .B1(new_n935), .B2(new_n662), .ZN(new_n1082));
  NAND4_X1  g0882(.A1(new_n709), .A2(new_n711), .A3(G330), .A4(new_n807), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1083), .A2(new_n896), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1081), .A2(new_n1082), .A3(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(new_n849), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1084), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n935), .A2(new_n662), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n803), .B1(new_n719), .B2(new_n809), .ZN(new_n1089));
  OR3_X1    g0889(.A1(new_n1087), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1086), .A2(new_n1090), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n922), .B(new_n924), .C1(new_n926), .C2(new_n897), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n920), .A2(new_n886), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n926), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n1089), .A2(new_n854), .B1(KEYINPUT121), .B2(new_n1094), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n1093), .B(new_n1095), .C1(KEYINPUT121), .C2(new_n1094), .ZN(new_n1096));
  AND3_X1   g0896(.A1(new_n1092), .A2(new_n1096), .A3(new_n1088), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1098), .B1(new_n1092), .B2(new_n1096), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n1079), .B(new_n1091), .C1(new_n1097), .C2(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1099), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1091), .A2(new_n1079), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1092), .A2(new_n1096), .A3(new_n1088), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1101), .A2(new_n1102), .A3(new_n1103), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1100), .A2(new_n1104), .A3(new_n691), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n925), .A2(new_n846), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(G68), .A2(new_n767), .B1(new_n759), .B2(G97), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1107), .B1(new_n770), .B2(new_n750), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1108), .B1(G116), .B2(new_n772), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n824), .A2(new_n252), .B1(new_n755), .B2(new_n831), .ZN(new_n1110));
  AOI211_X1 g0910(.A(new_n261), .B(new_n1110), .C1(G77), .C2(new_n745), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n1109), .B(new_n1111), .C1(new_n232), .C2(new_n741), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n261), .B1(new_n824), .B2(new_n1010), .ZN(new_n1113));
  INV_X1    g0913(.A(G128), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n755), .A2(new_n1114), .B1(new_n744), .B2(new_n751), .ZN(new_n1115));
  AOI211_X1 g0915(.A(new_n1113), .B(new_n1115), .C1(G132), .C2(new_n772), .ZN(new_n1116));
  XOR2_X1   g0916(.A(KEYINPUT54), .B(G143), .Z(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(G125), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n1118), .A2(new_n758), .B1(new_n1119), .B2(new_n750), .ZN(new_n1120));
  INV_X1    g0920(.A(KEYINPUT53), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1121), .B1(new_n741), .B2(new_n326), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n817), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1120), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n1116), .B(new_n1124), .C1(new_n1012), .C2(new_n736), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n733), .B1(new_n1112), .B2(new_n1125), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n845), .A2(new_n432), .ZN(new_n1127));
  NOR4_X1   g0927(.A1(new_n1106), .A2(new_n727), .A3(new_n1126), .A4(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1128), .B1(new_n1129), .B2(new_n993), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1105), .A2(new_n1130), .ZN(G378));
  NOR2_X1   g0931(.A1(new_n341), .A2(new_n669), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1132), .ZN(new_n1133));
  AND3_X1   g0933(.A1(new_n345), .A2(new_n351), .A3(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1133), .B1(new_n345), .B2(new_n351), .ZN(new_n1135));
  NOR3_X1   g0935(.A1(new_n1134), .A2(new_n1135), .A3(KEYINPUT55), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  OAI21_X1  g0937(.A(KEYINPUT55), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1138));
  AND3_X1   g0938(.A1(new_n1137), .A2(KEYINPUT56), .A3(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(KEYINPUT56), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  AND3_X1   g0941(.A1(new_n937), .A2(G330), .A3(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1141), .B1(new_n937), .B2(G330), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n928), .A2(new_n929), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(KEYINPUT111), .ZN(new_n1145));
  AOI211_X1 g0945(.A(KEYINPUT109), .B(new_n894), .C1(new_n923), .C2(new_n897), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n901), .B1(new_n900), .B2(new_n893), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1094), .B1(new_n922), .B2(new_n924), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1145), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n937), .A2(G330), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1141), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n903), .A2(new_n927), .A3(KEYINPUT111), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n937), .A2(G330), .A3(new_n1141), .ZN(new_n1155));
  NAND4_X1  g0955(.A1(new_n1150), .A2(new_n1153), .A3(new_n1154), .A4(new_n1155), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1144), .A2(new_n1156), .A3(KEYINPUT123), .ZN(new_n1157));
  INV_X1    g0957(.A(KEYINPUT123), .ZN(new_n1158));
  OAI221_X1 g0958(.A(new_n1158), .B1(new_n1142), .B2(new_n1143), .C1(new_n928), .C2(new_n929), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1100), .A2(new_n1079), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1157), .A2(new_n1159), .A3(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(KEYINPUT57), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n1144), .A2(new_n1156), .B1(new_n1100), .B2(new_n1079), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n692), .B1(new_n1164), .B2(KEYINPUT57), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1163), .A2(new_n1165), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1157), .A2(new_n993), .A3(new_n1159), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1141), .A2(new_n790), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n844), .A2(new_n1012), .ZN(new_n1169));
  OAI221_X1 g0969(.A(new_n1007), .B1(new_n824), .B2(new_n266), .C1(new_n254), .C2(new_n755), .ZN(new_n1170));
  NOR4_X1   g0970(.A1(new_n1170), .A2(G41), .A3(new_n261), .A4(new_n1045), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n356), .A2(new_n758), .B1(new_n736), .B2(new_n230), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1172), .B1(G107), .B2(new_n772), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n1171), .B(new_n1173), .C1(new_n831), .C2(new_n750), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(new_n1174), .B(KEYINPUT58), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n740), .A2(new_n1114), .B1(new_n758), .B2(new_n1010), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1176), .B1(new_n817), .B2(new_n1117), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n748), .A2(G132), .B1(new_n754), .B2(G125), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n1177), .B(new_n1178), .C1(new_n326), .C2(new_n744), .ZN(new_n1179));
  XOR2_X1   g0979(.A(new_n1179), .B(KEYINPUT59), .Z(new_n1180));
  AOI21_X1  g0980(.A(G41), .B1(new_n828), .B2(G124), .ZN(new_n1181));
  AOI21_X1  g0981(.A(G33), .B1(new_n767), .B2(G159), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1180), .A2(new_n1181), .A3(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(G41), .B1(KEYINPUT3), .B2(G33), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n1175), .B(new_n1183), .C1(G50), .C2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n727), .B1(new_n1185), .B2(new_n842), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1168), .A2(new_n1169), .A3(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1167), .A2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1166), .A2(new_n1189), .ZN(G375));
  OR2_X1    g0990(.A1(new_n1091), .A2(new_n1079), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1191), .A2(new_n977), .A3(new_n1102), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n740), .A2(new_n831), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n741), .A2(new_n266), .B1(new_n758), .B2(new_n252), .ZN(new_n1194));
  AOI211_X1 g0994(.A(new_n1193), .B(new_n1194), .C1(G303), .C2(new_n828), .ZN(new_n1195));
  OAI22_X1  g0995(.A1(new_n824), .A2(new_n254), .B1(new_n755), .B2(new_n770), .ZN(new_n1196));
  NOR3_X1   g0996(.A1(new_n1196), .A2(new_n261), .A3(new_n1046), .ZN(new_n1197));
  OAI211_X1 g0997(.A(new_n1195), .B(new_n1197), .C1(new_n298), .C2(new_n736), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(G159), .A2(new_n817), .B1(new_n828), .B2(G128), .ZN(new_n1199));
  OAI221_X1 g0999(.A(new_n1199), .B1(new_n230), .B2(new_n736), .C1(new_n326), .C2(new_n758), .ZN(new_n1200));
  AOI211_X1 g1000(.A(new_n372), .B(new_n1200), .C1(G50), .C2(new_n745), .ZN(new_n1201));
  INV_X1    g1001(.A(KEYINPUT124), .ZN(new_n1202));
  OR2_X1    g1002(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n1117), .A2(new_n748), .B1(G132), .B2(new_n754), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1203), .A2(new_n1204), .A3(new_n1205), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n740), .A2(new_n1010), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1198), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1208), .A2(new_n842), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1209), .B1(G68), .B2(new_n845), .ZN(new_n1210));
  AOI211_X1 g1010(.A(new_n727), .B(new_n1210), .C1(new_n790), .C2(new_n896), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1211), .B1(new_n1091), .B2(new_n993), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1192), .A2(new_n1212), .ZN(G381));
  NAND2_X1  g1013(.A1(G378), .A2(KEYINPUT125), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT125), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1105), .A2(new_n1130), .A3(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1214), .A2(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1217), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(G375), .A2(new_n1218), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(G387), .A2(G381), .ZN(new_n1220));
  INV_X1    g1020(.A(G396), .ZN(new_n1221));
  NAND4_X1  g1021(.A1(new_n1023), .A2(new_n1221), .A3(new_n1024), .A4(new_n1054), .ZN(new_n1222));
  NOR3_X1   g1022(.A1(G390), .A2(new_n1222), .A3(G384), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1219), .A2(new_n1220), .A3(new_n1223), .ZN(G407));
  INV_X1    g1024(.A(G213), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1225), .B1(new_n1219), .B2(new_n670), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1226), .A2(G407), .ZN(G409));
  NAND2_X1  g1027(.A1(G393), .A2(G396), .ZN(new_n1228));
  AND2_X1   g1028(.A1(new_n1228), .A2(new_n1222), .ZN(new_n1229));
  AND3_X1   g1029(.A1(new_n994), .A2(new_n1020), .A3(G390), .ZN(new_n1230));
  AOI21_X1  g1030(.A(G390), .B1(new_n994), .B2(new_n1020), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1229), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(G390), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(G387), .A2(new_n1233), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n994), .A2(new_n1020), .A3(G390), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT126), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1236), .B1(new_n1228), .B2(new_n1222), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1234), .A2(new_n1235), .A3(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1231), .A2(new_n1236), .ZN(new_n1239));
  AND3_X1   g1039(.A1(new_n1232), .A2(new_n1238), .A3(new_n1239), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1240), .A2(KEYINPUT61), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1225), .A2(G343), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1166), .A2(G378), .A3(new_n1189), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1157), .A2(new_n977), .A3(new_n1159), .A4(new_n1160), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1187), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1144), .A2(new_n1156), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1245), .B1(new_n1246), .B2(new_n993), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(new_n1214), .A2(new_n1216), .B1(new_n1244), .B2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1248), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1242), .B1(new_n1243), .B2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT60), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n692), .B1(new_n1191), .B2(new_n1251), .ZN(new_n1252));
  OAI211_X1 g1052(.A(new_n1252), .B(new_n1102), .C1(new_n1251), .C2(new_n1191), .ZN(new_n1253));
  AOI21_X1  g1053(.A(G384), .B1(new_n1253), .B2(new_n1212), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1253), .A2(G384), .A3(new_n1212), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1250), .A2(KEYINPUT63), .A3(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT63), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1243), .A2(new_n1249), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1242), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1256), .ZN(new_n1264));
  OAI211_X1 g1064(.A(G2897), .B(new_n1242), .C1(new_n1264), .C2(new_n1254), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1242), .A2(G2897), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1255), .A2(new_n1256), .A3(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1265), .A2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1260), .B1(new_n1263), .B2(new_n1269), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1263), .A2(new_n1257), .ZN(new_n1271));
  OAI211_X1 g1071(.A(new_n1241), .B(new_n1259), .C1(new_n1270), .C2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT61), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1273), .B1(new_n1250), .B2(new_n1268), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1188), .B1(new_n1163), .B2(new_n1165), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1248), .B1(new_n1275), .B2(G378), .ZN(new_n1276));
  NOR4_X1   g1076(.A1(new_n1276), .A2(KEYINPUT62), .A3(new_n1242), .A4(new_n1257), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT62), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1278), .B1(new_n1250), .B2(new_n1258), .ZN(new_n1279));
  NOR3_X1   g1079(.A1(new_n1274), .A2(new_n1277), .A3(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1240), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1272), .B1(new_n1280), .B2(new_n1281), .ZN(G405));
  INV_X1    g1082(.A(new_n1243), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1275), .A2(new_n1218), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1258), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1285));
  OAI211_X1 g1085(.A(new_n1243), .B(new_n1257), .C1(new_n1275), .C2(new_n1218), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1285), .A2(new_n1240), .A3(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1287), .A2(KEYINPUT127), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1289), .A2(new_n1281), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT127), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1285), .A2(new_n1240), .A3(new_n1291), .A4(new_n1286), .ZN(new_n1292));
  AND3_X1   g1092(.A1(new_n1288), .A2(new_n1290), .A3(new_n1292), .ZN(G402));
endmodule


