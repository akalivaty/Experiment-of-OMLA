//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 0 0 0 0 0 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 1 0 1 0 0 1 1 1 1 0 1 0 1 1 0 1 0 1 1 0 1 0 0 0 0 0 0 0 1 1 1 0 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:17 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n450, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n561, new_n563, new_n564, new_n565,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n581,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n626, new_n627, new_n628, new_n631, new_n632,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n836,
    new_n837, new_n838, new_n839, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1163, new_n1164;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT64), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  XOR2_X1   g031(.A(G325), .B(KEYINPUT65), .Z(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT66), .Z(new_n459));
  INV_X1    g034(.A(G567), .ZN(new_n460));
  OAI21_X1  g035(.A(new_n459), .B1(new_n460), .B2(new_n454), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  NAND4_X1  g042(.A1(new_n464), .A2(new_n466), .A3(G137), .A4(new_n467), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n463), .A2(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G101), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  AND3_X1   g046(.A1(KEYINPUT67), .A2(G113), .A3(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(KEYINPUT67), .B1(G113), .B2(G2104), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n464), .A2(new_n466), .A3(G125), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n471), .B1(G2105), .B2(new_n476), .ZN(G160));
  NAND2_X1  g052(.A1(new_n464), .A2(new_n466), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n478), .A2(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G136), .ZN(new_n480));
  OR2_X1    g055(.A1(new_n480), .A2(KEYINPUT68), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n480), .A2(KEYINPUT68), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n478), .A2(new_n467), .ZN(new_n483));
  AOI22_X1  g058(.A1(new_n481), .A2(new_n482), .B1(G124), .B2(new_n483), .ZN(new_n484));
  OR2_X1    g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G112), .C2(new_n467), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  NAND4_X1  g063(.A1(new_n464), .A2(new_n466), .A3(G138), .A4(new_n467), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT69), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  XNOR2_X1  g066(.A(KEYINPUT3), .B(G2104), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n492), .A2(KEYINPUT69), .A3(G138), .A4(new_n467), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n491), .A2(new_n493), .A3(KEYINPUT4), .ZN(new_n494));
  AND2_X1   g069(.A1(new_n469), .A2(G102), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n464), .A2(new_n466), .A3(G126), .ZN(new_n496));
  NAND2_X1  g071(.A1(G114), .A2(G2104), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n495), .B1(new_n498), .B2(G2105), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n489), .A2(new_n490), .A3(new_n500), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n494), .A2(new_n499), .A3(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(G164));
  INV_X1    g078(.A(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(KEYINPUT5), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT5), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(G62), .ZN(new_n509));
  OAI21_X1  g084(.A(KEYINPUT71), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(G75), .A2(G543), .ZN(new_n511));
  XNOR2_X1  g086(.A(KEYINPUT5), .B(G543), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT71), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n512), .A2(new_n513), .A3(G62), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n510), .A2(new_n511), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G651), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT72), .ZN(new_n517));
  XNOR2_X1  g092(.A(new_n516), .B(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(G651), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(KEYINPUT6), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT6), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G651), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n523), .A2(new_n504), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G50), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT70), .ZN(new_n526));
  NOR3_X1   g101(.A1(new_n523), .A2(new_n508), .A3(new_n526), .ZN(new_n527));
  XNOR2_X1  g102(.A(KEYINPUT6), .B(G651), .ZN(new_n528));
  AOI21_X1  g103(.A(KEYINPUT70), .B1(new_n528), .B2(new_n512), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(G88), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n518), .A2(new_n525), .A3(new_n531), .ZN(G303));
  INV_X1    g107(.A(G303), .ZN(G166));
  AND2_X1   g108(.A1(new_n530), .A2(G89), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT7), .ZN(new_n535));
  NAND2_X1  g110(.A1(G76), .A2(G543), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n535), .B1(new_n536), .B2(new_n519), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n536), .A2(new_n535), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n538), .B1(new_n512), .B2(G63), .ZN(new_n539));
  INV_X1    g114(.A(new_n524), .ZN(new_n540));
  XNOR2_X1  g115(.A(KEYINPUT73), .B(G51), .ZN(new_n541));
  OAI221_X1 g116(.A(new_n537), .B1(new_n539), .B2(new_n519), .C1(new_n540), .C2(new_n541), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n534), .A2(new_n542), .ZN(G168));
  NAND2_X1  g118(.A1(new_n530), .A2(G90), .ZN(new_n544));
  NAND2_X1  g119(.A1(G77), .A2(G543), .ZN(new_n545));
  INV_X1    g120(.A(G64), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n545), .B1(new_n508), .B2(new_n546), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n547), .A2(G651), .B1(new_n524), .B2(G52), .ZN(new_n548));
  AND2_X1   g123(.A1(new_n544), .A2(new_n548), .ZN(G171));
  NAND2_X1  g124(.A1(G68), .A2(G543), .ZN(new_n550));
  INV_X1    g125(.A(G56), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n550), .B1(new_n508), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G651), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT74), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n553), .B(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n530), .A2(G81), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n524), .A2(G43), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n555), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT75), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G860), .ZN(G153));
  AND3_X1   g135(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G36), .ZN(G176));
  XOR2_X1   g137(.A(KEYINPUT76), .B(KEYINPUT8), .Z(new_n563));
  NAND2_X1  g138(.A1(G1), .A2(G3), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n563), .B(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n561), .A2(new_n565), .ZN(G188));
  INV_X1    g141(.A(KEYINPUT77), .ZN(new_n567));
  NOR3_X1   g142(.A1(new_n527), .A2(new_n529), .A3(new_n567), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n526), .B1(new_n523), .B2(new_n508), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n528), .A2(new_n512), .A3(KEYINPUT70), .ZN(new_n570));
  AOI21_X1  g145(.A(KEYINPUT77), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  OAI21_X1  g146(.A(G91), .B1(new_n568), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n512), .A2(G65), .ZN(new_n573));
  NAND2_X1  g148(.A1(G78), .A2(G543), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n519), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n524), .A2(G53), .ZN(new_n577));
  XNOR2_X1  g152(.A(new_n577), .B(KEYINPUT9), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n572), .A2(new_n576), .A3(new_n578), .ZN(new_n579));
  XNOR2_X1  g154(.A(new_n579), .B(KEYINPUT78), .ZN(G299));
  XOR2_X1   g155(.A(G171), .B(KEYINPUT79), .Z(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(G301));
  INV_X1    g157(.A(G168), .ZN(G286));
  OAI21_X1  g158(.A(new_n567), .B1(new_n527), .B2(new_n529), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n569), .A2(KEYINPUT77), .A3(new_n570), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n586), .A2(G87), .ZN(new_n587));
  OR2_X1    g162(.A1(new_n512), .A2(G74), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n588), .A2(G651), .B1(new_n524), .B2(G49), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n587), .A2(new_n589), .ZN(G288));
  INV_X1    g165(.A(KEYINPUT80), .ZN(new_n591));
  INV_X1    g166(.A(G61), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n508), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(G73), .A2(G543), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n512), .A2(KEYINPUT80), .A3(G61), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n596), .A2(G651), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n598), .A2(KEYINPUT81), .B1(G48), .B2(new_n524), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n586), .A2(G86), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT81), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n597), .A2(new_n601), .ZN(new_n602));
  AND3_X1   g177(.A1(new_n599), .A2(new_n600), .A3(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(G305));
  XNOR2_X1  g179(.A(KEYINPUT82), .B(G85), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n530), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(G72), .A2(G543), .ZN(new_n607));
  INV_X1    g182(.A(G60), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n508), .B2(new_n608), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n609), .A2(G651), .B1(new_n524), .B2(G47), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n606), .A2(new_n610), .ZN(G290));
  NAND2_X1  g186(.A1(new_n512), .A2(G66), .ZN(new_n612));
  NAND2_X1  g187(.A1(G79), .A2(G543), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n519), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n586), .A2(G92), .ZN(new_n615));
  INV_X1    g190(.A(KEYINPUT10), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n586), .A2(KEYINPUT10), .A3(G92), .ZN(new_n618));
  AOI21_X1  g193(.A(new_n614), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n524), .A2(G54), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g196(.A(G868), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(new_n622), .B2(new_n581), .ZN(G284));
  OAI21_X1  g199(.A(new_n623), .B1(new_n622), .B2(new_n581), .ZN(G321));
  OAI21_X1  g200(.A(KEYINPUT83), .B1(G168), .B2(new_n622), .ZN(new_n626));
  OR3_X1    g201(.A1(G168), .A2(KEYINPUT83), .A3(new_n622), .ZN(new_n627));
  INV_X1    g202(.A(G299), .ZN(new_n628));
  OAI211_X1 g203(.A(new_n626), .B(new_n627), .C1(new_n628), .C2(G868), .ZN(G297));
  OAI211_X1 g204(.A(new_n626), .B(new_n627), .C1(new_n628), .C2(G868), .ZN(G280));
  INV_X1    g205(.A(new_n621), .ZN(new_n631));
  INV_X1    g206(.A(G559), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n631), .B1(new_n632), .B2(G860), .ZN(G148));
  NOR2_X1   g208(.A1(new_n621), .A2(G559), .ZN(new_n634));
  NOR2_X1   g209(.A1(new_n634), .A2(new_n622), .ZN(new_n635));
  INV_X1    g210(.A(new_n635), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n636), .B1(G868), .B2(new_n559), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n637), .A2(KEYINPUT84), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n638), .B1(KEYINPUT84), .B2(new_n635), .ZN(G323));
  XNOR2_X1  g214(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g215(.A1(new_n492), .A2(new_n469), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT12), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT13), .ZN(new_n643));
  INV_X1    g218(.A(G2100), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n644), .A2(KEYINPUT85), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n643), .B(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n479), .A2(G135), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n483), .A2(G123), .ZN(new_n648));
  NOR2_X1   g223(.A1(G99), .A2(G2105), .ZN(new_n649));
  OAI21_X1  g224(.A(G2104), .B1(new_n467), .B2(G111), .ZN(new_n650));
  OAI211_X1 g225(.A(new_n647), .B(new_n648), .C1(new_n649), .C2(new_n650), .ZN(new_n651));
  INV_X1    g226(.A(G2096), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  OAI211_X1 g228(.A(new_n646), .B(new_n653), .C1(KEYINPUT85), .C2(new_n644), .ZN(G156));
  XNOR2_X1  g229(.A(G2451), .B(G2454), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT16), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2443), .B(G2446), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1341), .B(G1348), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n658), .B(new_n659), .Z(new_n660));
  XNOR2_X1  g235(.A(KEYINPUT15), .B(G2430), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(G2435), .ZN(new_n662));
  XOR2_X1   g237(.A(G2427), .B(G2438), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n664), .A2(KEYINPUT14), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n660), .B(new_n665), .ZN(new_n666));
  AND2_X1   g241(.A1(new_n666), .A2(G14), .ZN(G401));
  XOR2_X1   g242(.A(G2084), .B(G2090), .Z(new_n668));
  XNOR2_X1  g243(.A(G2067), .B(G2678), .ZN(new_n669));
  XNOR2_X1  g244(.A(G2072), .B(G2078), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n668), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n671), .B(KEYINPUT18), .Z(new_n672));
  XOR2_X1   g247(.A(new_n669), .B(KEYINPUT86), .Z(new_n673));
  OAI21_X1  g248(.A(KEYINPUT17), .B1(new_n673), .B2(new_n668), .ZN(new_n674));
  XOR2_X1   g249(.A(new_n674), .B(new_n670), .Z(new_n675));
  AND2_X1   g250(.A1(new_n673), .A2(new_n668), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n672), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(new_n652), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(G2100), .ZN(G227));
  XNOR2_X1  g254(.A(G1956), .B(G2474), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT87), .ZN(new_n681));
  XOR2_X1   g256(.A(G1961), .B(G1966), .Z(new_n682));
  NAND2_X1  g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1971), .B(G1976), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT19), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT88), .ZN(new_n687));
  OR2_X1    g262(.A1(new_n687), .A2(KEYINPUT20), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n687), .A2(KEYINPUT20), .ZN(new_n689));
  INV_X1    g264(.A(new_n683), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n681), .A2(new_n682), .ZN(new_n691));
  INV_X1    g266(.A(new_n685), .ZN(new_n692));
  OR3_X1    g267(.A1(new_n690), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n691), .A2(new_n692), .ZN(new_n694));
  NAND4_X1  g269(.A1(new_n688), .A2(new_n689), .A3(new_n693), .A4(new_n694), .ZN(new_n695));
  XOR2_X1   g270(.A(G1991), .B(G1996), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1981), .B(G1986), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(G229));
  NAND2_X1  g277(.A1(G168), .A2(G16), .ZN(new_n703));
  OAI211_X1 g278(.A(new_n703), .B(KEYINPUT101), .C1(G16), .C2(G21), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(KEYINPUT101), .B2(new_n703), .ZN(new_n705));
  OR2_X1    g280(.A1(new_n705), .A2(G1966), .ZN(new_n706));
  INV_X1    g281(.A(G29), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n707), .A2(G27), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(G164), .B2(new_n707), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(G2078), .ZN(new_n710));
  AND2_X1   g285(.A1(new_n707), .A2(G35), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n711), .B1(new_n487), .B2(G29), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT29), .ZN(new_n713));
  INV_X1    g288(.A(G2090), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT31), .B(G11), .ZN(new_n716));
  INV_X1    g291(.A(KEYINPUT30), .ZN(new_n717));
  OR2_X1    g292(.A1(new_n717), .A2(G28), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n717), .A2(G28), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n718), .A2(new_n719), .A3(new_n707), .ZN(new_n720));
  OAI211_X1 g295(.A(new_n716), .B(new_n720), .C1(new_n651), .C2(new_n707), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT102), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n479), .A2(G141), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n483), .A2(G129), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n469), .A2(G105), .ZN(new_n725));
  NAND3_X1  g300(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n726));
  XOR2_X1   g301(.A(new_n726), .B(KEYINPUT26), .Z(new_n727));
  NAND4_X1  g302(.A1(new_n723), .A2(new_n724), .A3(new_n725), .A4(new_n727), .ZN(new_n728));
  MUX2_X1   g303(.A(G32), .B(new_n728), .S(G29), .Z(new_n729));
  XOR2_X1   g304(.A(KEYINPUT27), .B(G1996), .Z(new_n730));
  AOI21_X1  g305(.A(new_n722), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(G16), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n732), .A2(G5), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(G171), .B2(new_n732), .ZN(new_n734));
  INV_X1    g309(.A(G1961), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n734), .B(new_n735), .ZN(new_n736));
  AND2_X1   g311(.A1(new_n731), .A2(new_n736), .ZN(new_n737));
  OR2_X1    g312(.A1(KEYINPUT24), .A2(G34), .ZN(new_n738));
  NAND2_X1  g313(.A1(KEYINPUT24), .A2(G34), .ZN(new_n739));
  NAND3_X1  g314(.A1(new_n738), .A2(new_n707), .A3(new_n739), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(G160), .B2(new_n707), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n741), .A2(G2084), .ZN(new_n742));
  XNOR2_X1  g317(.A(KEYINPUT91), .B(G16), .ZN(new_n743));
  INV_X1    g318(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n744), .A2(G19), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(new_n559), .B2(new_n744), .ZN(new_n746));
  XNOR2_X1  g321(.A(KEYINPUT94), .B(G1341), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND4_X1  g323(.A1(new_n715), .A2(new_n737), .A3(new_n742), .A4(new_n748), .ZN(new_n749));
  XNOR2_X1  g324(.A(KEYINPUT97), .B(KEYINPUT28), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT98), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n707), .A2(G26), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n483), .A2(G128), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT96), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n479), .A2(G140), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT95), .ZN(new_n757));
  OR2_X1    g332(.A1(G104), .A2(G2105), .ZN(new_n758));
  OAI211_X1 g333(.A(new_n758), .B(G2104), .C1(G116), .C2(new_n467), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n755), .A2(new_n757), .A3(new_n759), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n753), .B1(new_n760), .B2(G29), .ZN(new_n761));
  XOR2_X1   g336(.A(KEYINPUT99), .B(G2067), .Z(new_n762));
  XNOR2_X1  g337(.A(new_n761), .B(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n705), .A2(G1966), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(new_n746), .B2(new_n747), .ZN(new_n765));
  OR4_X1    g340(.A1(new_n710), .A2(new_n749), .A3(new_n763), .A4(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n469), .A2(G103), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT25), .Z(new_n768));
  NAND2_X1  g343(.A1(new_n479), .A2(G139), .ZN(new_n769));
  AOI22_X1  g344(.A1(new_n492), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n770));
  OAI211_X1 g345(.A(new_n768), .B(new_n769), .C1(new_n467), .C2(new_n770), .ZN(new_n771));
  MUX2_X1   g346(.A(G33), .B(new_n771), .S(G29), .Z(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(G2072), .Z(new_n773));
  NAND2_X1  g348(.A1(new_n741), .A2(G2084), .ZN(new_n774));
  OAI211_X1 g349(.A(new_n773), .B(new_n774), .C1(new_n729), .C2(new_n730), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT100), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n713), .A2(new_n714), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT103), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n732), .A2(G4), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(new_n631), .B2(new_n732), .ZN(new_n781));
  XNOR2_X1  g356(.A(KEYINPUT93), .B(G1348), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n781), .B(new_n782), .Z(new_n783));
  NAND3_X1  g358(.A1(new_n744), .A2(KEYINPUT23), .A3(G20), .ZN(new_n784));
  INV_X1    g359(.A(KEYINPUT23), .ZN(new_n785));
  INV_X1    g360(.A(G20), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n785), .B1(new_n743), .B2(new_n786), .ZN(new_n787));
  OAI211_X1 g362(.A(new_n784), .B(new_n787), .C1(new_n628), .C2(new_n732), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(G1956), .ZN(new_n789));
  NOR4_X1   g364(.A1(new_n766), .A2(new_n779), .A3(new_n783), .A4(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n732), .A2(G23), .ZN(new_n791));
  AND2_X1   g366(.A1(new_n587), .A2(new_n589), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n791), .B1(new_n792), .B2(new_n732), .ZN(new_n793));
  OR2_X1    g368(.A1(new_n793), .A2(KEYINPUT33), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n793), .A2(KEYINPUT33), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  INV_X1    g371(.A(G1976), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n794), .A2(G1976), .A3(new_n795), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n732), .A2(G6), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(new_n603), .B2(new_n732), .ZN(new_n802));
  XOR2_X1   g377(.A(KEYINPUT32), .B(G1981), .Z(new_n803));
  INV_X1    g378(.A(new_n803), .ZN(new_n804));
  OR2_X1    g379(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  OR2_X1    g380(.A1(new_n743), .A2(G22), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(G303), .B2(new_n744), .ZN(new_n807));
  INV_X1    g382(.A(G1971), .ZN(new_n808));
  OR2_X1    g383(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n807), .A2(new_n808), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n802), .A2(new_n804), .ZN(new_n811));
  NAND4_X1  g386(.A1(new_n805), .A2(new_n809), .A3(new_n810), .A4(new_n811), .ZN(new_n812));
  OR3_X1    g387(.A1(new_n800), .A2(KEYINPUT34), .A3(new_n812), .ZN(new_n813));
  OAI21_X1  g388(.A(KEYINPUT34), .B1(new_n800), .B2(new_n812), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n744), .A2(G24), .ZN(new_n815));
  INV_X1    g390(.A(G290), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n815), .B1(new_n816), .B2(new_n744), .ZN(new_n817));
  XNOR2_X1  g392(.A(KEYINPUT92), .B(G1986), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  NOR2_X1   g394(.A1(G25), .A2(G29), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n479), .A2(G131), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT89), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n483), .A2(G119), .ZN(new_n823));
  NOR2_X1   g398(.A1(G95), .A2(G2105), .ZN(new_n824));
  OAI21_X1  g399(.A(G2104), .B1(new_n467), .B2(G107), .ZN(new_n825));
  OAI211_X1 g400(.A(new_n822), .B(new_n823), .C1(new_n824), .C2(new_n825), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT90), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n820), .B1(new_n827), .B2(G29), .ZN(new_n828));
  XOR2_X1   g403(.A(KEYINPUT35), .B(G1991), .Z(new_n829));
  XNOR2_X1  g404(.A(new_n828), .B(new_n829), .ZN(new_n830));
  NAND4_X1  g405(.A1(new_n813), .A2(new_n814), .A3(new_n819), .A4(new_n830), .ZN(new_n831));
  AND2_X1   g406(.A1(new_n831), .A2(KEYINPUT36), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n831), .A2(KEYINPUT36), .ZN(new_n833));
  OAI211_X1 g408(.A(new_n706), .B(new_n790), .C1(new_n832), .C2(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(new_n834), .ZN(G311));
  NAND2_X1  g410(.A1(new_n834), .A2(KEYINPUT104), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n831), .B(KEYINPUT36), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT104), .ZN(new_n838));
  NAND4_X1  g413(.A1(new_n837), .A2(new_n838), .A3(new_n706), .A4(new_n790), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n836), .A2(new_n839), .ZN(G150));
  NAND2_X1  g415(.A1(new_n530), .A2(G93), .ZN(new_n841));
  NAND2_X1  g416(.A1(G80), .A2(G543), .ZN(new_n842));
  INV_X1    g417(.A(G67), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n842), .B1(new_n508), .B2(new_n843), .ZN(new_n844));
  XOR2_X1   g419(.A(KEYINPUT105), .B(G55), .Z(new_n845));
  AOI22_X1  g420(.A1(new_n844), .A2(G651), .B1(new_n524), .B2(new_n845), .ZN(new_n846));
  AND2_X1   g421(.A1(new_n841), .A2(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(G860), .ZN(new_n849));
  XOR2_X1   g424(.A(new_n849), .B(KEYINPUT37), .Z(new_n850));
  NOR2_X1   g425(.A1(new_n621), .A2(new_n632), .ZN(new_n851));
  XNOR2_X1  g426(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n851), .B(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n558), .A2(new_n847), .ZN(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n855), .B1(new_n559), .B2(new_n848), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n853), .B(new_n856), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n850), .B1(new_n857), .B2(G860), .ZN(G145));
  XNOR2_X1  g433(.A(new_n651), .B(G160), .ZN(new_n859));
  XOR2_X1   g434(.A(new_n859), .B(new_n826), .Z(new_n860));
  NAND2_X1  g435(.A1(new_n479), .A2(G142), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n483), .A2(G130), .ZN(new_n862));
  NOR2_X1   g437(.A1(G106), .A2(G2105), .ZN(new_n863));
  OAI21_X1  g438(.A(G2104), .B1(new_n467), .B2(G118), .ZN(new_n864));
  OAI211_X1 g439(.A(new_n861), .B(new_n862), .C1(new_n863), .C2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(new_n642), .ZN(new_n866));
  XOR2_X1   g441(.A(new_n860), .B(new_n866), .Z(new_n867));
  XNOR2_X1  g442(.A(new_n760), .B(new_n502), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(new_n728), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n771), .B(KEYINPUT106), .ZN(new_n870));
  OR2_X1    g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT106), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n869), .B1(new_n872), .B2(new_n771), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n871), .A2(new_n487), .A3(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n487), .B1(new_n871), .B2(new_n873), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n867), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n876), .ZN(new_n878));
  INV_X1    g453(.A(new_n867), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n878), .A2(new_n874), .A3(new_n879), .ZN(new_n880));
  XOR2_X1   g455(.A(KEYINPUT107), .B(G37), .Z(new_n881));
  NAND3_X1  g456(.A1(new_n877), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g458(.A(new_n634), .ZN(new_n884));
  OR2_X1    g459(.A1(new_n884), .A2(new_n856), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n856), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n628), .A2(new_n631), .ZN(new_n888));
  NAND2_X1  g463(.A1(G299), .A2(new_n621), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n887), .A2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT41), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n890), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n888), .A2(new_n889), .A3(KEYINPUT41), .ZN(new_n895));
  NAND4_X1  g470(.A1(new_n894), .A2(new_n885), .A3(new_n886), .A4(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n892), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(G303), .A2(new_n792), .ZN(new_n898));
  NAND4_X1  g473(.A1(G288), .A2(new_n518), .A3(new_n525), .A4(new_n531), .ZN(new_n899));
  NAND3_X1  g474(.A1(G305), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(G305), .B1(new_n898), .B2(new_n899), .ZN(new_n902));
  OAI21_X1  g477(.A(G290), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n898), .A2(new_n899), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(new_n603), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n905), .A2(new_n816), .A3(new_n900), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n903), .A2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT108), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(KEYINPUT42), .ZN(new_n909));
  OR2_X1    g484(.A1(new_n908), .A2(KEYINPUT42), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n907), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  NAND4_X1  g486(.A1(new_n903), .A2(new_n906), .A3(new_n908), .A4(KEYINPUT42), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n897), .A2(new_n913), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n892), .A2(new_n911), .A3(new_n896), .A4(new_n912), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n914), .A2(KEYINPUT109), .A3(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT109), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n897), .A2(new_n913), .A3(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n622), .B1(new_n916), .B2(new_n918), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n848), .A2(G868), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n919), .A2(new_n920), .ZN(G295));
  INV_X1    g496(.A(KEYINPUT110), .ZN(new_n922));
  INV_X1    g497(.A(new_n920), .ZN(new_n923));
  AND2_X1   g498(.A1(new_n916), .A2(new_n918), .ZN(new_n924));
  OAI211_X1 g499(.A(new_n922), .B(new_n923), .C1(new_n924), .C2(new_n622), .ZN(new_n925));
  OAI21_X1  g500(.A(KEYINPUT110), .B1(new_n919), .B2(new_n920), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(G331));
  INV_X1    g502(.A(KEYINPUT44), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n894), .A2(new_n895), .ZN(new_n929));
  INV_X1    g504(.A(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(G286), .A2(G171), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n931), .B1(new_n581), .B2(G286), .ZN(new_n932));
  OR2_X1    g507(.A1(new_n932), .A2(new_n856), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n856), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n930), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n891), .B1(new_n933), .B2(new_n934), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n907), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(new_n935), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n937), .B1(new_n929), .B2(new_n939), .ZN(new_n940));
  XNOR2_X1  g515(.A(new_n907), .B(KEYINPUT111), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT43), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n938), .A2(new_n942), .A3(new_n943), .A4(new_n881), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(G37), .B1(new_n940), .B2(new_n941), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n943), .B1(new_n946), .B2(new_n938), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n928), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  AND4_X1   g523(.A1(KEYINPUT43), .A2(new_n938), .A3(new_n881), .A4(new_n942), .ZN(new_n949));
  AOI21_X1  g524(.A(KEYINPUT43), .B1(new_n946), .B2(new_n938), .ZN(new_n950));
  OAI21_X1  g525(.A(KEYINPUT44), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n948), .A2(new_n951), .ZN(G397));
  INV_X1    g527(.A(G1384), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n502), .A2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT45), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n476), .A2(G2105), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n958), .A2(G40), .A3(new_n470), .A4(new_n468), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(KEYINPUT112), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT112), .ZN(new_n961));
  NAND3_X1  g536(.A1(G160), .A2(new_n961), .A3(G40), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n957), .A2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(new_n964), .ZN(new_n965));
  XNOR2_X1  g540(.A(new_n760), .B(G2067), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n965), .B1(new_n966), .B2(new_n728), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT46), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n968), .B1(new_n964), .B2(G1996), .ZN(new_n969));
  INV_X1    g544(.A(G1996), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n965), .A2(KEYINPUT46), .A3(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n967), .A2(new_n969), .A3(new_n971), .ZN(new_n972));
  XNOR2_X1  g547(.A(new_n972), .B(KEYINPUT126), .ZN(new_n973));
  XNOR2_X1  g548(.A(new_n973), .B(KEYINPUT47), .ZN(new_n974));
  XNOR2_X1  g549(.A(new_n728), .B(G1996), .ZN(new_n975));
  OR2_X1    g550(.A1(new_n966), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n827), .A2(new_n829), .ZN(new_n977));
  OAI22_X1  g552(.A1(new_n976), .A2(new_n977), .B1(G2067), .B2(new_n760), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(new_n965), .ZN(new_n979));
  NOR3_X1   g554(.A1(new_n964), .A2(G1986), .A3(G290), .ZN(new_n980));
  XNOR2_X1  g555(.A(KEYINPUT127), .B(KEYINPUT48), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n980), .B(new_n981), .ZN(new_n982));
  XOR2_X1   g557(.A(new_n826), .B(new_n829), .Z(new_n983));
  NOR2_X1   g558(.A1(new_n976), .A2(new_n983), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n982), .B1(new_n964), .B2(new_n984), .ZN(new_n985));
  AND3_X1   g560(.A1(new_n974), .A2(new_n979), .A3(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(KEYINPUT114), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT55), .ZN(new_n989));
  INV_X1    g564(.A(G8), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n989), .B1(G166), .B2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT114), .ZN(new_n992));
  NAND4_X1  g567(.A1(G303), .A2(new_n992), .A3(KEYINPUT55), .A4(G8), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n988), .A2(new_n991), .A3(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n502), .A2(KEYINPUT45), .A3(new_n953), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n956), .A2(new_n963), .A3(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT113), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  AOI22_X1  g573(.A1(new_n954), .A2(new_n955), .B1(new_n960), .B2(new_n962), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n999), .A2(KEYINPUT113), .A3(new_n995), .ZN(new_n1000));
  AOI21_X1  g575(.A(G1971), .B1(new_n998), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT50), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n954), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n502), .A2(KEYINPUT50), .A3(new_n953), .ZN(new_n1004));
  AOI22_X1  g579(.A1(new_n1003), .A2(new_n1004), .B1(new_n960), .B2(new_n962), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(new_n714), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1006), .ZN(new_n1007));
  OAI211_X1 g582(.A(new_n994), .B(G8), .C1(new_n1001), .C2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n963), .A2(new_n953), .A3(new_n502), .ZN(new_n1010));
  OAI211_X1 g585(.A(new_n1010), .B(G8), .C1(G288), .C2(new_n797), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT52), .ZN(new_n1012));
  OR2_X1    g587(.A1(new_n1012), .A2(KEYINPUT115), .ZN(new_n1013));
  OR2_X1    g588(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g589(.A1(G288), .A2(new_n1012), .A3(new_n797), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1014), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(G1981), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n599), .A2(new_n1018), .A3(new_n600), .A4(new_n602), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n530), .A2(G86), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n524), .A2(G48), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1020), .A2(new_n597), .A3(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(G1981), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1019), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT49), .ZN(new_n1025));
  OAI21_X1  g600(.A(KEYINPUT116), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1027));
  AND2_X1   g602(.A1(new_n1010), .A2(G8), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT116), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1019), .A2(new_n1029), .A3(KEYINPUT49), .A4(new_n1023), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1026), .A2(new_n1027), .A3(new_n1028), .A4(new_n1030), .ZN(new_n1031));
  AND2_X1   g606(.A1(new_n1017), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1009), .A2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1031), .A2(new_n797), .A3(new_n792), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(new_n1019), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT117), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1034), .A2(KEYINPUT117), .A3(new_n1019), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1037), .A2(new_n1028), .A3(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(G8), .B1(new_n1001), .B2(new_n1007), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1040), .A2(new_n991), .A3(new_n988), .A4(new_n993), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1032), .A2(new_n1008), .A3(new_n1041), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1042), .A2(G286), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n502), .A2(KEYINPUT118), .A3(KEYINPUT45), .A4(new_n953), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT118), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n995), .A2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n999), .A2(new_n1044), .A3(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(G1966), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT119), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1004), .ZN(new_n1052));
  AOI21_X1  g627(.A(KEYINPUT50), .B1(new_n502), .B2(new_n953), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n963), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  OR2_X1    g629(.A1(new_n1054), .A2(G2084), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1047), .A2(KEYINPUT119), .A3(new_n1048), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1051), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(G8), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(KEYINPUT63), .B1(new_n1043), .B2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT63), .ZN(new_n1061));
  NOR4_X1   g636(.A1(new_n1042), .A2(new_n1061), .A3(G286), .A4(new_n1058), .ZN(new_n1062));
  OAI211_X1 g637(.A(new_n1033), .B(new_n1039), .C1(new_n1060), .C2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n572), .A2(KEYINPUT120), .A3(new_n576), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT57), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n579), .A2(new_n1064), .A3(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n575), .B1(new_n586), .B2(G91), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n1067), .B(new_n578), .C1(KEYINPUT120), .C2(KEYINPUT57), .ZN(new_n1068));
  AND2_X1   g643(.A1(new_n1066), .A2(new_n1068), .ZN(new_n1069));
  XNOR2_X1  g644(.A(KEYINPUT56), .B(G2072), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n956), .A2(new_n963), .A3(new_n995), .A4(new_n1070), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1071), .B1(new_n1005), .B2(G1956), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1069), .A2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT61), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1066), .A2(new_n1068), .ZN(new_n1075));
  INV_X1    g650(.A(G1956), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1054), .A2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1075), .A2(new_n1077), .A3(new_n1071), .ZN(new_n1078));
  AND3_X1   g653(.A1(new_n1073), .A2(new_n1074), .A3(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1074), .B1(new_n1073), .B2(new_n1078), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n956), .A2(new_n963), .A3(new_n970), .A4(new_n995), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT122), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n999), .A2(KEYINPUT122), .A3(new_n970), .A4(new_n995), .ZN(new_n1084));
  XOR2_X1   g659(.A(KEYINPUT58), .B(G1341), .Z(new_n1085));
  NAND2_X1  g660(.A1(new_n1010), .A2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1083), .A2(new_n1084), .A3(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT59), .ZN(new_n1088));
  AND3_X1   g663(.A1(new_n1087), .A2(new_n1088), .A3(new_n559), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1088), .B1(new_n1087), .B2(new_n559), .ZN(new_n1090));
  OAI22_X1  g665(.A1(new_n1079), .A2(new_n1080), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(KEYINPUT123), .ZN(new_n1092));
  OAI22_X1  g667(.A1(new_n1005), .A2(G1348), .B1(G2067), .B2(new_n1010), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(KEYINPUT121), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT121), .ZN(new_n1095));
  OAI221_X1 g670(.A(new_n1095), .B1(new_n1010), .B2(G2067), .C1(new_n1005), .C2(G1348), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n621), .B1(new_n1097), .B2(KEYINPUT60), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT60), .ZN(new_n1099));
  AOI211_X1 g674(.A(new_n1099), .B(new_n631), .C1(new_n1094), .C2(new_n1096), .ZN(new_n1100));
  OAI22_X1  g675(.A1(new_n1098), .A2(new_n1100), .B1(KEYINPUT60), .B2(new_n1097), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT123), .ZN(new_n1102));
  OAI221_X1 g677(.A(new_n1102), .B1(new_n1089), .B2(new_n1090), .C1(new_n1079), .C2(new_n1080), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1092), .A2(new_n1101), .A3(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1097), .ZN(new_n1105));
  AND2_X1   g680(.A1(new_n1078), .A2(new_n631), .ZN(new_n1106));
  AOI22_X1  g681(.A1(new_n1105), .A2(new_n1106), .B1(new_n1069), .B2(new_n1072), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1104), .A2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(G2078), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n998), .A2(new_n1109), .A3(new_n1000), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT124), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT53), .ZN(new_n1112));
  AND3_X1   g687(.A1(new_n1110), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1111), .B1(new_n1110), .B2(new_n1112), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1005), .A2(G1961), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT125), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1118), .B1(new_n957), .B2(new_n959), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n956), .A2(KEYINPUT125), .A3(G40), .A4(G160), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1112), .A2(G2078), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1119), .A2(new_n995), .A3(new_n1120), .A4(new_n1121), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1115), .A2(G301), .A3(new_n1117), .A4(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(KEYINPUT124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1110), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1126));
  NOR3_X1   g701(.A1(new_n1047), .A2(new_n1112), .A3(G2078), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1127), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1125), .A2(new_n1117), .A3(new_n1126), .A4(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(new_n581), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT54), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1123), .A2(new_n1130), .A3(new_n1131), .ZN(new_n1132));
  NOR4_X1   g707(.A1(new_n1113), .A2(new_n1114), .A3(new_n1116), .A4(new_n1127), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1125), .A2(new_n1117), .A3(new_n1126), .A4(new_n1122), .ZN(new_n1134));
  AOI22_X1  g709(.A1(new_n1133), .A2(G301), .B1(G171), .B2(new_n1134), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1132), .B1(new_n1135), .B2(new_n1131), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT51), .ZN(new_n1137));
  NOR2_X1   g712(.A1(G168), .A2(new_n990), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1138), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1058), .A2(new_n1137), .A3(new_n1139), .ZN(new_n1140));
  OAI211_X1 g715(.A(KEYINPUT51), .B(G8), .C1(new_n1057), .C2(G286), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1057), .A2(new_n1138), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1108), .A2(new_n1136), .A3(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1144), .A2(KEYINPUT62), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT62), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1142), .A2(new_n1147), .A3(new_n1143), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1146), .A2(new_n581), .A3(new_n1129), .A4(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1145), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1042), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1063), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  XOR2_X1   g727(.A(G290), .B(G1986), .Z(new_n1153));
  AOI21_X1  g728(.A(new_n964), .B1(new_n984), .B2(new_n1153), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n986), .B1(new_n1152), .B2(new_n1154), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g730(.A1(G227), .A2(G401), .ZN(new_n1157));
  NAND2_X1  g731(.A1(new_n882), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g732(.A1(new_n701), .A2(G319), .ZN(new_n1159));
  NAND2_X1  g733(.A1(new_n946), .A2(new_n938), .ZN(new_n1160));
  NAND2_X1  g734(.A1(new_n1160), .A2(KEYINPUT43), .ZN(new_n1161));
  AOI211_X1 g735(.A(new_n1158), .B(new_n1159), .C1(new_n1161), .C2(new_n944), .ZN(G308));
  AOI21_X1  g736(.A(new_n1159), .B1(new_n1161), .B2(new_n944), .ZN(new_n1163));
  INV_X1    g737(.A(new_n1158), .ZN(new_n1164));
  NAND2_X1  g738(.A1(new_n1163), .A2(new_n1164), .ZN(G225));
endmodule


