

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U549 ( .A1(n695), .A2(n593), .ZN(n651) );
  INV_X1 U550 ( .A(n651), .ZN(n634) );
  NOR2_X2 U551 ( .A1(G164), .A2(G1384), .ZN(n695) );
  NOR2_X2 U552 ( .A1(n527), .A2(n526), .ZN(G164) );
  NOR2_X2 U553 ( .A1(G2105), .A2(G2104), .ZN(n518) );
  AND2_X1 U554 ( .A1(n535), .A2(n534), .ZN(G160) );
  OR2_X1 U555 ( .A1(G301), .A2(n642), .ZN(n514) );
  XOR2_X1 U556 ( .A(KEYINPUT90), .B(KEYINPUT29), .Z(n515) );
  AND2_X1 U557 ( .A1(n735), .A2(n728), .ZN(n516) );
  AND2_X1 U558 ( .A1(n727), .A2(n726), .ZN(n517) );
  NOR2_X1 U559 ( .A1(n609), .A2(n1000), .ZN(n610) );
  NOR2_X1 U560 ( .A1(G1966), .A2(n650), .ZN(n664) );
  NAND2_X1 U561 ( .A1(G8), .A2(n651), .ZN(n650) );
  AND2_X1 U562 ( .A1(n725), .A2(n516), .ZN(n726) );
  NOR2_X1 U563 ( .A1(G651), .A2(n563), .ZN(n767) );
  XNOR2_X1 U564 ( .A(KEYINPUT69), .B(n608), .ZN(n1000) );
  XOR2_X2 U565 ( .A(KEYINPUT17), .B(n518), .Z(n857) );
  NAND2_X1 U566 ( .A1(G138), .A2(n857), .ZN(n521) );
  INV_X1 U567 ( .A(G2104), .ZN(n523) );
  NOR2_X1 U568 ( .A1(n523), .A2(G2105), .ZN(n519) );
  XNOR2_X2 U569 ( .A(n519), .B(KEYINPUT64), .ZN(n858) );
  NAND2_X1 U570 ( .A1(G102), .A2(n858), .ZN(n520) );
  NAND2_X1 U571 ( .A1(n521), .A2(n520), .ZN(n522) );
  XNOR2_X1 U572 ( .A(n522), .B(KEYINPUT82), .ZN(n527) );
  AND2_X1 U573 ( .A1(n523), .A2(G2105), .ZN(n862) );
  NAND2_X1 U574 ( .A1(G126), .A2(n862), .ZN(n525) );
  AND2_X1 U575 ( .A1(G2105), .A2(G2104), .ZN(n863) );
  NAND2_X1 U576 ( .A1(G114), .A2(n863), .ZN(n524) );
  NAND2_X1 U577 ( .A1(n525), .A2(n524), .ZN(n526) );
  NAND2_X1 U578 ( .A1(n858), .A2(G101), .ZN(n528) );
  XOR2_X1 U579 ( .A(n528), .B(KEYINPUT23), .Z(n535) );
  NAND2_X1 U580 ( .A1(G113), .A2(n863), .ZN(n529) );
  XNOR2_X1 U581 ( .A(KEYINPUT65), .B(n529), .ZN(n533) );
  NAND2_X1 U582 ( .A1(G137), .A2(n857), .ZN(n531) );
  NAND2_X1 U583 ( .A1(G125), .A2(n862), .ZN(n530) );
  NAND2_X1 U584 ( .A1(n531), .A2(n530), .ZN(n532) );
  NOR2_X1 U585 ( .A1(n533), .A2(n532), .ZN(n534) );
  XOR2_X1 U586 ( .A(KEYINPUT0), .B(G543), .Z(n563) );
  NAND2_X1 U587 ( .A1(G52), .A2(n767), .ZN(n538) );
  INV_X1 U588 ( .A(G651), .ZN(n539) );
  NOR2_X1 U589 ( .A1(G543), .A2(n539), .ZN(n536) );
  XOR2_X1 U590 ( .A(KEYINPUT1), .B(n536), .Z(n768) );
  NAND2_X1 U591 ( .A1(G64), .A2(n768), .ZN(n537) );
  NAND2_X1 U592 ( .A1(n538), .A2(n537), .ZN(n544) );
  NOR2_X1 U593 ( .A1(G651), .A2(G543), .ZN(n771) );
  NAND2_X1 U594 ( .A1(G90), .A2(n771), .ZN(n541) );
  NOR2_X2 U595 ( .A1(n563), .A2(n539), .ZN(n772) );
  NAND2_X1 U596 ( .A1(G77), .A2(n772), .ZN(n540) );
  NAND2_X1 U597 ( .A1(n541), .A2(n540), .ZN(n542) );
  XOR2_X1 U598 ( .A(KEYINPUT9), .B(n542), .Z(n543) );
  NOR2_X1 U599 ( .A1(n544), .A2(n543), .ZN(G171) );
  INV_X1 U600 ( .A(G171), .ZN(G301) );
  NAND2_X1 U601 ( .A1(G89), .A2(n771), .ZN(n545) );
  XNOR2_X1 U602 ( .A(n545), .B(KEYINPUT4), .ZN(n546) );
  XNOR2_X1 U603 ( .A(n546), .B(KEYINPUT70), .ZN(n548) );
  NAND2_X1 U604 ( .A1(G76), .A2(n772), .ZN(n547) );
  NAND2_X1 U605 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U606 ( .A(n549), .B(KEYINPUT5), .ZN(n554) );
  NAND2_X1 U607 ( .A1(G51), .A2(n767), .ZN(n551) );
  NAND2_X1 U608 ( .A1(G63), .A2(n768), .ZN(n550) );
  NAND2_X1 U609 ( .A1(n551), .A2(n550), .ZN(n552) );
  XOR2_X1 U610 ( .A(KEYINPUT6), .B(n552), .Z(n553) );
  NAND2_X1 U611 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U612 ( .A(n555), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U613 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U614 ( .A1(G88), .A2(n771), .ZN(n557) );
  NAND2_X1 U615 ( .A1(G75), .A2(n772), .ZN(n556) );
  NAND2_X1 U616 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U617 ( .A(KEYINPUT77), .B(n558), .ZN(n562) );
  NAND2_X1 U618 ( .A1(G50), .A2(n767), .ZN(n560) );
  NAND2_X1 U619 ( .A1(G62), .A2(n768), .ZN(n559) );
  AND2_X1 U620 ( .A1(n560), .A2(n559), .ZN(n561) );
  NAND2_X1 U621 ( .A1(n562), .A2(n561), .ZN(G303) );
  NAND2_X1 U622 ( .A1(G49), .A2(n767), .ZN(n565) );
  NAND2_X1 U623 ( .A1(G87), .A2(n563), .ZN(n564) );
  NAND2_X1 U624 ( .A1(n565), .A2(n564), .ZN(n566) );
  NOR2_X1 U625 ( .A1(n768), .A2(n566), .ZN(n568) );
  NAND2_X1 U626 ( .A1(G651), .A2(G74), .ZN(n567) );
  NAND2_X1 U627 ( .A1(n568), .A2(n567), .ZN(G288) );
  XOR2_X1 U628 ( .A(KEYINPUT76), .B(KEYINPUT2), .Z(n570) );
  NAND2_X1 U629 ( .A1(G73), .A2(n772), .ZN(n569) );
  XNOR2_X1 U630 ( .A(n570), .B(n569), .ZN(n576) );
  NAND2_X1 U631 ( .A1(n771), .A2(G86), .ZN(n571) );
  XNOR2_X1 U632 ( .A(n571), .B(KEYINPUT74), .ZN(n573) );
  NAND2_X1 U633 ( .A1(G61), .A2(n768), .ZN(n572) );
  NAND2_X1 U634 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U635 ( .A(KEYINPUT75), .B(n574), .Z(n575) );
  NOR2_X1 U636 ( .A1(n576), .A2(n575), .ZN(n578) );
  NAND2_X1 U637 ( .A1(n767), .A2(G48), .ZN(n577) );
  NAND2_X1 U638 ( .A1(n578), .A2(n577), .ZN(G305) );
  NAND2_X1 U639 ( .A1(G47), .A2(n767), .ZN(n580) );
  NAND2_X1 U640 ( .A1(G60), .A2(n768), .ZN(n579) );
  NAND2_X1 U641 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U642 ( .A(KEYINPUT66), .B(n581), .Z(n585) );
  NAND2_X1 U643 ( .A1(G85), .A2(n771), .ZN(n583) );
  NAND2_X1 U644 ( .A1(G72), .A2(n772), .ZN(n582) );
  AND2_X1 U645 ( .A1(n583), .A2(n582), .ZN(n584) );
  NAND2_X1 U646 ( .A1(n585), .A2(n584), .ZN(G290) );
  NAND2_X1 U647 ( .A1(G92), .A2(n771), .ZN(n587) );
  NAND2_X1 U648 ( .A1(G79), .A2(n772), .ZN(n586) );
  NAND2_X1 U649 ( .A1(n587), .A2(n586), .ZN(n591) );
  NAND2_X1 U650 ( .A1(G54), .A2(n767), .ZN(n589) );
  NAND2_X1 U651 ( .A1(G66), .A2(n768), .ZN(n588) );
  NAND2_X1 U652 ( .A1(n589), .A2(n588), .ZN(n590) );
  NOR2_X1 U653 ( .A1(n591), .A2(n590), .ZN(n592) );
  XOR2_X1 U654 ( .A(KEYINPUT15), .B(n592), .Z(n877) );
  NAND2_X1 U655 ( .A1(G160), .A2(G40), .ZN(n696) );
  INV_X1 U656 ( .A(n696), .ZN(n593) );
  INV_X1 U657 ( .A(G1996), .ZN(n933) );
  NOR2_X1 U658 ( .A1(n651), .A2(n933), .ZN(n595) );
  INV_X1 U659 ( .A(KEYINPUT26), .ZN(n594) );
  XNOR2_X1 U660 ( .A(n595), .B(n594), .ZN(n597) );
  NAND2_X1 U661 ( .A1(n651), .A2(G1341), .ZN(n596) );
  NAND2_X1 U662 ( .A1(n597), .A2(n596), .ZN(n609) );
  NAND2_X1 U663 ( .A1(n772), .A2(G68), .ZN(n598) );
  XNOR2_X1 U664 ( .A(KEYINPUT68), .B(n598), .ZN(n601) );
  NAND2_X1 U665 ( .A1(n771), .A2(G81), .ZN(n599) );
  XNOR2_X1 U666 ( .A(KEYINPUT12), .B(n599), .ZN(n600) );
  NAND2_X1 U667 ( .A1(n601), .A2(n600), .ZN(n602) );
  XNOR2_X1 U668 ( .A(n602), .B(KEYINPUT13), .ZN(n604) );
  NAND2_X1 U669 ( .A1(G43), .A2(n767), .ZN(n603) );
  NAND2_X1 U670 ( .A1(n604), .A2(n603), .ZN(n607) );
  NAND2_X1 U671 ( .A1(n768), .A2(G56), .ZN(n605) );
  XOR2_X1 U672 ( .A(KEYINPUT14), .B(n605), .Z(n606) );
  NOR2_X1 U673 ( .A1(n607), .A2(n606), .ZN(n608) );
  OR2_X1 U674 ( .A1(n877), .A2(n610), .ZN(n617) );
  NAND2_X1 U675 ( .A1(n877), .A2(n610), .ZN(n615) );
  AND2_X1 U676 ( .A1(n634), .A2(G2067), .ZN(n611) );
  XNOR2_X1 U677 ( .A(n611), .B(KEYINPUT89), .ZN(n613) );
  NAND2_X1 U678 ( .A1(n651), .A2(G1348), .ZN(n612) );
  NAND2_X1 U679 ( .A1(n613), .A2(n612), .ZN(n614) );
  NAND2_X1 U680 ( .A1(n615), .A2(n614), .ZN(n616) );
  NAND2_X1 U681 ( .A1(n617), .A2(n616), .ZN(n628) );
  NAND2_X1 U682 ( .A1(G53), .A2(n767), .ZN(n619) );
  NAND2_X1 U683 ( .A1(G65), .A2(n768), .ZN(n618) );
  NAND2_X1 U684 ( .A1(n619), .A2(n618), .ZN(n623) );
  NAND2_X1 U685 ( .A1(G91), .A2(n771), .ZN(n621) );
  NAND2_X1 U686 ( .A1(G78), .A2(n772), .ZN(n620) );
  NAND2_X1 U687 ( .A1(n621), .A2(n620), .ZN(n622) );
  NOR2_X1 U688 ( .A1(n623), .A2(n622), .ZN(n985) );
  NAND2_X1 U689 ( .A1(n634), .A2(G2072), .ZN(n624) );
  XNOR2_X1 U690 ( .A(n624), .B(KEYINPUT27), .ZN(n626) );
  INV_X1 U691 ( .A(G1956), .ZN(n960) );
  NOR2_X1 U692 ( .A1(n960), .A2(n634), .ZN(n625) );
  NOR2_X1 U693 ( .A1(n626), .A2(n625), .ZN(n629) );
  NAND2_X1 U694 ( .A1(n985), .A2(n629), .ZN(n627) );
  NAND2_X1 U695 ( .A1(n628), .A2(n627), .ZN(n632) );
  NOR2_X1 U696 ( .A1(n985), .A2(n629), .ZN(n630) );
  XOR2_X1 U697 ( .A(n630), .B(KEYINPUT28), .Z(n631) );
  NAND2_X1 U698 ( .A1(n632), .A2(n631), .ZN(n633) );
  XNOR2_X1 U699 ( .A(n633), .B(n515), .ZN(n637) );
  NAND2_X1 U700 ( .A1(G1961), .A2(n651), .ZN(n636) );
  XOR2_X1 U701 ( .A(G2078), .B(KEYINPUT25), .Z(n931) );
  NAND2_X1 U702 ( .A1(n634), .A2(n931), .ZN(n635) );
  NAND2_X1 U703 ( .A1(n636), .A2(n635), .ZN(n642) );
  AND2_X1 U704 ( .A1(n637), .A2(n514), .ZN(n648) );
  NOR2_X1 U705 ( .A1(G2084), .A2(n651), .ZN(n661) );
  NOR2_X1 U706 ( .A1(n664), .A2(n661), .ZN(n638) );
  XOR2_X1 U707 ( .A(KEYINPUT91), .B(n638), .Z(n639) );
  NAND2_X1 U708 ( .A1(n639), .A2(G8), .ZN(n640) );
  XNOR2_X1 U709 ( .A(n640), .B(KEYINPUT30), .ZN(n641) );
  NOR2_X1 U710 ( .A1(n641), .A2(G168), .ZN(n645) );
  NAND2_X1 U711 ( .A1(G301), .A2(n642), .ZN(n643) );
  XOR2_X1 U712 ( .A(KEYINPUT92), .B(n643), .Z(n644) );
  NOR2_X1 U713 ( .A1(n645), .A2(n644), .ZN(n646) );
  XNOR2_X1 U714 ( .A(n646), .B(KEYINPUT31), .ZN(n647) );
  NOR2_X1 U715 ( .A1(n648), .A2(n647), .ZN(n649) );
  XNOR2_X1 U716 ( .A(n649), .B(KEYINPUT93), .ZN(n662) );
  NAND2_X1 U717 ( .A1(n662), .A2(G286), .ZN(n659) );
  INV_X1 U718 ( .A(G8), .ZN(n657) );
  INV_X1 U719 ( .A(n650), .ZN(n673) );
  INV_X1 U720 ( .A(n673), .ZN(n691) );
  NOR2_X1 U721 ( .A1(G1971), .A2(n691), .ZN(n653) );
  NOR2_X1 U722 ( .A1(G2090), .A2(n651), .ZN(n652) );
  NOR2_X1 U723 ( .A1(n653), .A2(n652), .ZN(n654) );
  NAND2_X1 U724 ( .A1(n654), .A2(G303), .ZN(n655) );
  XNOR2_X1 U725 ( .A(n655), .B(KEYINPUT94), .ZN(n656) );
  OR2_X1 U726 ( .A1(n657), .A2(n656), .ZN(n658) );
  AND2_X1 U727 ( .A1(n659), .A2(n658), .ZN(n660) );
  XNOR2_X1 U728 ( .A(n660), .B(KEYINPUT32), .ZN(n668) );
  NAND2_X1 U729 ( .A1(G8), .A2(n661), .ZN(n666) );
  INV_X1 U730 ( .A(n662), .ZN(n663) );
  NOR2_X1 U731 ( .A1(n664), .A2(n663), .ZN(n665) );
  NAND2_X1 U732 ( .A1(n666), .A2(n665), .ZN(n667) );
  NAND2_X1 U733 ( .A1(n668), .A2(n667), .ZN(n689) );
  NOR2_X1 U734 ( .A1(G1976), .A2(G288), .ZN(n989) );
  NOR2_X1 U735 ( .A1(G1971), .A2(G303), .ZN(n669) );
  NOR2_X1 U736 ( .A1(n989), .A2(n669), .ZN(n671) );
  INV_X1 U737 ( .A(KEYINPUT33), .ZN(n670) );
  AND2_X1 U738 ( .A1(n671), .A2(n670), .ZN(n672) );
  NAND2_X1 U739 ( .A1(n689), .A2(n672), .ZN(n679) );
  NAND2_X1 U740 ( .A1(G1976), .A2(G288), .ZN(n986) );
  AND2_X1 U741 ( .A1(n673), .A2(n986), .ZN(n674) );
  NOR2_X1 U742 ( .A1(KEYINPUT33), .A2(n674), .ZN(n677) );
  NAND2_X1 U743 ( .A1(n989), .A2(KEYINPUT33), .ZN(n675) );
  NOR2_X1 U744 ( .A1(n675), .A2(n691), .ZN(n676) );
  NOR2_X1 U745 ( .A1(n677), .A2(n676), .ZN(n678) );
  AND2_X1 U746 ( .A1(n679), .A2(n678), .ZN(n680) );
  XOR2_X1 U747 ( .A(G1981), .B(G305), .Z(n1003) );
  NAND2_X1 U748 ( .A1(n680), .A2(n1003), .ZN(n681) );
  XNOR2_X1 U749 ( .A(n681), .B(KEYINPUT95), .ZN(n686) );
  NOR2_X1 U750 ( .A1(G1981), .A2(G305), .ZN(n682) );
  XOR2_X1 U751 ( .A(n682), .B(KEYINPUT24), .Z(n683) );
  XNOR2_X1 U752 ( .A(KEYINPUT88), .B(n683), .ZN(n684) );
  NOR2_X1 U753 ( .A1(n691), .A2(n684), .ZN(n685) );
  NOR2_X1 U754 ( .A1(n686), .A2(n685), .ZN(n694) );
  NOR2_X1 U755 ( .A1(G2090), .A2(G303), .ZN(n687) );
  NAND2_X1 U756 ( .A1(G8), .A2(n687), .ZN(n688) );
  XNOR2_X1 U757 ( .A(n688), .B(KEYINPUT96), .ZN(n690) );
  NAND2_X1 U758 ( .A1(n690), .A2(n689), .ZN(n692) );
  NAND2_X1 U759 ( .A1(n692), .A2(n691), .ZN(n693) );
  NAND2_X1 U760 ( .A1(n694), .A2(n693), .ZN(n727) );
  XNOR2_X1 U761 ( .A(G1986), .B(G290), .ZN(n992) );
  NOR2_X1 U762 ( .A1(n696), .A2(n695), .ZN(n740) );
  NAND2_X1 U763 ( .A1(n992), .A2(n740), .ZN(n697) );
  XOR2_X1 U764 ( .A(KEYINPUT83), .B(n697), .Z(n725) );
  NAND2_X1 U765 ( .A1(G140), .A2(n857), .ZN(n699) );
  NAND2_X1 U766 ( .A1(G104), .A2(n858), .ZN(n698) );
  NAND2_X1 U767 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U768 ( .A(KEYINPUT34), .B(n700), .ZN(n706) );
  NAND2_X1 U769 ( .A1(n862), .A2(G128), .ZN(n701) );
  XNOR2_X1 U770 ( .A(n701), .B(KEYINPUT84), .ZN(n703) );
  NAND2_X1 U771 ( .A1(G116), .A2(n863), .ZN(n702) );
  NAND2_X1 U772 ( .A1(n703), .A2(n702), .ZN(n704) );
  XOR2_X1 U773 ( .A(n704), .B(KEYINPUT35), .Z(n705) );
  NOR2_X1 U774 ( .A1(n706), .A2(n705), .ZN(n707) );
  XOR2_X1 U775 ( .A(KEYINPUT36), .B(n707), .Z(n708) );
  XNOR2_X1 U776 ( .A(KEYINPUT85), .B(n708), .ZN(n874) );
  XNOR2_X1 U777 ( .A(G2067), .B(KEYINPUT37), .ZN(n737) );
  NOR2_X1 U778 ( .A1(n874), .A2(n737), .ZN(n912) );
  NAND2_X1 U779 ( .A1(n740), .A2(n912), .ZN(n735) );
  XOR2_X1 U780 ( .A(KEYINPUT87), .B(G1991), .Z(n937) );
  NAND2_X1 U781 ( .A1(G119), .A2(n862), .ZN(n710) );
  NAND2_X1 U782 ( .A1(G107), .A2(n863), .ZN(n709) );
  NAND2_X1 U783 ( .A1(n710), .A2(n709), .ZN(n713) );
  NAND2_X1 U784 ( .A1(n858), .A2(G95), .ZN(n711) );
  XOR2_X1 U785 ( .A(KEYINPUT86), .B(n711), .Z(n712) );
  NOR2_X1 U786 ( .A1(n713), .A2(n712), .ZN(n715) );
  NAND2_X1 U787 ( .A1(n857), .A2(G131), .ZN(n714) );
  NAND2_X1 U788 ( .A1(n715), .A2(n714), .ZN(n851) );
  NAND2_X1 U789 ( .A1(n937), .A2(n851), .ZN(n724) );
  NAND2_X1 U790 ( .A1(G129), .A2(n862), .ZN(n717) );
  NAND2_X1 U791 ( .A1(G117), .A2(n863), .ZN(n716) );
  NAND2_X1 U792 ( .A1(n717), .A2(n716), .ZN(n720) );
  NAND2_X1 U793 ( .A1(n858), .A2(G105), .ZN(n718) );
  XOR2_X1 U794 ( .A(KEYINPUT38), .B(n718), .Z(n719) );
  NOR2_X1 U795 ( .A1(n720), .A2(n719), .ZN(n722) );
  NAND2_X1 U796 ( .A1(n857), .A2(G141), .ZN(n721) );
  NAND2_X1 U797 ( .A1(n722), .A2(n721), .ZN(n850) );
  NAND2_X1 U798 ( .A1(G1996), .A2(n850), .ZN(n723) );
  NAND2_X1 U799 ( .A1(n724), .A2(n723), .ZN(n905) );
  NAND2_X1 U800 ( .A1(n740), .A2(n905), .ZN(n728) );
  XNOR2_X1 U801 ( .A(n517), .B(KEYINPUT97), .ZN(n742) );
  NOR2_X1 U802 ( .A1(G1996), .A2(n850), .ZN(n902) );
  INV_X1 U803 ( .A(n728), .ZN(n731) );
  NOR2_X1 U804 ( .A1(n937), .A2(n851), .ZN(n909) );
  NOR2_X1 U805 ( .A1(G1986), .A2(G290), .ZN(n729) );
  NOR2_X1 U806 ( .A1(n909), .A2(n729), .ZN(n730) );
  NOR2_X1 U807 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U808 ( .A(n732), .B(KEYINPUT98), .ZN(n733) );
  NOR2_X1 U809 ( .A1(n902), .A2(n733), .ZN(n734) );
  XNOR2_X1 U810 ( .A(n734), .B(KEYINPUT39), .ZN(n736) );
  NAND2_X1 U811 ( .A1(n736), .A2(n735), .ZN(n738) );
  NAND2_X1 U812 ( .A1(n874), .A2(n737), .ZN(n920) );
  NAND2_X1 U813 ( .A1(n738), .A2(n920), .ZN(n739) );
  NAND2_X1 U814 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U815 ( .A1(n742), .A2(n741), .ZN(n743) );
  XNOR2_X1 U816 ( .A(n743), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U817 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U818 ( .A1(G123), .A2(n862), .ZN(n744) );
  XNOR2_X1 U819 ( .A(n744), .B(KEYINPUT18), .ZN(n751) );
  NAND2_X1 U820 ( .A1(G135), .A2(n857), .ZN(n746) );
  NAND2_X1 U821 ( .A1(G111), .A2(n863), .ZN(n745) );
  NAND2_X1 U822 ( .A1(n746), .A2(n745), .ZN(n749) );
  NAND2_X1 U823 ( .A1(G99), .A2(n858), .ZN(n747) );
  XNOR2_X1 U824 ( .A(KEYINPUT71), .B(n747), .ZN(n748) );
  NOR2_X1 U825 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U826 ( .A1(n751), .A2(n750), .ZN(n752) );
  XNOR2_X1 U827 ( .A(KEYINPUT72), .B(n752), .ZN(n906) );
  XNOR2_X1 U828 ( .A(n906), .B(G2096), .ZN(n753) );
  OR2_X1 U829 ( .A1(G2100), .A2(n753), .ZN(G156) );
  INV_X1 U830 ( .A(G57), .ZN(G237) );
  INV_X1 U831 ( .A(G120), .ZN(G236) );
  NAND2_X1 U832 ( .A1(G7), .A2(G661), .ZN(n754) );
  XNOR2_X1 U833 ( .A(n754), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U834 ( .A(G223), .ZN(n807) );
  NAND2_X1 U835 ( .A1(n807), .A2(G567), .ZN(n755) );
  XOR2_X1 U836 ( .A(KEYINPUT11), .B(n755), .Z(G234) );
  INV_X1 U837 ( .A(n1000), .ZN(n756) );
  NAND2_X1 U838 ( .A1(n756), .A2(G860), .ZN(G153) );
  NAND2_X1 U839 ( .A1(G868), .A2(G301), .ZN(n758) );
  INV_X1 U840 ( .A(n877), .ZN(n990) );
  INV_X1 U841 ( .A(G868), .ZN(n788) );
  NAND2_X1 U842 ( .A1(n990), .A2(n788), .ZN(n757) );
  NAND2_X1 U843 ( .A1(n758), .A2(n757), .ZN(G284) );
  XNOR2_X1 U844 ( .A(n985), .B(KEYINPUT67), .ZN(G299) );
  NAND2_X1 U845 ( .A1(G286), .A2(G868), .ZN(n760) );
  NAND2_X1 U846 ( .A1(G299), .A2(n788), .ZN(n759) );
  NAND2_X1 U847 ( .A1(n760), .A2(n759), .ZN(G297) );
  INV_X1 U848 ( .A(G559), .ZN(n763) );
  NOR2_X1 U849 ( .A1(G860), .A2(n763), .ZN(n761) );
  NOR2_X1 U850 ( .A1(n990), .A2(n761), .ZN(n762) );
  XOR2_X1 U851 ( .A(KEYINPUT16), .B(n762), .Z(G148) );
  NAND2_X1 U852 ( .A1(n763), .A2(n877), .ZN(n764) );
  NAND2_X1 U853 ( .A1(n764), .A2(G868), .ZN(n766) );
  NAND2_X1 U854 ( .A1(n1000), .A2(n788), .ZN(n765) );
  NAND2_X1 U855 ( .A1(n766), .A2(n765), .ZN(G282) );
  NAND2_X1 U856 ( .A1(G55), .A2(n767), .ZN(n770) );
  NAND2_X1 U857 ( .A1(G67), .A2(n768), .ZN(n769) );
  NAND2_X1 U858 ( .A1(n770), .A2(n769), .ZN(n776) );
  NAND2_X1 U859 ( .A1(G93), .A2(n771), .ZN(n774) );
  NAND2_X1 U860 ( .A1(G80), .A2(n772), .ZN(n773) );
  NAND2_X1 U861 ( .A1(n774), .A2(n773), .ZN(n775) );
  NOR2_X1 U862 ( .A1(n776), .A2(n775), .ZN(n787) );
  NAND2_X1 U863 ( .A1(G559), .A2(n877), .ZN(n777) );
  XNOR2_X1 U864 ( .A(n777), .B(n1000), .ZN(n785) );
  NOR2_X1 U865 ( .A1(G860), .A2(n785), .ZN(n778) );
  XOR2_X1 U866 ( .A(KEYINPUT73), .B(n778), .Z(n779) );
  XNOR2_X1 U867 ( .A(n787), .B(n779), .ZN(G145) );
  INV_X1 U868 ( .A(G303), .ZN(G166) );
  XNOR2_X1 U869 ( .A(n787), .B(G299), .ZN(n782) );
  XNOR2_X1 U870 ( .A(G166), .B(KEYINPUT19), .ZN(n780) );
  XNOR2_X1 U871 ( .A(n780), .B(G288), .ZN(n781) );
  XNOR2_X1 U872 ( .A(n782), .B(n781), .ZN(n783) );
  XNOR2_X1 U873 ( .A(n783), .B(G290), .ZN(n784) );
  XNOR2_X1 U874 ( .A(n784), .B(G305), .ZN(n880) );
  XNOR2_X1 U875 ( .A(n785), .B(n880), .ZN(n786) );
  NAND2_X1 U876 ( .A1(n786), .A2(G868), .ZN(n790) );
  NAND2_X1 U877 ( .A1(n788), .A2(n787), .ZN(n789) );
  NAND2_X1 U878 ( .A1(n790), .A2(n789), .ZN(n791) );
  XOR2_X1 U879 ( .A(KEYINPUT78), .B(n791), .Z(G295) );
  NAND2_X1 U880 ( .A1(G2078), .A2(G2084), .ZN(n792) );
  XNOR2_X1 U881 ( .A(n792), .B(KEYINPUT20), .ZN(n793) );
  XNOR2_X1 U882 ( .A(n793), .B(KEYINPUT79), .ZN(n794) );
  NAND2_X1 U883 ( .A1(n794), .A2(G2090), .ZN(n795) );
  XNOR2_X1 U884 ( .A(KEYINPUT21), .B(n795), .ZN(n796) );
  NAND2_X1 U885 ( .A1(n796), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U886 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U887 ( .A1(G236), .A2(G237), .ZN(n797) );
  NAND2_X1 U888 ( .A1(G69), .A2(n797), .ZN(n798) );
  XNOR2_X1 U889 ( .A(KEYINPUT81), .B(n798), .ZN(n799) );
  NAND2_X1 U890 ( .A1(n799), .A2(G108), .ZN(n812) );
  NAND2_X1 U891 ( .A1(G567), .A2(n812), .ZN(n805) );
  NAND2_X1 U892 ( .A1(G132), .A2(G82), .ZN(n800) );
  XNOR2_X1 U893 ( .A(n800), .B(KEYINPUT22), .ZN(n801) );
  XNOR2_X1 U894 ( .A(n801), .B(KEYINPUT80), .ZN(n802) );
  NOR2_X1 U895 ( .A1(G218), .A2(n802), .ZN(n803) );
  NAND2_X1 U896 ( .A1(G96), .A2(n803), .ZN(n813) );
  NAND2_X1 U897 ( .A1(G2106), .A2(n813), .ZN(n804) );
  NAND2_X1 U898 ( .A1(n805), .A2(n804), .ZN(n814) );
  NAND2_X1 U899 ( .A1(G483), .A2(G661), .ZN(n806) );
  NOR2_X1 U900 ( .A1(n814), .A2(n806), .ZN(n810) );
  NAND2_X1 U901 ( .A1(n810), .A2(G36), .ZN(G176) );
  NAND2_X1 U902 ( .A1(G2106), .A2(n807), .ZN(G217) );
  AND2_X1 U903 ( .A1(G15), .A2(G2), .ZN(n808) );
  NAND2_X1 U904 ( .A1(G661), .A2(n808), .ZN(G259) );
  NAND2_X1 U905 ( .A1(G3), .A2(G1), .ZN(n809) );
  XNOR2_X1 U906 ( .A(KEYINPUT100), .B(n809), .ZN(n811) );
  NAND2_X1 U907 ( .A1(n811), .A2(n810), .ZN(G188) );
  INV_X1 U909 ( .A(G132), .ZN(G219) );
  INV_X1 U910 ( .A(G108), .ZN(G238) );
  INV_X1 U911 ( .A(G82), .ZN(G220) );
  NOR2_X1 U912 ( .A1(n813), .A2(n812), .ZN(G325) );
  INV_X1 U913 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U914 ( .A(KEYINPUT101), .B(n814), .ZN(G319) );
  XOR2_X1 U915 ( .A(G2100), .B(G2096), .Z(n816) );
  XNOR2_X1 U916 ( .A(KEYINPUT42), .B(G2678), .ZN(n815) );
  XNOR2_X1 U917 ( .A(n816), .B(n815), .ZN(n820) );
  XOR2_X1 U918 ( .A(KEYINPUT43), .B(G2090), .Z(n818) );
  XNOR2_X1 U919 ( .A(G2067), .B(G2072), .ZN(n817) );
  XNOR2_X1 U920 ( .A(n818), .B(n817), .ZN(n819) );
  XOR2_X1 U921 ( .A(n820), .B(n819), .Z(n822) );
  XNOR2_X1 U922 ( .A(G2078), .B(G2084), .ZN(n821) );
  XNOR2_X1 U923 ( .A(n822), .B(n821), .ZN(G227) );
  XOR2_X1 U924 ( .A(KEYINPUT41), .B(G1976), .Z(n824) );
  XNOR2_X1 U925 ( .A(G1961), .B(G1956), .ZN(n823) );
  XNOR2_X1 U926 ( .A(n824), .B(n823), .ZN(n825) );
  XOR2_X1 U927 ( .A(n825), .B(G2474), .Z(n827) );
  XNOR2_X1 U928 ( .A(G1996), .B(G1991), .ZN(n826) );
  XNOR2_X1 U929 ( .A(n827), .B(n826), .ZN(n831) );
  XOR2_X1 U930 ( .A(G1981), .B(G1971), .Z(n829) );
  XNOR2_X1 U931 ( .A(G1986), .B(G1966), .ZN(n828) );
  XNOR2_X1 U932 ( .A(n829), .B(n828), .ZN(n830) );
  XOR2_X1 U933 ( .A(n831), .B(n830), .Z(n833) );
  XNOR2_X1 U934 ( .A(KEYINPUT102), .B(KEYINPUT103), .ZN(n832) );
  XNOR2_X1 U935 ( .A(n833), .B(n832), .ZN(G229) );
  NAND2_X1 U936 ( .A1(n862), .A2(G124), .ZN(n834) );
  XNOR2_X1 U937 ( .A(n834), .B(KEYINPUT44), .ZN(n836) );
  NAND2_X1 U938 ( .A1(G112), .A2(n863), .ZN(n835) );
  NAND2_X1 U939 ( .A1(n836), .A2(n835), .ZN(n840) );
  NAND2_X1 U940 ( .A1(G136), .A2(n857), .ZN(n838) );
  NAND2_X1 U941 ( .A1(G100), .A2(n858), .ZN(n837) );
  NAND2_X1 U942 ( .A1(n838), .A2(n837), .ZN(n839) );
  NOR2_X1 U943 ( .A1(n840), .A2(n839), .ZN(G162) );
  NAND2_X1 U944 ( .A1(n857), .A2(G142), .ZN(n841) );
  XOR2_X1 U945 ( .A(KEYINPUT105), .B(n841), .Z(n843) );
  NAND2_X1 U946 ( .A1(G106), .A2(n858), .ZN(n842) );
  NAND2_X1 U947 ( .A1(n843), .A2(n842), .ZN(n844) );
  XNOR2_X1 U948 ( .A(n844), .B(KEYINPUT45), .ZN(n846) );
  NAND2_X1 U949 ( .A1(G118), .A2(n863), .ZN(n845) );
  NAND2_X1 U950 ( .A1(n846), .A2(n845), .ZN(n849) );
  NAND2_X1 U951 ( .A1(n862), .A2(G130), .ZN(n847) );
  XOR2_X1 U952 ( .A(KEYINPUT104), .B(n847), .Z(n848) );
  NOR2_X1 U953 ( .A1(n849), .A2(n848), .ZN(n854) );
  XNOR2_X1 U954 ( .A(n906), .B(n850), .ZN(n852) );
  XNOR2_X1 U955 ( .A(n852), .B(n851), .ZN(n853) );
  XNOR2_X1 U956 ( .A(n854), .B(n853), .ZN(n873) );
  XOR2_X1 U957 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n856) );
  XNOR2_X1 U958 ( .A(G162), .B(KEYINPUT106), .ZN(n855) );
  XNOR2_X1 U959 ( .A(n856), .B(n855), .ZN(n869) );
  NAND2_X1 U960 ( .A1(G139), .A2(n857), .ZN(n860) );
  NAND2_X1 U961 ( .A1(G103), .A2(n858), .ZN(n859) );
  NAND2_X1 U962 ( .A1(n860), .A2(n859), .ZN(n861) );
  XOR2_X1 U963 ( .A(KEYINPUT107), .B(n861), .Z(n868) );
  NAND2_X1 U964 ( .A1(G127), .A2(n862), .ZN(n865) );
  NAND2_X1 U965 ( .A1(G115), .A2(n863), .ZN(n864) );
  NAND2_X1 U966 ( .A1(n865), .A2(n864), .ZN(n866) );
  XOR2_X1 U967 ( .A(KEYINPUT47), .B(n866), .Z(n867) );
  NOR2_X1 U968 ( .A1(n868), .A2(n867), .ZN(n916) );
  XOR2_X1 U969 ( .A(n869), .B(n916), .Z(n871) );
  XNOR2_X1 U970 ( .A(G160), .B(G164), .ZN(n870) );
  XNOR2_X1 U971 ( .A(n871), .B(n870), .ZN(n872) );
  XNOR2_X1 U972 ( .A(n873), .B(n872), .ZN(n875) );
  XOR2_X1 U973 ( .A(n875), .B(n874), .Z(n876) );
  NOR2_X1 U974 ( .A1(G37), .A2(n876), .ZN(G395) );
  XNOR2_X1 U975 ( .A(n1000), .B(G286), .ZN(n879) );
  XNOR2_X1 U976 ( .A(G171), .B(n877), .ZN(n878) );
  XNOR2_X1 U977 ( .A(n879), .B(n878), .ZN(n881) );
  XNOR2_X1 U978 ( .A(n881), .B(n880), .ZN(n882) );
  NOR2_X1 U979 ( .A1(G37), .A2(n882), .ZN(n883) );
  XNOR2_X1 U980 ( .A(KEYINPUT108), .B(n883), .ZN(G397) );
  XOR2_X1 U981 ( .A(G2454), .B(G2435), .Z(n885) );
  XNOR2_X1 U982 ( .A(G2438), .B(G2427), .ZN(n884) );
  XNOR2_X1 U983 ( .A(n885), .B(n884), .ZN(n892) );
  XOR2_X1 U984 ( .A(KEYINPUT99), .B(G2446), .Z(n887) );
  XNOR2_X1 U985 ( .A(G2443), .B(G2430), .ZN(n886) );
  XNOR2_X1 U986 ( .A(n887), .B(n886), .ZN(n888) );
  XOR2_X1 U987 ( .A(n888), .B(G2451), .Z(n890) );
  XNOR2_X1 U988 ( .A(G1341), .B(G1348), .ZN(n889) );
  XNOR2_X1 U989 ( .A(n890), .B(n889), .ZN(n891) );
  XNOR2_X1 U990 ( .A(n892), .B(n891), .ZN(n893) );
  NAND2_X1 U991 ( .A1(n893), .A2(G14), .ZN(n899) );
  NAND2_X1 U992 ( .A1(G319), .A2(n899), .ZN(n896) );
  NOR2_X1 U993 ( .A1(G227), .A2(G229), .ZN(n894) );
  XNOR2_X1 U994 ( .A(KEYINPUT49), .B(n894), .ZN(n895) );
  NOR2_X1 U995 ( .A1(n896), .A2(n895), .ZN(n898) );
  NOR2_X1 U996 ( .A1(G395), .A2(G397), .ZN(n897) );
  NAND2_X1 U997 ( .A1(n898), .A2(n897), .ZN(G225) );
  INV_X1 U998 ( .A(G225), .ZN(G308) );
  INV_X1 U999 ( .A(G96), .ZN(G221) );
  INV_X1 U1000 ( .A(G69), .ZN(G235) );
  INV_X1 U1001 ( .A(n899), .ZN(G401) );
  XNOR2_X1 U1002 ( .A(G2090), .B(G162), .ZN(n900) );
  XNOR2_X1 U1003 ( .A(n900), .B(KEYINPUT111), .ZN(n901) );
  NOR2_X1 U1004 ( .A1(n902), .A2(n901), .ZN(n903) );
  XNOR2_X1 U1005 ( .A(KEYINPUT51), .B(n903), .ZN(n904) );
  NOR2_X1 U1006 ( .A1(n905), .A2(n904), .ZN(n915) );
  XNOR2_X1 U1007 ( .A(G160), .B(G2084), .ZN(n907) );
  NAND2_X1 U1008 ( .A1(n907), .A2(n906), .ZN(n908) );
  NOR2_X1 U1009 ( .A1(n909), .A2(n908), .ZN(n910) );
  XNOR2_X1 U1010 ( .A(KEYINPUT109), .B(n910), .ZN(n911) );
  NOR2_X1 U1011 ( .A1(n912), .A2(n911), .ZN(n913) );
  XNOR2_X1 U1012 ( .A(n913), .B(KEYINPUT110), .ZN(n914) );
  NAND2_X1 U1013 ( .A1(n915), .A2(n914), .ZN(n923) );
  XOR2_X1 U1014 ( .A(G2072), .B(n916), .Z(n918) );
  XOR2_X1 U1015 ( .A(G164), .B(G2078), .Z(n917) );
  NOR2_X1 U1016 ( .A1(n918), .A2(n917), .ZN(n919) );
  XNOR2_X1 U1017 ( .A(n919), .B(KEYINPUT50), .ZN(n921) );
  NAND2_X1 U1018 ( .A1(n921), .A2(n920), .ZN(n922) );
  NOR2_X1 U1019 ( .A1(n923), .A2(n922), .ZN(n924) );
  XOR2_X1 U1020 ( .A(KEYINPUT52), .B(n924), .Z(n925) );
  NOR2_X1 U1021 ( .A1(KEYINPUT55), .A2(n925), .ZN(n926) );
  XOR2_X1 U1022 ( .A(KEYINPUT112), .B(n926), .Z(n927) );
  NAND2_X1 U1023 ( .A1(G29), .A2(n927), .ZN(n1015) );
  XOR2_X1 U1024 ( .A(G2090), .B(G35), .Z(n930) );
  XOR2_X1 U1025 ( .A(KEYINPUT54), .B(G34), .Z(n928) );
  XNOR2_X1 U1026 ( .A(G2084), .B(n928), .ZN(n929) );
  NAND2_X1 U1027 ( .A1(n930), .A2(n929), .ZN(n947) );
  XOR2_X1 U1028 ( .A(n931), .B(G27), .Z(n932) );
  NAND2_X1 U1029 ( .A1(n932), .A2(G28), .ZN(n936) );
  XOR2_X1 U1030 ( .A(KEYINPUT114), .B(n933), .Z(n934) );
  XNOR2_X1 U1031 ( .A(G32), .B(n934), .ZN(n935) );
  NOR2_X1 U1032 ( .A1(n936), .A2(n935), .ZN(n944) );
  XNOR2_X1 U1033 ( .A(n937), .B(G25), .ZN(n942) );
  XNOR2_X1 U1034 ( .A(G2067), .B(G26), .ZN(n939) );
  XNOR2_X1 U1035 ( .A(G2072), .B(G33), .ZN(n938) );
  NOR2_X1 U1036 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1037 ( .A(KEYINPUT113), .B(n940), .ZN(n941) );
  NOR2_X1 U1038 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1039 ( .A1(n944), .A2(n943), .ZN(n945) );
  XOR2_X1 U1040 ( .A(n945), .B(KEYINPUT53), .Z(n946) );
  NOR2_X1 U1041 ( .A1(n947), .A2(n946), .ZN(n948) );
  XOR2_X1 U1042 ( .A(KEYINPUT116), .B(n948), .Z(n950) );
  XOR2_X1 U1043 ( .A(KEYINPUT55), .B(KEYINPUT115), .Z(n949) );
  XNOR2_X1 U1044 ( .A(n950), .B(n949), .ZN(n951) );
  OR2_X1 U1045 ( .A1(G29), .A2(n951), .ZN(n952) );
  NAND2_X1 U1046 ( .A1(G11), .A2(n952), .ZN(n1013) );
  XNOR2_X1 U1047 ( .A(KEYINPUT119), .B(G16), .ZN(n983) );
  XOR2_X1 U1048 ( .A(KEYINPUT126), .B(KEYINPUT127), .Z(n981) );
  XNOR2_X1 U1049 ( .A(G1966), .B(G21), .ZN(n954) );
  XNOR2_X1 U1050 ( .A(G5), .B(G1961), .ZN(n953) );
  NOR2_X1 U1051 ( .A1(n954), .A2(n953), .ZN(n969) );
  XNOR2_X1 U1052 ( .A(KEYINPUT60), .B(KEYINPUT123), .ZN(n967) );
  XNOR2_X1 U1053 ( .A(G1341), .B(G19), .ZN(n955) );
  XNOR2_X1 U1054 ( .A(n955), .B(KEYINPUT120), .ZN(n958) );
  XOR2_X1 U1055 ( .A(G1981), .B(G6), .Z(n956) );
  XNOR2_X1 U1056 ( .A(KEYINPUT121), .B(n956), .ZN(n957) );
  NOR2_X1 U1057 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1058 ( .A(KEYINPUT122), .B(n959), .ZN(n962) );
  XNOR2_X1 U1059 ( .A(n960), .B(G20), .ZN(n961) );
  NAND2_X1 U1060 ( .A1(n962), .A2(n961), .ZN(n965) );
  XOR2_X1 U1061 ( .A(G1348), .B(KEYINPUT59), .Z(n963) );
  XNOR2_X1 U1062 ( .A(G4), .B(n963), .ZN(n964) );
  NOR2_X1 U1063 ( .A1(n965), .A2(n964), .ZN(n966) );
  XOR2_X1 U1064 ( .A(n967), .B(n966), .Z(n968) );
  NAND2_X1 U1065 ( .A1(n969), .A2(n968), .ZN(n978) );
  XOR2_X1 U1066 ( .A(G1986), .B(G24), .Z(n974) );
  XNOR2_X1 U1067 ( .A(G1971), .B(G22), .ZN(n971) );
  XNOR2_X1 U1068 ( .A(G1976), .B(G23), .ZN(n970) );
  NOR2_X1 U1069 ( .A1(n971), .A2(n970), .ZN(n972) );
  XNOR2_X1 U1070 ( .A(n972), .B(KEYINPUT124), .ZN(n973) );
  NAND2_X1 U1071 ( .A1(n974), .A2(n973), .ZN(n975) );
  XOR2_X1 U1072 ( .A(KEYINPUT125), .B(n975), .Z(n976) );
  XNOR2_X1 U1073 ( .A(KEYINPUT58), .B(n976), .ZN(n977) );
  NOR2_X1 U1074 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1075 ( .A(n979), .B(KEYINPUT61), .ZN(n980) );
  XNOR2_X1 U1076 ( .A(n981), .B(n980), .ZN(n982) );
  NAND2_X1 U1077 ( .A1(n983), .A2(n982), .ZN(n1011) );
  XNOR2_X1 U1078 ( .A(KEYINPUT56), .B(G16), .ZN(n1009) );
  XNOR2_X1 U1079 ( .A(G1971), .B(G166), .ZN(n984) );
  XNOR2_X1 U1080 ( .A(n984), .B(KEYINPUT118), .ZN(n999) );
  XNOR2_X1 U1081 ( .A(n985), .B(G1956), .ZN(n987) );
  NAND2_X1 U1082 ( .A1(n987), .A2(n986), .ZN(n988) );
  NOR2_X1 U1083 ( .A1(n989), .A2(n988), .ZN(n994) );
  XNOR2_X1 U1084 ( .A(G1348), .B(n990), .ZN(n991) );
  NOR2_X1 U1085 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1086 ( .A1(n994), .A2(n993), .ZN(n997) );
  XOR2_X1 U1087 ( .A(G1961), .B(G301), .Z(n995) );
  XNOR2_X1 U1088 ( .A(KEYINPUT117), .B(n995), .ZN(n996) );
  NOR2_X1 U1089 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1090 ( .A1(n999), .A2(n998), .ZN(n1002) );
  XNOR2_X1 U1091 ( .A(G1341), .B(n1000), .ZN(n1001) );
  NOR2_X1 U1092 ( .A1(n1002), .A2(n1001), .ZN(n1007) );
  XNOR2_X1 U1093 ( .A(G1966), .B(G168), .ZN(n1004) );
  NAND2_X1 U1094 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1095 ( .A(n1005), .B(KEYINPUT57), .ZN(n1006) );
  NAND2_X1 U1096 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1098 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NOR2_X1 U1099 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1100 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XOR2_X1 U1101 ( .A(KEYINPUT62), .B(n1016), .Z(G311) );
  INV_X1 U1102 ( .A(G311), .ZN(G150) );
endmodule

