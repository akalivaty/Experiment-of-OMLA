

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578;

  XOR2_X1 U321 ( .A(KEYINPUT41), .B(n567), .Z(n550) );
  XNOR2_X1 U322 ( .A(n403), .B(n295), .ZN(n296) );
  XNOR2_X1 U323 ( .A(n371), .B(KEYINPUT48), .ZN(n372) );
  XNOR2_X1 U324 ( .A(n382), .B(n296), .ZN(n297) );
  XNOR2_X1 U325 ( .A(n373), .B(n372), .ZN(n532) );
  XNOR2_X1 U326 ( .A(G169GAT), .B(KEYINPUT119), .ZN(n445) );
  XNOR2_X1 U327 ( .A(n446), .B(n445), .ZN(G1348GAT) );
  XOR2_X1 U328 ( .A(KEYINPUT33), .B(KEYINPUT73), .Z(n290) );
  XNOR2_X1 U329 ( .A(G120GAT), .B(KEYINPUT74), .ZN(n289) );
  XNOR2_X1 U330 ( .A(n290), .B(n289), .ZN(n305) );
  XOR2_X1 U331 ( .A(KEYINPUT13), .B(KEYINPUT31), .Z(n292) );
  XNOR2_X1 U332 ( .A(KEYINPUT71), .B(KEYINPUT32), .ZN(n291) );
  XNOR2_X1 U333 ( .A(n292), .B(n291), .ZN(n298) );
  XOR2_X1 U334 ( .A(G64GAT), .B(KEYINPUT72), .Z(n294) );
  XNOR2_X1 U335 ( .A(G204GAT), .B(G92GAT), .ZN(n293) );
  XNOR2_X1 U336 ( .A(n294), .B(n293), .ZN(n382) );
  XOR2_X1 U337 ( .A(G85GAT), .B(G57GAT), .Z(n403) );
  AND2_X1 U338 ( .A1(G230GAT), .A2(G233GAT), .ZN(n295) );
  XOR2_X1 U339 ( .A(n298), .B(n297), .Z(n303) );
  XNOR2_X1 U340 ( .A(G99GAT), .B(G71GAT), .ZN(n299) );
  XNOR2_X1 U341 ( .A(n299), .B(G176GAT), .ZN(n435) );
  XOR2_X1 U342 ( .A(G78GAT), .B(G148GAT), .Z(n301) );
  XNOR2_X1 U343 ( .A(G106GAT), .B(KEYINPUT70), .ZN(n300) );
  XNOR2_X1 U344 ( .A(n301), .B(n300), .ZN(n415) );
  XNOR2_X1 U345 ( .A(n435), .B(n415), .ZN(n302) );
  XNOR2_X1 U346 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U347 ( .A(n305), .B(n304), .ZN(n567) );
  INV_X1 U348 ( .A(n550), .ZN(n538) );
  XOR2_X1 U349 ( .A(G29GAT), .B(G50GAT), .Z(n307) );
  XNOR2_X1 U350 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n306) );
  XNOR2_X1 U351 ( .A(n307), .B(n306), .ZN(n358) );
  XOR2_X1 U352 ( .A(G1GAT), .B(G8GAT), .Z(n309) );
  XNOR2_X1 U353 ( .A(G15GAT), .B(G22GAT), .ZN(n308) );
  XNOR2_X1 U354 ( .A(n309), .B(n308), .ZN(n341) );
  XNOR2_X1 U355 ( .A(n358), .B(n341), .ZN(n322) );
  XOR2_X1 U356 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n311) );
  NAND2_X1 U357 ( .A1(G229GAT), .A2(G233GAT), .ZN(n310) );
  XNOR2_X1 U358 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U359 ( .A(n312), .B(KEYINPUT67), .Z(n320) );
  XOR2_X1 U360 ( .A(G113GAT), .B(G43GAT), .Z(n314) );
  XNOR2_X1 U361 ( .A(G169GAT), .B(G36GAT), .ZN(n313) );
  XNOR2_X1 U362 ( .A(n314), .B(n313), .ZN(n318) );
  XOR2_X1 U363 ( .A(KEYINPUT68), .B(KEYINPUT69), .Z(n316) );
  XNOR2_X1 U364 ( .A(G197GAT), .B(G141GAT), .ZN(n315) );
  XNOR2_X1 U365 ( .A(n316), .B(n315), .ZN(n317) );
  XNOR2_X1 U366 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U367 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U368 ( .A(n322), .B(n321), .ZN(n564) );
  INV_X1 U369 ( .A(n564), .ZN(n536) );
  NAND2_X1 U370 ( .A1(n538), .A2(n536), .ZN(n325) );
  XOR2_X1 U371 ( .A(KEYINPUT46), .B(KEYINPUT110), .Z(n323) );
  XNOR2_X1 U372 ( .A(KEYINPUT109), .B(n323), .ZN(n324) );
  NAND2_X1 U373 ( .A1(n325), .A2(n324), .ZN(n327) );
  OR2_X1 U374 ( .A1(n325), .A2(n324), .ZN(n326) );
  NAND2_X1 U375 ( .A1(n327), .A2(n326), .ZN(n364) );
  XOR2_X1 U376 ( .A(KEYINPUT14), .B(G64GAT), .Z(n329) );
  XNOR2_X1 U377 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n328) );
  XNOR2_X1 U378 ( .A(n329), .B(n328), .ZN(n345) );
  XOR2_X1 U379 ( .A(KEYINPUT12), .B(KEYINPUT15), .Z(n331) );
  XNOR2_X1 U380 ( .A(KEYINPUT78), .B(KEYINPUT81), .ZN(n330) );
  XNOR2_X1 U381 ( .A(n331), .B(n330), .ZN(n339) );
  NAND2_X1 U382 ( .A1(G231GAT), .A2(G233GAT), .ZN(n337) );
  XOR2_X1 U383 ( .A(G78GAT), .B(G155GAT), .Z(n333) );
  XNOR2_X1 U384 ( .A(G71GAT), .B(G211GAT), .ZN(n332) );
  XNOR2_X1 U385 ( .A(n333), .B(n332), .ZN(n335) );
  XOR2_X1 U386 ( .A(G127GAT), .B(G183GAT), .Z(n334) );
  XNOR2_X1 U387 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U388 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U389 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U390 ( .A(n340), .B(KEYINPUT79), .Z(n343) );
  XNOR2_X1 U391 ( .A(n341), .B(KEYINPUT80), .ZN(n342) );
  XNOR2_X1 U392 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U393 ( .A(n345), .B(n344), .Z(n542) );
  XOR2_X1 U394 ( .A(KEYINPUT9), .B(G92GAT), .Z(n347) );
  XNOR2_X1 U395 ( .A(G99GAT), .B(G85GAT), .ZN(n346) );
  XNOR2_X1 U396 ( .A(n347), .B(n346), .ZN(n362) );
  XOR2_X1 U397 ( .A(G43GAT), .B(G134GAT), .Z(n432) );
  XOR2_X1 U398 ( .A(KEYINPUT75), .B(KEYINPUT77), .Z(n349) );
  XNOR2_X1 U399 ( .A(G218GAT), .B(KEYINPUT11), .ZN(n348) );
  XNOR2_X1 U400 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U401 ( .A(n432), .B(n350), .Z(n352) );
  NAND2_X1 U402 ( .A1(G232GAT), .A2(G233GAT), .ZN(n351) );
  XNOR2_X1 U403 ( .A(n352), .B(n351), .ZN(n356) );
  XOR2_X1 U404 ( .A(KEYINPUT10), .B(KEYINPUT66), .Z(n354) );
  XNOR2_X1 U405 ( .A(G162GAT), .B(G106GAT), .ZN(n353) );
  XNOR2_X1 U406 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U407 ( .A(n356), .B(n355), .Z(n360) );
  XNOR2_X1 U408 ( .A(G36GAT), .B(G190GAT), .ZN(n357) );
  XNOR2_X1 U409 ( .A(n357), .B(KEYINPUT76), .ZN(n380) );
  XNOR2_X1 U410 ( .A(n358), .B(n380), .ZN(n359) );
  XNOR2_X1 U411 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U412 ( .A(n362), .B(n361), .ZN(n557) );
  INV_X1 U413 ( .A(n557), .ZN(n545) );
  NOR2_X1 U414 ( .A1(n542), .A2(n545), .ZN(n363) );
  AND2_X1 U415 ( .A1(n364), .A2(n363), .ZN(n365) );
  XNOR2_X1 U416 ( .A(n365), .B(KEYINPUT47), .ZN(n370) );
  INV_X1 U417 ( .A(n567), .ZN(n447) );
  XNOR2_X1 U418 ( .A(KEYINPUT36), .B(n557), .ZN(n576) );
  INV_X1 U419 ( .A(n542), .ZN(n572) );
  NOR2_X1 U420 ( .A1(n576), .A2(n572), .ZN(n366) );
  XOR2_X1 U421 ( .A(KEYINPUT45), .B(n366), .Z(n367) );
  NOR2_X1 U422 ( .A1(n447), .A2(n367), .ZN(n368) );
  NAND2_X1 U423 ( .A1(n368), .A2(n564), .ZN(n369) );
  NAND2_X1 U424 ( .A1(n370), .A2(n369), .ZN(n373) );
  XNOR2_X1 U425 ( .A(KEYINPUT64), .B(KEYINPUT111), .ZN(n371) );
  XNOR2_X1 U426 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n374) );
  XNOR2_X1 U427 ( .A(n374), .B(KEYINPUT17), .ZN(n375) );
  XOR2_X1 U428 ( .A(n375), .B(KEYINPUT85), .Z(n377) );
  XNOR2_X1 U429 ( .A(G169GAT), .B(G183GAT), .ZN(n376) );
  XNOR2_X1 U430 ( .A(n377), .B(n376), .ZN(n440) );
  XOR2_X1 U431 ( .A(G176GAT), .B(KEYINPUT94), .Z(n379) );
  NAND2_X1 U432 ( .A1(G226GAT), .A2(G233GAT), .ZN(n378) );
  XNOR2_X1 U433 ( .A(n379), .B(n378), .ZN(n381) );
  XOR2_X1 U434 ( .A(n381), .B(n380), .Z(n384) );
  XNOR2_X1 U435 ( .A(G8GAT), .B(n382), .ZN(n383) );
  XNOR2_X1 U436 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U437 ( .A(n440), .B(n385), .ZN(n389) );
  XOR2_X1 U438 ( .A(KEYINPUT89), .B(G218GAT), .Z(n387) );
  XNOR2_X1 U439 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n386) );
  XNOR2_X1 U440 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U441 ( .A(G197GAT), .B(n388), .ZN(n425) );
  XNOR2_X1 U442 ( .A(n389), .B(n425), .ZN(n506) );
  NOR2_X1 U443 ( .A1(n532), .A2(n506), .ZN(n390) );
  XNOR2_X1 U444 ( .A(n390), .B(KEYINPUT54), .ZN(n413) );
  XOR2_X1 U445 ( .A(KEYINPUT0), .B(G127GAT), .Z(n392) );
  XNOR2_X1 U446 ( .A(KEYINPUT82), .B(G120GAT), .ZN(n391) );
  XNOR2_X1 U447 ( .A(n392), .B(n391), .ZN(n393) );
  XOR2_X1 U448 ( .A(G113GAT), .B(n393), .Z(n441) );
  XOR2_X1 U449 ( .A(G148GAT), .B(G134GAT), .Z(n395) );
  XNOR2_X1 U450 ( .A(G29GAT), .B(G1GAT), .ZN(n394) );
  XNOR2_X1 U451 ( .A(n395), .B(n394), .ZN(n399) );
  XOR2_X1 U452 ( .A(KEYINPUT6), .B(KEYINPUT5), .Z(n397) );
  XNOR2_X1 U453 ( .A(KEYINPUT91), .B(KEYINPUT92), .ZN(n396) );
  XNOR2_X1 U454 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U455 ( .A(n399), .B(n398), .Z(n405) );
  XOR2_X1 U456 ( .A(KEYINPUT4), .B(KEYINPUT1), .Z(n401) );
  NAND2_X1 U457 ( .A1(G225GAT), .A2(G233GAT), .ZN(n400) );
  XNOR2_X1 U458 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U459 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U460 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U461 ( .A(n441), .B(n406), .ZN(n412) );
  XNOR2_X1 U462 ( .A(G155GAT), .B(KEYINPUT2), .ZN(n407) );
  XNOR2_X1 U463 ( .A(n407), .B(KEYINPUT3), .ZN(n408) );
  XOR2_X1 U464 ( .A(n408), .B(KEYINPUT90), .Z(n410) );
  XNOR2_X1 U465 ( .A(G141GAT), .B(G162GAT), .ZN(n409) );
  XNOR2_X1 U466 ( .A(n410), .B(n409), .ZN(n422) );
  INV_X1 U467 ( .A(n422), .ZN(n411) );
  XNOR2_X1 U468 ( .A(n412), .B(n411), .ZN(n455) );
  XNOR2_X1 U469 ( .A(KEYINPUT93), .B(n455), .ZN(n503) );
  NAND2_X1 U470 ( .A1(n413), .A2(n503), .ZN(n414) );
  XNOR2_X1 U471 ( .A(n414), .B(KEYINPUT65), .ZN(n563) );
  XOR2_X1 U472 ( .A(n415), .B(G22GAT), .Z(n417) );
  NAND2_X1 U473 ( .A1(G228GAT), .A2(G233GAT), .ZN(n416) );
  XNOR2_X1 U474 ( .A(n417), .B(n416), .ZN(n421) );
  XOR2_X1 U475 ( .A(G204GAT), .B(KEYINPUT23), .Z(n419) );
  XNOR2_X1 U476 ( .A(KEYINPUT22), .B(KEYINPUT24), .ZN(n418) );
  XNOR2_X1 U477 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U478 ( .A(n421), .B(n420), .Z(n424) );
  XNOR2_X1 U479 ( .A(G50GAT), .B(n422), .ZN(n423) );
  XNOR2_X1 U480 ( .A(n424), .B(n423), .ZN(n426) );
  XNOR2_X1 U481 ( .A(n426), .B(n425), .ZN(n456) );
  NAND2_X1 U482 ( .A1(n563), .A2(n456), .ZN(n428) );
  XNOR2_X1 U483 ( .A(KEYINPUT55), .B(KEYINPUT118), .ZN(n427) );
  XNOR2_X1 U484 ( .A(n428), .B(n427), .ZN(n444) );
  XOR2_X1 U485 ( .A(KEYINPUT84), .B(KEYINPUT86), .Z(n430) );
  XNOR2_X1 U486 ( .A(KEYINPUT83), .B(KEYINPUT87), .ZN(n429) );
  XNOR2_X1 U487 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U488 ( .A(n431), .B(G190GAT), .Z(n434) );
  XNOR2_X1 U489 ( .A(G15GAT), .B(n432), .ZN(n433) );
  XNOR2_X1 U490 ( .A(n434), .B(n433), .ZN(n439) );
  XOR2_X1 U491 ( .A(n435), .B(KEYINPUT20), .Z(n437) );
  NAND2_X1 U492 ( .A1(G227GAT), .A2(G233GAT), .ZN(n436) );
  XNOR2_X1 U493 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U494 ( .A(n439), .B(n438), .Z(n443) );
  XNOR2_X1 U495 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U496 ( .A(n443), .B(n442), .ZN(n517) );
  NAND2_X1 U497 ( .A1(n444), .A2(n517), .ZN(n549) );
  NOR2_X1 U498 ( .A1(n549), .A2(n564), .ZN(n446) );
  NOR2_X1 U499 ( .A1(n564), .A2(n447), .ZN(n479) );
  INV_X1 U500 ( .A(n517), .ZN(n508) );
  OR2_X1 U501 ( .A1(n508), .A2(n506), .ZN(n448) );
  NAND2_X1 U502 ( .A1(n456), .A2(n448), .ZN(n449) );
  XOR2_X1 U503 ( .A(KEYINPUT25), .B(n449), .Z(n452) );
  NOR2_X1 U504 ( .A1(n456), .A2(n517), .ZN(n450) );
  XNOR2_X1 U505 ( .A(n450), .B(KEYINPUT26), .ZN(n562) );
  XNOR2_X1 U506 ( .A(KEYINPUT27), .B(KEYINPUT95), .ZN(n451) );
  XNOR2_X1 U507 ( .A(n451), .B(n506), .ZN(n457) );
  NAND2_X1 U508 ( .A1(n562), .A2(n457), .ZN(n531) );
  NAND2_X1 U509 ( .A1(n452), .A2(n531), .ZN(n453) );
  XOR2_X1 U510 ( .A(KEYINPUT98), .B(n453), .Z(n454) );
  NOR2_X1 U511 ( .A1(n455), .A2(n454), .ZN(n463) );
  INV_X1 U512 ( .A(n503), .ZN(n534) );
  XNOR2_X1 U513 ( .A(n456), .B(KEYINPUT28), .ZN(n511) );
  AND2_X1 U514 ( .A1(n534), .A2(n511), .ZN(n458) );
  NAND2_X1 U515 ( .A1(n458), .A2(n457), .ZN(n515) );
  XNOR2_X1 U516 ( .A(n515), .B(KEYINPUT96), .ZN(n460) );
  XNOR2_X1 U517 ( .A(n517), .B(KEYINPUT88), .ZN(n459) );
  NOR2_X1 U518 ( .A1(n460), .A2(n459), .ZN(n461) );
  XOR2_X1 U519 ( .A(KEYINPUT97), .B(n461), .Z(n462) );
  NOR2_X1 U520 ( .A1(n463), .A2(n462), .ZN(n476) );
  NOR2_X1 U521 ( .A1(n545), .A2(n572), .ZN(n464) );
  XOR2_X1 U522 ( .A(KEYINPUT16), .B(n464), .Z(n465) );
  NOR2_X1 U523 ( .A1(n476), .A2(n465), .ZN(n491) );
  NAND2_X1 U524 ( .A1(n479), .A2(n491), .ZN(n473) );
  NOR2_X1 U525 ( .A1(n503), .A2(n473), .ZN(n467) );
  XNOR2_X1 U526 ( .A(KEYINPUT99), .B(KEYINPUT34), .ZN(n466) );
  XNOR2_X1 U527 ( .A(n467), .B(n466), .ZN(n468) );
  XNOR2_X1 U528 ( .A(G1GAT), .B(n468), .ZN(G1324GAT) );
  NOR2_X1 U529 ( .A1(n506), .A2(n473), .ZN(n469) );
  XOR2_X1 U530 ( .A(G8GAT), .B(n469), .Z(G1325GAT) );
  NOR2_X1 U531 ( .A1(n508), .A2(n473), .ZN(n471) );
  XNOR2_X1 U532 ( .A(KEYINPUT100), .B(KEYINPUT35), .ZN(n470) );
  XNOR2_X1 U533 ( .A(n471), .B(n470), .ZN(n472) );
  XNOR2_X1 U534 ( .A(G15GAT), .B(n472), .ZN(G1326GAT) );
  NOR2_X1 U535 ( .A1(n511), .A2(n473), .ZN(n474) );
  XOR2_X1 U536 ( .A(G22GAT), .B(n474), .Z(G1327GAT) );
  XNOR2_X1 U537 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n475) );
  XNOR2_X1 U538 ( .A(n475), .B(KEYINPUT101), .ZN(n482) );
  NOR2_X1 U539 ( .A1(n576), .A2(n476), .ZN(n477) );
  NAND2_X1 U540 ( .A1(n572), .A2(n477), .ZN(n478) );
  XNOR2_X1 U541 ( .A(n478), .B(KEYINPUT37), .ZN(n502) );
  NAND2_X1 U542 ( .A1(n502), .A2(n479), .ZN(n480) );
  XNOR2_X1 U543 ( .A(KEYINPUT38), .B(n480), .ZN(n488) );
  NOR2_X1 U544 ( .A1(n503), .A2(n488), .ZN(n481) );
  XOR2_X1 U545 ( .A(n482), .B(n481), .Z(G1328GAT) );
  NOR2_X1 U546 ( .A1(n488), .A2(n506), .ZN(n483) );
  XOR2_X1 U547 ( .A(G36GAT), .B(n483), .Z(G1329GAT) );
  XOR2_X1 U548 ( .A(KEYINPUT40), .B(KEYINPUT103), .Z(n485) );
  XNOR2_X1 U549 ( .A(G43GAT), .B(KEYINPUT102), .ZN(n484) );
  XNOR2_X1 U550 ( .A(n485), .B(n484), .ZN(n487) );
  NOR2_X1 U551 ( .A1(n488), .A2(n508), .ZN(n486) );
  XOR2_X1 U552 ( .A(n487), .B(n486), .Z(G1330GAT) );
  NOR2_X1 U553 ( .A1(n488), .A2(n511), .ZN(n489) );
  XOR2_X1 U554 ( .A(KEYINPUT104), .B(n489), .Z(n490) );
  XNOR2_X1 U555 ( .A(G50GAT), .B(n490), .ZN(G1331GAT) );
  NOR2_X1 U556 ( .A1(n536), .A2(n550), .ZN(n501) );
  NAND2_X1 U557 ( .A1(n501), .A2(n491), .ZN(n497) );
  NOR2_X1 U558 ( .A1(n503), .A2(n497), .ZN(n492) );
  XOR2_X1 U559 ( .A(G57GAT), .B(n492), .Z(n493) );
  XNOR2_X1 U560 ( .A(KEYINPUT42), .B(n493), .ZN(G1332GAT) );
  NOR2_X1 U561 ( .A1(n506), .A2(n497), .ZN(n494) );
  XOR2_X1 U562 ( .A(G64GAT), .B(n494), .Z(G1333GAT) );
  NOR2_X1 U563 ( .A1(n508), .A2(n497), .ZN(n496) );
  XNOR2_X1 U564 ( .A(G71GAT), .B(KEYINPUT105), .ZN(n495) );
  XNOR2_X1 U565 ( .A(n496), .B(n495), .ZN(G1334GAT) );
  NOR2_X1 U566 ( .A1(n511), .A2(n497), .ZN(n499) );
  XNOR2_X1 U567 ( .A(KEYINPUT43), .B(KEYINPUT106), .ZN(n498) );
  XNOR2_X1 U568 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U569 ( .A(G78GAT), .B(n500), .ZN(G1335GAT) );
  NAND2_X1 U570 ( .A1(n502), .A2(n501), .ZN(n510) );
  NOR2_X1 U571 ( .A1(n503), .A2(n510), .ZN(n505) );
  XNOR2_X1 U572 ( .A(G85GAT), .B(KEYINPUT107), .ZN(n504) );
  XNOR2_X1 U573 ( .A(n505), .B(n504), .ZN(G1336GAT) );
  NOR2_X1 U574 ( .A1(n506), .A2(n510), .ZN(n507) );
  XOR2_X1 U575 ( .A(G92GAT), .B(n507), .Z(G1337GAT) );
  NOR2_X1 U576 ( .A1(n508), .A2(n510), .ZN(n509) );
  XOR2_X1 U577 ( .A(G99GAT), .B(n509), .Z(G1338GAT) );
  NOR2_X1 U578 ( .A1(n511), .A2(n510), .ZN(n513) );
  XNOR2_X1 U579 ( .A(KEYINPUT108), .B(KEYINPUT44), .ZN(n512) );
  XNOR2_X1 U580 ( .A(n513), .B(n512), .ZN(n514) );
  XOR2_X1 U581 ( .A(G106GAT), .B(n514), .Z(G1339GAT) );
  NOR2_X1 U582 ( .A1(n532), .A2(n515), .ZN(n516) );
  NAND2_X1 U583 ( .A1(n517), .A2(n516), .ZN(n527) );
  NOR2_X1 U584 ( .A1(n564), .A2(n527), .ZN(n519) );
  XNOR2_X1 U585 ( .A(KEYINPUT112), .B(KEYINPUT113), .ZN(n518) );
  XNOR2_X1 U586 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U587 ( .A(G113GAT), .B(n520), .ZN(G1340GAT) );
  NOR2_X1 U588 ( .A1(n550), .A2(n527), .ZN(n522) );
  XNOR2_X1 U589 ( .A(KEYINPUT114), .B(KEYINPUT49), .ZN(n521) );
  XNOR2_X1 U590 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U591 ( .A(G120GAT), .B(n523), .ZN(G1341GAT) );
  NOR2_X1 U592 ( .A1(n572), .A2(n527), .ZN(n525) );
  XNOR2_X1 U593 ( .A(KEYINPUT50), .B(KEYINPUT115), .ZN(n524) );
  XNOR2_X1 U594 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U595 ( .A(G127GAT), .B(n526), .ZN(G1342GAT) );
  NOR2_X1 U596 ( .A1(n557), .A2(n527), .ZN(n529) );
  XNOR2_X1 U597 ( .A(KEYINPUT116), .B(KEYINPUT51), .ZN(n528) );
  XNOR2_X1 U598 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U599 ( .A(G134GAT), .B(n530), .ZN(G1343GAT) );
  NOR2_X1 U600 ( .A1(n532), .A2(n531), .ZN(n533) );
  NAND2_X1 U601 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U602 ( .A(n535), .B(KEYINPUT117), .ZN(n544) );
  NAND2_X1 U603 ( .A1(n536), .A2(n544), .ZN(n537) );
  XNOR2_X1 U604 ( .A(n537), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n540) );
  NAND2_X1 U606 ( .A1(n544), .A2(n538), .ZN(n539) );
  XNOR2_X1 U607 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U608 ( .A(G148GAT), .B(n541), .ZN(G1345GAT) );
  NAND2_X1 U609 ( .A1(n544), .A2(n542), .ZN(n543) );
  XNOR2_X1 U610 ( .A(n543), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U611 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U612 ( .A(G162GAT), .B(n546), .ZN(G1347GAT) );
  XOR2_X1 U613 ( .A(KEYINPUT56), .B(KEYINPUT120), .Z(n548) );
  XNOR2_X1 U614 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n547) );
  XNOR2_X1 U615 ( .A(n548), .B(n547), .ZN(n552) );
  NOR2_X1 U616 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U617 ( .A(n552), .B(n551), .Z(G1349GAT) );
  NOR2_X1 U618 ( .A1(n572), .A2(n549), .ZN(n554) );
  XNOR2_X1 U619 ( .A(G183GAT), .B(KEYINPUT121), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n554), .B(n553), .ZN(G1350GAT) );
  XOR2_X1 U621 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n556) );
  XNOR2_X1 U622 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n555) );
  XNOR2_X1 U623 ( .A(n556), .B(n555), .ZN(n559) );
  NOR2_X1 U624 ( .A1(n557), .A2(n549), .ZN(n558) );
  XOR2_X1 U625 ( .A(n559), .B(n558), .Z(G1351GAT) );
  XOR2_X1 U626 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n561) );
  XNOR2_X1 U627 ( .A(G197GAT), .B(KEYINPUT124), .ZN(n560) );
  XNOR2_X1 U628 ( .A(n561), .B(n560), .ZN(n566) );
  NAND2_X1 U629 ( .A1(n563), .A2(n562), .ZN(n575) );
  NOR2_X1 U630 ( .A1(n564), .A2(n575), .ZN(n565) );
  XOR2_X1 U631 ( .A(n566), .B(n565), .Z(G1352GAT) );
  NOR2_X1 U632 ( .A1(n575), .A2(n567), .ZN(n571) );
  XOR2_X1 U633 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n569) );
  XNOR2_X1 U634 ( .A(G204GAT), .B(KEYINPUT126), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(G1353GAT) );
  NOR2_X1 U637 ( .A1(n572), .A2(n575), .ZN(n574) );
  XNOR2_X1 U638 ( .A(G211GAT), .B(KEYINPUT127), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(G1354GAT) );
  NOR2_X1 U640 ( .A1(n576), .A2(n575), .ZN(n577) );
  XOR2_X1 U641 ( .A(KEYINPUT62), .B(n577), .Z(n578) );
  XNOR2_X1 U642 ( .A(G218GAT), .B(n578), .ZN(G1355GAT) );
endmodule

