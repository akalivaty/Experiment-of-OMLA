

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751;

  NAND2_X1 U377 ( .A1(n610), .A2(n609), .ZN(n382) );
  XNOR2_X1 U378 ( .A(n354), .B(n408), .ZN(n605) );
  NAND2_X1 U379 ( .A1(n376), .A2(n667), .ZN(n354) );
  XNOR2_X1 U380 ( .A(n556), .B(n555), .ZN(n749) );
  BUF_X1 U381 ( .A(n651), .Z(n657) );
  NOR2_X1 U382 ( .A1(n680), .A2(n681), .ZN(n553) );
  XNOR2_X1 U383 ( .A(n392), .B(n478), .ZN(n734) );
  OR2_X1 U384 ( .A1(n611), .A2(G902), .ZN(n457) );
  NOR2_X2 U385 ( .A1(n628), .A2(n725), .ZN(n630) );
  NOR2_X2 U386 ( .A1(n620), .A2(n725), .ZN(n622) );
  NOR2_X1 U387 ( .A1(n658), .A2(n652), .ZN(n682) );
  INV_X1 U388 ( .A(G953), .ZN(n742) );
  INV_X1 U389 ( .A(n660), .ZN(n658) );
  XNOR2_X2 U390 ( .A(n606), .B(KEYINPUT84), .ZN(n741) );
  BUF_X1 U391 ( .A(n623), .Z(n721) );
  AND2_X1 U392 ( .A1(n670), .A2(n603), .ZN(n631) );
  NOR2_X1 U393 ( .A1(n404), .A2(n406), .ZN(n403) );
  AND2_X1 U394 ( .A1(n371), .A2(n398), .ZN(n370) );
  XNOR2_X1 U395 ( .A(n394), .B(n393), .ZN(n588) );
  XNOR2_X1 U396 ( .A(n362), .B(n420), .ZN(n506) );
  XNOR2_X1 U397 ( .A(n356), .B(n418), .ZN(n477) );
  XNOR2_X1 U398 ( .A(n419), .B(G128), .ZN(n362) );
  XNOR2_X2 U399 ( .A(n575), .B(KEYINPUT35), .ZN(n750) );
  AND2_X1 U400 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U401 ( .A(n405), .B(KEYINPUT79), .ZN(n404) );
  XNOR2_X1 U402 ( .A(n656), .B(n407), .ZN(n406) );
  NAND2_X1 U403 ( .A1(n380), .A2(n378), .ZN(n377) );
  XNOR2_X1 U404 ( .A(n559), .B(n379), .ZN(n378) );
  AND2_X1 U405 ( .A1(n551), .A2(n666), .ZN(n380) );
  INV_X1 U406 ( .A(KEYINPUT46), .ZN(n379) );
  XNOR2_X1 U407 ( .A(n413), .B(n412), .ZN(n633) );
  XNOR2_X1 U408 ( .A(n506), .B(n411), .ZN(n412) );
  XNOR2_X1 U409 ( .A(n477), .B(n414), .ZN(n413) );
  XNOR2_X1 U410 ( .A(n423), .B(n360), .ZN(n411) );
  INV_X1 U411 ( .A(KEYINPUT86), .ZN(n408) );
  XNOR2_X1 U412 ( .A(n377), .B(n361), .ZN(n376) );
  INV_X1 U413 ( .A(G143), .ZN(n419) );
  XNOR2_X1 U414 ( .A(n531), .B(KEYINPUT1), .ZN(n690) );
  AND2_X1 U415 ( .A1(n524), .A2(n692), .ZN(n374) );
  XNOR2_X1 U416 ( .A(n509), .B(n395), .ZN(n533) );
  INV_X1 U417 ( .A(KEYINPUT19), .ZN(n395) );
  XNOR2_X1 U418 ( .A(n435), .B(n441), .ZN(n739) );
  XNOR2_X1 U419 ( .A(n506), .B(n421), .ZN(n435) );
  XNOR2_X1 U420 ( .A(n734), .B(n384), .ZN(n624) );
  XNOR2_X1 U421 ( .A(n389), .B(n385), .ZN(n384) );
  XNOR2_X1 U422 ( .A(n391), .B(n390), .ZN(n389) );
  XNOR2_X1 U423 ( .A(n388), .B(n386), .ZN(n385) );
  XNOR2_X1 U424 ( .A(n482), .B(KEYINPUT39), .ZN(n523) );
  NOR2_X1 U425 ( .A1(n596), .A2(n545), .ZN(n546) );
  NAND2_X1 U426 ( .A1(n688), .A2(n400), .ZN(n371) );
  XNOR2_X1 U427 ( .A(n520), .B(n519), .ZN(n582) );
  XNOR2_X1 U428 ( .A(n518), .B(KEYINPUT70), .ZN(n519) );
  XNOR2_X1 U429 ( .A(n401), .B(KEYINPUT71), .ZN(n551) );
  NAND2_X1 U430 ( .A1(n403), .A2(n402), .ZN(n401) );
  XNOR2_X1 U431 ( .A(n415), .B(n421), .ZN(n414) );
  XNOR2_X1 U432 ( .A(n424), .B(n422), .ZN(n415) );
  XNOR2_X1 U433 ( .A(G116), .B(G146), .ZN(n424) );
  NOR2_X1 U434 ( .A1(G953), .A2(G237), .ZN(n489) );
  AND2_X1 U435 ( .A1(n367), .A2(n365), .ZN(n364) );
  AND2_X1 U436 ( .A1(n417), .A2(n366), .ZN(n365) );
  NOR2_X1 U437 ( .A1(n585), .A2(KEYINPUT44), .ZN(n368) );
  XNOR2_X1 U438 ( .A(n381), .B(KEYINPUT10), .ZN(n483) );
  XOR2_X1 U439 ( .A(KEYINPUT8), .B(KEYINPUT66), .Z(n446) );
  BUF_X1 U440 ( .A(n483), .Z(n740) );
  INV_X1 U441 ( .A(KEYINPUT18), .ZN(n387) );
  XNOR2_X1 U442 ( .A(n472), .B(n475), .ZN(n391) );
  XOR2_X1 U443 ( .A(KEYINPUT91), .B(KEYINPUT73), .Z(n475) );
  XNOR2_X1 U444 ( .A(n473), .B(n476), .ZN(n390) );
  OR2_X1 U445 ( .A1(n730), .A2(n601), .ZN(n670) );
  NAND2_X1 U446 ( .A1(G234), .A2(G237), .ZN(n462) );
  INV_X1 U447 ( .A(G134), .ZN(n420) );
  XOR2_X1 U448 ( .A(KEYINPUT69), .B(G110), .Z(n472) );
  XNOR2_X1 U449 ( .A(G101), .B(G146), .ZN(n429) );
  XOR2_X1 U450 ( .A(G107), .B(G104), .Z(n430) );
  INV_X1 U451 ( .A(KEYINPUT0), .ZN(n393) );
  NOR2_X1 U452 ( .A1(n533), .A2(n359), .ZN(n394) );
  AND2_X1 U453 ( .A1(n471), .A2(n470), .ZN(n541) );
  XNOR2_X1 U454 ( .A(n375), .B(n469), .ZN(n470) );
  OR2_X1 U455 ( .A1(n714), .A2(G902), .ZN(n372) );
  AND2_X1 U456 ( .A1(n595), .A2(n692), .ZN(n689) );
  XNOR2_X1 U457 ( .A(n477), .B(KEYINPUT16), .ZN(n392) );
  AND2_X1 U458 ( .A1(n614), .A2(G953), .ZN(n725) );
  XNOR2_X1 U459 ( .A(n410), .B(n355), .ZN(n558) );
  NOR2_X1 U460 ( .A1(n560), .A2(n563), .ZN(n549) );
  NAND2_X1 U461 ( .A1(n396), .A2(n370), .ZN(n399) );
  XNOR2_X1 U462 ( .A(n583), .B(KEYINPUT32), .ZN(n751) );
  XOR2_X1 U463 ( .A(KEYINPUT107), .B(KEYINPUT40), .Z(n355) );
  XOR2_X1 U464 ( .A(G101), .B(G113), .Z(n356) );
  XOR2_X1 U465 ( .A(KEYINPUT78), .B(n567), .Z(n357) );
  NAND2_X1 U466 ( .A1(n531), .A2(n689), .ZN(n358) );
  AND2_X1 U467 ( .A1(n513), .A2(n512), .ZN(n359) );
  AND2_X1 U468 ( .A1(n489), .A2(G210), .ZN(n360) );
  INV_X1 U469 ( .A(KEYINPUT34), .ZN(n400) );
  XOR2_X1 U470 ( .A(KEYINPUT88), .B(KEYINPUT48), .Z(n361) );
  XNOR2_X1 U471 ( .A(n362), .B(n474), .ZN(n388) );
  NAND2_X1 U472 ( .A1(n364), .A2(n363), .ZN(n383) );
  NAND2_X1 U473 ( .A1(n750), .A2(KEYINPUT44), .ZN(n363) );
  NAND2_X1 U474 ( .A1(n585), .A2(KEYINPUT44), .ZN(n366) );
  NAND2_X1 U475 ( .A1(n369), .A2(n368), .ZN(n367) );
  INV_X1 U476 ( .A(n750), .ZN(n369) );
  XNOR2_X2 U477 ( .A(n571), .B(KEYINPUT33), .ZN(n688) );
  INV_X1 U478 ( .A(n690), .ZN(n568) );
  XNOR2_X2 U479 ( .A(n372), .B(G469), .ZN(n531) );
  NAND2_X1 U480 ( .A1(n531), .A2(n373), .ZN(n375) );
  AND2_X1 U481 ( .A1(n595), .A2(n374), .ZN(n373) );
  XNOR2_X1 U482 ( .A(n381), .B(n387), .ZN(n386) );
  XNOR2_X2 U483 ( .A(G146), .B(G125), .ZN(n381) );
  AND2_X2 U484 ( .A1(n382), .A2(n631), .ZN(n623) );
  NAND2_X1 U485 ( .A1(n632), .A2(n382), .ZN(n637) );
  XNOR2_X2 U486 ( .A(n383), .B(n416), .ZN(n730) );
  OR2_X1 U487 ( .A1(n397), .A2(n688), .ZN(n396) );
  NAND2_X1 U488 ( .A1(n591), .A2(KEYINPUT34), .ZN(n397) );
  OR2_X1 U489 ( .A1(n591), .A2(KEYINPUT34), .ZN(n398) );
  NAND2_X1 U490 ( .A1(n399), .A2(n574), .ZN(n575) );
  NAND2_X1 U491 ( .A1(n536), .A2(n535), .ZN(n402) );
  NAND2_X1 U492 ( .A1(n682), .A2(KEYINPUT47), .ZN(n405) );
  INV_X1 U493 ( .A(KEYINPUT80), .ZN(n407) );
  NAND2_X1 U494 ( .A1(n605), .A2(n357), .ZN(n601) );
  NAND2_X1 U495 ( .A1(n624), .A2(n602), .ZN(n409) );
  XNOR2_X1 U496 ( .A(n537), .B(n481), .ZN(n678) );
  XNOR2_X2 U497 ( .A(n409), .B(n480), .ZN(n537) );
  INV_X1 U498 ( .A(n558), .ZN(n552) );
  NAND2_X1 U499 ( .A1(n523), .A2(n658), .ZN(n410) );
  XOR2_X1 U500 ( .A(n600), .B(KEYINPUT45), .Z(n416) );
  XNOR2_X1 U501 ( .A(n527), .B(KEYINPUT67), .ZN(n544) );
  AND2_X1 U502 ( .A1(n599), .A2(n642), .ZN(n417) );
  INV_X1 U503 ( .A(KEYINPUT47), .ZN(n534) );
  INV_X1 U504 ( .A(G137), .ZN(n422) );
  NAND2_X1 U505 ( .A1(n526), .A2(n525), .ZN(n527) );
  INV_X1 U506 ( .A(n730), .ZN(n607) );
  INV_X1 U507 ( .A(KEYINPUT2), .ZN(n609) );
  INV_X1 U508 ( .A(KEYINPUT94), .ZN(n572) );
  XNOR2_X1 U509 ( .A(n635), .B(n634), .ZN(n636) );
  BUF_X1 U510 ( .A(n526), .Z(n576) );
  XNOR2_X1 U511 ( .A(G119), .B(KEYINPUT3), .ZN(n418) );
  XNOR2_X1 U512 ( .A(KEYINPUT4), .B(G131), .ZN(n421) );
  XOR2_X1 U513 ( .A(KEYINPUT5), .B(KEYINPUT96), .Z(n423) );
  NOR2_X1 U514 ( .A1(G902), .A2(n633), .ZN(n426) );
  XNOR2_X1 U515 ( .A(G472), .B(KEYINPUT97), .ZN(n425) );
  XNOR2_X1 U516 ( .A(n426), .B(n425), .ZN(n542) );
  XNOR2_X1 U517 ( .A(n542), .B(KEYINPUT104), .ZN(n528) );
  OR2_X1 U518 ( .A1(G237), .A2(G902), .ZN(n479) );
  NAND2_X1 U519 ( .A1(G214), .A2(n479), .ZN(n677) );
  NAND2_X1 U520 ( .A1(n528), .A2(n677), .ZN(n428) );
  INV_X1 U521 ( .A(KEYINPUT30), .ZN(n427) );
  XNOR2_X1 U522 ( .A(n428), .B(n427), .ZN(n471) );
  XNOR2_X1 U523 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U524 ( .A(n472), .B(n431), .Z(n433) );
  NAND2_X1 U525 ( .A1(G227), .A2(n742), .ZN(n432) );
  XNOR2_X1 U526 ( .A(n433), .B(n432), .ZN(n436) );
  INV_X1 U527 ( .A(G140), .ZN(n434) );
  XNOR2_X1 U528 ( .A(n434), .B(G137), .ZN(n441) );
  XNOR2_X1 U529 ( .A(n436), .B(n739), .ZN(n714) );
  XNOR2_X1 U530 ( .A(G110), .B(KEYINPUT24), .ZN(n438) );
  XNOR2_X1 U531 ( .A(KEYINPUT68), .B(KEYINPUT95), .ZN(n437) );
  XNOR2_X1 U532 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U533 ( .A(n483), .B(n439), .ZN(n444) );
  XNOR2_X1 U534 ( .A(G128), .B(G119), .ZN(n440) );
  XNOR2_X1 U535 ( .A(n440), .B(KEYINPUT23), .ZN(n442) );
  XNOR2_X1 U536 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U537 ( .A(n444), .B(n443), .ZN(n450) );
  NAND2_X1 U538 ( .A1(G234), .A2(n742), .ZN(n445) );
  XNOR2_X1 U539 ( .A(n446), .B(n445), .ZN(n448) );
  INV_X1 U540 ( .A(KEYINPUT81), .ZN(n447) );
  XNOR2_X1 U541 ( .A(n448), .B(n447), .ZN(n499) );
  NAND2_X1 U542 ( .A1(n499), .A2(G221), .ZN(n449) );
  XNOR2_X1 U543 ( .A(n450), .B(n449), .ZN(n611) );
  XNOR2_X1 U544 ( .A(G902), .B(KEYINPUT15), .ZN(n602) );
  NAND2_X1 U545 ( .A1(n602), .A2(G234), .ZN(n452) );
  INV_X1 U546 ( .A(KEYINPUT20), .ZN(n451) );
  XNOR2_X1 U547 ( .A(n452), .B(n451), .ZN(n459) );
  INV_X1 U548 ( .A(G217), .ZN(n453) );
  OR2_X1 U549 ( .A1(n459), .A2(n453), .ZN(n455) );
  INV_X1 U550 ( .A(KEYINPUT25), .ZN(n454) );
  XNOR2_X1 U551 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X2 U552 ( .A(n457), .B(n456), .ZN(n595) );
  INV_X1 U553 ( .A(G221), .ZN(n458) );
  OR2_X1 U554 ( .A1(n459), .A2(n458), .ZN(n461) );
  INV_X1 U555 ( .A(KEYINPUT21), .ZN(n460) );
  XNOR2_X1 U556 ( .A(n461), .B(n460), .ZN(n692) );
  XNOR2_X1 U557 ( .A(KEYINPUT14), .B(n462), .ZN(n465) );
  NAND2_X1 U558 ( .A1(G952), .A2(n465), .ZN(n463) );
  XNOR2_X1 U559 ( .A(KEYINPUT92), .B(n463), .ZN(n706) );
  NOR2_X1 U560 ( .A1(n706), .A2(G953), .ZN(n464) );
  XNOR2_X1 U561 ( .A(n464), .B(KEYINPUT93), .ZN(n512) );
  NAND2_X1 U562 ( .A1(G902), .A2(n465), .ZN(n510) );
  NOR2_X1 U563 ( .A1(G900), .A2(n510), .ZN(n466) );
  NAND2_X1 U564 ( .A1(n466), .A2(G953), .ZN(n467) );
  AND2_X1 U565 ( .A1(n512), .A2(n467), .ZN(n468) );
  XNOR2_X1 U566 ( .A(n468), .B(KEYINPUT77), .ZN(n524) );
  INV_X1 U567 ( .A(KEYINPUT72), .ZN(n469) );
  AND2_X1 U568 ( .A1(G224), .A2(n742), .ZN(n473) );
  XNOR2_X1 U569 ( .A(KEYINPUT4), .B(KEYINPUT75), .ZN(n474) );
  XNOR2_X1 U570 ( .A(KEYINPUT74), .B(KEYINPUT17), .ZN(n476) );
  XOR2_X1 U571 ( .A(G116), .B(G107), .Z(n500) );
  XOR2_X1 U572 ( .A(G122), .B(G104), .Z(n493) );
  XOR2_X1 U573 ( .A(n500), .B(n493), .Z(n478) );
  AND2_X1 U574 ( .A1(G210), .A2(n479), .ZN(n480) );
  INV_X1 U575 ( .A(KEYINPUT38), .ZN(n481) );
  NAND2_X1 U576 ( .A1(n541), .A2(n678), .ZN(n482) );
  XOR2_X1 U577 ( .A(KEYINPUT12), .B(KEYINPUT99), .Z(n485) );
  XNOR2_X1 U578 ( .A(G131), .B(G140), .ZN(n484) );
  XNOR2_X1 U579 ( .A(n485), .B(n484), .ZN(n487) );
  XNOR2_X1 U580 ( .A(G113), .B(G143), .ZN(n486) );
  XNOR2_X1 U581 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U582 ( .A(n740), .B(n488), .ZN(n495) );
  XOR2_X1 U583 ( .A(KEYINPUT11), .B(KEYINPUT100), .Z(n491) );
  NAND2_X1 U584 ( .A1(G214), .A2(n489), .ZN(n490) );
  XNOR2_X1 U585 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U586 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U587 ( .A(n495), .B(n494), .ZN(n617) );
  INV_X1 U588 ( .A(G902), .ZN(n496) );
  NAND2_X1 U589 ( .A1(n617), .A2(n496), .ZN(n498) );
  XNOR2_X1 U590 ( .A(KEYINPUT13), .B(G475), .ZN(n497) );
  XNOR2_X1 U591 ( .A(n498), .B(n497), .ZN(n539) );
  XOR2_X1 U592 ( .A(KEYINPUT101), .B(G478), .Z(n508) );
  NAND2_X1 U593 ( .A1(n499), .A2(G217), .ZN(n504) );
  XOR2_X1 U594 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n502) );
  XNOR2_X1 U595 ( .A(G122), .B(n500), .ZN(n501) );
  XNOR2_X1 U596 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U597 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U598 ( .A(n506), .B(n505), .ZN(n722) );
  NOR2_X1 U599 ( .A1(G902), .A2(n722), .ZN(n507) );
  XNOR2_X1 U600 ( .A(n508), .B(n507), .ZN(n538) );
  INV_X1 U601 ( .A(n538), .ZN(n522) );
  NAND2_X1 U602 ( .A1(n539), .A2(n522), .ZN(n663) );
  INV_X1 U603 ( .A(n663), .ZN(n652) );
  AND2_X1 U604 ( .A1(n523), .A2(n652), .ZN(n566) );
  XOR2_X1 U605 ( .A(G134), .B(n566), .Z(G36) );
  INV_X1 U606 ( .A(n595), .ZN(n526) );
  NAND2_X1 U607 ( .A1(n677), .A2(n537), .ZN(n509) );
  NOR2_X1 U608 ( .A1(G898), .A2(n742), .ZN(n736) );
  INV_X1 U609 ( .A(n510), .ZN(n511) );
  NAND2_X1 U610 ( .A1(n736), .A2(n511), .ZN(n513) );
  INV_X1 U611 ( .A(n588), .ZN(n517) );
  INV_X1 U612 ( .A(n692), .ZN(n514) );
  NAND2_X1 U613 ( .A1(n539), .A2(n538), .ZN(n680) );
  NOR2_X1 U614 ( .A1(n514), .A2(n680), .ZN(n515) );
  XNOR2_X1 U615 ( .A(KEYINPUT102), .B(n515), .ZN(n516) );
  NAND2_X1 U616 ( .A1(n517), .A2(n516), .ZN(n520) );
  XOR2_X1 U617 ( .A(KEYINPUT22), .B(KEYINPUT64), .Z(n518) );
  NAND2_X1 U618 ( .A1(n568), .A2(n582), .ZN(n598) );
  NOR2_X1 U619 ( .A1(n528), .A2(n598), .ZN(n521) );
  NAND2_X1 U620 ( .A1(n576), .A2(n521), .ZN(n584) );
  XNOR2_X1 U621 ( .A(n584), .B(G110), .ZN(G12) );
  OR2_X1 U622 ( .A1(n539), .A2(n522), .ZN(n660) );
  XOR2_X1 U623 ( .A(G131), .B(n552), .Z(G33) );
  AND2_X1 U624 ( .A1(n524), .A2(n692), .ZN(n525) );
  NAND2_X1 U625 ( .A1(n544), .A2(n528), .ZN(n530) );
  INV_X1 U626 ( .A(KEYINPUT28), .ZN(n529) );
  XNOR2_X1 U627 ( .A(n530), .B(n529), .ZN(n532) );
  NAND2_X1 U628 ( .A1(n532), .A2(n531), .ZN(n554) );
  NOR2_X2 U629 ( .A1(n554), .A2(n533), .ZN(n651) );
  XNOR2_X1 U630 ( .A(n651), .B(n534), .ZN(n536) );
  NAND2_X1 U631 ( .A1(n657), .A2(n682), .ZN(n535) );
  INV_X1 U632 ( .A(n537), .ZN(n563) );
  OR2_X1 U633 ( .A1(n539), .A2(n538), .ZN(n573) );
  NOR2_X1 U634 ( .A1(n563), .A2(n573), .ZN(n540) );
  NAND2_X1 U635 ( .A1(n541), .A2(n540), .ZN(n656) );
  INV_X1 U636 ( .A(n542), .ZN(n543) );
  INV_X2 U637 ( .A(n543), .ZN(n695) );
  XNOR2_X2 U638 ( .A(KEYINPUT6), .B(n695), .ZN(n596) );
  INV_X1 U639 ( .A(n544), .ZN(n545) );
  XOR2_X1 U640 ( .A(KEYINPUT106), .B(n546), .Z(n547) );
  NOR2_X1 U641 ( .A1(n660), .A2(n547), .ZN(n548) );
  NAND2_X1 U642 ( .A1(n548), .A2(n677), .ZN(n560) );
  XNOR2_X1 U643 ( .A(n549), .B(KEYINPUT36), .ZN(n550) );
  XNOR2_X1 U644 ( .A(n568), .B(KEYINPUT89), .ZN(n577) );
  NAND2_X1 U645 ( .A1(n550), .A2(n577), .ZN(n666) );
  NAND2_X1 U646 ( .A1(n678), .A2(n677), .ZN(n681) );
  XNOR2_X1 U647 ( .A(KEYINPUT41), .B(n553), .ZN(n702) );
  NOR2_X1 U648 ( .A1(n702), .A2(n554), .ZN(n556) );
  XNOR2_X1 U649 ( .A(KEYINPUT108), .B(KEYINPUT42), .ZN(n555) );
  INV_X1 U650 ( .A(n749), .ZN(n557) );
  NAND2_X1 U651 ( .A1(n558), .A2(n557), .ZN(n559) );
  INV_X1 U652 ( .A(n560), .ZN(n561) );
  NAND2_X1 U653 ( .A1(n568), .A2(n561), .ZN(n562) );
  XNOR2_X1 U654 ( .A(n562), .B(KEYINPUT43), .ZN(n564) );
  NAND2_X1 U655 ( .A1(n564), .A2(n563), .ZN(n667) );
  INV_X1 U656 ( .A(n566), .ZN(n604) );
  NAND2_X1 U657 ( .A1(n604), .A2(KEYINPUT2), .ZN(n567) );
  NAND2_X1 U658 ( .A1(n690), .A2(n689), .ZN(n586) );
  XNOR2_X1 U659 ( .A(n586), .B(KEYINPUT105), .ZN(n570) );
  INV_X1 U660 ( .A(n596), .ZN(n569) );
  XNOR2_X1 U661 ( .A(n588), .B(n572), .ZN(n591) );
  INV_X1 U662 ( .A(n573), .ZN(n574) );
  XNOR2_X1 U663 ( .A(n596), .B(KEYINPUT76), .ZN(n580) );
  NAND2_X1 U664 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U665 ( .A(KEYINPUT103), .B(n578), .ZN(n579) );
  AND2_X1 U666 ( .A1(n580), .A2(n579), .ZN(n581) );
  NAND2_X1 U667 ( .A1(n582), .A2(n581), .ZN(n583) );
  NAND2_X1 U668 ( .A1(n751), .A2(n584), .ZN(n585) );
  INV_X1 U669 ( .A(n586), .ZN(n587) );
  NAND2_X1 U670 ( .A1(n587), .A2(n695), .ZN(n698) );
  NOR2_X1 U671 ( .A1(n698), .A2(n588), .ZN(n589) );
  XNOR2_X1 U672 ( .A(n589), .B(KEYINPUT31), .ZN(n662) );
  NOR2_X1 U673 ( .A1(n358), .A2(n695), .ZN(n590) );
  NAND2_X1 U674 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U675 ( .A(KEYINPUT98), .B(n592), .ZN(n648) );
  NAND2_X1 U676 ( .A1(n662), .A2(n648), .ZN(n594) );
  INV_X1 U677 ( .A(n682), .ZN(n593) );
  NAND2_X1 U678 ( .A1(n594), .A2(n593), .ZN(n599) );
  NAND2_X1 U679 ( .A1(n596), .A2(n595), .ZN(n597) );
  OR2_X1 U680 ( .A1(n598), .A2(n597), .ZN(n642) );
  INV_X1 U681 ( .A(KEYINPUT85), .ZN(n600) );
  INV_X1 U682 ( .A(n602), .ZN(n603) );
  NAND2_X1 U683 ( .A1(n605), .A2(n604), .ZN(n606) );
  INV_X1 U684 ( .A(n741), .ZN(n608) );
  NAND2_X1 U685 ( .A1(n608), .A2(n607), .ZN(n610) );
  NAND2_X1 U686 ( .A1(n721), .A2(G217), .ZN(n613) );
  XNOR2_X1 U687 ( .A(n611), .B(KEYINPUT124), .ZN(n612) );
  XNOR2_X1 U688 ( .A(n613), .B(n612), .ZN(n615) );
  INV_X1 U689 ( .A(G952), .ZN(n614) );
  NOR2_X1 U690 ( .A1(n615), .A2(n725), .ZN(G66) );
  NAND2_X1 U691 ( .A1(n623), .A2(G475), .ZN(n619) );
  XOR2_X1 U692 ( .A(KEYINPUT65), .B(KEYINPUT59), .Z(n616) );
  XNOR2_X1 U693 ( .A(n617), .B(n616), .ZN(n618) );
  XNOR2_X1 U694 ( .A(n619), .B(n618), .ZN(n620) );
  XOR2_X1 U695 ( .A(KEYINPUT123), .B(KEYINPUT60), .Z(n621) );
  XNOR2_X1 U696 ( .A(n622), .B(n621), .ZN(G60) );
  NAND2_X1 U697 ( .A1(n623), .A2(G210), .ZN(n627) );
  XNOR2_X1 U698 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n625) );
  XNOR2_X1 U699 ( .A(n624), .B(n625), .ZN(n626) );
  XNOR2_X1 U700 ( .A(n627), .B(n626), .ZN(n628) );
  XOR2_X1 U701 ( .A(KEYINPUT87), .B(KEYINPUT56), .Z(n629) );
  XNOR2_X1 U702 ( .A(n630), .B(n629), .ZN(G51) );
  AND2_X1 U703 ( .A1(n631), .A2(G472), .ZN(n632) );
  XNOR2_X1 U704 ( .A(n633), .B(KEYINPUT109), .ZN(n635) );
  XOR2_X1 U705 ( .A(KEYINPUT62), .B(KEYINPUT110), .Z(n634) );
  XNOR2_X1 U706 ( .A(n637), .B(n636), .ZN(n638) );
  NOR2_X1 U707 ( .A1(n725), .A2(n638), .ZN(n641) );
  XNOR2_X1 U708 ( .A(KEYINPUT90), .B(KEYINPUT111), .ZN(n639) );
  XNOR2_X1 U709 ( .A(n639), .B(KEYINPUT63), .ZN(n640) );
  XNOR2_X1 U710 ( .A(n641), .B(n640), .ZN(G57) );
  XNOR2_X1 U711 ( .A(G101), .B(KEYINPUT112), .ZN(n643) );
  XNOR2_X1 U712 ( .A(n643), .B(n642), .ZN(G3) );
  NOR2_X1 U713 ( .A1(n648), .A2(n660), .ZN(n645) );
  XNOR2_X1 U714 ( .A(G104), .B(KEYINPUT113), .ZN(n644) );
  XNOR2_X1 U715 ( .A(n645), .B(n644), .ZN(G6) );
  XOR2_X1 U716 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n647) );
  XNOR2_X1 U717 ( .A(G107), .B(KEYINPUT114), .ZN(n646) );
  XNOR2_X1 U718 ( .A(n647), .B(n646), .ZN(n650) );
  NOR2_X1 U719 ( .A1(n648), .A2(n663), .ZN(n649) );
  XOR2_X1 U720 ( .A(n650), .B(n649), .Z(G9) );
  XOR2_X1 U721 ( .A(G128), .B(KEYINPUT29), .Z(n654) );
  NAND2_X1 U722 ( .A1(n657), .A2(n652), .ZN(n653) );
  XNOR2_X1 U723 ( .A(n654), .B(n653), .ZN(G30) );
  XOR2_X1 U724 ( .A(G143), .B(KEYINPUT115), .Z(n655) );
  XNOR2_X1 U725 ( .A(n656), .B(n655), .ZN(G45) );
  NAND2_X1 U726 ( .A1(n658), .A2(n657), .ZN(n659) );
  XNOR2_X1 U727 ( .A(G146), .B(n659), .ZN(G48) );
  NOR2_X1 U728 ( .A1(n660), .A2(n662), .ZN(n661) );
  XOR2_X1 U729 ( .A(G113), .B(n661), .Z(G15) );
  NOR2_X1 U730 ( .A1(n663), .A2(n662), .ZN(n664) );
  XOR2_X1 U731 ( .A(G116), .B(n664), .Z(G18) );
  XOR2_X1 U732 ( .A(G125), .B(KEYINPUT37), .Z(n665) );
  XNOR2_X1 U733 ( .A(n666), .B(n665), .ZN(G27) );
  XNOR2_X1 U734 ( .A(G140), .B(n667), .ZN(G42) );
  NAND2_X1 U735 ( .A1(n609), .A2(n730), .ZN(n668) );
  XNOR2_X1 U736 ( .A(n668), .B(KEYINPUT82), .ZN(n669) );
  NAND2_X1 U737 ( .A1(n670), .A2(n669), .ZN(n673) );
  NAND2_X1 U738 ( .A1(n741), .A2(n609), .ZN(n671) );
  XNOR2_X1 U739 ( .A(n671), .B(KEYINPUT83), .ZN(n672) );
  NOR2_X1 U740 ( .A1(n673), .A2(n672), .ZN(n676) );
  NOR2_X1 U741 ( .A1(n688), .A2(n702), .ZN(n674) );
  XOR2_X1 U742 ( .A(KEYINPUT119), .B(n674), .Z(n675) );
  NOR2_X1 U743 ( .A1(n676), .A2(n675), .ZN(n710) );
  NOR2_X1 U744 ( .A1(n678), .A2(n677), .ZN(n679) );
  NOR2_X1 U745 ( .A1(n680), .A2(n679), .ZN(n685) );
  NOR2_X1 U746 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U747 ( .A(n683), .B(KEYINPUT116), .ZN(n684) );
  NOR2_X1 U748 ( .A1(n685), .A2(n684), .ZN(n686) );
  XOR2_X1 U749 ( .A(KEYINPUT117), .B(n686), .Z(n687) );
  NOR2_X1 U750 ( .A1(n688), .A2(n687), .ZN(n704) );
  NOR2_X1 U751 ( .A1(n690), .A2(n689), .ZN(n691) );
  XOR2_X1 U752 ( .A(KEYINPUT50), .B(n691), .Z(n697) );
  NOR2_X1 U753 ( .A1(n595), .A2(n692), .ZN(n693) );
  XOR2_X1 U754 ( .A(KEYINPUT49), .B(n693), .Z(n694) );
  NOR2_X1 U755 ( .A1(n695), .A2(n694), .ZN(n696) );
  NAND2_X1 U756 ( .A1(n697), .A2(n696), .ZN(n699) );
  NAND2_X1 U757 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U758 ( .A(KEYINPUT51), .B(n700), .ZN(n701) );
  NOR2_X1 U759 ( .A1(n702), .A2(n701), .ZN(n703) );
  NOR2_X1 U760 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U761 ( .A(KEYINPUT52), .B(n705), .ZN(n707) );
  NOR2_X1 U762 ( .A1(n707), .A2(n706), .ZN(n708) );
  XOR2_X1 U763 ( .A(KEYINPUT118), .B(n708), .Z(n709) );
  NAND2_X1 U764 ( .A1(n710), .A2(n709), .ZN(n711) );
  NOR2_X1 U765 ( .A1(G953), .A2(n711), .ZN(n713) );
  XNOR2_X1 U766 ( .A(KEYINPUT53), .B(KEYINPUT120), .ZN(n712) );
  XNOR2_X1 U767 ( .A(n713), .B(n712), .ZN(G75) );
  NAND2_X1 U768 ( .A1(n721), .A2(G469), .ZN(n719) );
  XOR2_X1 U769 ( .A(KEYINPUT122), .B(KEYINPUT121), .Z(n716) );
  XNOR2_X1 U770 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n715) );
  XNOR2_X1 U771 ( .A(n716), .B(n715), .ZN(n717) );
  XOR2_X1 U772 ( .A(n714), .B(n717), .Z(n718) );
  XNOR2_X1 U773 ( .A(n719), .B(n718), .ZN(n720) );
  NOR2_X1 U774 ( .A1(n725), .A2(n720), .ZN(G54) );
  NAND2_X1 U775 ( .A1(n721), .A2(G478), .ZN(n723) );
  XNOR2_X1 U776 ( .A(n723), .B(n722), .ZN(n724) );
  NOR2_X1 U777 ( .A1(n725), .A2(n724), .ZN(G63) );
  XOR2_X1 U778 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n727) );
  NAND2_X1 U779 ( .A1(G224), .A2(G953), .ZN(n726) );
  XNOR2_X1 U780 ( .A(n727), .B(n726), .ZN(n728) );
  NAND2_X1 U781 ( .A1(G898), .A2(n728), .ZN(n729) );
  XOR2_X1 U782 ( .A(KEYINPUT126), .B(n729), .Z(n732) );
  NOR2_X1 U783 ( .A1(G953), .A2(n730), .ZN(n731) );
  NOR2_X1 U784 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U785 ( .A(n733), .B(KEYINPUT127), .ZN(n738) );
  XNOR2_X1 U786 ( .A(n734), .B(G110), .ZN(n735) );
  NOR2_X1 U787 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U788 ( .A(n738), .B(n737), .ZN(G69) );
  XNOR2_X1 U789 ( .A(n740), .B(n739), .ZN(n744) );
  XNOR2_X1 U790 ( .A(n741), .B(n744), .ZN(n743) );
  NAND2_X1 U791 ( .A1(n743), .A2(n742), .ZN(n748) );
  XNOR2_X1 U792 ( .A(n744), .B(G227), .ZN(n745) );
  NAND2_X1 U793 ( .A1(n745), .A2(G900), .ZN(n746) );
  NAND2_X1 U794 ( .A1(n746), .A2(G953), .ZN(n747) );
  NAND2_X1 U795 ( .A1(n748), .A2(n747), .ZN(G72) );
  XOR2_X1 U796 ( .A(n749), .B(G137), .Z(G39) );
  XOR2_X1 U797 ( .A(n750), .B(G122), .Z(G24) );
  XNOR2_X1 U798 ( .A(G119), .B(n751), .ZN(G21) );
endmodule

