//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 1 0 0 0 1 0 1 0 1 1 1 1 0 0 0 1 0 1 1 0 1 1 1 1 0 1 0 1 0 0 1 1 1 0 0 0 1 1 0 1 0 0 0 0 1 0 1 0 1 0 0 1 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n694, new_n695, new_n696, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n771, new_n772, new_n773, new_n774, new_n776, new_n777, new_n778,
    new_n779, new_n781, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n880, new_n881, new_n882, new_n883,
    new_n885, new_n886, new_n887, new_n889, new_n890, new_n891, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n941, new_n942, new_n943, new_n945,
    new_n946, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n958, new_n959, new_n960, new_n962, new_n963,
    new_n964, new_n965, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n993, new_n994;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G169gat), .B(G197gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(KEYINPUT89), .B(KEYINPUT11), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  XOR2_X1   g005(.A(new_n206), .B(KEYINPUT12), .Z(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(G15gat), .B(G22gat), .ZN(new_n209));
  OR2_X1    g008(.A1(new_n209), .A2(G1gat), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT93), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT16), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n209), .B1(new_n212), .B2(G1gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n210), .A2(new_n211), .A3(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(G8gat), .ZN(new_n215));
  INV_X1    g014(.A(G8gat), .ZN(new_n216));
  NAND4_X1  g015(.A1(new_n210), .A2(new_n213), .A3(new_n211), .A4(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT14), .ZN(new_n219));
  NOR3_X1   g018(.A1(new_n219), .A2(G29gat), .A3(G36gat), .ZN(new_n220));
  INV_X1    g019(.A(G29gat), .ZN(new_n221));
  INV_X1    g020(.A(G36gat), .ZN(new_n222));
  AOI21_X1  g021(.A(KEYINPUT14), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  OAI21_X1  g022(.A(KEYINPUT90), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n221), .A2(new_n222), .A3(KEYINPUT14), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n219), .B1(G29gat), .B2(G36gat), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT90), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  AND2_X1   g027(.A1(KEYINPUT91), .A2(G36gat), .ZN(new_n229));
  NOR2_X1   g028(.A1(KEYINPUT91), .A2(G36gat), .ZN(new_n230));
  OAI21_X1  g029(.A(G29gat), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n224), .A2(new_n228), .A3(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT15), .ZN(new_n233));
  INV_X1    g032(.A(G43gat), .ZN(new_n234));
  INV_X1    g033(.A(G50gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(G43gat), .A2(G50gat), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n233), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n232), .A2(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n236), .A2(new_n233), .A3(new_n237), .ZN(new_n240));
  AND2_X1   g039(.A1(new_n231), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n226), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n238), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n239), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n218), .A2(new_n245), .ZN(new_n246));
  AOI22_X1  g045(.A1(new_n232), .A2(new_n238), .B1(new_n243), .B2(new_n241), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n247), .A2(new_n215), .A3(new_n217), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(G229gat), .A2(G233gat), .ZN(new_n250));
  XOR2_X1   g049(.A(new_n250), .B(KEYINPUT13), .Z(new_n251));
  NAND2_X1  g050(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT17), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT92), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n253), .B1(new_n247), .B2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(new_n238), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n227), .B1(new_n225), .B2(new_n226), .ZN(new_n257));
  INV_X1    g056(.A(new_n230), .ZN(new_n258));
  NAND2_X1  g057(.A1(KEYINPUT91), .A2(G36gat), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n221), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n257), .A2(new_n260), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n256), .B1(new_n261), .B2(new_n228), .ZN(new_n262));
  AND2_X1   g061(.A1(new_n241), .A2(new_n243), .ZN(new_n263));
  OAI211_X1 g062(.A(KEYINPUT92), .B(KEYINPUT17), .C1(new_n262), .C2(new_n263), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n218), .B1(new_n255), .B2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(new_n250), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n247), .B1(new_n215), .B2(new_n217), .ZN(new_n267));
  NOR3_X1   g066(.A1(new_n265), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n252), .B1(new_n268), .B2(KEYINPUT18), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT18), .ZN(new_n270));
  NOR4_X1   g069(.A1(new_n265), .A2(new_n270), .A3(new_n266), .A4(new_n267), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n208), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n255), .A2(new_n264), .ZN(new_n273));
  INV_X1    g072(.A(new_n218), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n275), .A2(new_n250), .A3(new_n246), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(new_n270), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n268), .A2(KEYINPUT18), .ZN(new_n278));
  NAND4_X1  g077(.A1(new_n277), .A2(new_n278), .A3(new_n252), .A4(new_n207), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n272), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT72), .ZN(new_n282));
  INV_X1    g081(.A(G169gat), .ZN(new_n283));
  INV_X1    g082(.A(G176gat), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT26), .ZN(new_n286));
  NOR2_X1   g085(.A1(G169gat), .A2(G176gat), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n285), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n288), .B1(new_n286), .B2(new_n287), .ZN(new_n289));
  NAND2_X1  g088(.A1(G183gat), .A2(G190gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  XNOR2_X1  g091(.A(KEYINPUT27), .B(G183gat), .ZN(new_n293));
  INV_X1    g092(.A(G190gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT28), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n295), .B(new_n296), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n292), .A2(KEYINPUT66), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n299));
  MUX2_X1   g098(.A(G183gat), .B(new_n299), .S(G190gat), .Z(new_n300));
  INV_X1    g099(.A(KEYINPUT24), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n290), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n285), .B1(KEYINPUT23), .B2(new_n287), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n283), .A2(new_n284), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT23), .ZN(new_n306));
  AOI21_X1  g105(.A(KEYINPUT64), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT64), .ZN(new_n308));
  NOR3_X1   g107(.A1(new_n287), .A2(new_n308), .A3(KEYINPUT23), .ZN(new_n309));
  OAI211_X1 g108(.A(new_n303), .B(new_n304), .C1(new_n307), .C2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT25), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  AND2_X1   g111(.A1(new_n302), .A2(KEYINPUT65), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n302), .A2(KEYINPUT65), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n300), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  OR2_X1    g114(.A1(new_n307), .A2(new_n309), .ZN(new_n316));
  NAND4_X1  g115(.A1(new_n315), .A2(new_n316), .A3(KEYINPUT25), .A4(new_n304), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n312), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT66), .ZN(new_n319));
  XNOR2_X1  g118(.A(new_n295), .B(KEYINPUT28), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n319), .B1(new_n320), .B2(new_n291), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n298), .A2(new_n318), .A3(new_n321), .ZN(new_n322));
  XNOR2_X1  g121(.A(KEYINPUT67), .B(G127gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(G134gat), .ZN(new_n324));
  OR2_X1    g123(.A1(G127gat), .A2(G134gat), .ZN(new_n325));
  AOI21_X1  g124(.A(KEYINPUT68), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(G113gat), .B(G120gat), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n327), .A2(KEYINPUT1), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n324), .A2(KEYINPUT68), .A3(new_n325), .ZN(new_n330));
  XOR2_X1   g129(.A(new_n327), .B(KEYINPUT69), .Z(new_n331));
  NAND2_X1  g130(.A1(G127gat), .A2(G134gat), .ZN(new_n332));
  AOI21_X1  g131(.A(KEYINPUT1), .B1(new_n325), .B2(new_n332), .ZN(new_n333));
  AOI22_X1  g132(.A1(new_n329), .A2(new_n330), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n322), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n329), .A2(new_n330), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n331), .A2(new_n333), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND4_X1  g137(.A1(new_n338), .A2(new_n298), .A3(new_n318), .A4(new_n321), .ZN(new_n339));
  NAND4_X1  g138(.A1(new_n335), .A2(G227gat), .A3(G233gat), .A4(new_n339), .ZN(new_n340));
  XNOR2_X1  g139(.A(G15gat), .B(G43gat), .ZN(new_n341));
  XNOR2_X1  g140(.A(G71gat), .B(G99gat), .ZN(new_n342));
  XNOR2_X1  g141(.A(new_n341), .B(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT33), .ZN(new_n344));
  OR2_X1    g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n340), .A2(KEYINPUT32), .A3(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT70), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND4_X1  g147(.A1(new_n340), .A2(KEYINPUT70), .A3(KEYINPUT32), .A4(new_n345), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n343), .B1(new_n340), .B2(KEYINPUT32), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n340), .A2(new_n344), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n350), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n335), .A2(new_n339), .ZN(new_n355));
  NAND2_X1  g154(.A1(G227gat), .A2(G233gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  OAI21_X1  g156(.A(KEYINPUT71), .B1(new_n357), .B2(KEYINPUT34), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT71), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT34), .ZN(new_n360));
  NAND4_X1  g159(.A1(new_n355), .A2(new_n359), .A3(new_n360), .A4(new_n356), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n357), .A2(KEYINPUT34), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n358), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n282), .B1(new_n354), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n354), .A2(new_n363), .ZN(new_n365));
  AOI22_X1  g164(.A1(new_n348), .A2(new_n349), .B1(new_n352), .B2(new_n351), .ZN(new_n366));
  AND2_X1   g165(.A1(new_n358), .A2(new_n362), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n366), .A2(new_n361), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n365), .A2(new_n368), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n364), .B1(new_n369), .B2(new_n282), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT36), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n369), .A2(KEYINPUT36), .ZN(new_n373));
  AND2_X1   g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  XNOR2_X1  g173(.A(KEYINPUT81), .B(KEYINPUT6), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT2), .ZN(new_n377));
  INV_X1    g176(.A(G148gat), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n378), .A2(G141gat), .ZN(new_n379));
  INV_X1    g178(.A(G141gat), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n380), .A2(G148gat), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n377), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(G155gat), .A2(G162gat), .ZN(new_n383));
  INV_X1    g182(.A(G155gat), .ZN(new_n384));
  INV_X1    g183(.A(G162gat), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n384), .A2(new_n385), .A3(KEYINPUT77), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n384), .A2(new_n385), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT77), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND4_X1  g188(.A1(new_n382), .A2(new_n383), .A3(new_n386), .A4(new_n389), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n383), .B1(new_n387), .B2(KEYINPUT2), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n380), .A2(KEYINPUT78), .A3(G148gat), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n392), .B1(new_n380), .B2(G148gat), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n379), .A2(KEYINPUT78), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n391), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  AND2_X1   g194(.A1(new_n395), .A2(KEYINPUT79), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n395), .A2(KEYINPUT79), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n390), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT4), .ZN(new_n399));
  NOR3_X1   g198(.A1(new_n338), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n390), .ZN(new_n401));
  INV_X1    g200(.A(new_n397), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n395), .A2(KEYINPUT79), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n401), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  AOI21_X1  g203(.A(KEYINPUT4), .B1(new_n404), .B2(new_n334), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n400), .A2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT80), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n398), .A2(new_n407), .ZN(new_n408));
  OAI211_X1 g207(.A(KEYINPUT80), .B(new_n390), .C1(new_n396), .C2(new_n397), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n408), .A2(KEYINPUT3), .A3(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT3), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n334), .B1(new_n404), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(G225gat), .A2(G233gat), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n406), .A2(new_n413), .A3(KEYINPUT5), .A4(new_n414), .ZN(new_n415));
  AND3_X1   g214(.A1(new_n406), .A2(new_n413), .A3(new_n414), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT5), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n408), .A2(new_n409), .A3(new_n338), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n404), .A2(new_n334), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(new_n414), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n417), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n415), .B1(new_n416), .B2(new_n422), .ZN(new_n423));
  XNOR2_X1  g222(.A(G1gat), .B(G29gat), .ZN(new_n424));
  XNOR2_X1  g223(.A(new_n424), .B(KEYINPUT0), .ZN(new_n425));
  XNOR2_X1  g224(.A(G57gat), .B(G85gat), .ZN(new_n426));
  XOR2_X1   g225(.A(new_n425), .B(new_n426), .Z(new_n427));
  AOI21_X1  g226(.A(new_n376), .B1(new_n423), .B2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n427), .ZN(new_n429));
  OAI211_X1 g228(.A(new_n429), .B(new_n415), .C1(new_n416), .C2(new_n422), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n430), .A2(new_n375), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(G226gat), .A2(G233gat), .ZN(new_n435));
  XOR2_X1   g234(.A(new_n435), .B(KEYINPUT75), .Z(new_n436));
  INV_X1    g235(.A(KEYINPUT29), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n436), .B1(new_n322), .B2(new_n437), .ZN(new_n438));
  AOI22_X1  g237(.A1(new_n312), .A2(new_n317), .B1(new_n292), .B2(new_n297), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n439), .A2(new_n435), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  XNOR2_X1  g241(.A(G197gat), .B(G204gat), .ZN(new_n443));
  INV_X1    g242(.A(G211gat), .ZN(new_n444));
  INV_X1    g243(.A(G218gat), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n443), .B1(KEYINPUT22), .B2(new_n446), .ZN(new_n447));
  XNOR2_X1  g246(.A(G211gat), .B(G218gat), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  OR2_X1    g249(.A1(new_n450), .A2(KEYINPUT73), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT74), .ZN(new_n452));
  OAI211_X1 g251(.A(new_n448), .B(new_n443), .C1(KEYINPUT22), .C2(new_n446), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n450), .A2(KEYINPUT73), .A3(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n451), .A2(new_n452), .A3(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n452), .B1(new_n451), .B2(new_n454), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n458), .ZN(new_n459));
  XNOR2_X1  g258(.A(G8gat), .B(G36gat), .ZN(new_n460));
  XNOR2_X1  g259(.A(new_n460), .B(KEYINPUT76), .ZN(new_n461));
  XNOR2_X1  g260(.A(G64gat), .B(G92gat), .ZN(new_n462));
  XOR2_X1   g261(.A(new_n461), .B(new_n462), .Z(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(new_n458), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n322), .A2(new_n436), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n435), .B1(new_n439), .B2(KEYINPUT29), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n459), .A2(KEYINPUT30), .A3(new_n464), .A4(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT30), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n468), .B1(new_n441), .B2(new_n465), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n470), .B1(new_n471), .B2(new_n463), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n463), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n469), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n434), .A2(new_n475), .ZN(new_n476));
  XNOR2_X1  g275(.A(G78gat), .B(G106gat), .ZN(new_n477));
  XNOR2_X1  g276(.A(KEYINPUT31), .B(G50gat), .ZN(new_n478));
  XOR2_X1   g277(.A(new_n477), .B(new_n478), .Z(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n437), .B1(new_n398), .B2(KEYINPUT3), .ZN(new_n481));
  INV_X1    g280(.A(new_n457), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n481), .A2(new_n482), .A3(new_n455), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n451), .A2(new_n437), .A3(new_n454), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(new_n411), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n485), .A2(new_n408), .A3(new_n409), .ZN(new_n486));
  NAND2_X1  g285(.A1(G228gat), .A2(G233gat), .ZN(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n483), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(G22gat), .ZN(new_n490));
  AOI21_X1  g289(.A(KEYINPUT29), .B1(new_n450), .B2(new_n453), .ZN(new_n491));
  OR2_X1    g290(.A1(new_n491), .A2(KEYINPUT3), .ZN(new_n492));
  AOI22_X1  g291(.A1(new_n458), .A2(new_n481), .B1(new_n398), .B2(new_n492), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n489), .B(new_n490), .C1(new_n493), .C2(new_n488), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT82), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AND3_X1   g295(.A1(new_n483), .A2(new_n486), .A3(new_n488), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n492), .A2(new_n398), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n488), .B1(new_n483), .B2(new_n498), .ZN(new_n499));
  OAI21_X1  g298(.A(G22gat), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n496), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n483), .A2(new_n498), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(new_n487), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n490), .B1(new_n503), .B2(new_n489), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n504), .A2(new_n495), .A3(new_n494), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n480), .B1(new_n501), .B2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT83), .ZN(new_n507));
  OAI211_X1 g306(.A(new_n507), .B(G22gat), .C1(new_n497), .C2(new_n499), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n508), .A2(new_n480), .A3(new_n494), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n504), .A2(new_n507), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n506), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n476), .A2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT85), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n423), .A2(new_n514), .ZN(new_n515));
  OAI211_X1 g314(.A(KEYINPUT85), .B(new_n415), .C1(new_n416), .C2(new_n422), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n515), .A2(new_n429), .A3(new_n516), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n432), .B1(new_n517), .B2(new_n428), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n471), .A2(new_n463), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n471), .A2(KEYINPUT37), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n520), .A2(new_n464), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT37), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n522), .B1(new_n442), .B2(new_n465), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n467), .A2(new_n466), .A3(new_n458), .ZN(new_n524));
  AOI21_X1  g323(.A(KEYINPUT38), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n519), .B1(new_n521), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n518), .A2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT86), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n518), .A2(KEYINPUT86), .A3(new_n526), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n471), .A2(KEYINPUT37), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n521), .A2(new_n531), .ZN(new_n532));
  AOI22_X1  g331(.A1(new_n529), .A2(new_n530), .B1(KEYINPUT38), .B2(new_n532), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n504), .B1(new_n495), .B2(new_n494), .ZN(new_n534));
  AOI211_X1 g333(.A(KEYINPUT82), .B(new_n490), .C1(new_n503), .C2(new_n489), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n479), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  OR2_X1    g335(.A1(new_n509), .A2(new_n510), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n406), .A2(new_n413), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(new_n421), .ZN(new_n540));
  OAI211_X1 g339(.A(new_n540), .B(KEYINPUT39), .C1(new_n421), .C2(new_n420), .ZN(new_n541));
  OR2_X1    g340(.A1(new_n540), .A2(KEYINPUT39), .ZN(new_n542));
  AND3_X1   g341(.A1(new_n542), .A2(KEYINPUT84), .A3(new_n427), .ZN(new_n543));
  AOI21_X1  g342(.A(KEYINPUT84), .B1(new_n542), .B2(new_n427), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n541), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT40), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  OAI211_X1 g347(.A(KEYINPUT40), .B(new_n541), .C1(new_n543), .C2(new_n544), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n549), .A2(new_n517), .A3(new_n474), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n538), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  OAI211_X1 g350(.A(new_n374), .B(new_n513), .C1(new_n533), .C2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT87), .ZN(new_n553));
  AND2_X1   g352(.A1(new_n517), .A2(new_n428), .ZN(new_n554));
  OAI211_X1 g353(.A(new_n553), .B(new_n475), .C1(new_n554), .C2(new_n432), .ZN(new_n555));
  OAI21_X1  g354(.A(KEYINPUT87), .B1(new_n518), .B2(new_n474), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n512), .A2(KEYINPUT35), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n555), .A2(new_n556), .A3(new_n370), .A4(new_n557), .ZN(new_n558));
  OAI211_X1 g357(.A(new_n365), .B(new_n368), .C1(new_n506), .C2(new_n511), .ZN(new_n559));
  OAI211_X1 g358(.A(KEYINPUT88), .B(KEYINPUT35), .C1(new_n476), .C2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n474), .B1(new_n431), .B2(new_n433), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n366), .B(new_n363), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n562), .A2(new_n538), .A3(new_n563), .ZN(new_n564));
  AOI21_X1  g363(.A(KEYINPUT88), .B1(new_n564), .B2(KEYINPUT35), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n558), .B1(new_n561), .B2(new_n565), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n281), .B1(new_n552), .B2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT97), .ZN(new_n568));
  XNOR2_X1  g367(.A(G57gat), .B(G64gat), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  OR2_X1    g369(.A1(G71gat), .A2(G78gat), .ZN(new_n571));
  NAND2_X1  g370(.A1(G71gat), .A2(G78gat), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT9), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n570), .A2(new_n573), .A3(new_n575), .ZN(new_n576));
  OAI211_X1 g375(.A(new_n572), .B(new_n571), .C1(new_n569), .C2(new_n574), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(G99gat), .B(G106gat), .ZN(new_n579));
  NAND2_X1  g378(.A1(G85gat), .A2(G92gat), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT95), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT7), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(G99gat), .A2(G106gat), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n584), .A2(KEYINPUT8), .ZN(new_n585));
  INV_X1    g384(.A(G85gat), .ZN(new_n586));
  INV_X1    g385(.A(G92gat), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AND3_X1   g387(.A1(new_n583), .A2(new_n585), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n580), .A2(new_n581), .ZN(new_n590));
  NAND3_X1  g389(.A1(KEYINPUT95), .A2(G85gat), .A3(G92gat), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n590), .A2(KEYINPUT7), .A3(new_n591), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n579), .B1(new_n589), .B2(new_n592), .ZN(new_n593));
  AOI22_X1  g392(.A1(KEYINPUT8), .A2(new_n584), .B1(new_n586), .B2(new_n587), .ZN(new_n594));
  AND4_X1   g393(.A1(new_n579), .A2(new_n592), .A3(new_n583), .A4(new_n594), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n578), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n592), .A2(new_n583), .A3(new_n594), .ZN(new_n597));
  INV_X1    g396(.A(new_n579), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND4_X1  g398(.A1(new_n592), .A2(new_n579), .A3(new_n583), .A4(new_n594), .ZN(new_n600));
  NAND4_X1  g399(.A1(new_n599), .A2(new_n577), .A3(new_n576), .A4(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT10), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n596), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n578), .ZN(new_n604));
  NAND4_X1  g403(.A1(new_n604), .A2(KEYINPUT10), .A3(new_n600), .A4(new_n599), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(G230gat), .A2(G233gat), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n568), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n607), .ZN(new_n609));
  AOI211_X1 g408(.A(KEYINPUT97), .B(new_n609), .C1(new_n603), .C2(new_n605), .ZN(new_n610));
  XNOR2_X1  g409(.A(G120gat), .B(G148gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(G176gat), .B(G204gat), .ZN(new_n612));
  XOR2_X1   g411(.A(new_n611), .B(new_n612), .Z(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n607), .B1(new_n596), .B2(new_n601), .ZN(new_n615));
  NOR4_X1   g414(.A1(new_n608), .A2(new_n610), .A3(new_n614), .A4(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n615), .ZN(new_n618));
  AOI21_X1  g417(.A(KEYINPUT98), .B1(new_n606), .B2(new_n607), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT98), .ZN(new_n620));
  AOI211_X1 g419(.A(new_n620), .B(new_n609), .C1(new_n603), .C2(new_n605), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n618), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT99), .ZN(new_n623));
  AND3_X1   g422(.A1(new_n622), .A2(new_n623), .A3(new_n614), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n623), .B1(new_n622), .B2(new_n614), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n617), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT100), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT21), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n578), .A2(new_n629), .ZN(new_n630));
  AND2_X1   g429(.A1(G231gat), .A2(G233gat), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n630), .A2(new_n631), .ZN(new_n634));
  OAI21_X1  g433(.A(G127gat), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n634), .ZN(new_n636));
  INV_X1    g435(.A(G127gat), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n636), .A2(new_n637), .A3(new_n632), .ZN(new_n638));
  XOR2_X1   g437(.A(G183gat), .B(G211gat), .Z(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n635), .A2(new_n638), .A3(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n640), .B1(new_n635), .B2(new_n638), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n578), .A2(new_n629), .ZN(new_n644));
  OR3_X1    g443(.A1(new_n218), .A2(KEYINPUT94), .A3(new_n644), .ZN(new_n645));
  OAI21_X1  g444(.A(KEYINPUT94), .B1(new_n218), .B2(new_n644), .ZN(new_n646));
  XNOR2_X1  g445(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(new_n384), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  AND3_X1   g448(.A1(new_n645), .A2(new_n646), .A3(new_n649), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n649), .B1(new_n645), .B2(new_n646), .ZN(new_n651));
  OAI22_X1  g450(.A1(new_n642), .A2(new_n643), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n635), .A2(new_n638), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n653), .A2(new_n639), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n645), .A2(new_n646), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n655), .A2(new_n648), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n645), .A2(new_n646), .A3(new_n649), .ZN(new_n657));
  NAND4_X1  g456(.A1(new_n654), .A2(new_n656), .A3(new_n641), .A4(new_n657), .ZN(new_n658));
  AND2_X1   g457(.A1(new_n652), .A2(new_n658), .ZN(new_n659));
  AOI21_X1  g458(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  NAND3_X1  g460(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n599), .A2(new_n600), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n662), .B1(new_n247), .B2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT96), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n273), .A2(new_n663), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n661), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n666), .A2(new_n667), .A3(new_n661), .ZN(new_n670));
  XNOR2_X1  g469(.A(G190gat), .B(G218gat), .ZN(new_n671));
  XNOR2_X1  g470(.A(G134gat), .B(G162gat), .ZN(new_n672));
  XOR2_X1   g471(.A(new_n671), .B(new_n672), .Z(new_n673));
  NAND3_X1  g472(.A1(new_n669), .A2(new_n670), .A3(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n673), .ZN(new_n675));
  INV_X1    g474(.A(new_n670), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n675), .B1(new_n676), .B2(new_n668), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n659), .B1(new_n674), .B2(new_n677), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n627), .A2(new_n628), .A3(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n677), .A2(new_n674), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n652), .A2(new_n658), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  OAI21_X1  g481(.A(KEYINPUT100), .B1(new_n682), .B2(new_n626), .ZN(new_n683));
  AND2_X1   g482(.A1(new_n679), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n567), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n685), .A2(new_n434), .ZN(new_n686));
  XOR2_X1   g485(.A(new_n686), .B(G1gat), .Z(G1324gat));
  NOR2_X1   g486(.A1(new_n685), .A2(new_n475), .ZN(new_n688));
  XOR2_X1   g487(.A(KEYINPUT16), .B(G8gat), .Z(new_n689));
  AND2_X1   g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  OR2_X1    g489(.A1(new_n690), .A2(KEYINPUT42), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(KEYINPUT42), .ZN(new_n692));
  OAI211_X1 g491(.A(new_n691), .B(new_n692), .C1(new_n216), .C2(new_n688), .ZN(G1325gat));
  OAI21_X1  g492(.A(G15gat), .B1(new_n685), .B2(new_n374), .ZN(new_n694));
  INV_X1    g493(.A(new_n370), .ZN(new_n695));
  OR2_X1    g494(.A1(new_n695), .A2(G15gat), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n694), .B1(new_n685), .B2(new_n696), .ZN(G1326gat));
  NAND3_X1  g496(.A1(new_n567), .A2(new_n512), .A3(new_n684), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(KEYINPUT101), .ZN(new_n699));
  XNOR2_X1  g498(.A(KEYINPUT43), .B(G22gat), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n699), .B(new_n700), .ZN(G1327gat));
  AND2_X1   g500(.A1(new_n677), .A2(new_n674), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT44), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT104), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n566), .A2(new_n705), .ZN(new_n706));
  OAI211_X1 g505(.A(new_n558), .B(KEYINPUT104), .C1(new_n561), .C2(new_n565), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n704), .B1(new_n708), .B2(new_n552), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n552), .A2(new_n566), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n703), .B1(new_n710), .B2(new_n702), .ZN(new_n711));
  OR2_X1    g510(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n626), .B(KEYINPUT103), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n681), .B(KEYINPUT102), .ZN(new_n714));
  AND3_X1   g513(.A1(new_n713), .A2(new_n280), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n712), .A2(new_n715), .ZN(new_n716));
  OAI21_X1  g515(.A(G29gat), .B1(new_n716), .B2(new_n434), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n680), .A2(new_n681), .ZN(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n719), .A2(new_n626), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  AOI211_X1 g520(.A(new_n281), .B(new_n721), .C1(new_n552), .C2(new_n566), .ZN(new_n722));
  INV_X1    g521(.A(new_n434), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n722), .A2(new_n221), .A3(new_n723), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n724), .B(KEYINPUT45), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n717), .A2(new_n725), .ZN(G1328gat));
  NAND2_X1  g525(.A1(new_n258), .A2(new_n259), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n727), .B1(new_n716), .B2(new_n475), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n567), .A2(new_n720), .ZN(new_n729));
  NOR3_X1   g528(.A1(new_n729), .A2(new_n475), .A3(new_n727), .ZN(new_n730));
  XNOR2_X1  g529(.A(KEYINPUT105), .B(KEYINPUT46), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n730), .B(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n728), .A2(new_n732), .ZN(G1329gat));
  NAND2_X1  g532(.A1(new_n372), .A2(new_n373), .ZN(new_n734));
  OAI211_X1 g533(.A(new_n734), .B(new_n715), .C1(new_n709), .C2(new_n711), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(G43gat), .ZN(new_n736));
  NOR3_X1   g535(.A1(new_n729), .A2(G43gat), .A3(new_n695), .ZN(new_n737));
  INV_X1    g536(.A(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  AOI21_X1  g538(.A(KEYINPUT47), .B1(new_n739), .B2(KEYINPUT106), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n737), .B1(new_n735), .B2(G43gat), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT106), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT47), .ZN(new_n743));
  NOR3_X1   g542(.A1(new_n741), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n740), .A2(new_n744), .ZN(G1330gat));
  INV_X1    g544(.A(KEYINPUT107), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n538), .A2(G50gat), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n746), .B1(new_n722), .B2(new_n747), .ZN(new_n748));
  OAI21_X1  g547(.A(KEYINPUT108), .B1(new_n748), .B2(KEYINPUT48), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n567), .A2(new_n720), .A3(new_n747), .ZN(new_n750));
  AOI21_X1  g549(.A(KEYINPUT48), .B1(new_n750), .B2(KEYINPUT107), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT108), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n749), .A2(new_n753), .ZN(new_n754));
  OAI211_X1 g553(.A(new_n512), .B(new_n715), .C1(new_n709), .C2(new_n711), .ZN(new_n755));
  AOI22_X1  g554(.A1(new_n755), .A2(G50gat), .B1(new_n722), .B2(new_n747), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n754), .B(new_n756), .ZN(G1331gat));
  NAND3_X1  g556(.A1(new_n372), .A2(new_n513), .A3(new_n373), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n529), .A2(new_n530), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n532), .A2(KEYINPUT38), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(new_n550), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n512), .B1(new_n762), .B2(new_n547), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n758), .B1(new_n761), .B2(new_n763), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n764), .B1(new_n706), .B2(new_n707), .ZN(new_n765));
  NOR3_X1   g564(.A1(new_n713), .A2(new_n280), .A3(new_n682), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(KEYINPUT109), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(new_n723), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n769), .B(G57gat), .ZN(G1332gat));
  INV_X1    g569(.A(KEYINPUT49), .ZN(new_n771));
  INV_X1    g570(.A(G64gat), .ZN(new_n772));
  OAI211_X1 g571(.A(new_n768), .B(new_n474), .C1(new_n771), .C2(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n771), .A2(new_n772), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n773), .B(new_n774), .ZN(G1333gat));
  INV_X1    g574(.A(G71gat), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n768), .A2(new_n776), .A3(new_n370), .ZN(new_n777));
  NOR3_X1   g576(.A1(new_n765), .A2(new_n374), .A3(new_n767), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n777), .B1(new_n778), .B2(new_n776), .ZN(new_n779));
  XOR2_X1   g578(.A(new_n779), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g579(.A1(new_n768), .A2(new_n512), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n781), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g581(.A1(new_n627), .A2(new_n280), .A3(new_n681), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n712), .A2(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(G85gat), .B1(new_n784), .B2(new_n434), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT51), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n719), .A2(new_n280), .ZN(new_n787));
  INV_X1    g586(.A(new_n787), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n786), .B1(new_n765), .B2(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(new_n707), .ZN(new_n790));
  OAI21_X1  g589(.A(KEYINPUT35), .B1(new_n476), .B2(new_n559), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT88), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(new_n560), .ZN(new_n794));
  AOI21_X1  g593(.A(KEYINPUT104), .B1(new_n794), .B2(new_n558), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n552), .B1(new_n790), .B2(new_n795), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n796), .A2(KEYINPUT51), .A3(new_n787), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n789), .A2(new_n797), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n798), .A2(new_n586), .A3(new_n723), .A4(new_n626), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n785), .A2(new_n799), .ZN(G1336gat));
  XNOR2_X1  g599(.A(KEYINPUT110), .B(KEYINPUT52), .ZN(new_n801));
  INV_X1    g600(.A(new_n801), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n709), .A2(new_n711), .ZN(new_n803));
  INV_X1    g602(.A(new_n783), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n587), .B1(new_n805), .B2(new_n474), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n713), .B1(new_n789), .B2(new_n797), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n475), .A2(G92gat), .ZN(new_n808));
  AND2_X1   g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n802), .B1(new_n806), .B2(new_n809), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n712), .A2(new_n474), .A3(new_n783), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(G92gat), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n807), .A2(new_n808), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n812), .A2(new_n813), .A3(new_n801), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n810), .A2(new_n814), .ZN(G1337gat));
  OAI21_X1  g614(.A(KEYINPUT111), .B1(new_n784), .B2(new_n374), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT111), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n805), .A2(new_n817), .A3(new_n734), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n816), .A2(G99gat), .A3(new_n818), .ZN(new_n819));
  NOR3_X1   g618(.A1(new_n695), .A2(G99gat), .A3(new_n627), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n798), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n819), .A2(new_n821), .ZN(G1338gat));
  OR2_X1    g621(.A1(KEYINPUT112), .A2(KEYINPUT53), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n538), .A2(G106gat), .ZN(new_n824));
  AOI22_X1  g623(.A1(new_n807), .A2(new_n824), .B1(KEYINPUT112), .B2(KEYINPUT53), .ZN(new_n825));
  OAI211_X1 g624(.A(new_n512), .B(new_n783), .C1(new_n709), .C2(new_n711), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(G106gat), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n823), .B1(new_n825), .B2(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(new_n713), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n798), .A2(new_n829), .A3(new_n824), .ZN(new_n830));
  NAND2_X1  g629(.A1(KEYINPUT112), .A2(KEYINPUT53), .ZN(new_n831));
  AND4_X1   g630(.A1(new_n827), .A2(new_n830), .A3(new_n831), .A4(new_n823), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n828), .A2(new_n832), .ZN(G1339gat));
  INV_X1    g632(.A(new_n251), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n246), .A2(new_n248), .A3(new_n834), .ZN(new_n835));
  XNOR2_X1  g634(.A(new_n835), .B(KEYINPUT113), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n266), .B1(new_n265), .B2(new_n267), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n206), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n269), .A2(new_n271), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n838), .B1(new_n839), .B2(new_n207), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n626), .A2(new_n840), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n619), .A2(new_n621), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT54), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n613), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT55), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n608), .A2(new_n610), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n603), .A2(new_n609), .A3(new_n605), .ZN(new_n847));
  AND2_X1   g646(.A1(new_n847), .A2(KEYINPUT54), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n845), .B1(new_n846), .B2(new_n848), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n616), .B1(new_n844), .B2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(new_n619), .ZN(new_n851));
  INV_X1    g650(.A(new_n621), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n851), .A2(new_n852), .A3(new_n843), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n606), .A2(new_n607), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(KEYINPUT97), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n606), .A2(new_n568), .A3(new_n607), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n855), .A2(new_n848), .A3(new_n856), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n853), .A2(new_n857), .A3(new_n614), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(new_n845), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n280), .A2(new_n850), .A3(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n702), .B1(new_n841), .B2(new_n860), .ZN(new_n861));
  AND4_X1   g660(.A1(new_n702), .A2(new_n840), .A3(new_n859), .A4(new_n850), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n714), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n678), .A2(new_n281), .A3(new_n627), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n512), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  XNOR2_X1  g664(.A(new_n865), .B(KEYINPUT114), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n866), .A2(new_n695), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n723), .A2(new_n475), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  OR2_X1    g669(.A1(new_n870), .A2(KEYINPUT115), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(KEYINPUT115), .ZN(new_n872));
  NAND4_X1  g671(.A1(new_n871), .A2(G113gat), .A3(new_n280), .A4(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(G113gat), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n434), .B1(new_n863), .B2(new_n864), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n559), .A2(new_n474), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n874), .B1(new_n877), .B2(new_n281), .ZN(new_n878));
  AND2_X1   g677(.A1(new_n873), .A2(new_n878), .ZN(G1340gat));
  OR3_X1    g678(.A1(new_n877), .A2(G120gat), .A3(new_n627), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n871), .A2(new_n829), .A3(new_n872), .ZN(new_n881));
  AND3_X1   g680(.A1(new_n881), .A2(KEYINPUT116), .A3(G120gat), .ZN(new_n882));
  AOI21_X1  g681(.A(KEYINPUT116), .B1(new_n881), .B2(G120gat), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n880), .B1(new_n882), .B2(new_n883), .ZN(G1341gat));
  NAND2_X1  g683(.A1(new_n871), .A2(new_n872), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n323), .B1(new_n885), .B2(new_n714), .ZN(new_n886));
  OR2_X1    g685(.A1(new_n659), .A2(new_n323), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n886), .B1(new_n877), .B2(new_n887), .ZN(G1342gat));
  OAI21_X1  g687(.A(G134gat), .B1(new_n885), .B2(new_n680), .ZN(new_n889));
  NOR3_X1   g688(.A1(new_n877), .A2(G134gat), .A3(new_n680), .ZN(new_n890));
  XNOR2_X1  g689(.A(new_n890), .B(KEYINPUT56), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n889), .A2(new_n891), .ZN(G1343gat));
  NOR3_X1   g691(.A1(new_n734), .A2(new_n538), .A3(new_n474), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(new_n875), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n380), .B1(new_n894), .B2(new_n281), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n734), .A2(new_n868), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n512), .A2(KEYINPUT57), .ZN(new_n897));
  INV_X1    g696(.A(new_n862), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n898), .B1(new_n861), .B2(KEYINPUT117), .ZN(new_n899));
  AND2_X1   g698(.A1(new_n861), .A2(KEYINPUT117), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n659), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n897), .B1(new_n901), .B2(new_n864), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT118), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n538), .B1(new_n863), .B2(new_n864), .ZN(new_n904));
  OAI22_X1  g703(.A1(new_n902), .A2(new_n903), .B1(KEYINPUT57), .B2(new_n904), .ZN(new_n905));
  AND2_X1   g704(.A1(new_n902), .A2(new_n903), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n896), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n280), .A2(G141gat), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n895), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  XOR2_X1   g708(.A(new_n909), .B(KEYINPUT58), .Z(G1344gat));
  OAI211_X1 g709(.A(new_n626), .B(new_n896), .C1(new_n905), .C2(new_n906), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n378), .A2(KEYINPUT59), .ZN(new_n912));
  AND2_X1   g711(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NOR3_X1   g712(.A1(new_n734), .A2(new_n627), .A3(new_n868), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT119), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n897), .B1(new_n863), .B2(new_n864), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n659), .B1(new_n861), .B2(new_n862), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n679), .A2(new_n683), .A3(new_n281), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n538), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  OAI22_X1  g718(.A1(new_n915), .A2(new_n916), .B1(new_n919), .B2(KEYINPUT57), .ZN(new_n920));
  AND2_X1   g719(.A1(new_n916), .A2(new_n915), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n914), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT120), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  OAI211_X1 g723(.A(KEYINPUT120), .B(new_n914), .C1(new_n920), .C2(new_n921), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n924), .A2(G148gat), .A3(new_n925), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n926), .A2(KEYINPUT59), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT121), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n926), .A2(KEYINPUT121), .A3(KEYINPUT59), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n913), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NOR3_X1   g730(.A1(new_n894), .A2(G148gat), .A3(new_n627), .ZN(new_n932));
  OAI21_X1  g731(.A(KEYINPUT122), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT122), .ZN(new_n934));
  INV_X1    g733(.A(new_n932), .ZN(new_n935));
  AND3_X1   g734(.A1(new_n926), .A2(KEYINPUT121), .A3(KEYINPUT59), .ZN(new_n936));
  AOI21_X1  g735(.A(KEYINPUT121), .B1(new_n926), .B2(KEYINPUT59), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  OAI211_X1 g737(.A(new_n934), .B(new_n935), .C1(new_n938), .C2(new_n913), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n933), .A2(new_n939), .ZN(G1345gat));
  OAI21_X1  g739(.A(G155gat), .B1(new_n907), .B2(new_n714), .ZN(new_n941));
  INV_X1    g740(.A(new_n894), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n942), .A2(new_n384), .A3(new_n681), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n941), .A2(new_n943), .ZN(G1346gat));
  OR3_X1    g743(.A1(new_n907), .A2(new_n385), .A3(new_n680), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n385), .B1(new_n894), .B2(new_n680), .ZN(new_n946));
  AND2_X1   g745(.A1(new_n945), .A2(new_n946), .ZN(G1347gat));
  NAND3_X1  g746(.A1(new_n867), .A2(new_n434), .A3(new_n474), .ZN(new_n948));
  NOR3_X1   g747(.A1(new_n948), .A2(new_n283), .A3(new_n281), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n723), .B1(new_n863), .B2(new_n864), .ZN(new_n950));
  NAND4_X1  g749(.A1(new_n950), .A2(new_n538), .A3(new_n474), .A4(new_n563), .ZN(new_n951));
  INV_X1    g750(.A(new_n951), .ZN(new_n952));
  AOI21_X1  g751(.A(G169gat), .B1(new_n952), .B2(new_n280), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n949), .A2(new_n953), .ZN(G1348gat));
  OAI21_X1  g753(.A(G176gat), .B1(new_n948), .B2(new_n713), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n952), .A2(new_n284), .A3(new_n626), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n955), .A2(new_n956), .ZN(G1349gat));
  OAI21_X1  g756(.A(G183gat), .B1(new_n948), .B2(new_n714), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n952), .A2(new_n293), .A3(new_n681), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  XNOR2_X1  g759(.A(new_n960), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g760(.A(G190gat), .B1(new_n948), .B2(new_n680), .ZN(new_n962));
  XOR2_X1   g761(.A(KEYINPUT123), .B(KEYINPUT61), .Z(new_n963));
  XNOR2_X1  g762(.A(new_n962), .B(new_n963), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n952), .A2(new_n294), .A3(new_n702), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n964), .A2(new_n965), .ZN(G1351gat));
  AND4_X1   g765(.A1(new_n512), .A2(new_n374), .A3(new_n474), .A4(new_n950), .ZN(new_n967));
  AOI21_X1  g766(.A(G197gat), .B1(new_n967), .B2(new_n280), .ZN(new_n968));
  OR2_X1    g767(.A1(new_n920), .A2(new_n921), .ZN(new_n969));
  NOR3_X1   g768(.A1(new_n734), .A2(new_n723), .A3(new_n475), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g770(.A(new_n971), .ZN(new_n972));
  AND2_X1   g771(.A1(new_n280), .A2(G197gat), .ZN(new_n973));
  AOI21_X1  g772(.A(new_n968), .B1(new_n972), .B2(new_n973), .ZN(G1352gat));
  XOR2_X1   g773(.A(KEYINPUT124), .B(G204gat), .Z(new_n975));
  NOR2_X1   g774(.A1(new_n627), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n967), .A2(new_n976), .ZN(new_n977));
  XOR2_X1   g776(.A(new_n977), .B(KEYINPUT62), .Z(new_n978));
  OAI21_X1  g777(.A(new_n975), .B1(new_n971), .B2(new_n713), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  XOR2_X1   g779(.A(new_n980), .B(KEYINPUT125), .Z(G1353gat));
  NAND3_X1  g780(.A1(new_n972), .A2(KEYINPUT126), .A3(new_n681), .ZN(new_n982));
  INV_X1    g781(.A(KEYINPUT126), .ZN(new_n983));
  OAI21_X1  g782(.A(new_n983), .B1(new_n971), .B2(new_n659), .ZN(new_n984));
  INV_X1    g783(.A(KEYINPUT63), .ZN(new_n985));
  AOI21_X1  g784(.A(new_n444), .B1(KEYINPUT127), .B2(new_n985), .ZN(new_n986));
  NAND3_X1  g785(.A1(new_n982), .A2(new_n984), .A3(new_n986), .ZN(new_n987));
  NOR2_X1   g786(.A1(new_n985), .A2(KEYINPUT127), .ZN(new_n988));
  OR2_X1    g787(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n967), .A2(new_n444), .A3(new_n681), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n987), .A2(new_n988), .ZN(new_n991));
  NAND3_X1  g790(.A1(new_n989), .A2(new_n990), .A3(new_n991), .ZN(G1354gat));
  OAI21_X1  g791(.A(G218gat), .B1(new_n971), .B2(new_n680), .ZN(new_n993));
  NAND3_X1  g792(.A1(new_n967), .A2(new_n445), .A3(new_n702), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n993), .A2(new_n994), .ZN(G1355gat));
endmodule


