

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715;

  INV_X1 U367 ( .A(G953), .ZN(n702) );
  NOR2_X2 U368 ( .A1(n681), .A2(n589), .ZN(n592) );
  NOR2_X2 U369 ( .A1(n681), .A2(n675), .ZN(n676) );
  XNOR2_X2 U370 ( .A(n385), .B(G143), .ZN(n378) );
  AND2_X1 U371 ( .A1(n507), .A2(n506), .ZN(n508) );
  NOR2_X1 U372 ( .A1(n538), .A2(n537), .ZN(n539) );
  AND2_X1 U373 ( .A1(n359), .A2(n358), .ZN(n596) );
  BUF_X1 U374 ( .A(n668), .Z(n671) );
  AND2_X2 U375 ( .A1(n668), .A2(n669), .ZN(n677) );
  NAND2_X1 U376 ( .A1(n580), .A2(n579), .ZN(n668) );
  XNOR2_X1 U377 ( .A(n392), .B(n391), .ZN(n711) );
  NOR2_X1 U378 ( .A1(n513), .A2(n528), .ZN(n497) );
  XNOR2_X1 U379 ( .A(n569), .B(n438), .ZN(n561) );
  NOR2_X1 U380 ( .A1(G902), .A2(n594), .ZN(n486) );
  XNOR2_X1 U381 ( .A(n672), .B(n350), .ZN(n673) );
  XNOR2_X2 U382 ( .A(G128), .B(KEYINPUT78), .ZN(n385) );
  XNOR2_X2 U383 ( .A(n698), .B(G146), .ZN(n484) );
  XNOR2_X2 U384 ( .A(n406), .B(n394), .ZN(n698) );
  XNOR2_X2 U385 ( .A(n636), .B(KEYINPUT6), .ZN(n528) );
  XNOR2_X1 U386 ( .A(n429), .B(n355), .ZN(n431) );
  XNOR2_X1 U387 ( .A(n430), .B(n448), .ZN(n355) );
  NOR2_X1 U388 ( .A1(n561), .A2(n445), .ZN(n447) );
  XOR2_X1 U389 ( .A(G125), .B(G146), .Z(n448) );
  XNOR2_X1 U390 ( .A(n396), .B(G131), .ZN(n449) );
  INV_X1 U391 ( .A(KEYINPUT67), .ZN(n396) );
  XOR2_X1 U392 ( .A(KEYINPUT10), .B(n448), .Z(n468) );
  XNOR2_X1 U393 ( .A(n682), .B(n413), .ZN(n429) );
  XNOR2_X1 U394 ( .A(n484), .B(n483), .ZN(n594) );
  XNOR2_X1 U395 ( .A(n366), .B(n365), .ZN(n364) );
  XNOR2_X1 U396 ( .A(G128), .B(G110), .ZN(n365) );
  XNOR2_X1 U397 ( .A(n367), .B(G119), .ZN(n366) );
  XNOR2_X1 U398 ( .A(n363), .B(n362), .ZN(n361) );
  XNOR2_X1 U399 ( .A(KEYINPUT88), .B(KEYINPUT24), .ZN(n363) );
  XNOR2_X1 U400 ( .A(KEYINPUT23), .B(KEYINPUT89), .ZN(n362) );
  XNOR2_X1 U401 ( .A(n436), .B(n388), .ZN(n535) );
  XNOR2_X1 U402 ( .A(n435), .B(KEYINPUT84), .ZN(n388) );
  XNOR2_X1 U403 ( .A(n434), .B(n433), .ZN(n435) );
  NAND2_X1 U404 ( .A1(n535), .A2(n642), .ZN(n569) );
  AND2_X1 U405 ( .A1(n658), .A2(KEYINPUT34), .ZN(n383) );
  XNOR2_X1 U406 ( .A(n356), .B(n347), .ZN(n490) );
  AND2_X1 U407 ( .A1(n542), .A2(n344), .ZN(n357) );
  NOR2_X1 U408 ( .A1(G902), .A2(n581), .ZN(n464) );
  NAND2_X1 U409 ( .A1(n677), .A2(G472), .ZN(n360) );
  XNOR2_X1 U410 ( .A(n427), .B(n387), .ZN(n386) );
  INV_X1 U411 ( .A(KEYINPUT18), .ZN(n387) );
  NOR2_X1 U412 ( .A1(n566), .A2(n623), .ZN(n373) );
  AND2_X1 U413 ( .A1(n377), .A2(n376), .ZN(n375) );
  NOR2_X1 U414 ( .A1(n393), .A2(n573), .ZN(n376) );
  XNOR2_X1 U415 ( .A(n449), .B(n395), .ZN(n394) );
  XNOR2_X1 U416 ( .A(n367), .B(KEYINPUT4), .ZN(n395) );
  XNOR2_X1 U417 ( .A(G116), .B(KEYINPUT3), .ZN(n424) );
  XOR2_X1 U418 ( .A(G140), .B(KEYINPUT68), .Z(n466) );
  NAND2_X1 U419 ( .A1(G237), .A2(G234), .ZN(n439) );
  XNOR2_X1 U420 ( .A(KEYINPUT38), .B(n557), .ZN(n641) );
  AND2_X1 U421 ( .A1(n344), .A2(n522), .ZN(n627) );
  XNOR2_X1 U422 ( .A(n412), .B(n411), .ZN(n682) );
  XNOR2_X1 U423 ( .A(G107), .B(G110), .ZN(n411) );
  XNOR2_X1 U424 ( .A(n478), .B(n426), .ZN(n683) );
  XNOR2_X1 U425 ( .A(n425), .B(G122), .ZN(n426) );
  XOR2_X1 U426 ( .A(KEYINPUT73), .B(KEYINPUT16), .Z(n425) );
  XNOR2_X1 U427 ( .A(n378), .B(n397), .ZN(n406) );
  INV_X1 U428 ( .A(G134), .ZN(n397) );
  XOR2_X1 U429 ( .A(KEYINPUT7), .B(G116), .Z(n402) );
  XNOR2_X1 U430 ( .A(G104), .B(G113), .ZN(n450) );
  NOR2_X1 U431 ( .A1(n531), .A2(n530), .ZN(n567) );
  XNOR2_X1 U432 ( .A(n498), .B(KEYINPUT100), .ZN(n556) );
  INV_X1 U433 ( .A(n535), .ZN(n557) );
  INV_X1 U434 ( .A(KEYINPUT19), .ZN(n438) );
  NAND2_X1 U435 ( .A1(n540), .A2(n627), .ZN(n547) );
  XNOR2_X1 U436 ( .A(n364), .B(n361), .ZN(n471) );
  XNOR2_X1 U437 ( .A(n390), .B(n389), .ZN(n714) );
  INV_X1 U438 ( .A(KEYINPUT42), .ZN(n389) );
  OR2_X1 U439 ( .A1(n659), .A2(n562), .ZN(n390) );
  INV_X1 U440 ( .A(KEYINPUT40), .ZN(n391) );
  XNOR2_X1 U441 ( .A(n379), .B(KEYINPUT35), .ZN(n713) );
  NAND2_X1 U442 ( .A1(n343), .A2(n496), .ZN(n382) );
  AND2_X1 U443 ( .A1(n490), .A2(n489), .ZN(n493) );
  XNOR2_X1 U444 ( .A(n360), .B(n348), .ZN(n359) );
  XNOR2_X1 U445 ( .A(n351), .B(n581), .ZN(n582) );
  NAND2_X1 U446 ( .A1(n677), .A2(G478), .ZN(n351) );
  INV_X1 U447 ( .A(KEYINPUT116), .ZN(n352) );
  NOR2_X1 U448 ( .A1(n658), .A2(KEYINPUT34), .ZN(n343) );
  XOR2_X1 U449 ( .A(n630), .B(KEYINPUT92), .Z(n344) );
  XOR2_X1 U450 ( .A(G113), .B(G119), .Z(n345) );
  INV_X1 U451 ( .A(G137), .ZN(n367) );
  XOR2_X1 U452 ( .A(n556), .B(KEYINPUT76), .Z(n346) );
  XOR2_X1 U453 ( .A(KEYINPUT22), .B(KEYINPUT72), .Z(n347) );
  XOR2_X1 U454 ( .A(n594), .B(n593), .Z(n348) );
  XOR2_X1 U455 ( .A(n664), .B(n665), .Z(n349) );
  INV_X1 U456 ( .A(n572), .ZN(n573) );
  XNOR2_X1 U457 ( .A(KEYINPUT48), .B(KEYINPUT80), .ZN(n572) );
  XNOR2_X1 U458 ( .A(KEYINPUT59), .B(KEYINPUT117), .ZN(n350) );
  NOR2_X1 U459 ( .A1(G952), .A2(n702), .ZN(n681) );
  INV_X1 U460 ( .A(n681), .ZN(n358) );
  AND2_X2 U461 ( .A1(n559), .A2(n641), .ZN(n554) );
  NOR2_X2 U462 ( .A1(n552), .A2(n551), .ZN(n559) );
  NAND2_X1 U463 ( .A1(n473), .A2(G221), .ZN(n423) );
  XNOR2_X1 U464 ( .A(n422), .B(KEYINPUT90), .ZN(n473) );
  NOR2_X1 U465 ( .A1(n547), .A2(n546), .ZN(n549) );
  NOR2_X1 U466 ( .A1(n623), .A2(n572), .ZN(n369) );
  NOR2_X1 U467 ( .A1(n383), .A2(n381), .ZN(n380) );
  XNOR2_X1 U468 ( .A(n353), .B(n352), .ZN(G54) );
  NAND2_X1 U469 ( .A1(n667), .A2(n358), .ZN(n353) );
  NAND2_X1 U470 ( .A1(n518), .A2(n354), .ZN(n521) );
  AND2_X1 U471 ( .A1(n517), .A2(n519), .ZN(n354) );
  NAND2_X1 U472 ( .A1(n496), .A2(n357), .ZN(n356) );
  INV_X1 U473 ( .A(n522), .ZN(n631) );
  XNOR2_X2 U474 ( .A(n477), .B(n476), .ZN(n522) );
  NAND2_X1 U475 ( .A1(n371), .A2(n368), .ZN(n370) );
  INV_X1 U476 ( .A(n566), .ZN(n368) );
  NOR2_X1 U477 ( .A1(n565), .A2(n393), .ZN(n371) );
  NAND2_X1 U478 ( .A1(n370), .A2(n369), .ZN(n374) );
  NAND2_X1 U479 ( .A1(n374), .A2(n372), .ZN(n576) );
  NAND2_X1 U480 ( .A1(n373), .A2(n375), .ZN(n372) );
  INV_X1 U481 ( .A(n565), .ZN(n377) );
  XNOR2_X1 U482 ( .A(n378), .B(n386), .ZN(n428) );
  NAND2_X1 U483 ( .A1(n380), .A2(n382), .ZN(n379) );
  NAND2_X1 U484 ( .A1(n384), .A2(n346), .ZN(n381) );
  XNOR2_X2 U485 ( .A(n540), .B(KEYINPUT1), .ZN(n626) );
  NAND2_X1 U486 ( .A1(n510), .A2(KEYINPUT34), .ZN(n384) );
  XNOR2_X1 U487 ( .A(n544), .B(n543), .ZN(n659) );
  NOR2_X2 U488 ( .A1(n711), .A2(n714), .ZN(n555) );
  NAND2_X1 U489 ( .A1(n575), .A2(n613), .ZN(n392) );
  XNOR2_X2 U490 ( .A(n554), .B(n553), .ZN(n575) );
  INV_X1 U491 ( .A(n620), .ZN(n393) );
  XNOR2_X1 U492 ( .A(n588), .B(n398), .ZN(n589) );
  XNOR2_X1 U493 ( .A(n666), .B(n349), .ZN(n667) );
  XOR2_X2 U494 ( .A(G902), .B(KEYINPUT15), .Z(n577) );
  XOR2_X1 U495 ( .A(n587), .B(n586), .Z(n398) );
  XNOR2_X1 U496 ( .A(n499), .B(KEYINPUT82), .ZN(n494) );
  XNOR2_X1 U497 ( .A(KEYINPUT0), .B(KEYINPUT66), .ZN(n446) );
  XNOR2_X1 U498 ( .A(n484), .B(n417), .ZN(n664) );
  XNOR2_X1 U499 ( .A(n447), .B(n446), .ZN(n496) );
  XNOR2_X1 U500 ( .A(n478), .B(n482), .ZN(n483) );
  XNOR2_X1 U501 ( .A(n402), .B(G107), .ZN(n403) );
  BUF_X1 U502 ( .A(n624), .Z(n625) );
  INV_X1 U503 ( .A(KEYINPUT74), .ZN(n548) );
  XOR2_X1 U504 ( .A(n464), .B(G478), .Z(n507) );
  XNOR2_X1 U505 ( .A(n674), .B(n673), .ZN(n675) );
  XNOR2_X1 U506 ( .A(n592), .B(n591), .ZN(G51) );
  XOR2_X1 U507 ( .A(G122), .B(KEYINPUT9), .Z(n401) );
  NAND2_X1 U508 ( .A1(G234), .A2(n702), .ZN(n399) );
  XOR2_X1 U509 ( .A(KEYINPUT8), .B(n399), .Z(n469) );
  NAND2_X1 U510 ( .A1(G217), .A2(n469), .ZN(n400) );
  XNOR2_X1 U511 ( .A(n401), .B(n400), .ZN(n405) );
  XNOR2_X1 U512 ( .A(n406), .B(n403), .ZN(n404) );
  XOR2_X1 U513 ( .A(n405), .B(n404), .Z(n581) );
  INV_X1 U514 ( .A(KEYINPUT70), .ZN(n413) );
  INV_X1 U515 ( .A(G104), .ZN(n407) );
  NAND2_X1 U516 ( .A1(G101), .A2(n407), .ZN(n410) );
  INV_X1 U517 ( .A(G101), .ZN(n408) );
  NAND2_X1 U518 ( .A1(n408), .A2(G104), .ZN(n409) );
  NAND2_X1 U519 ( .A1(n410), .A2(n409), .ZN(n412) );
  XOR2_X1 U520 ( .A(n466), .B(KEYINPUT75), .Z(n415) );
  NAND2_X1 U521 ( .A1(G227), .A2(n702), .ZN(n414) );
  XNOR2_X1 U522 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U523 ( .A(n429), .B(n416), .ZN(n417) );
  NOR2_X1 U524 ( .A1(G902), .A2(n664), .ZN(n419) );
  XNOR2_X1 U525 ( .A(KEYINPUT69), .B(G469), .ZN(n418) );
  XNOR2_X2 U526 ( .A(n419), .B(n418), .ZN(n540) );
  INV_X1 U527 ( .A(n626), .ZN(n465) );
  INV_X1 U528 ( .A(n577), .ZN(n420) );
  NAND2_X1 U529 ( .A1(n420), .A2(G234), .ZN(n421) );
  XNOR2_X1 U530 ( .A(n421), .B(KEYINPUT20), .ZN(n422) );
  XNOR2_X1 U531 ( .A(n423), .B(KEYINPUT21), .ZN(n630) );
  XNOR2_X1 U532 ( .A(n345), .B(n424), .ZN(n478) );
  NAND2_X1 U533 ( .A1(G224), .A2(n702), .ZN(n427) );
  XNOR2_X1 U534 ( .A(n683), .B(n428), .ZN(n432) );
  XOR2_X1 U535 ( .A(KEYINPUT17), .B(KEYINPUT4), .Z(n430) );
  XNOR2_X1 U536 ( .A(n432), .B(n431), .ZN(n585) );
  NOR2_X1 U537 ( .A1(n577), .A2(n585), .ZN(n436) );
  OR2_X1 U538 ( .A1(G902), .A2(G237), .ZN(n437) );
  AND2_X1 U539 ( .A1(G210), .A2(n437), .ZN(n434) );
  XOR2_X1 U540 ( .A(KEYINPUT85), .B(KEYINPUT79), .Z(n433) );
  NAND2_X1 U541 ( .A1(G214), .A2(n437), .ZN(n642) );
  XNOR2_X1 U542 ( .A(n439), .B(KEYINPUT14), .ZN(n441) );
  NAND2_X1 U543 ( .A1(G952), .A2(n441), .ZN(n440) );
  XOR2_X1 U544 ( .A(KEYINPUT86), .B(n440), .Z(n654) );
  NAND2_X1 U545 ( .A1(n702), .A2(n654), .ZN(n526) );
  INV_X1 U546 ( .A(n526), .ZN(n444) );
  NAND2_X1 U547 ( .A1(G902), .A2(n441), .ZN(n523) );
  NOR2_X1 U548 ( .A1(G898), .A2(n702), .ZN(n442) );
  XNOR2_X1 U549 ( .A(KEYINPUT87), .B(n442), .ZN(n684) );
  NOR2_X1 U550 ( .A1(n523), .A2(n684), .ZN(n443) );
  NOR2_X1 U551 ( .A1(n444), .A2(n443), .ZN(n445) );
  XNOR2_X1 U552 ( .A(n450), .B(n449), .ZN(n451) );
  XOR2_X1 U553 ( .A(n468), .B(n451), .Z(n453) );
  NOR2_X1 U554 ( .A1(G953), .A2(G237), .ZN(n479) );
  NAND2_X1 U555 ( .A1(n479), .A2(G214), .ZN(n452) );
  XNOR2_X1 U556 ( .A(n453), .B(n452), .ZN(n461) );
  XOR2_X1 U557 ( .A(KEYINPUT95), .B(KEYINPUT96), .Z(n455) );
  XNOR2_X1 U558 ( .A(G143), .B(G122), .ZN(n454) );
  XNOR2_X1 U559 ( .A(n455), .B(n454), .ZN(n459) );
  XOR2_X1 U560 ( .A(G140), .B(KEYINPUT12), .Z(n457) );
  XNOR2_X1 U561 ( .A(KEYINPUT94), .B(KEYINPUT11), .ZN(n456) );
  XNOR2_X1 U562 ( .A(n457), .B(n456), .ZN(n458) );
  XOR2_X1 U563 ( .A(n459), .B(n458), .Z(n460) );
  XNOR2_X1 U564 ( .A(n461), .B(n460), .ZN(n672) );
  NOR2_X1 U565 ( .A1(G902), .A2(n672), .ZN(n463) );
  XNOR2_X1 U566 ( .A(KEYINPUT13), .B(G475), .ZN(n462) );
  XNOR2_X1 U567 ( .A(n463), .B(n462), .ZN(n505) );
  NOR2_X1 U568 ( .A1(n505), .A2(n507), .ZN(n542) );
  NAND2_X1 U569 ( .A1(n465), .A2(n490), .ZN(n504) );
  INV_X1 U570 ( .A(n466), .ZN(n467) );
  XNOR2_X1 U571 ( .A(n468), .B(n467), .ZN(n697) );
  NAND2_X1 U572 ( .A1(G221), .A2(n469), .ZN(n470) );
  XNOR2_X1 U573 ( .A(n471), .B(n470), .ZN(n472) );
  XNOR2_X1 U574 ( .A(n697), .B(n472), .ZN(n679) );
  NOR2_X1 U575 ( .A1(n679), .A2(G902), .ZN(n477) );
  XOR2_X1 U576 ( .A(KEYINPUT91), .B(KEYINPUT25), .Z(n475) );
  NAND2_X1 U577 ( .A1(G217), .A2(n473), .ZN(n474) );
  XNOR2_X1 U578 ( .A(n475), .B(n474), .ZN(n476) );
  XOR2_X1 U579 ( .A(G101), .B(KEYINPUT5), .Z(n481) );
  NAND2_X1 U580 ( .A1(n479), .A2(G210), .ZN(n480) );
  XNOR2_X1 U581 ( .A(n481), .B(n480), .ZN(n482) );
  INV_X1 U582 ( .A(G472), .ZN(n485) );
  XNOR2_X2 U583 ( .A(n486), .B(n485), .ZN(n636) );
  INV_X1 U584 ( .A(n636), .ZN(n538) );
  NAND2_X1 U585 ( .A1(n631), .A2(n538), .ZN(n487) );
  NOR2_X1 U586 ( .A1(n504), .A2(n487), .ZN(n606) );
  AND2_X1 U587 ( .A1(n626), .A2(n528), .ZN(n488) );
  AND2_X1 U588 ( .A1(n631), .A2(n488), .ZN(n489) );
  XOR2_X1 U589 ( .A(KEYINPUT32), .B(KEYINPUT77), .Z(n491) );
  XNOR2_X1 U590 ( .A(KEYINPUT64), .B(n491), .ZN(n492) );
  XNOR2_X1 U591 ( .A(n493), .B(n492), .ZN(n712) );
  NOR2_X1 U592 ( .A1(n606), .A2(n712), .ZN(n495) );
  INV_X1 U593 ( .A(KEYINPUT44), .ZN(n499) );
  XNOR2_X1 U594 ( .A(n495), .B(n494), .ZN(n501) );
  INV_X1 U595 ( .A(n496), .ZN(n510) );
  NAND2_X1 U596 ( .A1(n627), .A2(n626), .ZN(n513) );
  XNOR2_X1 U597 ( .A(n497), .B(KEYINPUT33), .ZN(n658) );
  NAND2_X1 U598 ( .A1(n507), .A2(n505), .ZN(n498) );
  NAND2_X1 U599 ( .A1(n499), .A2(n713), .ZN(n500) );
  NAND2_X1 U600 ( .A1(n501), .A2(n500), .ZN(n519) );
  NAND2_X1 U601 ( .A1(n713), .A2(KEYINPUT44), .ZN(n502) );
  XOR2_X1 U602 ( .A(KEYINPUT81), .B(n502), .Z(n518) );
  NAND2_X1 U603 ( .A1(n522), .A2(n528), .ZN(n503) );
  NOR2_X1 U604 ( .A1(n504), .A2(n503), .ZN(n597) );
  INV_X1 U605 ( .A(n505), .ZN(n506) );
  NOR2_X1 U606 ( .A1(n506), .A2(n507), .ZN(n613) );
  XOR2_X2 U607 ( .A(n508), .B(KEYINPUT97), .Z(n616) );
  XNOR2_X1 U608 ( .A(KEYINPUT98), .B(n616), .ZN(n574) );
  OR2_X1 U609 ( .A1(n613), .A2(n574), .ZN(n509) );
  XOR2_X1 U610 ( .A(KEYINPUT99), .B(n509), .Z(n563) );
  INV_X1 U611 ( .A(n563), .ZN(n646) );
  NOR2_X1 U612 ( .A1(n547), .A2(n510), .ZN(n511) );
  NAND2_X1 U613 ( .A1(n511), .A2(n538), .ZN(n512) );
  XNOR2_X1 U614 ( .A(KEYINPUT93), .B(n512), .ZN(n601) );
  NOR2_X1 U615 ( .A1(n538), .A2(n513), .ZN(n638) );
  NAND2_X1 U616 ( .A1(n496), .A2(n638), .ZN(n514) );
  XNOR2_X1 U617 ( .A(KEYINPUT31), .B(n514), .ZN(n617) );
  NOR2_X1 U618 ( .A1(n601), .A2(n617), .ZN(n515) );
  NOR2_X1 U619 ( .A1(n646), .A2(n515), .ZN(n516) );
  NOR2_X1 U620 ( .A1(n597), .A2(n516), .ZN(n517) );
  INV_X1 U621 ( .A(KEYINPUT45), .ZN(n520) );
  XNOR2_X1 U622 ( .A(n521), .B(n520), .ZN(n688) );
  INV_X1 U623 ( .A(n613), .ZN(n531) );
  NOR2_X1 U624 ( .A1(n630), .A2(n522), .ZN(n527) );
  NOR2_X1 U625 ( .A1(G900), .A2(n523), .ZN(n524) );
  NAND2_X1 U626 ( .A1(G953), .A2(n524), .ZN(n525) );
  NAND2_X1 U627 ( .A1(n526), .A2(n525), .ZN(n545) );
  NAND2_X1 U628 ( .A1(n527), .A2(n545), .ZN(n537) );
  NOR2_X1 U629 ( .A1(n537), .A2(n528), .ZN(n529) );
  XNOR2_X1 U630 ( .A(n529), .B(KEYINPUT101), .ZN(n530) );
  NAND2_X1 U631 ( .A1(n567), .A2(n642), .ZN(n532) );
  NOR2_X1 U632 ( .A1(n626), .A2(n532), .ZN(n534) );
  XNOR2_X1 U633 ( .A(KEYINPUT43), .B(KEYINPUT102), .ZN(n533) );
  XNOR2_X1 U634 ( .A(n534), .B(n533), .ZN(n536) );
  NOR2_X1 U635 ( .A1(n536), .A2(n535), .ZN(n623) );
  XNOR2_X1 U636 ( .A(KEYINPUT28), .B(n539), .ZN(n541) );
  NAND2_X1 U637 ( .A1(n541), .A2(n540), .ZN(n562) );
  NAND2_X1 U638 ( .A1(n642), .A2(n641), .ZN(n645) );
  INV_X1 U639 ( .A(n542), .ZN(n644) );
  NOR2_X1 U640 ( .A1(n645), .A2(n644), .ZN(n544) );
  XOR2_X1 U641 ( .A(KEYINPUT41), .B(KEYINPUT103), .Z(n543) );
  INV_X1 U642 ( .A(n545), .ZN(n546) );
  XNOR2_X1 U643 ( .A(n549), .B(n548), .ZN(n552) );
  NAND2_X1 U644 ( .A1(n636), .A2(n642), .ZN(n550) );
  XNOR2_X1 U645 ( .A(KEYINPUT30), .B(n550), .ZN(n551) );
  XNOR2_X1 U646 ( .A(KEYINPUT39), .B(KEYINPUT71), .ZN(n553) );
  XNOR2_X1 U647 ( .A(n555), .B(KEYINPUT46), .ZN(n560) );
  NOR2_X1 U648 ( .A1(n557), .A2(n556), .ZN(n558) );
  NAND2_X1 U649 ( .A1(n559), .A2(n558), .ZN(n610) );
  NAND2_X1 U650 ( .A1(n560), .A2(n610), .ZN(n566) );
  NOR2_X1 U651 ( .A1(n562), .A2(n561), .ZN(n611) );
  NAND2_X1 U652 ( .A1(n563), .A2(n611), .ZN(n564) );
  XNOR2_X1 U653 ( .A(n564), .B(KEYINPUT47), .ZN(n565) );
  XOR2_X1 U654 ( .A(KEYINPUT104), .B(n567), .Z(n568) );
  NOR2_X1 U655 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U656 ( .A(n570), .B(KEYINPUT36), .ZN(n571) );
  NAND2_X1 U657 ( .A1(n571), .A2(n626), .ZN(n620) );
  NAND2_X1 U658 ( .A1(n575), .A2(n574), .ZN(n622) );
  NAND2_X1 U659 ( .A1(n576), .A2(n622), .ZN(n696) );
  NOR2_X2 U660 ( .A1(n688), .A2(n696), .ZN(n624) );
  NAND2_X1 U661 ( .A1(n624), .A2(n577), .ZN(n580) );
  NAND2_X1 U662 ( .A1(n577), .A2(KEYINPUT2), .ZN(n578) );
  XOR2_X1 U663 ( .A(KEYINPUT65), .B(n578), .Z(n579) );
  NAND2_X1 U664 ( .A1(KEYINPUT2), .A2(n624), .ZN(n669) );
  NOR2_X2 U665 ( .A1(n582), .A2(n681), .ZN(n583) );
  XNOR2_X1 U666 ( .A(n583), .B(KEYINPUT118), .ZN(G63) );
  AND2_X1 U667 ( .A1(G210), .A2(n669), .ZN(n584) );
  NAND2_X1 U668 ( .A1(n584), .A2(n671), .ZN(n588) );
  XOR2_X1 U669 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n587) );
  XNOR2_X1 U670 ( .A(n585), .B(KEYINPUT83), .ZN(n586) );
  INV_X1 U671 ( .A(KEYINPUT115), .ZN(n590) );
  XNOR2_X1 U672 ( .A(n590), .B(KEYINPUT56), .ZN(n591) );
  XOR2_X1 U673 ( .A(KEYINPUT105), .B(KEYINPUT62), .Z(n593) );
  XOR2_X1 U674 ( .A(KEYINPUT63), .B(KEYINPUT106), .Z(n595) );
  XNOR2_X1 U675 ( .A(n596), .B(n595), .ZN(G57) );
  XOR2_X1 U676 ( .A(G101), .B(n597), .Z(G3) );
  XOR2_X1 U677 ( .A(KEYINPUT107), .B(KEYINPUT108), .Z(n599) );
  NAND2_X1 U678 ( .A1(n601), .A2(n613), .ZN(n598) );
  XNOR2_X1 U679 ( .A(n599), .B(n598), .ZN(n600) );
  XNOR2_X1 U680 ( .A(G104), .B(n600), .ZN(G6) );
  XOR2_X1 U681 ( .A(G107), .B(KEYINPUT109), .Z(n603) );
  NAND2_X1 U682 ( .A1(n601), .A2(n616), .ZN(n602) );
  XNOR2_X1 U683 ( .A(n603), .B(n602), .ZN(n605) );
  XOR2_X1 U684 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n604) );
  XNOR2_X1 U685 ( .A(n605), .B(n604), .ZN(G9) );
  XOR2_X1 U686 ( .A(G110), .B(n606), .Z(G12) );
  XOR2_X1 U687 ( .A(KEYINPUT110), .B(KEYINPUT29), .Z(n608) );
  NAND2_X1 U688 ( .A1(n611), .A2(n616), .ZN(n607) );
  XNOR2_X1 U689 ( .A(n608), .B(n607), .ZN(n609) );
  XNOR2_X1 U690 ( .A(G128), .B(n609), .ZN(G30) );
  XNOR2_X1 U691 ( .A(G143), .B(n610), .ZN(G45) );
  NAND2_X1 U692 ( .A1(n611), .A2(n613), .ZN(n612) );
  XNOR2_X1 U693 ( .A(n612), .B(G146), .ZN(G48) );
  XOR2_X1 U694 ( .A(G113), .B(KEYINPUT111), .Z(n615) );
  NAND2_X1 U695 ( .A1(n617), .A2(n613), .ZN(n614) );
  XNOR2_X1 U696 ( .A(n615), .B(n614), .ZN(G15) );
  NAND2_X1 U697 ( .A1(n617), .A2(n616), .ZN(n618) );
  XNOR2_X1 U698 ( .A(n618), .B(G116), .ZN(G18) );
  XOR2_X1 U699 ( .A(KEYINPUT112), .B(KEYINPUT37), .Z(n619) );
  XNOR2_X1 U700 ( .A(n620), .B(n619), .ZN(n621) );
  XNOR2_X1 U701 ( .A(G125), .B(n621), .ZN(G27) );
  XNOR2_X1 U702 ( .A(G134), .B(n622), .ZN(G36) );
  XOR2_X1 U703 ( .A(G140), .B(n623), .Z(G42) );
  XNOR2_X1 U704 ( .A(KEYINPUT2), .B(n625), .ZN(n657) );
  NOR2_X1 U705 ( .A1(n627), .A2(n626), .ZN(n629) );
  XNOR2_X1 U706 ( .A(KEYINPUT50), .B(KEYINPUT113), .ZN(n628) );
  XNOR2_X1 U707 ( .A(n629), .B(n628), .ZN(n634) );
  NAND2_X1 U708 ( .A1(n631), .A2(n630), .ZN(n632) );
  XOR2_X1 U709 ( .A(KEYINPUT49), .B(n632), .Z(n633) );
  NAND2_X1 U710 ( .A1(n634), .A2(n633), .ZN(n635) );
  NOR2_X1 U711 ( .A1(n636), .A2(n635), .ZN(n637) );
  NOR2_X1 U712 ( .A1(n638), .A2(n637), .ZN(n639) );
  XOR2_X1 U713 ( .A(KEYINPUT51), .B(n639), .Z(n640) );
  NOR2_X1 U714 ( .A1(n659), .A2(n640), .ZN(n652) );
  NOR2_X1 U715 ( .A1(n642), .A2(n641), .ZN(n643) );
  NOR2_X1 U716 ( .A1(n644), .A2(n643), .ZN(n649) );
  NOR2_X1 U717 ( .A1(n646), .A2(n645), .ZN(n647) );
  XNOR2_X1 U718 ( .A(n647), .B(KEYINPUT114), .ZN(n648) );
  NOR2_X1 U719 ( .A1(n649), .A2(n648), .ZN(n650) );
  NOR2_X1 U720 ( .A1(n650), .A2(n658), .ZN(n651) );
  NOR2_X1 U721 ( .A1(n652), .A2(n651), .ZN(n653) );
  XOR2_X1 U722 ( .A(KEYINPUT52), .B(n653), .Z(n655) );
  NAND2_X1 U723 ( .A1(n655), .A2(n654), .ZN(n656) );
  NAND2_X1 U724 ( .A1(n657), .A2(n656), .ZN(n661) );
  NOR2_X1 U725 ( .A1(n659), .A2(n658), .ZN(n660) );
  NOR2_X1 U726 ( .A1(n661), .A2(n660), .ZN(n662) );
  NAND2_X1 U727 ( .A1(n702), .A2(n662), .ZN(n663) );
  XOR2_X1 U728 ( .A(KEYINPUT53), .B(n663), .Z(G75) );
  NAND2_X1 U729 ( .A1(n677), .A2(G469), .ZN(n666) );
  XOR2_X1 U730 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n665) );
  AND2_X1 U731 ( .A1(n669), .A2(G475), .ZN(n670) );
  NAND2_X1 U732 ( .A1(n671), .A2(n670), .ZN(n674) );
  XNOR2_X1 U733 ( .A(KEYINPUT60), .B(n676), .ZN(G60) );
  NAND2_X1 U734 ( .A1(G217), .A2(n677), .ZN(n678) );
  XNOR2_X1 U735 ( .A(n679), .B(n678), .ZN(n680) );
  NOR2_X1 U736 ( .A1(n681), .A2(n680), .ZN(G66) );
  XOR2_X1 U737 ( .A(KEYINPUT121), .B(KEYINPUT120), .Z(n687) );
  XOR2_X1 U738 ( .A(n683), .B(n682), .Z(n685) );
  NAND2_X1 U739 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U740 ( .A(n687), .B(n686), .ZN(n695) );
  NOR2_X1 U741 ( .A1(G953), .A2(n688), .ZN(n689) );
  XNOR2_X1 U742 ( .A(n689), .B(KEYINPUT119), .ZN(n693) );
  NAND2_X1 U743 ( .A1(G953), .A2(G224), .ZN(n690) );
  XNOR2_X1 U744 ( .A(KEYINPUT61), .B(n690), .ZN(n691) );
  NAND2_X1 U745 ( .A1(n691), .A2(G898), .ZN(n692) );
  NAND2_X1 U746 ( .A1(n693), .A2(n692), .ZN(n694) );
  XOR2_X1 U747 ( .A(n695), .B(n694), .Z(G69) );
  XNOR2_X1 U748 ( .A(KEYINPUT123), .B(n696), .ZN(n701) );
  XOR2_X1 U749 ( .A(n698), .B(n697), .Z(n699) );
  XNOR2_X1 U750 ( .A(KEYINPUT122), .B(n699), .ZN(n704) );
  INV_X1 U751 ( .A(n704), .ZN(n700) );
  XNOR2_X1 U752 ( .A(n701), .B(n700), .ZN(n703) );
  NAND2_X1 U753 ( .A1(n703), .A2(n702), .ZN(n709) );
  XNOR2_X1 U754 ( .A(n704), .B(G227), .ZN(n705) );
  XNOR2_X1 U755 ( .A(n705), .B(KEYINPUT124), .ZN(n706) );
  NAND2_X1 U756 ( .A1(n706), .A2(G900), .ZN(n707) );
  NAND2_X1 U757 ( .A1(n707), .A2(G953), .ZN(n708) );
  NAND2_X1 U758 ( .A1(n709), .A2(n708), .ZN(G72) );
  XOR2_X1 U759 ( .A(G131), .B(KEYINPUT126), .Z(n710) );
  XNOR2_X1 U760 ( .A(n711), .B(n710), .ZN(G33) );
  XOR2_X1 U761 ( .A(n712), .B(G119), .Z(G21) );
  XOR2_X1 U762 ( .A(n713), .B(G122), .Z(G24) );
  XNOR2_X1 U763 ( .A(G137), .B(KEYINPUT125), .ZN(n715) );
  XNOR2_X1 U764 ( .A(n715), .B(n714), .ZN(G39) );
endmodule

