//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 0 0 0 1 0 1 0 0 1 1 1 1 0 1 1 0 1 1 0 1 0 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 1 1 1 1 1 1 0 0 1 0 0 0 0 0 1 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n785, new_n786, new_n787, new_n788, new_n790, new_n791, new_n792,
    new_n793, new_n795, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n825, new_n826, new_n827, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n875, new_n876,
    new_n878, new_n879, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n941, new_n942, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1017, new_n1018, new_n1019, new_n1020;
  XOR2_X1   g000(.A(KEYINPUT78), .B(KEYINPUT0), .Z(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT79), .ZN(new_n203));
  XNOR2_X1  g002(.A(G1gat), .B(G29gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(G57gat), .B(G85gat), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n205), .B(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  OAI21_X1  g007(.A(KEYINPUT76), .B1(G155gat), .B2(G162gat), .ZN(new_n209));
  XNOR2_X1  g008(.A(G141gat), .B(G148gat), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT2), .ZN(new_n211));
  AOI21_X1  g010(.A(new_n211), .B1(G155gat), .B2(G162gat), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n209), .B1(new_n210), .B2(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(G155gat), .B(G162gat), .ZN(new_n214));
  INV_X1    g013(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(G155gat), .ZN(new_n217));
  INV_X1    g016(.A(G162gat), .ZN(new_n218));
  OAI21_X1  g017(.A(KEYINPUT2), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(G141gat), .ZN(new_n220));
  INV_X1    g019(.A(G148gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(G141gat), .A2(G148gat), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n219), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n224), .A2(new_n214), .A3(new_n209), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n216), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(G134gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(G127gat), .ZN(new_n228));
  INV_X1    g027(.A(G127gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(G134gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  XNOR2_X1  g030(.A(G113gat), .B(G120gat), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n231), .B1(new_n232), .B2(KEYINPUT1), .ZN(new_n233));
  INV_X1    g032(.A(G120gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(G113gat), .ZN(new_n235));
  INV_X1    g034(.A(G113gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(G120gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(G127gat), .B(G134gat), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT1), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n238), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n233), .A2(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n226), .B(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(G225gat), .A2(G233gat), .ZN(new_n244));
  OAI21_X1  g043(.A(KEYINPUT5), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  AND3_X1   g044(.A1(new_n233), .A2(new_n241), .A3(KEYINPUT67), .ZN(new_n246));
  AOI21_X1  g045(.A(KEYINPUT67), .B1(new_n233), .B2(new_n241), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n226), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT77), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n248), .A2(new_n249), .A3(KEYINPUT4), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT3), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n226), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n216), .A2(KEYINPUT3), .A3(new_n225), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n252), .A2(new_n242), .A3(new_n253), .ZN(new_n254));
  AND3_X1   g053(.A1(new_n250), .A2(new_n244), .A3(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT4), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT67), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n242), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n233), .A2(new_n241), .A3(KEYINPUT67), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n256), .B1(new_n260), .B2(new_n226), .ZN(new_n261));
  INV_X1    g060(.A(new_n242), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n226), .A2(new_n262), .A3(new_n256), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(KEYINPUT77), .ZN(new_n264));
  OR2_X1    g063(.A1(new_n261), .A2(new_n264), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n245), .B1(new_n255), .B2(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n260), .A2(new_n256), .A3(new_n226), .ZN(new_n267));
  INV_X1    g066(.A(new_n226), .ZN(new_n268));
  OAI21_X1  g067(.A(KEYINPUT4), .B1(new_n268), .B2(new_n242), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT5), .ZN(new_n271));
  NAND4_X1  g070(.A1(new_n270), .A2(new_n271), .A3(new_n244), .A4(new_n254), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n208), .B1(new_n266), .B2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT6), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n250), .A2(new_n244), .A3(new_n254), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n261), .A2(new_n264), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  OAI211_X1 g077(.A(new_n207), .B(new_n272), .C1(new_n278), .C2(new_n245), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n274), .A2(new_n275), .A3(new_n279), .ZN(new_n280));
  OAI211_X1 g079(.A(KEYINPUT6), .B(new_n208), .C1(new_n266), .C2(new_n273), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT91), .ZN(new_n284));
  XOR2_X1   g083(.A(G15gat), .B(G43gat), .Z(new_n285));
  XNOR2_X1  g084(.A(G71gat), .B(G99gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n285), .B(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(G227gat), .A2(G233gat), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(G169gat), .ZN(new_n291));
  INV_X1    g090(.A(G176gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT26), .ZN(new_n294));
  NAND2_X1  g093(.A1(G169gat), .A2(G176gat), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n293), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(G183gat), .A2(G190gat), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n291), .A2(new_n292), .A3(KEYINPUT26), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n296), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(G190gat), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT27), .ZN(new_n301));
  OAI211_X1 g100(.A(KEYINPUT66), .B(new_n300), .C1(new_n301), .C2(G183gat), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT28), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n300), .B1(new_n301), .B2(G183gat), .ZN(new_n304));
  INV_X1    g103(.A(G183gat), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n305), .A2(KEYINPUT27), .ZN(new_n306));
  OAI211_X1 g105(.A(new_n302), .B(new_n303), .C1(new_n304), .C2(new_n306), .ZN(new_n307));
  AOI21_X1  g106(.A(G190gat), .B1(new_n305), .B2(KEYINPUT27), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n301), .A2(G183gat), .ZN(new_n309));
  OAI211_X1 g108(.A(new_n308), .B(new_n309), .C1(KEYINPUT66), .C2(KEYINPUT28), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n299), .B1(new_n307), .B2(new_n310), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n291), .A2(new_n292), .A3(KEYINPUT23), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT23), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n313), .B1(G169gat), .B2(G176gat), .ZN(new_n314));
  NAND4_X1  g113(.A1(new_n312), .A2(new_n314), .A3(KEYINPUT25), .A4(new_n295), .ZN(new_n315));
  AND3_X1   g114(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n316));
  NOR2_X1   g115(.A1(G183gat), .A2(G190gat), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT24), .ZN(new_n319));
  AOI22_X1  g118(.A1(new_n319), .A2(KEYINPUT64), .B1(G183gat), .B2(G190gat), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n320), .B1(KEYINPUT64), .B2(new_n319), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n315), .B1(new_n318), .B2(new_n321), .ZN(new_n322));
  AND3_X1   g121(.A1(new_n312), .A2(new_n314), .A3(new_n295), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n297), .A2(new_n319), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n305), .A2(new_n300), .ZN(new_n325));
  NAND3_X1  g124(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n324), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  AOI21_X1  g126(.A(KEYINPUT25), .B1(new_n323), .B2(new_n327), .ZN(new_n328));
  OAI21_X1  g127(.A(KEYINPUT65), .B1(new_n322), .B2(new_n328), .ZN(new_n329));
  AND4_X1   g128(.A1(KEYINPUT25), .A2(new_n312), .A3(new_n314), .A4(new_n295), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT64), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n297), .B1(new_n331), .B2(KEYINPUT24), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n319), .A2(KEYINPUT64), .ZN(new_n333));
  OAI211_X1 g132(.A(new_n325), .B(new_n326), .C1(new_n332), .C2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n330), .A2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT25), .ZN(new_n336));
  AOI21_X1  g135(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n337));
  NOR3_X1   g136(.A1(new_n316), .A2(new_n337), .A3(new_n317), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n312), .A2(new_n314), .A3(new_n295), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n336), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT65), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n335), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n311), .B1(new_n329), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n260), .A2(KEYINPUT68), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT68), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n258), .A2(new_n345), .A3(new_n259), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n343), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n343), .A2(new_n346), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n290), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT33), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n288), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n344), .A2(new_n346), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n329), .A2(new_n342), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n307), .A2(new_n310), .ZN(new_n355));
  AND3_X1   g154(.A1(new_n296), .A2(new_n297), .A3(new_n298), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n354), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n353), .A2(new_n358), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n359), .A2(new_n289), .A3(new_n348), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(KEYINPUT34), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT34), .ZN(new_n362));
  NAND4_X1  g161(.A1(new_n359), .A2(new_n362), .A3(new_n289), .A4(new_n348), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n352), .A2(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n289), .B1(new_n359), .B2(new_n348), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n287), .B1(new_n366), .B2(KEYINPUT33), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n367), .A2(new_n361), .A3(new_n363), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n365), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n350), .A2(KEYINPUT32), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n365), .A2(new_n368), .A3(KEYINPUT32), .A4(new_n350), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  XNOR2_X1  g172(.A(KEYINPUT31), .B(G50gat), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT22), .ZN(new_n375));
  INV_X1    g174(.A(G211gat), .ZN(new_n376));
  INV_X1    g175(.A(G218gat), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n375), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  OR2_X1    g177(.A1(KEYINPUT69), .A2(G197gat), .ZN(new_n379));
  NAND2_X1  g178(.A1(KEYINPUT69), .A2(G197gat), .ZN(new_n380));
  AND3_X1   g179(.A1(new_n379), .A2(G204gat), .A3(new_n380), .ZN(new_n381));
  AOI21_X1  g180(.A(G204gat), .B1(new_n379), .B2(new_n380), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n378), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  XOR2_X1   g182(.A(G211gat), .B(G218gat), .Z(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT70), .ZN(new_n386));
  INV_X1    g185(.A(new_n384), .ZN(new_n387));
  OAI211_X1 g186(.A(new_n387), .B(new_n378), .C1(new_n381), .C2(new_n382), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n385), .A2(new_n386), .A3(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n383), .A2(KEYINPUT70), .A3(new_n384), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  AOI21_X1  g191(.A(KEYINPUT29), .B1(new_n226), .B2(new_n251), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT29), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n389), .A2(new_n395), .A3(new_n390), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n226), .B1(new_n396), .B2(new_n251), .ZN(new_n397));
  OAI211_X1 g196(.A(G228gat), .B(G233gat), .C1(new_n394), .C2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT80), .ZN(new_n399));
  AOI21_X1  g198(.A(KEYINPUT29), .B1(new_n385), .B2(new_n388), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n268), .B1(new_n400), .B2(KEYINPUT3), .ZN(new_n401));
  NAND2_X1  g200(.A1(G228gat), .A2(G233gat), .ZN(new_n402));
  OAI211_X1 g201(.A(new_n401), .B(new_n402), .C1(new_n392), .C2(new_n393), .ZN(new_n403));
  AND3_X1   g202(.A1(new_n398), .A2(new_n399), .A3(new_n403), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n399), .B1(new_n398), .B2(new_n403), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n374), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n398), .A2(new_n403), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(KEYINPUT80), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n398), .A2(new_n399), .A3(new_n403), .ZN(new_n409));
  INV_X1    g208(.A(new_n374), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n408), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  XNOR2_X1  g210(.A(G78gat), .B(G106gat), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n412), .B(G22gat), .ZN(new_n413));
  AND3_X1   g212(.A1(new_n406), .A2(new_n411), .A3(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n413), .B1(new_n406), .B2(new_n411), .ZN(new_n415));
  NOR3_X1   g214(.A1(new_n373), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT35), .ZN(new_n417));
  NAND2_X1  g216(.A1(G226gat), .A2(G233gat), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n418), .B1(new_n343), .B2(KEYINPUT29), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(KEYINPUT71), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT72), .ZN(new_n421));
  AND2_X1   g220(.A1(G169gat), .A2(G176gat), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n422), .B1(new_n293), .B2(new_n313), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n423), .A2(new_n327), .A3(new_n312), .ZN(new_n424));
  AOI22_X1  g223(.A1(new_n424), .A2(new_n336), .B1(new_n330), .B2(new_n334), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n421), .B1(new_n425), .B2(new_n311), .ZN(new_n426));
  INV_X1    g225(.A(new_n418), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n335), .A2(new_n340), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n428), .A2(KEYINPUT72), .A3(new_n357), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n426), .A2(new_n427), .A3(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT73), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND4_X1  g231(.A1(new_n426), .A2(new_n429), .A3(KEYINPUT73), .A4(new_n427), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT71), .ZN(new_n435));
  OAI211_X1 g234(.A(new_n435), .B(new_n418), .C1(new_n343), .C2(KEYINPUT29), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n420), .A2(new_n434), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(new_n391), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n343), .A2(new_n427), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n426), .A2(new_n429), .A3(new_n395), .A4(new_n418), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n391), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n438), .A2(new_n442), .ZN(new_n443));
  XNOR2_X1  g242(.A(G8gat), .B(G36gat), .ZN(new_n444));
  XNOR2_X1  g243(.A(G64gat), .B(G92gat), .ZN(new_n445));
  XOR2_X1   g244(.A(new_n444), .B(new_n445), .Z(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n443), .A2(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n441), .B1(new_n437), .B2(new_n391), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n449), .A2(KEYINPUT30), .A3(new_n446), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n438), .A2(new_n446), .A3(new_n442), .ZN(new_n452));
  XOR2_X1   g251(.A(KEYINPUT74), .B(KEYINPUT30), .Z(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT75), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n452), .A2(KEYINPUT75), .A3(new_n453), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n451), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n416), .A2(new_n417), .A3(new_n282), .A4(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n282), .ZN(new_n460));
  INV_X1    g259(.A(new_n413), .ZN(new_n461));
  NOR3_X1   g260(.A1(new_n404), .A2(new_n405), .A3(new_n374), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n410), .B1(new_n408), .B2(new_n409), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n461), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n406), .A2(new_n411), .A3(new_n413), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n464), .A2(new_n465), .A3(new_n372), .A4(new_n371), .ZN(new_n466));
  OAI21_X1  g265(.A(KEYINPUT35), .B1(new_n460), .B2(new_n466), .ZN(new_n467));
  AND2_X1   g266(.A1(new_n459), .A2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT84), .ZN(new_n469));
  AND3_X1   g268(.A1(new_n280), .A2(new_n452), .A3(new_n281), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT83), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT37), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n446), .B1(new_n449), .B2(new_n472), .ZN(new_n473));
  XOR2_X1   g272(.A(KEYINPUT82), .B(KEYINPUT38), .Z(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n437), .A2(new_n392), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n439), .A2(new_n440), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n472), .B1(new_n477), .B2(new_n391), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n475), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n473), .A2(new_n479), .ZN(new_n480));
  AND3_X1   g279(.A1(new_n470), .A2(new_n471), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n471), .B1(new_n470), .B2(new_n480), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n443), .A2(KEYINPUT37), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n474), .B1(new_n483), .B2(new_n473), .ZN(new_n484));
  NOR3_X1   g283(.A1(new_n481), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n414), .A2(new_n415), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n244), .B1(new_n270), .B2(new_n254), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT81), .ZN(new_n488));
  OR2_X1    g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n487), .A2(new_n488), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT39), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n491), .B1(new_n243), .B2(new_n244), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n489), .A2(new_n490), .A3(new_n492), .ZN(new_n493));
  XNOR2_X1  g292(.A(new_n487), .B(KEYINPUT81), .ZN(new_n494));
  OAI211_X1 g293(.A(new_n493), .B(new_n207), .C1(KEYINPUT39), .C2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT40), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n489), .A2(new_n490), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n208), .B1(new_n498), .B2(new_n491), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n499), .A2(KEYINPUT40), .A3(new_n493), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n497), .A2(new_n500), .A3(new_n274), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n486), .B1(new_n458), .B2(new_n501), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n469), .B1(new_n485), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n464), .A2(new_n465), .ZN(new_n504));
  AND3_X1   g303(.A1(new_n497), .A2(new_n274), .A3(new_n500), .ZN(new_n505));
  INV_X1    g304(.A(new_n457), .ZN(new_n506));
  AOI21_X1  g305(.A(KEYINPUT75), .B1(new_n452), .B2(new_n453), .ZN(new_n507));
  OAI211_X1 g306(.A(new_n448), .B(new_n450), .C1(new_n506), .C2(new_n507), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n504), .B1(new_n505), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n470), .A2(new_n480), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(KEYINPUT83), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n470), .A2(new_n480), .A3(new_n471), .ZN(new_n512));
  INV_X1    g311(.A(new_n484), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n511), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n509), .A2(new_n514), .A3(KEYINPUT84), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n503), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n460), .A2(new_n504), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT36), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n373), .B(new_n518), .ZN(new_n519));
  AND2_X1   g318(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n468), .B1(new_n516), .B2(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(G15gat), .B(G22gat), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT16), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n522), .B1(new_n523), .B2(G1gat), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n524), .B1(G1gat), .B2(new_n522), .ZN(new_n525));
  XOR2_X1   g324(.A(new_n525), .B(G8gat), .Z(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  NOR2_X1   g326(.A1(G29gat), .A2(G36gat), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT14), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n528), .B(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(KEYINPUT86), .B(G29gat), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(G36gat), .ZN(new_n532));
  AND2_X1   g331(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(G50gat), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n534), .A2(G43gat), .ZN(new_n535));
  INV_X1    g334(.A(G43gat), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(G50gat), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT15), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  OAI21_X1  g339(.A(KEYINPUT87), .B1(new_n538), .B2(new_n539), .ZN(new_n541));
  OR3_X1    g340(.A1(new_n538), .A2(KEYINPUT87), .A3(new_n539), .ZN(new_n542));
  NAND4_X1  g341(.A1(new_n533), .A2(new_n540), .A3(new_n541), .A4(new_n542), .ZN(new_n543));
  NOR2_X1   g342(.A1(new_n538), .A2(new_n539), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n528), .B(KEYINPUT14), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n532), .B1(new_n545), .B2(KEYINPUT85), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT85), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n530), .A2(new_n547), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n544), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n543), .A2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT88), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n543), .A2(new_n549), .A3(KEYINPUT88), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n527), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(G229gat), .A2(G233gat), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT17), .ZN(new_n556));
  AND3_X1   g355(.A1(new_n552), .A2(new_n556), .A3(new_n553), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n543), .A2(new_n549), .A3(KEYINPUT17), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n526), .A2(new_n558), .ZN(new_n559));
  OAI211_X1 g358(.A(new_n554), .B(new_n555), .C1(new_n557), .C2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(KEYINPUT89), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT18), .ZN(new_n562));
  INV_X1    g361(.A(new_n559), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n552), .A2(new_n553), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n563), .B1(new_n564), .B2(KEYINPUT17), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT89), .ZN(new_n566));
  NAND4_X1  g365(.A1(new_n565), .A2(new_n566), .A3(new_n554), .A4(new_n555), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n561), .A2(new_n562), .A3(new_n567), .ZN(new_n568));
  NAND4_X1  g367(.A1(new_n565), .A2(KEYINPUT18), .A3(new_n554), .A4(new_n555), .ZN(new_n569));
  XOR2_X1   g368(.A(new_n555), .B(KEYINPUT13), .Z(new_n570));
  INV_X1    g369(.A(new_n554), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n527), .B1(new_n552), .B2(new_n553), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  AND2_X1   g372(.A1(new_n569), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n568), .A2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT90), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(G113gat), .B(G141gat), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n578), .B(G197gat), .ZN(new_n579));
  XOR2_X1   g378(.A(KEYINPUT11), .B(G169gat), .Z(new_n580));
  XNOR2_X1  g379(.A(new_n579), .B(new_n580), .ZN(new_n581));
  XOR2_X1   g380(.A(new_n581), .B(KEYINPUT12), .Z(new_n582));
  NAND3_X1  g381(.A1(new_n575), .A2(new_n577), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n569), .A2(new_n573), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n582), .B1(new_n584), .B2(KEYINPUT90), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n585), .A2(new_n574), .A3(new_n568), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n284), .B1(new_n521), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n517), .A2(new_n519), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n590), .B1(new_n503), .B2(new_n515), .ZN(new_n591));
  OAI211_X1 g390(.A(KEYINPUT91), .B(new_n587), .C1(new_n591), .C2(new_n468), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(G85gat), .A2(G92gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n594), .B(KEYINPUT7), .ZN(new_n595));
  NAND2_X1  g394(.A1(G99gat), .A2(G106gat), .ZN(new_n596));
  INV_X1    g395(.A(G85gat), .ZN(new_n597));
  INV_X1    g396(.A(G92gat), .ZN(new_n598));
  AOI22_X1  g397(.A1(KEYINPUT8), .A2(new_n596), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(G99gat), .B(G106gat), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n595), .A2(new_n601), .A3(new_n599), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n603), .A2(KEYINPUT95), .A3(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT95), .ZN(new_n606));
  NAND4_X1  g405(.A1(new_n595), .A2(new_n606), .A3(new_n601), .A4(new_n599), .ZN(new_n607));
  AND3_X1   g406(.A1(new_n605), .A2(new_n607), .A3(KEYINPUT96), .ZN(new_n608));
  AOI21_X1  g407(.A(KEYINPUT96), .B1(new_n605), .B2(new_n607), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n564), .A2(new_n610), .ZN(new_n611));
  AND2_X1   g410(.A1(G232gat), .A2(G233gat), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n611), .B1(KEYINPUT41), .B2(new_n612), .ZN(new_n613));
  OAI211_X1 g412(.A(new_n558), .B(new_n610), .C1(new_n564), .C2(KEYINPUT17), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  XOR2_X1   g414(.A(G190gat), .B(G218gat), .Z(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n616), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n613), .A2(new_n614), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n612), .A2(KEYINPUT41), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(KEYINPUT94), .ZN(new_n622));
  XOR2_X1   g421(.A(G134gat), .B(G162gat), .Z(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(KEYINPUT97), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n620), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT97), .ZN(new_n627));
  NAND4_X1  g426(.A1(new_n617), .A2(new_n627), .A3(new_n624), .A4(new_n619), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(G57gat), .B(G64gat), .ZN(new_n631));
  AOI21_X1  g430(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  AOI22_X1  g432(.A1(KEYINPUT92), .A2(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n634), .B1(G71gat), .B2(G78gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n633), .B(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT21), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(G231gat), .A2(G233gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(G127gat), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n526), .B1(new_n637), .B2(new_n636), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(G183gat), .B(G211gat), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n644), .B(KEYINPUT93), .ZN(new_n645));
  XNOR2_X1  g444(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n646), .B(new_n217), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n645), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n643), .B(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n630), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(G230gat), .A2(G233gat), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n605), .A2(new_n607), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n653), .A2(new_n636), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT98), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n604), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n656), .A2(new_n603), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n600), .A2(new_n655), .A3(new_n602), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  XOR2_X1   g458(.A(new_n633), .B(new_n635), .Z(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  AOI21_X1  g460(.A(KEYINPUT10), .B1(new_n654), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n660), .A2(KEYINPUT10), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT96), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n653), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n605), .A2(new_n607), .A3(KEYINPUT96), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n663), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n652), .B1(new_n662), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n668), .A2(KEYINPUT99), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n660), .B1(new_n607), .B2(new_n605), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n636), .B1(new_n657), .B2(new_n658), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n652), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  XNOR2_X1  g474(.A(G120gat), .B(G148gat), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(KEYINPUT100), .ZN(new_n677));
  XNOR2_X1  g476(.A(G176gat), .B(G204gat), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n677), .B(new_n678), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n675), .A2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT99), .ZN(new_n681));
  OAI211_X1 g480(.A(new_n681), .B(new_n652), .C1(new_n662), .C2(new_n667), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n669), .A2(new_n680), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(KEYINPUT101), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT101), .ZN(new_n685));
  NAND4_X1  g484(.A1(new_n669), .A2(new_n680), .A3(new_n685), .A4(new_n682), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n679), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n688), .B1(new_n668), .B2(new_n674), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  AOI21_X1  g489(.A(KEYINPUT102), .B1(new_n687), .B2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT102), .ZN(new_n692));
  AOI211_X1 g491(.A(new_n692), .B(new_n689), .C1(new_n684), .C2(new_n686), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n651), .A2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT103), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n651), .A2(KEYINPUT103), .A3(new_n694), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  AOI21_X1  g499(.A(KEYINPUT104), .B1(new_n593), .B2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT104), .ZN(new_n702));
  AOI211_X1 g501(.A(new_n702), .B(new_n699), .C1(new_n589), .C2(new_n592), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n283), .B1(new_n701), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(G1gat), .ZN(new_n705));
  INV_X1    g504(.A(G1gat), .ZN(new_n706));
  OAI211_X1 g505(.A(new_n706), .B(new_n283), .C1(new_n701), .C2(new_n703), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n705), .A2(new_n707), .ZN(G1324gat));
  XOR2_X1   g507(.A(KEYINPUT16), .B(G8gat), .Z(new_n709));
  OAI211_X1 g508(.A(new_n508), .B(new_n709), .C1(new_n701), .C2(new_n703), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT42), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  AND2_X1   g511(.A1(new_n709), .A2(KEYINPUT42), .ZN(new_n713));
  OAI211_X1 g512(.A(new_n508), .B(new_n713), .C1(new_n701), .C2(new_n703), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n508), .B1(new_n701), .B2(new_n703), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(G8gat), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n712), .A2(new_n714), .A3(new_n716), .ZN(G1325gat));
  OR2_X1    g516(.A1(new_n701), .A2(new_n703), .ZN(new_n718));
  INV_X1    g517(.A(new_n519), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(G15gat), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(KEYINPUT105), .ZN(new_n721));
  INV_X1    g520(.A(new_n373), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n722), .B1(new_n701), .B2(new_n703), .ZN(new_n723));
  INV_X1    g522(.A(G15gat), .ZN(new_n724));
  AOI22_X1  g523(.A1(new_n718), .A2(new_n721), .B1(new_n723), .B2(new_n724), .ZN(G1326gat));
  OAI21_X1  g524(.A(new_n504), .B1(new_n701), .B2(new_n703), .ZN(new_n726));
  XNOR2_X1  g525(.A(KEYINPUT43), .B(G22gat), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(new_n727), .ZN(new_n729));
  OAI211_X1 g528(.A(new_n504), .B(new_n729), .C1(new_n701), .C2(new_n703), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n728), .A2(new_n730), .ZN(G1327gat));
  INV_X1    g530(.A(new_n694), .ZN(new_n732));
  NOR3_X1   g531(.A1(new_n732), .A2(new_n649), .A3(new_n629), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n282), .A2(new_n531), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n593), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT45), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NOR3_X1   g536(.A1(new_n485), .A2(new_n502), .A3(new_n469), .ZN(new_n738));
  AOI21_X1  g537(.A(KEYINPUT84), .B1(new_n509), .B2(new_n514), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n520), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(new_n468), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n629), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(KEYINPUT44), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n630), .B1(new_n591), .B2(new_n468), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT44), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NOR3_X1   g545(.A1(new_n732), .A2(new_n588), .A3(new_n649), .ZN(new_n747));
  NAND4_X1  g546(.A1(new_n743), .A2(new_n746), .A3(new_n283), .A4(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(new_n531), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n593), .A2(KEYINPUT45), .A3(new_n733), .A4(new_n734), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n737), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(KEYINPUT106), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT106), .ZN(new_n753));
  NAND4_X1  g552(.A1(new_n737), .A2(new_n749), .A3(new_n753), .A4(new_n750), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n752), .A2(new_n754), .ZN(G1328gat));
  AND2_X1   g554(.A1(new_n593), .A2(new_n733), .ZN(new_n756));
  INV_X1    g555(.A(G36gat), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n756), .A2(new_n757), .A3(new_n508), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(KEYINPUT46), .ZN(new_n759));
  AND2_X1   g558(.A1(new_n743), .A2(new_n746), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(new_n747), .ZN(new_n761));
  OAI21_X1  g560(.A(G36gat), .B1(new_n761), .B2(new_n458), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT46), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n756), .A2(new_n763), .A3(new_n757), .A4(new_n508), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n759), .A2(new_n762), .A3(new_n764), .ZN(G1329gat));
  NAND3_X1  g564(.A1(new_n593), .A2(new_n722), .A3(new_n733), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(new_n536), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n519), .A2(new_n536), .ZN(new_n768));
  INV_X1    g567(.A(new_n768), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n767), .B1(new_n761), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(KEYINPUT47), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT47), .ZN(new_n772));
  OAI211_X1 g571(.A(new_n767), .B(new_n772), .C1(new_n761), .C2(new_n769), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n771), .A2(new_n773), .ZN(G1330gat));
  NAND4_X1  g573(.A1(new_n743), .A2(new_n746), .A3(new_n504), .A4(new_n747), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(G50gat), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n593), .A2(new_n534), .A3(new_n504), .A4(new_n733), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT48), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n778), .B(new_n779), .ZN(G1331gat));
  NAND3_X1  g579(.A1(new_n651), .A2(new_n732), .A3(new_n588), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n521), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(new_n283), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n783), .B(G57gat), .ZN(G1332gat));
  INV_X1    g583(.A(KEYINPUT49), .ZN(new_n785));
  INV_X1    g584(.A(G64gat), .ZN(new_n786));
  OAI211_X1 g585(.A(new_n782), .B(new_n508), .C1(new_n785), .C2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n785), .A2(new_n786), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n787), .B(new_n788), .ZN(G1333gat));
  NAND2_X1  g588(.A1(new_n782), .A2(new_n719), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n373), .A2(G71gat), .ZN(new_n791));
  AOI22_X1  g590(.A1(new_n790), .A2(G71gat), .B1(new_n782), .B2(new_n791), .ZN(new_n792));
  XNOR2_X1  g591(.A(KEYINPUT107), .B(KEYINPUT50), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n792), .B(new_n793), .ZN(G1334gat));
  NAND2_X1  g593(.A1(new_n782), .A2(new_n504), .ZN(new_n795));
  XNOR2_X1  g594(.A(new_n795), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g595(.A1(new_n588), .A2(new_n650), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n797), .A2(new_n694), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n760), .A2(new_n798), .ZN(new_n799));
  OAI21_X1  g598(.A(G85gat), .B1(new_n799), .B2(new_n282), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT51), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n801), .B1(new_n744), .B2(new_n797), .ZN(new_n802));
  INV_X1    g601(.A(new_n802), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n797), .A2(new_n801), .ZN(new_n804));
  INV_X1    g603(.A(new_n804), .ZN(new_n805));
  OAI21_X1  g604(.A(KEYINPUT108), .B1(new_n744), .B2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT108), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n742), .A2(new_n807), .A3(new_n804), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(KEYINPUT109), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT109), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n806), .A2(new_n808), .A3(new_n811), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n803), .B1(new_n810), .B2(new_n812), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n732), .A2(new_n597), .A3(new_n283), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n800), .B1(new_n813), .B2(new_n814), .ZN(G1336gat));
  NAND4_X1  g614(.A1(new_n743), .A2(new_n746), .A3(new_n508), .A4(new_n798), .ZN(new_n816));
  AOI21_X1  g615(.A(KEYINPUT52), .B1(new_n816), .B2(G92gat), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n732), .A2(new_n598), .A3(new_n508), .ZN(new_n818));
  XNOR2_X1  g617(.A(new_n818), .B(KEYINPUT110), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n817), .B1(new_n813), .B2(new_n819), .ZN(new_n820));
  AND2_X1   g619(.A1(new_n816), .A2(G92gat), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n819), .B1(new_n809), .B2(new_n802), .ZN(new_n822));
  OAI21_X1  g621(.A(KEYINPUT52), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n820), .A2(new_n823), .ZN(G1337gat));
  OAI21_X1  g623(.A(G99gat), .B1(new_n799), .B2(new_n519), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n694), .A2(G99gat), .A3(new_n373), .ZN(new_n826));
  XOR2_X1   g625(.A(new_n826), .B(KEYINPUT111), .Z(new_n827));
  OAI21_X1  g626(.A(new_n825), .B1(new_n813), .B2(new_n827), .ZN(G1338gat));
  NAND4_X1  g627(.A1(new_n743), .A2(new_n746), .A3(new_n504), .A4(new_n798), .ZN(new_n829));
  AOI21_X1  g628(.A(KEYINPUT53), .B1(new_n829), .B2(G106gat), .ZN(new_n830));
  OR3_X1    g629(.A1(new_n694), .A2(G106gat), .A3(new_n486), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n830), .B1(new_n813), .B2(new_n831), .ZN(new_n832));
  AND2_X1   g631(.A1(new_n829), .A2(G106gat), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n831), .B1(new_n809), .B2(new_n802), .ZN(new_n834));
  OAI21_X1  g633(.A(KEYINPUT53), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n832), .A2(new_n835), .ZN(G1339gat));
  NAND3_X1  g635(.A1(new_n651), .A2(new_n588), .A3(new_n694), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n555), .B1(new_n565), .B2(new_n554), .ZN(new_n838));
  NOR3_X1   g637(.A1(new_n571), .A2(new_n572), .A3(new_n570), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n581), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(new_n582), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n568), .A2(new_n574), .A3(new_n841), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n626), .A2(new_n628), .A3(new_n840), .A4(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT54), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n662), .A2(new_n667), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n844), .B1(new_n845), .B2(new_n673), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n846), .A2(new_n669), .A3(new_n682), .ZN(new_n847));
  INV_X1    g646(.A(new_n668), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n688), .B1(new_n848), .B2(new_n844), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT55), .ZN(new_n851));
  AND3_X1   g650(.A1(new_n850), .A2(KEYINPUT112), .A3(new_n851), .ZN(new_n852));
  AOI21_X1  g651(.A(KEYINPUT112), .B1(new_n850), .B2(new_n851), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n847), .A2(new_n849), .A3(KEYINPUT55), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n687), .A2(new_n855), .ZN(new_n856));
  NOR3_X1   g655(.A1(new_n843), .A2(new_n854), .A3(new_n856), .ZN(new_n857));
  AND2_X1   g656(.A1(new_n687), .A2(new_n855), .ZN(new_n858));
  OAI211_X1 g657(.A(new_n587), .B(new_n858), .C1(new_n852), .C2(new_n853), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n842), .A2(new_n840), .ZN(new_n860));
  INV_X1    g659(.A(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n861), .B1(new_n691), .B2(new_n693), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n859), .A2(new_n862), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n857), .B1(new_n863), .B2(new_n629), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n837), .B1(new_n864), .B2(new_n649), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n508), .A2(new_n282), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n865), .A2(new_n486), .A3(new_n722), .A4(new_n866), .ZN(new_n867));
  NOR3_X1   g666(.A1(new_n867), .A2(new_n236), .A3(new_n588), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n865), .A2(new_n283), .A3(new_n416), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT113), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n508), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND4_X1  g670(.A1(new_n865), .A2(KEYINPUT113), .A3(new_n283), .A4(new_n416), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n871), .A2(new_n587), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n868), .B1(new_n873), .B2(new_n236), .ZN(G1340gat));
  NOR3_X1   g673(.A1(new_n867), .A2(new_n234), .A3(new_n694), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n871), .A2(new_n732), .A3(new_n872), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n875), .B1(new_n876), .B2(new_n234), .ZN(G1341gat));
  NAND4_X1  g676(.A1(new_n871), .A2(new_n229), .A3(new_n649), .A4(new_n872), .ZN(new_n878));
  OAI21_X1  g677(.A(G127gat), .B1(new_n867), .B2(new_n650), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(G1342gat));
  NOR2_X1   g679(.A1(new_n629), .A2(G134gat), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n871), .A2(new_n872), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(KEYINPUT56), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT56), .ZN(new_n884));
  NAND4_X1  g683(.A1(new_n871), .A2(new_n884), .A3(new_n872), .A4(new_n881), .ZN(new_n885));
  OAI21_X1  g684(.A(G134gat), .B1(new_n867), .B2(new_n629), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n883), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n887), .A2(KEYINPUT114), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT114), .ZN(new_n889));
  NAND4_X1  g688(.A1(new_n883), .A2(new_n889), .A3(new_n885), .A4(new_n886), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n888), .A2(new_n890), .ZN(G1343gat));
  INV_X1    g690(.A(new_n865), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n892), .A2(new_n282), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n719), .A2(new_n486), .A3(new_n508), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(new_n895), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n896), .A2(new_n220), .A3(new_n587), .ZN(new_n897));
  INV_X1    g696(.A(new_n866), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n719), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g698(.A(KEYINPUT57), .B1(new_n865), .B2(new_n504), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n504), .A2(KEYINPUT57), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n850), .A2(new_n851), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n587), .A2(new_n858), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n630), .B1(new_n862), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n650), .B1(new_n904), .B2(new_n857), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n901), .B1(new_n905), .B2(new_n837), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n899), .B1(new_n900), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g706(.A(G141gat), .B1(new_n907), .B2(new_n588), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n897), .A2(new_n908), .ZN(new_n909));
  XOR2_X1   g708(.A(KEYINPUT115), .B(KEYINPUT58), .Z(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(new_n910), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n897), .A2(new_n912), .A3(new_n908), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n911), .A2(new_n913), .ZN(G1344gat));
  OAI21_X1  g713(.A(KEYINPUT59), .B1(new_n895), .B2(new_n694), .ZN(new_n915));
  INV_X1    g714(.A(new_n907), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n694), .A2(KEYINPUT59), .ZN(new_n917));
  AOI22_X1  g716(.A1(new_n915), .A2(new_n221), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n862), .A2(new_n903), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(new_n629), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT116), .ZN(new_n921));
  INV_X1    g720(.A(new_n857), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n920), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  OAI21_X1  g722(.A(KEYINPUT116), .B1(new_n904), .B2(new_n857), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n923), .A2(new_n924), .A3(new_n650), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n697), .A2(new_n588), .A3(new_n698), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g726(.A(KEYINPUT57), .B1(new_n927), .B2(new_n504), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n892), .A2(new_n901), .ZN(new_n929));
  OR2_X1    g728(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  AND3_X1   g729(.A1(new_n930), .A2(new_n732), .A3(new_n899), .ZN(new_n931));
  NAND2_X1  g730(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n918), .B1(new_n931), .B2(new_n932), .ZN(G1345gat));
  NAND3_X1  g732(.A1(new_n896), .A2(new_n217), .A3(new_n649), .ZN(new_n934));
  OAI21_X1  g733(.A(G155gat), .B1(new_n907), .B2(new_n650), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT117), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n934), .A2(KEYINPUT117), .A3(new_n935), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n938), .A2(new_n939), .ZN(G1346gat));
  AOI21_X1  g739(.A(G162gat), .B1(new_n896), .B2(new_n630), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n629), .A2(new_n218), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n941), .B1(new_n916), .B2(new_n942), .ZN(G1347gat));
  NOR2_X1   g742(.A1(new_n892), .A2(new_n283), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n466), .A2(new_n458), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NOR3_X1   g745(.A1(new_n946), .A2(G169gat), .A3(new_n588), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n947), .B(KEYINPUT118), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n458), .A2(new_n283), .ZN(new_n949));
  NAND4_X1  g748(.A1(new_n865), .A2(new_n486), .A3(new_n722), .A4(new_n949), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT119), .ZN(new_n951));
  XNOR2_X1  g750(.A(new_n950), .B(new_n951), .ZN(new_n952));
  OAI21_X1  g751(.A(G169gat), .B1(new_n952), .B2(new_n588), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n948), .A2(new_n953), .ZN(G1348gat));
  NAND3_X1  g753(.A1(new_n944), .A2(new_n732), .A3(new_n945), .ZN(new_n955));
  AND3_X1   g754(.A1(new_n955), .A2(KEYINPUT120), .A3(new_n292), .ZN(new_n956));
  AOI21_X1  g755(.A(KEYINPUT120), .B1(new_n955), .B2(new_n292), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT121), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n732), .A2(G176gat), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n959), .B1(new_n952), .B2(new_n960), .ZN(new_n961));
  XNOR2_X1  g760(.A(new_n950), .B(KEYINPUT119), .ZN(new_n962));
  NAND4_X1  g761(.A1(new_n962), .A2(KEYINPUT121), .A3(G176gat), .A4(new_n732), .ZN(new_n963));
  AND3_X1   g762(.A1(new_n958), .A2(new_n961), .A3(new_n963), .ZN(G1349gat));
  AOI21_X1  g763(.A(new_n305), .B1(new_n962), .B2(new_n649), .ZN(new_n965));
  INV_X1    g764(.A(new_n946), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n301), .A2(G183gat), .ZN(new_n967));
  NOR3_X1   g766(.A1(new_n650), .A2(new_n967), .A3(new_n306), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  INV_X1    g768(.A(new_n969), .ZN(new_n970));
  OAI21_X1  g769(.A(KEYINPUT60), .B1(new_n965), .B2(new_n970), .ZN(new_n971));
  OAI21_X1  g770(.A(G183gat), .B1(new_n952), .B2(new_n650), .ZN(new_n972));
  INV_X1    g771(.A(KEYINPUT60), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n972), .A2(new_n973), .A3(new_n969), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n971), .A2(new_n974), .ZN(G1350gat));
  NAND3_X1  g774(.A1(new_n966), .A2(new_n300), .A3(new_n630), .ZN(new_n976));
  INV_X1    g775(.A(KEYINPUT61), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n962), .A2(new_n630), .ZN(new_n978));
  AOI21_X1  g777(.A(new_n977), .B1(new_n978), .B2(G190gat), .ZN(new_n979));
  AOI211_X1 g778(.A(KEYINPUT61), .B(new_n300), .C1(new_n962), .C2(new_n630), .ZN(new_n980));
  OAI21_X1  g779(.A(new_n976), .B1(new_n979), .B2(new_n980), .ZN(G1351gat));
  AND2_X1   g780(.A1(new_n519), .A2(new_n949), .ZN(new_n982));
  OAI211_X1 g781(.A(new_n587), .B(new_n982), .C1(new_n928), .C2(new_n929), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n983), .A2(G197gat), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n519), .A2(new_n504), .A3(new_n508), .ZN(new_n985));
  XNOR2_X1  g784(.A(new_n985), .B(KEYINPUT122), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n944), .A2(new_n986), .ZN(new_n987));
  OR3_X1    g786(.A1(new_n987), .A2(G197gat), .A3(new_n588), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n984), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n989), .A2(KEYINPUT123), .ZN(new_n990));
  INV_X1    g789(.A(KEYINPUT123), .ZN(new_n991));
  NAND3_X1  g790(.A1(new_n984), .A2(new_n988), .A3(new_n991), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n990), .A2(new_n992), .ZN(G1352gat));
  NAND2_X1  g792(.A1(new_n930), .A2(new_n982), .ZN(new_n994));
  OAI21_X1  g793(.A(G204gat), .B1(new_n994), .B2(new_n694), .ZN(new_n995));
  INV_X1    g794(.A(KEYINPUT124), .ZN(new_n996));
  NOR2_X1   g795(.A1(new_n694), .A2(G204gat), .ZN(new_n997));
  INV_X1    g796(.A(new_n997), .ZN(new_n998));
  OAI21_X1  g797(.A(new_n996), .B1(new_n987), .B2(new_n998), .ZN(new_n999));
  NAND4_X1  g798(.A1(new_n944), .A2(KEYINPUT124), .A3(new_n986), .A4(new_n997), .ZN(new_n1000));
  NAND2_X1  g799(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n1001));
  NAND3_X1  g800(.A1(new_n999), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  INV_X1    g801(.A(KEYINPUT125), .ZN(new_n1003));
  INV_X1    g802(.A(KEYINPUT62), .ZN(new_n1004));
  NAND2_X1  g803(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n1002), .A2(new_n1005), .ZN(new_n1006));
  NAND4_X1  g805(.A1(new_n999), .A2(new_n1003), .A3(new_n1004), .A4(new_n1000), .ZN(new_n1007));
  NAND3_X1  g806(.A1(new_n995), .A2(new_n1006), .A3(new_n1007), .ZN(G1353gat));
  OAI211_X1 g807(.A(new_n649), .B(new_n982), .C1(new_n928), .C2(new_n929), .ZN(new_n1009));
  NAND2_X1  g808(.A1(new_n1009), .A2(G211gat), .ZN(new_n1010));
  NAND2_X1  g809(.A1(new_n1010), .A2(KEYINPUT63), .ZN(new_n1011));
  INV_X1    g810(.A(KEYINPUT63), .ZN(new_n1012));
  NAND3_X1  g811(.A1(new_n1009), .A2(new_n1012), .A3(G211gat), .ZN(new_n1013));
  NAND4_X1  g812(.A1(new_n944), .A2(new_n376), .A3(new_n649), .A4(new_n986), .ZN(new_n1014));
  XNOR2_X1  g813(.A(new_n1014), .B(KEYINPUT126), .ZN(new_n1015));
  NAND3_X1  g814(.A1(new_n1011), .A2(new_n1013), .A3(new_n1015), .ZN(G1354gat));
  NOR3_X1   g815(.A1(new_n994), .A2(new_n377), .A3(new_n629), .ZN(new_n1017));
  NAND3_X1  g816(.A1(new_n944), .A2(new_n630), .A3(new_n986), .ZN(new_n1018));
  NAND2_X1  g817(.A1(new_n1018), .A2(new_n377), .ZN(new_n1019));
  XNOR2_X1  g818(.A(new_n1019), .B(KEYINPUT127), .ZN(new_n1020));
  NOR2_X1   g819(.A1(new_n1017), .A2(new_n1020), .ZN(G1355gat));
endmodule


