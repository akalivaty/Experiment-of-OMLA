//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1 0 0 1 1 0 0 1 1 1 1 0 0 1 1 0 0 1 0 0 0 0 1 1 1 1 0 1 1 0 0 0 1 1 1 1 0 0 1 1 0 1 0 0 0 1 0 1 1 0 0 0 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n714, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n751, new_n752, new_n753, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n761, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n787, new_n788, new_n789,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n839, new_n840, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n873, new_n874,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n896, new_n897, new_n898,
    new_n900, new_n901, new_n902, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n935, new_n936, new_n937, new_n938,
    new_n940, new_n941;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT90), .B(G197gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(KEYINPUT11), .B(G169gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  XOR2_X1   g005(.A(new_n206), .B(KEYINPUT12), .Z(new_n207));
  XNOR2_X1  g006(.A(G15gat), .B(G22gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT16), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n208), .B1(new_n209), .B2(G1gat), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n210), .B1(G1gat), .B2(new_n208), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n211), .A2(G8gat), .ZN(new_n212));
  XNOR2_X1  g011(.A(new_n212), .B(KEYINPUT95), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n211), .A2(G8gat), .ZN(new_n214));
  XNOR2_X1  g013(.A(new_n214), .B(KEYINPUT94), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(new_n216), .ZN(new_n217));
  XOR2_X1   g016(.A(G43gat), .B(G50gat), .Z(new_n218));
  INV_X1    g017(.A(KEYINPUT15), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  XOR2_X1   g019(.A(KEYINPUT92), .B(G36gat), .Z(new_n221));
  INV_X1    g020(.A(G29gat), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NOR2_X1   g022(.A1(G29gat), .A2(G36gat), .ZN(new_n224));
  XNOR2_X1  g023(.A(new_n224), .B(KEYINPUT14), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n220), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n226), .B(KEYINPUT93), .ZN(new_n227));
  AND2_X1   g026(.A1(new_n218), .A2(new_n219), .ZN(new_n228));
  OR4_X1    g027(.A1(new_n220), .A2(new_n228), .A3(new_n223), .A4(new_n225), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n227), .A2(KEYINPUT17), .A3(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n227), .A2(new_n229), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT17), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n217), .A2(new_n230), .A3(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n216), .A2(new_n231), .ZN(new_n235));
  AND2_X1   g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(G229gat), .A2(G233gat), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n236), .A2(KEYINPUT18), .A3(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n216), .B(new_n231), .ZN(new_n239));
  XOR2_X1   g038(.A(new_n237), .B(KEYINPUT13), .Z(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n234), .A2(new_n237), .A3(new_n235), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT18), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n238), .A2(new_n241), .A3(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT91), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n207), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n207), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n245), .A2(KEYINPUT91), .A3(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT30), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT76), .ZN(new_n254));
  AND2_X1   g053(.A1(G211gat), .A2(G218gat), .ZN(new_n255));
  NOR2_X1   g054(.A1(G211gat), .A2(G218gat), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  OR2_X1    g056(.A1(new_n257), .A2(KEYINPUT75), .ZN(new_n258));
  AND2_X1   g057(.A1(KEYINPUT74), .A2(G197gat), .ZN(new_n259));
  NOR2_X1   g058(.A1(KEYINPUT74), .A2(G197gat), .ZN(new_n260));
  OAI21_X1  g059(.A(G204gat), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT74), .ZN(new_n262));
  INV_X1    g061(.A(G197gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(G204gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(KEYINPUT74), .A2(G197gat), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n264), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  AND2_X1   g066(.A1(new_n261), .A2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT22), .ZN(new_n269));
  NAND2_X1  g068(.A1(G211gat), .A2(G218gat), .ZN(new_n270));
  AOI22_X1  g069(.A1(new_n257), .A2(KEYINPUT75), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n258), .B1(new_n268), .B2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(G211gat), .ZN(new_n273));
  INV_X1    g072(.A(G218gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n275), .A2(KEYINPUT75), .A3(new_n270), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n270), .A2(new_n269), .ZN(new_n277));
  NAND4_X1  g076(.A1(new_n276), .A2(new_n261), .A3(new_n267), .A4(new_n277), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n257), .A2(KEYINPUT75), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n254), .B1(new_n272), .B2(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n268), .A2(new_n258), .A3(new_n271), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n278), .A2(new_n279), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n282), .A2(new_n283), .A3(KEYINPUT76), .ZN(new_n284));
  AND2_X1   g083(.A1(new_n281), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(G226gat), .ZN(new_n287));
  INV_X1    g086(.A(G233gat), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n289), .A2(KEYINPUT29), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT23), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n292), .A2(G169gat), .ZN(new_n293));
  INV_X1    g092(.A(G176gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(KEYINPUT66), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT66), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(G176gat), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n293), .A2(new_n295), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(G169gat), .A2(G176gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(KEYINPUT23), .ZN(new_n300));
  INV_X1    g099(.A(G169gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(new_n294), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n298), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT67), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n298), .A2(new_n303), .A3(KEYINPUT67), .ZN(new_n307));
  AOI21_X1  g106(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n308));
  OR2_X1    g107(.A1(new_n308), .A2(KEYINPUT65), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(KEYINPUT65), .ZN(new_n310));
  INV_X1    g109(.A(G183gat), .ZN(new_n311));
  INV_X1    g110(.A(G190gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g112(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n314));
  NAND4_X1  g113(.A1(new_n309), .A2(new_n310), .A3(new_n313), .A4(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n306), .A2(new_n307), .A3(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT25), .ZN(new_n317));
  AND3_X1   g116(.A1(new_n316), .A2(KEYINPUT68), .A3(new_n317), .ZN(new_n318));
  AOI21_X1  g117(.A(KEYINPUT68), .B1(new_n316), .B2(new_n317), .ZN(new_n319));
  INV_X1    g118(.A(new_n308), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n320), .A2(new_n313), .A3(new_n314), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n317), .B1(new_n293), .B2(new_n294), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n321), .A2(new_n303), .A3(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  NOR3_X1   g123(.A1(new_n318), .A2(new_n319), .A3(new_n324), .ZN(new_n325));
  XNOR2_X1  g124(.A(KEYINPUT27), .B(G183gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(new_n312), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT28), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(KEYINPUT69), .ZN(new_n329));
  XOR2_X1   g128(.A(new_n327), .B(new_n329), .Z(new_n330));
  NAND2_X1  g129(.A1(G183gat), .A2(G190gat), .ZN(new_n331));
  OR2_X1    g130(.A1(new_n302), .A2(KEYINPUT26), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n302), .A2(KEYINPUT26), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n332), .A2(new_n333), .A3(new_n299), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n330), .A2(new_n331), .A3(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  OAI21_X1  g135(.A(KEYINPUT77), .B1(new_n325), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n316), .A2(new_n317), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT68), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n316), .A2(KEYINPUT68), .A3(new_n317), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n340), .A2(new_n341), .A3(new_n323), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT77), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n342), .A2(new_n343), .A3(new_n335), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n291), .B1(new_n337), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n342), .A2(new_n335), .ZN(new_n346));
  NOR3_X1   g145(.A1(new_n346), .A2(new_n287), .A3(new_n288), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n286), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n337), .A2(new_n289), .A3(new_n344), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n346), .A2(new_n290), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n349), .A2(new_n285), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n348), .A2(new_n351), .ZN(new_n352));
  XNOR2_X1  g151(.A(G8gat), .B(G36gat), .ZN(new_n353));
  XNOR2_X1  g152(.A(G64gat), .B(G92gat), .ZN(new_n354));
  XOR2_X1   g153(.A(new_n353), .B(new_n354), .Z(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n253), .B1(new_n352), .B2(new_n356), .ZN(new_n357));
  NAND4_X1  g156(.A1(new_n348), .A2(new_n351), .A3(KEYINPUT30), .A4(new_n355), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n344), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n343), .B1(new_n342), .B2(new_n335), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n290), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n347), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n285), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  AND3_X1   g163(.A1(new_n349), .A2(new_n285), .A3(new_n350), .ZN(new_n365));
  OAI21_X1  g164(.A(KEYINPUT78), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT78), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n348), .A2(new_n367), .A3(new_n351), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n355), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  OAI21_X1  g168(.A(KEYINPUT85), .B1(new_n359), .B2(new_n369), .ZN(new_n370));
  AND3_X1   g169(.A1(new_n348), .A2(new_n367), .A3(new_n351), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n367), .B1(new_n348), .B2(new_n351), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n356), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT85), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n373), .A2(new_n374), .A3(new_n357), .A4(new_n358), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n370), .A2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(G120gat), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n377), .A2(G113gat), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT70), .ZN(new_n379));
  INV_X1    g178(.A(G113gat), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n380), .A2(G120gat), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n378), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  OAI21_X1  g181(.A(KEYINPUT70), .B1(new_n380), .B2(G120gat), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  XOR2_X1   g183(.A(G127gat), .B(G134gat), .Z(new_n385));
  NOR2_X1   g184(.A1(new_n385), .A2(KEYINPUT1), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n381), .A2(new_n378), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n385), .B1(new_n388), .B2(KEYINPUT1), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(KEYINPUT71), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT71), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n390), .A2(new_n393), .ZN(new_n394));
  OAI211_X1 g193(.A(new_n392), .B(new_n394), .C1(new_n325), .C2(new_n336), .ZN(new_n395));
  NAND4_X1  g194(.A1(new_n342), .A2(new_n393), .A3(new_n390), .A4(new_n335), .ZN(new_n396));
  NAND2_X1  g195(.A1(G227gat), .A2(G233gat), .ZN(new_n397));
  XOR2_X1   g196(.A(new_n397), .B(KEYINPUT64), .Z(new_n398));
  NAND3_X1  g197(.A1(new_n395), .A2(new_n396), .A3(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT32), .ZN(new_n400));
  XNOR2_X1  g199(.A(G15gat), .B(G43gat), .ZN(new_n401));
  XNOR2_X1  g200(.A(G71gat), .B(G99gat), .ZN(new_n402));
  XNOR2_X1  g201(.A(new_n401), .B(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n400), .B1(new_n404), .B2(KEYINPUT33), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n399), .A2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT72), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n400), .A2(KEYINPUT33), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n399), .A2(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n407), .B1(new_n409), .B2(new_n404), .ZN(new_n410));
  AOI211_X1 g209(.A(KEYINPUT72), .B(new_n403), .C1(new_n399), .C2(new_n408), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n406), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  OR2_X1    g211(.A1(new_n398), .A2(KEYINPUT34), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n413), .B1(new_n395), .B2(new_n396), .ZN(new_n414));
  INV_X1    g213(.A(new_n395), .ZN(new_n415));
  INV_X1    g214(.A(new_n396), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n397), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n414), .B1(new_n417), .B2(KEYINPUT34), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n412), .A2(new_n419), .ZN(new_n420));
  OAI211_X1 g219(.A(new_n418), .B(new_n406), .C1(new_n410), .C2(new_n411), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT29), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n282), .A2(new_n283), .A3(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT83), .ZN(new_n425));
  AOI21_X1  g224(.A(KEYINPUT3), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n426), .B1(new_n425), .B2(new_n424), .ZN(new_n427));
  NAND2_X1  g226(.A1(G155gat), .A2(G162gat), .ZN(new_n428));
  INV_X1    g227(.A(G155gat), .ZN(new_n429));
  INV_X1    g228(.A(G162gat), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n428), .B1(new_n431), .B2(KEYINPUT2), .ZN(new_n432));
  INV_X1    g231(.A(G141gat), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n433), .A2(KEYINPUT79), .A3(G148gat), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n434), .B1(new_n433), .B2(G148gat), .ZN(new_n435));
  INV_X1    g234(.A(G148gat), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n436), .A2(G141gat), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n437), .A2(KEYINPUT79), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n432), .B1(new_n435), .B2(new_n438), .ZN(new_n439));
  XNOR2_X1  g238(.A(G141gat), .B(G148gat), .ZN(new_n440));
  OAI211_X1 g239(.A(new_n428), .B(new_n431), .C1(new_n440), .C2(KEYINPUT2), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n427), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(G228gat), .A2(G233gat), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n423), .B1(new_n442), .B2(KEYINPUT3), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n444), .B1(new_n285), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n443), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT82), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT3), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n424), .A2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT80), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n442), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n439), .A2(KEYINPUT80), .A3(new_n441), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n450), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n281), .A2(new_n284), .A3(new_n445), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  XOR2_X1   g256(.A(new_n444), .B(KEYINPUT81), .Z(new_n458));
  AOI21_X1  g257(.A(new_n448), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(new_n458), .ZN(new_n460));
  AOI211_X1 g259(.A(KEYINPUT82), .B(new_n460), .C1(new_n455), .C2(new_n456), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n447), .B1(new_n459), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(G22gat), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT84), .ZN(new_n464));
  INV_X1    g263(.A(G22gat), .ZN(new_n465));
  OAI211_X1 g264(.A(new_n447), .B(new_n465), .C1(new_n459), .C2(new_n461), .ZN(new_n466));
  XNOR2_X1  g265(.A(G78gat), .B(G106gat), .ZN(new_n467));
  XNOR2_X1  g266(.A(KEYINPUT31), .B(G50gat), .ZN(new_n468));
  XOR2_X1   g267(.A(new_n467), .B(new_n468), .Z(new_n469));
  NAND4_X1  g268(.A1(new_n463), .A2(new_n464), .A3(new_n466), .A4(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n463), .A2(new_n464), .A3(new_n466), .ZN(new_n471));
  INV_X1    g270(.A(new_n469), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n464), .B1(new_n463), .B2(new_n466), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n470), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n422), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n391), .B1(KEYINPUT3), .B2(new_n442), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n477), .B1(KEYINPUT3), .B2(new_n442), .ZN(new_n478));
  NAND2_X1  g277(.A1(G225gat), .A2(G233gat), .ZN(new_n479));
  INV_X1    g278(.A(new_n454), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n480), .A2(KEYINPUT4), .A3(new_n391), .ZN(new_n481));
  OR2_X1    g280(.A1(new_n390), .A2(new_n442), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT4), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n478), .A2(new_n479), .A3(new_n481), .A4(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT5), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n390), .B(new_n442), .ZN(new_n487));
  INV_X1    g286(.A(new_n479), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n486), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n485), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n480), .A2(new_n483), .A3(new_n391), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n482), .A2(KEYINPUT4), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n493), .A2(new_n486), .A3(new_n479), .A4(new_n478), .ZN(new_n494));
  XNOR2_X1  g293(.A(G1gat), .B(G29gat), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n495), .B(KEYINPUT0), .ZN(new_n496));
  XNOR2_X1  g295(.A(G57gat), .B(G85gat), .ZN(new_n497));
  XOR2_X1   g296(.A(new_n496), .B(new_n497), .Z(new_n498));
  NAND3_X1  g297(.A1(new_n490), .A2(new_n494), .A3(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT6), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n490), .A2(new_n494), .ZN(new_n502));
  INV_X1    g301(.A(new_n498), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  XNOR2_X1  g303(.A(new_n501), .B(new_n504), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n505), .A2(KEYINPUT35), .ZN(new_n506));
  AND3_X1   g305(.A1(new_n376), .A2(new_n476), .A3(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT73), .ZN(new_n508));
  INV_X1    g307(.A(new_n406), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n409), .A2(new_n404), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(KEYINPUT72), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n409), .A2(new_n407), .A3(new_n404), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n509), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n508), .B1(new_n513), .B2(new_n418), .ZN(new_n514));
  INV_X1    g313(.A(new_n470), .ZN(new_n515));
  AND2_X1   g314(.A1(new_n471), .A2(new_n472), .ZN(new_n516));
  INV_X1    g315(.A(new_n474), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n412), .A2(KEYINPUT73), .A3(new_n419), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n514), .A2(new_n518), .A3(new_n421), .A4(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT89), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NOR3_X1   g321(.A1(new_n359), .A2(new_n505), .A3(new_n369), .ZN(new_n523));
  INV_X1    g322(.A(new_n421), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n475), .A2(new_n524), .ZN(new_n525));
  NAND4_X1  g324(.A1(new_n525), .A2(KEYINPUT89), .A3(new_n514), .A4(new_n519), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n522), .A2(new_n523), .A3(new_n526), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n507), .B1(new_n527), .B2(KEYINPUT35), .ZN(new_n528));
  AND3_X1   g327(.A1(new_n412), .A2(KEYINPUT73), .A3(new_n419), .ZN(new_n529));
  AOI21_X1  g328(.A(KEYINPUT73), .B1(new_n412), .B2(new_n419), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n421), .A2(KEYINPUT36), .ZN(new_n531));
  NOR3_X1   g330(.A1(new_n529), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  AOI21_X1  g331(.A(KEYINPUT36), .B1(new_n420), .B2(new_n421), .ZN(new_n533));
  OAI22_X1  g332(.A1(new_n532), .A2(new_n533), .B1(new_n518), .B2(new_n523), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n479), .B1(new_n493), .B2(new_n478), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT39), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  OAI21_X1  g336(.A(KEYINPUT39), .B1(new_n487), .B2(new_n488), .ZN(new_n538));
  OAI211_X1 g337(.A(new_n537), .B(new_n498), .C1(new_n535), .C2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT40), .ZN(new_n540));
  OR2_X1    g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n539), .A2(new_n540), .ZN(new_n542));
  AND3_X1   g341(.A1(new_n541), .A2(new_n504), .A3(new_n542), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n370), .A2(new_n543), .A3(new_n375), .ZN(new_n544));
  AND2_X1   g343(.A1(new_n544), .A2(new_n518), .ZN(new_n545));
  XNOR2_X1  g344(.A(KEYINPUT86), .B(KEYINPUT38), .ZN(new_n546));
  OAI21_X1  g345(.A(KEYINPUT87), .B1(new_n352), .B2(KEYINPUT37), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT87), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT37), .ZN(new_n549));
  NAND4_X1  g348(.A1(new_n348), .A2(new_n351), .A3(new_n548), .A4(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n547), .A2(new_n550), .A3(new_n356), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n549), .B1(new_n366), .B2(new_n368), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n546), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n553), .A2(KEYINPUT88), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT88), .ZN(new_n555));
  OAI211_X1 g354(.A(new_n555), .B(new_n546), .C1(new_n551), .C2(new_n552), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n362), .A2(new_n363), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n549), .B1(new_n557), .B2(new_n285), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n349), .A2(new_n286), .A3(new_n350), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n546), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND4_X1  g359(.A1(new_n560), .A2(new_n547), .A3(new_n550), .A4(new_n356), .ZN(new_n561));
  INV_X1    g360(.A(new_n505), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n352), .A2(new_n356), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND4_X1  g363(.A1(new_n554), .A2(new_n556), .A3(new_n561), .A4(new_n564), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n534), .B1(new_n545), .B2(new_n565), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n252), .B1(new_n528), .B2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT96), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  OAI211_X1 g368(.A(KEYINPUT96), .B(new_n252), .C1(new_n528), .C2(new_n566), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  XOR2_X1   g370(.A(G57gat), .B(G64gat), .Z(new_n572));
  AOI21_X1  g371(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n572), .B1(KEYINPUT97), .B2(new_n573), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n574), .B1(KEYINPUT97), .B2(new_n573), .ZN(new_n575));
  XNOR2_X1  g374(.A(G71gat), .B(G78gat), .ZN(new_n576));
  OR2_X1    g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n575), .A2(new_n576), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT21), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(G231gat), .A2(G233gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n581), .B(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(G127gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n583), .B(new_n584), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n217), .B1(new_n580), .B2(new_n579), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n583), .B(G127gat), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(new_n586), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n592), .B(new_n429), .ZN(new_n593));
  XNOR2_X1  g392(.A(G183gat), .B(G211gat), .ZN(new_n594));
  XOR2_X1   g393(.A(new_n593), .B(new_n594), .Z(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n591), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n588), .A2(new_n590), .A3(new_n595), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(KEYINPUT100), .A2(KEYINPUT7), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n601), .A2(G85gat), .A3(G92gat), .ZN(new_n602));
  NOR2_X1   g401(.A1(KEYINPUT100), .A2(KEYINPUT7), .ZN(new_n603));
  OR2_X1    g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n602), .A2(new_n603), .ZN(new_n605));
  NAND2_X1  g404(.A1(G99gat), .A2(G106gat), .ZN(new_n606));
  INV_X1    g405(.A(G85gat), .ZN(new_n607));
  INV_X1    g406(.A(G92gat), .ZN(new_n608));
  AOI22_X1  g407(.A1(KEYINPUT8), .A2(new_n606), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n604), .A2(new_n605), .A3(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(KEYINPUT101), .ZN(new_n611));
  XOR2_X1   g410(.A(G99gat), .B(G106gat), .Z(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n611), .A2(new_n613), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n618), .A2(new_n231), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n617), .A2(new_n230), .A3(new_n233), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT41), .ZN(new_n621));
  NAND2_X1  g420(.A1(G232gat), .A2(G233gat), .ZN(new_n622));
  XOR2_X1   g421(.A(new_n622), .B(KEYINPUT98), .Z(new_n623));
  OAI211_X1 g422(.A(new_n619), .B(new_n620), .C1(new_n621), .C2(new_n623), .ZN(new_n624));
  XOR2_X1   g423(.A(G190gat), .B(G218gat), .Z(new_n625));
  XNOR2_X1  g424(.A(new_n625), .B(KEYINPUT102), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  AND2_X1   g426(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n624), .A2(new_n627), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  AOI21_X1  g429(.A(KEYINPUT103), .B1(new_n624), .B2(new_n627), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n623), .A2(new_n621), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(KEYINPUT99), .ZN(new_n633));
  XNOR2_X1  g432(.A(G134gat), .B(G162gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n633), .B(new_n634), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n631), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n630), .A2(new_n636), .ZN(new_n637));
  OAI22_X1  g436(.A1(new_n628), .A2(new_n629), .B1(new_n631), .B2(new_n635), .ZN(new_n638));
  AND2_X1   g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(G230gat), .A2(G233gat), .ZN(new_n640));
  INV_X1    g439(.A(new_n610), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n641), .A2(KEYINPUT104), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n579), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n616), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n643), .A2(new_n644), .A3(new_n614), .ZN(new_n645));
  OAI22_X1  g444(.A1(new_n615), .A2(new_n616), .B1(new_n579), .B2(new_n642), .ZN(new_n646));
  AOI21_X1  g445(.A(KEYINPUT10), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT10), .ZN(new_n648));
  NOR3_X1   g447(.A1(new_n617), .A2(new_n648), .A3(new_n579), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n640), .B1(new_n647), .B2(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(G120gat), .B(G148gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(KEYINPUT105), .ZN(new_n652));
  XNOR2_X1  g451(.A(G176gat), .B(G204gat), .ZN(new_n653));
  XOR2_X1   g452(.A(new_n652), .B(new_n653), .Z(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n645), .A2(new_n646), .ZN(new_n656));
  OAI211_X1 g455(.A(new_n650), .B(new_n655), .C1(new_n640), .C2(new_n656), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n656), .A2(new_n640), .ZN(new_n658));
  INV_X1    g457(.A(new_n647), .ZN(new_n659));
  INV_X1    g458(.A(new_n649), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n640), .B(KEYINPUT106), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n658), .B1(new_n661), .B2(new_n663), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n657), .B1(new_n664), .B2(new_n655), .ZN(new_n665));
  NOR3_X1   g464(.A1(new_n600), .A2(new_n639), .A3(new_n665), .ZN(new_n666));
  AND2_X1   g465(.A1(new_n571), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n667), .A2(new_n505), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(G1gat), .ZN(G1324gat));
  INV_X1    g468(.A(new_n376), .ZN(new_n670));
  XOR2_X1   g469(.A(KEYINPUT16), .B(G8gat), .Z(new_n671));
  NAND3_X1  g470(.A1(new_n667), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT42), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND4_X1  g473(.A1(new_n667), .A2(KEYINPUT42), .A3(new_n670), .A4(new_n671), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n667), .A2(new_n670), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n676), .A2(G8gat), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n674), .A2(new_n675), .A3(new_n677), .ZN(G1325gat));
  INV_X1    g477(.A(G15gat), .ZN(new_n679));
  INV_X1    g478(.A(new_n422), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n667), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n532), .ZN(new_n682));
  INV_X1    g481(.A(new_n533), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  AND2_X1   g484(.A1(new_n667), .A2(new_n685), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n681), .B1(new_n686), .B2(new_n679), .ZN(G1326gat));
  NAND2_X1  g486(.A1(new_n667), .A2(new_n475), .ZN(new_n688));
  XNOR2_X1  g487(.A(KEYINPUT43), .B(G22gat), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n688), .B(new_n689), .ZN(G1327gat));
  OAI21_X1  g489(.A(new_n639), .B1(new_n528), .B2(new_n566), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT44), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  OAI211_X1 g492(.A(KEYINPUT44), .B(new_n639), .C1(new_n528), .C2(new_n566), .ZN(new_n694));
  AND2_X1   g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n599), .A2(new_n665), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(new_n252), .ZN(new_n697));
  XOR2_X1   g496(.A(new_n697), .B(KEYINPUT108), .Z(new_n698));
  NAND3_X1  g497(.A1(new_n695), .A2(new_n505), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(G29gat), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n696), .A2(new_n639), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n701), .B1(new_n569), .B2(new_n570), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT107), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n562), .A2(G29gat), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n702), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n703), .B1(new_n702), .B2(new_n704), .ZN(new_n707));
  NOR3_X1   g506(.A1(new_n706), .A2(new_n707), .A3(KEYINPUT45), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT45), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n702), .A2(new_n704), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(KEYINPUT107), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n709), .B1(new_n711), .B2(new_n705), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n700), .B1(new_n708), .B2(new_n712), .ZN(G1328gat));
  NAND3_X1  g512(.A1(new_n702), .A2(new_n670), .A3(new_n221), .ZN(new_n714));
  OR2_X1    g513(.A1(new_n714), .A2(KEYINPUT46), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(KEYINPUT46), .ZN(new_n716));
  AND3_X1   g515(.A1(new_n695), .A2(new_n670), .A3(new_n698), .ZN(new_n717));
  OAI211_X1 g516(.A(new_n715), .B(new_n716), .C1(new_n221), .C2(new_n717), .ZN(G1329gat));
  NAND4_X1  g517(.A1(new_n693), .A2(new_n685), .A3(new_n694), .A4(new_n698), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(G43gat), .ZN(new_n720));
  INV_X1    g519(.A(new_n701), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n422), .A2(G43gat), .ZN(new_n722));
  AND4_X1   g521(.A1(KEYINPUT109), .A2(new_n571), .A3(new_n721), .A4(new_n722), .ZN(new_n723));
  AOI21_X1  g522(.A(KEYINPUT109), .B1(new_n702), .B2(new_n722), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n720), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT47), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  OAI211_X1 g526(.A(KEYINPUT47), .B(new_n720), .C1(new_n723), .C2(new_n724), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(G1330gat));
  XOR2_X1   g528(.A(KEYINPUT110), .B(KEYINPUT48), .Z(new_n730));
  NAND4_X1  g529(.A1(new_n693), .A2(new_n475), .A3(new_n694), .A4(new_n698), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(G50gat), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n518), .A2(G50gat), .ZN(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  AOI211_X1 g533(.A(new_n701), .B(new_n734), .C1(new_n569), .C2(new_n570), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT111), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n732), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n702), .A2(new_n733), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n738), .A2(KEYINPUT111), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n730), .B1(new_n737), .B2(new_n739), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n738), .A2(new_n732), .A3(KEYINPUT48), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(G1331gat));
  NOR2_X1   g541(.A1(new_n528), .A2(new_n566), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n637), .A2(new_n638), .ZN(new_n744));
  NAND4_X1  g543(.A1(new_n251), .A2(new_n599), .A3(new_n744), .A4(new_n665), .ZN(new_n745));
  XOR2_X1   g544(.A(new_n745), .B(KEYINPUT112), .Z(new_n746));
  NOR2_X1   g545(.A1(new_n743), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(new_n505), .ZN(new_n748));
  XOR2_X1   g547(.A(KEYINPUT113), .B(G57gat), .Z(new_n749));
  XNOR2_X1  g548(.A(new_n748), .B(new_n749), .ZN(G1332gat));
  NAND2_X1  g549(.A1(new_n747), .A2(new_n670), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n751), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n752));
  XOR2_X1   g551(.A(KEYINPUT49), .B(G64gat), .Z(new_n753));
  OAI21_X1  g552(.A(new_n752), .B1(new_n751), .B2(new_n753), .ZN(G1333gat));
  INV_X1    g553(.A(G71gat), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n747), .A2(new_n755), .A3(new_n680), .ZN(new_n756));
  INV_X1    g555(.A(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n747), .A2(new_n685), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n757), .B1(G71gat), .B2(new_n758), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n759), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g559(.A1(new_n747), .A2(new_n475), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g561(.A1(new_n252), .A2(new_n599), .ZN(new_n763));
  OAI211_X1 g562(.A(new_n639), .B(new_n763), .C1(new_n528), .C2(new_n566), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT51), .ZN(new_n765));
  AND2_X1   g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n764), .A2(new_n765), .ZN(new_n767));
  OR2_X1    g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n768), .A2(new_n607), .A3(new_n505), .A4(new_n665), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n763), .A2(new_n665), .ZN(new_n770));
  INV_X1    g569(.A(new_n770), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n693), .A2(new_n694), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(KEYINPUT114), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT114), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n693), .A2(new_n774), .A3(new_n694), .A4(new_n771), .ZN(new_n775));
  AND3_X1   g574(.A1(new_n773), .A2(new_n505), .A3(new_n775), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n769), .B1(new_n776), .B2(new_n607), .ZN(G1336gat));
  OAI21_X1  g576(.A(G92gat), .B1(new_n772), .B2(new_n376), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT52), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n766), .A2(new_n767), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n670), .A2(new_n608), .A3(new_n665), .ZN(new_n781));
  OAI211_X1 g580(.A(new_n778), .B(new_n779), .C1(new_n780), .C2(new_n781), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n780), .A2(new_n781), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n773), .A2(new_n670), .A3(new_n775), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n783), .B1(new_n784), .B2(G92gat), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n782), .B1(new_n785), .B2(new_n779), .ZN(G1337gat));
  INV_X1    g585(.A(G99gat), .ZN(new_n787));
  NAND4_X1  g586(.A1(new_n768), .A2(new_n787), .A3(new_n680), .A4(new_n665), .ZN(new_n788));
  AND3_X1   g587(.A1(new_n773), .A2(new_n685), .A3(new_n775), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n788), .B1(new_n789), .B2(new_n787), .ZN(G1338gat));
  NAND4_X1  g589(.A1(new_n695), .A2(KEYINPUT116), .A3(new_n475), .A4(new_n771), .ZN(new_n791));
  INV_X1    g590(.A(G106gat), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n693), .A2(new_n475), .A3(new_n694), .A4(new_n771), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT116), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n792), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n791), .A2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT115), .ZN(new_n797));
  AND3_X1   g596(.A1(new_n475), .A2(new_n792), .A3(new_n665), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n768), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n798), .B1(new_n766), .B2(new_n767), .ZN(new_n800));
  AOI21_X1  g599(.A(KEYINPUT53), .B1(new_n800), .B2(KEYINPUT115), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n796), .A2(new_n799), .A3(new_n801), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n773), .A2(new_n475), .A3(new_n775), .ZN(new_n803));
  AOI22_X1  g602(.A1(new_n803), .A2(G106gat), .B1(new_n768), .B2(new_n798), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT53), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n802), .B1(new_n804), .B2(new_n805), .ZN(G1339gat));
  OAI22_X1  g605(.A1(new_n236), .A2(new_n237), .B1(new_n239), .B2(new_n240), .ZN(new_n807));
  AOI22_X1  g606(.A1(new_n246), .A2(new_n249), .B1(new_n807), .B2(new_n206), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(new_n665), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT54), .ZN(new_n810));
  OAI211_X1 g609(.A(new_n810), .B(new_n663), .C1(new_n647), .C2(new_n649), .ZN(new_n811));
  AND2_X1   g610(.A1(new_n811), .A2(new_n654), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n659), .A2(new_n662), .A3(new_n660), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n813), .A2(new_n650), .A3(KEYINPUT54), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT55), .ZN(new_n815));
  AND3_X1   g614(.A1(new_n812), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n815), .B1(new_n812), .B2(new_n814), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n657), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  OAI211_X1 g617(.A(new_n744), .B(new_n809), .C1(new_n818), .C2(new_n251), .ZN(new_n819));
  INV_X1    g618(.A(new_n808), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n639), .B1(new_n818), .B2(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n819), .A2(new_n821), .A3(new_n600), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n666), .A2(new_n251), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n670), .A2(new_n562), .ZN(new_n825));
  AND2_X1   g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(new_n476), .ZN(new_n827));
  NOR3_X1   g626(.A1(new_n827), .A2(new_n380), .A3(new_n251), .ZN(new_n828));
  AND2_X1   g627(.A1(new_n522), .A2(new_n526), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n826), .A2(new_n829), .A3(new_n252), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n828), .B1(new_n380), .B2(new_n830), .ZN(G1340gat));
  NAND2_X1  g630(.A1(new_n826), .A2(new_n829), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n665), .A2(new_n377), .ZN(new_n833));
  XNOR2_X1  g632(.A(new_n833), .B(KEYINPUT117), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n826), .A2(new_n476), .A3(new_n665), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n835), .B1(new_n836), .B2(G120gat), .ZN(new_n837));
  XNOR2_X1  g636(.A(new_n837), .B(KEYINPUT118), .ZN(G1341gat));
  OAI21_X1  g637(.A(G127gat), .B1(new_n827), .B2(new_n600), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n599), .A2(new_n584), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n839), .B1(new_n832), .B2(new_n840), .ZN(G1342gat));
  NOR3_X1   g640(.A1(new_n832), .A2(G134gat), .A3(new_n744), .ZN(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  OR2_X1    g642(.A1(new_n843), .A2(KEYINPUT56), .ZN(new_n844));
  OAI21_X1  g643(.A(G134gat), .B1(new_n827), .B2(new_n744), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n843), .A2(KEYINPUT56), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n844), .A2(new_n845), .A3(new_n846), .ZN(G1343gat));
  AOI21_X1  g646(.A(new_n518), .B1(new_n822), .B2(new_n823), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n825), .A2(new_n684), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n433), .B1(new_n850), .B2(new_n251), .ZN(new_n851));
  OR2_X1    g650(.A1(new_n848), .A2(KEYINPUT57), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT119), .ZN(new_n853));
  OR2_X1    g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n848), .A2(KEYINPUT57), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n852), .A2(new_n853), .A3(new_n855), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n854), .A2(new_n849), .A3(new_n856), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n251), .A2(new_n433), .ZN(new_n858));
  INV_X1    g657(.A(new_n858), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n851), .B1(new_n857), .B2(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT58), .ZN(new_n861));
  XNOR2_X1  g660(.A(new_n860), .B(new_n861), .ZN(G1344gat));
  INV_X1    g661(.A(new_n850), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n863), .A2(new_n436), .A3(new_n665), .ZN(new_n864));
  XOR2_X1   g663(.A(new_n864), .B(KEYINPUT120), .Z(new_n865));
  NAND4_X1  g664(.A1(new_n854), .A2(new_n665), .A3(new_n849), .A4(new_n856), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT59), .ZN(new_n867));
  AND3_X1   g666(.A1(new_n866), .A2(new_n867), .A3(G148gat), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n855), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n869), .A2(new_n665), .A3(new_n849), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n867), .B1(new_n870), .B2(G148gat), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n865), .B1(new_n868), .B2(new_n871), .ZN(G1345gat));
  OAI21_X1  g671(.A(G155gat), .B1(new_n857), .B2(new_n600), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n863), .A2(new_n429), .A3(new_n599), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(G1346gat));
  OAI21_X1  g674(.A(new_n430), .B1(new_n850), .B2(new_n744), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n744), .A2(new_n430), .ZN(new_n877));
  INV_X1    g676(.A(new_n877), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n876), .B1(new_n857), .B2(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT121), .ZN(new_n880));
  XNOR2_X1  g679(.A(new_n879), .B(new_n880), .ZN(G1347gat));
  NOR2_X1   g680(.A1(new_n376), .A2(new_n505), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n824), .A2(new_n829), .A3(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(KEYINPUT122), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT122), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n883), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n885), .A2(new_n252), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(new_n301), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n824), .A2(new_n882), .ZN(new_n890));
  INV_X1    g689(.A(new_n476), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n892), .A2(G169gat), .A3(new_n252), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n889), .A2(new_n893), .ZN(new_n894));
  XOR2_X1   g693(.A(new_n894), .B(KEYINPUT123), .Z(G1348gat));
  NAND2_X1  g694(.A1(new_n295), .A2(new_n297), .ZN(new_n896));
  AND3_X1   g695(.A1(new_n892), .A2(new_n896), .A3(new_n665), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n885), .A2(new_n665), .A3(new_n887), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n897), .B1(new_n898), .B2(new_n294), .ZN(G1349gat));
  AOI21_X1  g698(.A(new_n311), .B1(new_n892), .B2(new_n599), .ZN(new_n900));
  AND2_X1   g699(.A1(new_n599), .A2(new_n326), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n900), .B1(new_n884), .B2(new_n901), .ZN(new_n902));
  XOR2_X1   g701(.A(new_n902), .B(KEYINPUT60), .Z(G1350gat));
  NOR2_X1   g702(.A1(new_n744), .A2(G190gat), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n885), .A2(new_n887), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(KEYINPUT124), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT124), .ZN(new_n907));
  NAND4_X1  g706(.A1(new_n885), .A2(new_n907), .A3(new_n887), .A4(new_n904), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  NOR3_X1   g708(.A1(new_n890), .A2(new_n891), .A3(new_n744), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n910), .A2(new_n312), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT61), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NOR3_X1   g712(.A1(new_n910), .A2(KEYINPUT61), .A3(new_n312), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  OAI21_X1  g714(.A(KEYINPUT125), .B1(new_n909), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n906), .A2(new_n908), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT125), .ZN(new_n918));
  OAI211_X1 g717(.A(new_n917), .B(new_n918), .C1(new_n913), .C2(new_n914), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n916), .A2(new_n919), .ZN(G1351gat));
  AND2_X1   g719(.A1(new_n684), .A2(new_n882), .ZN(new_n921));
  AND2_X1   g720(.A1(new_n848), .A2(new_n921), .ZN(new_n922));
  XNOR2_X1  g721(.A(new_n922), .B(KEYINPUT126), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n923), .A2(new_n263), .A3(new_n252), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n869), .A2(new_n921), .ZN(new_n925));
  OAI21_X1  g724(.A(G197gat), .B1(new_n925), .B2(new_n251), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n924), .A2(new_n926), .ZN(G1352gat));
  NAND3_X1  g726(.A1(new_n869), .A2(new_n665), .A3(new_n921), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(G204gat), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n922), .A2(new_n265), .A3(new_n665), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n930), .A2(KEYINPUT62), .ZN(new_n931));
  AND2_X1   g730(.A1(new_n931), .A2(KEYINPUT127), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n931), .A2(KEYINPUT127), .ZN(new_n933));
  OAI221_X1 g732(.A(new_n929), .B1(KEYINPUT62), .B2(new_n930), .C1(new_n932), .C2(new_n933), .ZN(G1353gat));
  NAND3_X1  g733(.A1(new_n923), .A2(new_n273), .A3(new_n599), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n869), .A2(new_n599), .A3(new_n921), .ZN(new_n936));
  AND3_X1   g735(.A1(new_n936), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n937));
  AOI21_X1  g736(.A(KEYINPUT63), .B1(new_n936), .B2(G211gat), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n935), .B1(new_n937), .B2(new_n938), .ZN(G1354gat));
  NAND3_X1  g738(.A1(new_n923), .A2(new_n274), .A3(new_n639), .ZN(new_n940));
  OAI21_X1  g739(.A(G218gat), .B1(new_n925), .B2(new_n744), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(new_n941), .ZN(G1355gat));
endmodule


