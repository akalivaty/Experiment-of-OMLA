//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 1 1 1 1 0 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 0 0 1 0 1 1 0 0 0 0 0 1 1 0 0 0 0 1 1 1 1 0 0 0 0 0 0 1 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:34 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1195,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1253, new_n1254, new_n1255;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XOR2_X1   g0010(.A(new_n210), .B(KEYINPUT0), .Z(new_n211));
  NAND2_X1  g0011(.A1(G107), .A2(G264), .ZN(new_n212));
  INV_X1    g0012(.A(G77), .ZN(new_n213));
  INV_X1    g0013(.A(G244), .ZN(new_n214));
  OAI21_X1  g0014(.A(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT64), .ZN(new_n217));
  AOI211_X1 g0017(.A(new_n215), .B(new_n217), .C1(G50), .C2(G226), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G116), .A2(G270), .ZN(new_n219));
  INV_X1    g0019(.A(G58), .ZN(new_n220));
  INV_X1    g0020(.A(G232), .ZN(new_n221));
  OAI211_X1 g0021(.A(new_n218), .B(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(G68), .ZN(new_n223));
  INV_X1    g0023(.A(G238), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n208), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT1), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  INV_X1    g0028(.A(G20), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g0030(.A(new_n201), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n231), .A2(G50), .ZN(new_n232));
  INV_X1    g0032(.A(new_n232), .ZN(new_n233));
  AOI211_X1 g0033(.A(new_n211), .B(new_n227), .C1(new_n230), .C2(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(new_n221), .ZN(new_n236));
  XOR2_X1   g0036(.A(KEYINPUT2), .B(G226), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G257), .ZN(new_n240));
  XOR2_X1   g0040(.A(KEYINPUT65), .B(G250), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n238), .B(new_n242), .Z(G358));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(G68), .B(G77), .Z(new_n247));
  XNOR2_X1  g0047(.A(G50), .B(G58), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  NAND3_X1  g0050(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n251));
  AND2_X1   g0051(.A1(new_n251), .A2(new_n228), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G1), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n253), .B1(new_n254), .B2(G20), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(G50), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n254), .A2(G13), .A3(G20), .ZN(new_n257));
  NOR2_X1   g0057(.A1(G20), .A2(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G150), .ZN(new_n259));
  XNOR2_X1  g0059(.A(KEYINPUT8), .B(G58), .ZN(new_n260));
  INV_X1    g0060(.A(G33), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n261), .A2(G20), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n259), .B1(new_n260), .B2(new_n263), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n264), .B1(G20), .B2(new_n203), .ZN(new_n265));
  OAI221_X1 g0065(.A(new_n256), .B1(G50), .B2(new_n257), .C1(new_n265), .C2(new_n252), .ZN(new_n266));
  XNOR2_X1  g0066(.A(new_n266), .B(KEYINPUT9), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT3), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(new_n261), .ZN(new_n269));
  NAND2_X1  g0069(.A1(KEYINPUT3), .A2(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NOR2_X1   g0071(.A1(G222), .A2(G1698), .ZN(new_n272));
  INV_X1    g0072(.A(G1698), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n273), .A2(G223), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n271), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n228), .B1(G33), .B2(G41), .ZN(new_n276));
  OAI211_X1 g0076(.A(new_n275), .B(new_n276), .C1(G77), .C2(new_n271), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n254), .B1(G41), .B2(G45), .ZN(new_n278));
  INV_X1    g0078(.A(G274), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G226), .ZN(new_n282));
  INV_X1    g0082(.A(G41), .ZN(new_n283));
  OAI211_X1 g0083(.A(G1), .B(G13), .C1(new_n261), .C2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(new_n278), .ZN(new_n285));
  OAI211_X1 g0085(.A(new_n277), .B(new_n281), .C1(new_n282), .C2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(G200), .ZN(new_n287));
  INV_X1    g0087(.A(G190), .ZN(new_n288));
  OAI211_X1 g0088(.A(new_n267), .B(new_n287), .C1(new_n288), .C2(new_n286), .ZN(new_n289));
  XNOR2_X1  g0089(.A(new_n289), .B(KEYINPUT10), .ZN(new_n290));
  OR2_X1    g0090(.A1(new_n286), .A2(G179), .ZN(new_n291));
  INV_X1    g0091(.A(G169), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n286), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n291), .A2(new_n266), .A3(new_n293), .ZN(new_n294));
  AND2_X1   g0094(.A1(new_n290), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n269), .A2(new_n229), .A3(new_n270), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(KEYINPUT7), .ZN(new_n297));
  XOR2_X1   g0097(.A(KEYINPUT68), .B(KEYINPUT7), .Z(new_n298));
  OAI211_X1 g0098(.A(new_n297), .B(G68), .C1(new_n296), .C2(new_n298), .ZN(new_n299));
  XNOR2_X1  g0099(.A(G58), .B(G68), .ZN(new_n300));
  AOI22_X1  g0100(.A1(new_n300), .A2(G20), .B1(G159), .B2(new_n258), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n299), .A2(KEYINPUT16), .A3(new_n301), .ZN(new_n302));
  AND2_X1   g0102(.A1(new_n302), .A2(new_n253), .ZN(new_n303));
  INV_X1    g0103(.A(new_n301), .ZN(new_n304));
  AND2_X1   g0104(.A1(KEYINPUT3), .A2(G33), .ZN(new_n305));
  NOR2_X1   g0105(.A1(KEYINPUT3), .A2(G33), .ZN(new_n306));
  NOR3_X1   g0106(.A1(new_n305), .A2(new_n306), .A3(G20), .ZN(new_n307));
  OAI21_X1  g0107(.A(KEYINPUT69), .B1(new_n307), .B2(new_n298), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT69), .ZN(new_n309));
  XNOR2_X1  g0109(.A(KEYINPUT68), .B(KEYINPUT7), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n296), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n308), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT7), .ZN(new_n313));
  OAI21_X1  g0113(.A(KEYINPUT70), .B1(new_n296), .B2(new_n313), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n305), .A2(new_n306), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT70), .ZN(new_n316));
  NAND4_X1  g0116(.A1(new_n315), .A2(new_n316), .A3(KEYINPUT7), .A4(new_n229), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n314), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n312), .A2(new_n318), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n304), .B1(new_n319), .B2(G68), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n303), .B1(new_n320), .B2(KEYINPUT16), .ZN(new_n321));
  INV_X1    g0121(.A(new_n260), .ZN(new_n322));
  INV_X1    g0122(.A(new_n257), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(new_n255), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n324), .B1(new_n325), .B2(new_n322), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n321), .A2(new_n327), .ZN(new_n328));
  OR2_X1    g0128(.A1(G223), .A2(G1698), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n282), .A2(G1698), .ZN(new_n330));
  OAI211_X1 g0130(.A(new_n329), .B(new_n330), .C1(new_n305), .C2(new_n306), .ZN(new_n331));
  NAND2_X1  g0131(.A1(G33), .A2(G87), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n284), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n333), .A2(new_n280), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n285), .A2(new_n221), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  AOI21_X1  g0136(.A(G169), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  NOR4_X1   g0137(.A1(new_n333), .A2(new_n335), .A3(G179), .A4(new_n280), .ZN(new_n338));
  OAI21_X1  g0138(.A(KEYINPUT71), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(G179), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n334), .A2(new_n340), .A3(new_n336), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT71), .ZN(new_n342));
  NOR3_X1   g0142(.A1(new_n333), .A2(new_n335), .A3(new_n280), .ZN(new_n343));
  OAI211_X1 g0143(.A(new_n341), .B(new_n342), .C1(G169), .C2(new_n343), .ZN(new_n344));
  AND2_X1   g0144(.A1(new_n339), .A2(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(KEYINPUT18), .B1(new_n328), .B2(new_n345), .ZN(new_n346));
  AOI22_X1  g0146(.A1(new_n308), .A2(new_n311), .B1(new_n314), .B2(new_n317), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n301), .B1(new_n347), .B2(new_n223), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT16), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n326), .B1(new_n350), .B2(new_n303), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n339), .A2(new_n344), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT18), .ZN(new_n353));
  NOR3_X1   g0153(.A1(new_n351), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n346), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n343), .A2(G190), .ZN(new_n356));
  INV_X1    g0156(.A(G200), .ZN(new_n357));
  OR2_X1    g0157(.A1(new_n343), .A2(new_n357), .ZN(new_n358));
  NAND4_X1  g0158(.A1(new_n321), .A2(new_n356), .A3(new_n327), .A4(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT17), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n351), .A2(KEYINPUT17), .A3(new_n356), .A4(new_n358), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n355), .A2(new_n363), .ZN(new_n364));
  AOI22_X1  g0164(.A1(new_n322), .A2(new_n258), .B1(G20), .B2(G77), .ZN(new_n365));
  XNOR2_X1  g0165(.A(KEYINPUT15), .B(G87), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT66), .ZN(new_n367));
  XNOR2_X1  g0167(.A(new_n366), .B(new_n367), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n365), .B1(new_n368), .B2(new_n263), .ZN(new_n369));
  AOI22_X1  g0169(.A1(new_n369), .A2(new_n253), .B1(new_n213), .B2(new_n323), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n255), .A2(G77), .ZN(new_n371));
  AND2_X1   g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n273), .B1(new_n269), .B2(new_n270), .ZN(new_n373));
  AOI22_X1  g0173(.A1(new_n373), .A2(G238), .B1(new_n315), .B2(G107), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n271), .A2(new_n273), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n374), .B1(new_n221), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(new_n276), .ZN(new_n377));
  OAI211_X1 g0177(.A(new_n377), .B(new_n281), .C1(new_n214), .C2(new_n285), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(G200), .ZN(new_n379));
  OAI211_X1 g0179(.A(new_n372), .B(new_n379), .C1(new_n288), .C2(new_n378), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n295), .A2(new_n364), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n258), .A2(G50), .ZN(new_n382));
  OAI221_X1 g0182(.A(new_n382), .B1(new_n229), .B2(G68), .C1(new_n213), .C2(new_n263), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(new_n253), .ZN(new_n384));
  XNOR2_X1  g0184(.A(new_n384), .B(KEYINPUT11), .ZN(new_n385));
  OAI21_X1  g0185(.A(KEYINPUT12), .B1(new_n257), .B2(G68), .ZN(new_n386));
  OR3_X1    g0186(.A1(new_n257), .A2(KEYINPUT12), .A3(G68), .ZN(new_n387));
  AOI22_X1  g0187(.A1(new_n255), .A2(G68), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n385), .A2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n282), .A2(new_n273), .ZN(new_n391));
  OAI211_X1 g0191(.A(new_n271), .B(new_n391), .C1(G232), .C2(new_n273), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT67), .ZN(new_n393));
  NAND2_X1  g0193(.A1(G33), .A2(G97), .ZN(new_n394));
  AND3_X1   g0194(.A1(new_n392), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n393), .B1(new_n392), .B2(new_n394), .ZN(new_n396));
  NOR3_X1   g0196(.A1(new_n395), .A2(new_n396), .A3(new_n284), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n281), .B1(new_n285), .B2(new_n224), .ZN(new_n398));
  OAI21_X1  g0198(.A(KEYINPUT13), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(new_n396), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n392), .A2(new_n393), .A3(new_n394), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n400), .A2(new_n276), .A3(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT13), .ZN(new_n403));
  INV_X1    g0203(.A(new_n398), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n402), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n292), .B1(new_n399), .B2(new_n405), .ZN(new_n406));
  XNOR2_X1  g0206(.A(new_n406), .B(KEYINPUT14), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n399), .A2(G179), .A3(new_n405), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n390), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  OR2_X1    g0210(.A1(new_n378), .A2(G179), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n370), .A2(new_n371), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n378), .A2(new_n292), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n399), .A2(new_n405), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n389), .B1(new_n415), .B2(G200), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n416), .B1(new_n288), .B2(new_n415), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n410), .A2(new_n414), .A3(new_n417), .ZN(new_n418));
  OR2_X1    g0218(.A1(new_n381), .A2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n258), .A2(G77), .ZN(new_n421));
  INV_X1    g0221(.A(G107), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n422), .A2(KEYINPUT6), .A3(G97), .ZN(new_n423));
  INV_X1    g0223(.A(G97), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n424), .A2(new_n422), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n425), .A2(new_n205), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n423), .B1(new_n426), .B2(KEYINPUT6), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(G20), .ZN(new_n428));
  OAI211_X1 g0228(.A(new_n421), .B(new_n428), .C1(new_n347), .C2(new_n422), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(new_n253), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n254), .A2(G33), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n252), .A2(new_n257), .A3(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT72), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n252), .A2(KEYINPUT72), .A3(new_n257), .A4(new_n431), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(G97), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n257), .A2(G97), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n430), .A2(new_n437), .A3(new_n439), .ZN(new_n440));
  AOI22_X1  g0240(.A1(new_n373), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT4), .ZN(new_n442));
  AOI21_X1  g0242(.A(G1698), .B1(new_n269), .B2(new_n270), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n442), .B1(new_n443), .B2(G244), .ZN(new_n444));
  OAI211_X1 g0244(.A(G244), .B(new_n273), .C1(new_n305), .C2(new_n306), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n445), .A2(KEYINPUT4), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n441), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(KEYINPUT73), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n445), .A2(KEYINPUT4), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n271), .A2(new_n442), .A3(G244), .A4(new_n273), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT73), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n451), .A2(new_n452), .A3(new_n441), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n448), .A2(new_n276), .A3(new_n453), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n254), .B(G45), .C1(new_n283), .C2(KEYINPUT5), .ZN(new_n455));
  AND2_X1   g0255(.A1(new_n283), .A2(KEYINPUT5), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n457), .A2(new_n276), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(G257), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n276), .A2(new_n456), .ZN(new_n460));
  INV_X1    g0260(.A(G45), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n461), .A2(G1), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT74), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n462), .B(new_n463), .C1(KEYINPUT5), .C2(new_n283), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n455), .A2(KEYINPUT74), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n460), .A2(new_n464), .A3(new_n465), .A4(G274), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n459), .A2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n454), .A2(new_n288), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n454), .A2(new_n468), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(new_n357), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n440), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  AND3_X1   g0272(.A1(new_n451), .A2(new_n452), .A3(new_n441), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n452), .B1(new_n451), .B2(new_n441), .ZN(new_n474));
  NOR3_X1   g0274(.A1(new_n473), .A2(new_n474), .A3(new_n284), .ZN(new_n475));
  OAI21_X1  g0275(.A(G169), .B1(new_n475), .B2(new_n467), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n454), .A2(G179), .A3(new_n468), .ZN(new_n477));
  INV_X1    g0277(.A(new_n437), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n478), .B1(new_n429), .B2(new_n253), .ZN(new_n479));
  AOI22_X1  g0279(.A1(new_n476), .A2(new_n477), .B1(new_n479), .B2(new_n439), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n472), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n373), .A2(KEYINPUT75), .A3(G264), .ZN(new_n482));
  OAI211_X1 g0282(.A(G264), .B(G1698), .C1(new_n305), .C2(new_n306), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT75), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n482), .A2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(G257), .ZN(new_n487));
  INV_X1    g0287(.A(G303), .ZN(new_n488));
  OAI22_X1  g0288(.A1(new_n375), .A2(new_n487), .B1(new_n488), .B2(new_n271), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n276), .B1(new_n486), .B2(new_n489), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n284), .B(G270), .C1(new_n455), .C2(new_n456), .ZN(new_n491));
  AND2_X1   g0291(.A1(new_n466), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n252), .A2(G116), .A3(new_n257), .A4(new_n431), .ZN(new_n494));
  INV_X1    g0294(.A(G116), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n323), .A2(new_n495), .ZN(new_n496));
  AND2_X1   g0296(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  AOI22_X1  g0297(.A1(new_n251), .A2(new_n228), .B1(G20), .B2(new_n495), .ZN(new_n498));
  NAND2_X1  g0298(.A1(G33), .A2(G283), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n499), .B(new_n229), .C1(G33), .C2(new_n424), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT20), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n498), .A2(KEYINPUT20), .A3(new_n500), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n292), .B1(new_n497), .B2(new_n505), .ZN(new_n506));
  AOI21_X1  g0306(.A(KEYINPUT21), .B1(new_n493), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n497), .A2(new_n505), .ZN(new_n508));
  AND4_X1   g0308(.A1(G179), .A2(new_n490), .A3(new_n508), .A4(new_n492), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n493), .A2(G200), .ZN(new_n511));
  INV_X1    g0311(.A(new_n508), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n511), .B(new_n512), .C1(new_n288), .C2(new_n493), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n493), .A2(KEYINPUT21), .A3(new_n506), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT76), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n493), .A2(new_n506), .A3(KEYINPUT76), .A4(KEYINPUT21), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n510), .A2(new_n513), .A3(new_n516), .A4(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n271), .A2(G257), .A3(G1698), .ZN(new_n520));
  XNOR2_X1  g0320(.A(KEYINPUT77), .B(G294), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(G33), .ZN(new_n522));
  OAI211_X1 g0322(.A(G250), .B(new_n273), .C1(new_n305), .C2(new_n306), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n520), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(new_n276), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n458), .A2(G264), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n525), .A2(new_n466), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(new_n357), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n528), .B1(G190), .B2(new_n527), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n436), .A2(G107), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n257), .A2(G107), .ZN(new_n531));
  XNOR2_X1  g0331(.A(new_n531), .B(KEYINPUT25), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n262), .A2(G116), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n229), .A2(G107), .ZN(new_n534));
  XNOR2_X1  g0334(.A(new_n534), .B(KEYINPUT23), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT22), .ZN(new_n536));
  AOI21_X1  g0336(.A(G20), .B1(new_n269), .B2(new_n270), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n536), .B1(new_n537), .B2(G87), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n229), .B(G87), .C1(new_n305), .C2(new_n306), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n539), .A2(KEYINPUT22), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n533), .B(new_n535), .C1(new_n538), .C2(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT24), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n537), .A2(new_n536), .A3(G87), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n539), .A2(KEYINPUT22), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n546), .A2(KEYINPUT24), .A3(new_n533), .A4(new_n535), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n543), .A2(new_n253), .A3(new_n547), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n529), .A2(new_n530), .A3(new_n532), .A4(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(new_n462), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n284), .A2(new_n550), .A3(G250), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n551), .B1(new_n279), .B2(new_n550), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n214), .A2(G1698), .ZN(new_n553));
  OAI221_X1 g0353(.A(new_n553), .B1(G238), .B2(G1698), .C1(new_n305), .C2(new_n306), .ZN(new_n554));
  NAND2_X1  g0354(.A1(G33), .A2(G116), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n284), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n552), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(G190), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n537), .A2(G68), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT19), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n560), .B1(new_n263), .B2(new_n424), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n229), .B1(new_n394), .B2(new_n560), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n562), .B1(G87), .B2(new_n206), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n559), .A2(new_n561), .A3(new_n563), .ZN(new_n564));
  AOI22_X1  g0364(.A1(new_n564), .A2(new_n253), .B1(new_n368), .B2(new_n323), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n436), .A2(G87), .ZN(new_n566));
  AND3_X1   g0366(.A1(new_n558), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(new_n557), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(G200), .ZN(new_n569));
  INV_X1    g0369(.A(new_n368), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n436), .A2(new_n570), .ZN(new_n571));
  AOI22_X1  g0371(.A1(new_n565), .A2(new_n571), .B1(new_n557), .B2(new_n340), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n568), .A2(new_n292), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n567), .A2(new_n569), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n548), .A2(new_n530), .A3(new_n532), .ZN(new_n575));
  AOI22_X1  g0375(.A1(new_n524), .A2(new_n276), .B1(new_n458), .B2(G264), .ZN(new_n576));
  AND3_X1   g0376(.A1(new_n576), .A2(new_n340), .A3(new_n466), .ZN(new_n577));
  AOI21_X1  g0377(.A(G169), .B1(new_n576), .B2(new_n466), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n575), .A2(new_n579), .ZN(new_n580));
  AND3_X1   g0380(.A1(new_n549), .A2(new_n574), .A3(new_n580), .ZN(new_n581));
  AND4_X1   g0381(.A1(new_n420), .A2(new_n481), .A3(new_n519), .A4(new_n581), .ZN(G372));
  INV_X1    g0382(.A(new_n552), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT78), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n556), .A2(new_n584), .ZN(new_n585));
  AOI211_X1 g0385(.A(KEYINPUT78), .B(new_n284), .C1(new_n554), .C2(new_n555), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n583), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(G200), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n292), .ZN(new_n589));
  AOI22_X1  g0389(.A1(new_n567), .A2(new_n588), .B1(new_n589), .B2(new_n572), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n580), .A2(new_n510), .A3(new_n516), .A4(new_n517), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n481), .A2(new_n549), .A3(new_n590), .A4(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT79), .ZN(new_n593));
  AND3_X1   g0393(.A1(new_n454), .A2(G179), .A3(new_n468), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n292), .B1(new_n454), .B2(new_n468), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n593), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n476), .A2(KEYINPUT79), .A3(new_n477), .ZN(new_n597));
  AND3_X1   g0397(.A1(new_n596), .A2(new_n440), .A3(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT26), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n598), .A2(new_n599), .A3(new_n590), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n480), .A2(new_n574), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(KEYINPUT26), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n589), .A2(new_n572), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n592), .A2(new_n600), .A3(new_n602), .A4(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n420), .A2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(new_n294), .ZN(new_n606));
  AND3_X1   g0406(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n417), .B1(new_n409), .B2(new_n607), .ZN(new_n608));
  OAI22_X1  g0408(.A1(new_n608), .A2(new_n363), .B1(new_n346), .B2(new_n354), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n606), .B1(new_n609), .B2(new_n290), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n605), .A2(new_n610), .ZN(G369));
  NAND3_X1  g0411(.A1(new_n510), .A2(new_n516), .A3(new_n517), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n254), .A2(new_n229), .A3(G13), .ZN(new_n613));
  XNOR2_X1  g0413(.A(new_n613), .B(KEYINPUT80), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT27), .ZN(new_n615));
  OR2_X1    g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n614), .A2(new_n615), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n616), .A2(new_n617), .A3(G213), .ZN(new_n618));
  INV_X1    g0418(.A(G343), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n621), .A2(new_n512), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n612), .A2(new_n622), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n623), .B1(new_n518), .B2(new_n622), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(G330), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n580), .A2(new_n620), .ZN(new_n627));
  INV_X1    g0427(.A(new_n575), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n549), .B1(new_n628), .B2(new_n621), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n627), .B1(new_n629), .B2(new_n580), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n626), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n612), .A2(new_n621), .ZN(new_n632));
  INV_X1    g0432(.A(new_n632), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n627), .B1(new_n630), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n631), .A2(new_n634), .ZN(G399));
  INV_X1    g0435(.A(new_n209), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n636), .A2(G41), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  NOR3_X1   g0438(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n638), .A2(G1), .A3(new_n639), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n640), .B1(new_n232), .B2(new_n638), .ZN(new_n641));
  XNOR2_X1  g0441(.A(new_n641), .B(KEYINPUT28), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT29), .ZN(new_n643));
  AOI211_X1 g0443(.A(new_n438), .B(new_n478), .C1(new_n253), .C2(new_n429), .ZN(new_n644));
  INV_X1    g0444(.A(new_n469), .ZN(new_n645));
  AOI21_X1  g0445(.A(G200), .B1(new_n454), .B2(new_n468), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n644), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n440), .B1(new_n594), .B2(new_n595), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n591), .A2(new_n647), .A3(new_n648), .A4(new_n549), .ZN(new_n649));
  INV_X1    g0449(.A(new_n590), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n603), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n596), .A2(new_n597), .A3(new_n440), .A4(new_n590), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(KEYINPUT26), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n480), .A2(new_n599), .A3(new_n574), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n621), .B1(new_n651), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(KEYINPUT82), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT82), .ZN(new_n658));
  OAI211_X1 g0458(.A(new_n658), .B(new_n621), .C1(new_n651), .C2(new_n655), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n643), .B1(new_n657), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(KEYINPUT83), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT83), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n604), .A2(new_n621), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n662), .B1(new_n663), .B2(new_n643), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n661), .B1(new_n664), .B2(new_n660), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT30), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(KEYINPUT81), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n490), .A2(new_n492), .A3(new_n557), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n594), .A2(new_n576), .A3(new_n667), .A4(new_n669), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n454), .A2(G179), .A3(new_n468), .A4(new_n576), .ZN(new_n671));
  OAI211_X1 g0471(.A(KEYINPUT81), .B(new_n666), .C1(new_n671), .C2(new_n668), .ZN(new_n672));
  AND2_X1   g0472(.A1(new_n493), .A2(new_n527), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n673), .A2(new_n470), .A3(new_n340), .A4(new_n587), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n670), .A2(new_n672), .A3(new_n674), .ZN(new_n675));
  AND2_X1   g0475(.A1(new_n675), .A2(new_n620), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n481), .A2(new_n519), .A3(new_n581), .A4(new_n621), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n676), .B1(new_n677), .B2(KEYINPUT31), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n675), .A2(KEYINPUT31), .A3(new_n620), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(G330), .B1(new_n678), .B2(new_n680), .ZN(new_n681));
  AND2_X1   g0481(.A1(new_n665), .A2(new_n681), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n642), .B1(new_n682), .B2(G1), .ZN(G364));
  NAND2_X1  g0483(.A1(new_n229), .A2(G13), .ZN(new_n684));
  XNOR2_X1  g0484(.A(new_n684), .B(KEYINPUT84), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(G45), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(G1), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n687), .A2(new_n637), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n626), .A2(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n689), .B1(G330), .B2(new_n624), .ZN(new_n690));
  INV_X1    g0490(.A(new_n688), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n233), .A2(new_n461), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n636), .A2(new_n271), .ZN(new_n693));
  OAI211_X1 g0493(.A(new_n692), .B(new_n693), .C1(new_n249), .C2(new_n461), .ZN(new_n694));
  NAND3_X1  g0494(.A1(G355), .A2(new_n271), .A3(new_n209), .ZN(new_n695));
  OAI211_X1 g0495(.A(new_n694), .B(new_n695), .C1(G116), .C2(new_n209), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n228), .B1(G20), .B2(new_n292), .ZN(new_n697));
  NOR3_X1   g0497(.A1(G13), .A2(G20), .A3(G33), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n229), .A2(G179), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n701), .A2(G190), .A3(G200), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n701), .A2(new_n288), .A3(G200), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  AOI22_X1  g0505(.A1(new_n703), .A2(G303), .B1(new_n705), .B2(G283), .ZN(new_n706));
  INV_X1    g0506(.A(G311), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n229), .A2(new_n340), .ZN(new_n708));
  NOR2_X1   g0508(.A1(G190), .A2(G200), .ZN(new_n709));
  AND3_X1   g0509(.A1(new_n708), .A2(KEYINPUT85), .A3(new_n709), .ZN(new_n710));
  AOI21_X1  g0510(.A(KEYINPUT85), .B1(new_n708), .B2(new_n709), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n706), .B1(new_n707), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n708), .A2(G200), .ZN(new_n714));
  XNOR2_X1  g0514(.A(new_n714), .B(KEYINPUT86), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n715), .A2(new_n288), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(G326), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n715), .A2(G190), .ZN(new_n718));
  XNOR2_X1  g0518(.A(KEYINPUT33), .B(G317), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n708), .ZN(new_n721));
  NOR3_X1   g0521(.A1(new_n721), .A2(new_n288), .A3(G200), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(G322), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n701), .A2(new_n709), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n271), .B1(new_n725), .B2(G329), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n717), .A2(new_n720), .A3(new_n723), .A4(new_n726), .ZN(new_n727));
  NOR3_X1   g0527(.A1(new_n288), .A2(G179), .A3(G200), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n728), .A2(new_n229), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  AOI211_X1 g0530(.A(new_n713), .B(new_n727), .C1(new_n521), .C2(new_n730), .ZN(new_n731));
  AOI22_X1  g0531(.A1(G50), .A2(new_n716), .B1(new_n718), .B2(G68), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n732), .B1(new_n213), .B2(new_n712), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n704), .A2(new_n422), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n734), .B1(G87), .B2(new_n703), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n315), .B1(new_n722), .B2(G58), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n730), .A2(G97), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n735), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n725), .A2(G159), .ZN(new_n739));
  XNOR2_X1  g0539(.A(new_n739), .B(KEYINPUT32), .ZN(new_n740));
  NOR3_X1   g0540(.A1(new_n733), .A2(new_n738), .A3(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n697), .B1(new_n731), .B2(new_n741), .ZN(new_n742));
  XOR2_X1   g0542(.A(new_n698), .B(KEYINPUT87), .Z(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  OAI211_X1 g0544(.A(new_n700), .B(new_n742), .C1(new_n624), .C2(new_n744), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n690), .B1(new_n691), .B2(new_n745), .ZN(G396));
  NAND2_X1  g0546(.A1(new_n412), .A2(new_n620), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n380), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(new_n414), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n607), .A2(new_n621), .ZN(new_n750));
  AND2_X1   g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  XOR2_X1   g0552(.A(new_n751), .B(KEYINPUT89), .Z(new_n753));
  MUX2_X1   g0553(.A(new_n752), .B(new_n753), .S(new_n663), .Z(new_n754));
  XNOR2_X1  g0554(.A(new_n754), .B(new_n681), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(new_n691), .ZN(new_n756));
  INV_X1    g0556(.A(G87), .ZN(new_n757));
  OAI221_X1 g0557(.A(new_n737), .B1(new_n757), .B2(new_n704), .C1(new_n422), .C2(new_n702), .ZN(new_n758));
  AOI211_X1 g0558(.A(new_n271), .B(new_n758), .C1(G311), .C2(new_n725), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n722), .A2(G294), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n716), .A2(G303), .ZN(new_n761));
  INV_X1    g0561(.A(new_n712), .ZN(new_n762));
  AOI22_X1  g0562(.A1(new_n718), .A2(G283), .B1(G116), .B2(new_n762), .ZN(new_n763));
  NAND4_X1  g0563(.A1(new_n759), .A2(new_n760), .A3(new_n761), .A4(new_n763), .ZN(new_n764));
  AOI22_X1  g0564(.A1(G137), .A2(new_n716), .B1(new_n718), .B2(G150), .ZN(new_n765));
  INV_X1    g0565(.A(G159), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n765), .B1(new_n766), .B2(new_n712), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n767), .B1(G143), .B2(new_n722), .ZN(new_n768));
  XOR2_X1   g0568(.A(new_n768), .B(KEYINPUT34), .Z(new_n769));
  OAI22_X1  g0569(.A1(new_n202), .A2(new_n702), .B1(new_n704), .B2(new_n223), .ZN(new_n770));
  XNOR2_X1  g0570(.A(new_n770), .B(KEYINPUT88), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n315), .B1(new_n730), .B2(G58), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n769), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  AND2_X1   g0573(.A1(new_n725), .A2(G132), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n764), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(new_n697), .ZN(new_n776));
  NOR2_X1   g0576(.A1(G13), .A2(G33), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n752), .A2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n697), .A2(new_n777), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(new_n213), .ZN(new_n780));
  NAND4_X1  g0580(.A1(new_n776), .A2(new_n778), .A3(new_n688), .A4(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n756), .A2(new_n781), .ZN(G384));
  INV_X1    g0582(.A(KEYINPUT93), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n679), .A2(new_n783), .ZN(new_n784));
  NAND4_X1  g0584(.A1(new_n675), .A2(KEYINPUT93), .A3(KEYINPUT31), .A4(new_n620), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n678), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n419), .A2(new_n786), .ZN(new_n787));
  XOR2_X1   g0587(.A(new_n787), .B(KEYINPUT96), .Z(new_n788));
  INV_X1    g0588(.A(KEYINPUT40), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n415), .A2(G169), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(KEYINPUT14), .ZN(new_n791));
  INV_X1    g0591(.A(KEYINPUT14), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n406), .A2(new_n792), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n791), .A2(new_n408), .A3(new_n793), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n794), .A2(new_n389), .A3(new_n621), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n389), .A2(new_n620), .ZN(new_n796));
  AND2_X1   g0596(.A1(new_n417), .A2(new_n796), .ZN(new_n797));
  OAI211_X1 g0597(.A(new_n751), .B(new_n795), .C1(new_n409), .C2(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n677), .A2(KEYINPUT31), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n675), .A2(new_n620), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n784), .A2(new_n785), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n798), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(KEYINPUT95), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n789), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n328), .A2(new_n345), .ZN(new_n806));
  INV_X1    g0606(.A(new_n618), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n328), .A2(new_n807), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n806), .A2(new_n808), .A3(new_n359), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(KEYINPUT37), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(KEYINPUT92), .ZN(new_n811));
  INV_X1    g0611(.A(KEYINPUT37), .ZN(new_n812));
  NAND4_X1  g0612(.A1(new_n806), .A2(new_n808), .A3(new_n812), .A4(new_n359), .ZN(new_n813));
  INV_X1    g0613(.A(KEYINPUT92), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n809), .A2(new_n814), .A3(KEYINPUT37), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n811), .A2(new_n813), .A3(new_n815), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n816), .B1(new_n364), .B2(new_n808), .ZN(new_n817));
  INV_X1    g0617(.A(KEYINPUT38), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n299), .A2(new_n301), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(new_n349), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n326), .B1(new_n303), .B2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  OAI211_X1 g0623(.A(new_n807), .B(new_n823), .C1(new_n355), .C2(new_n363), .ZN(new_n824));
  INV_X1    g0624(.A(new_n359), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n822), .B1(new_n352), .B2(new_n618), .ZN(new_n826));
  OAI21_X1  g0626(.A(KEYINPUT37), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n827), .A2(new_n813), .A3(KEYINPUT91), .ZN(new_n828));
  INV_X1    g0628(.A(KEYINPUT91), .ZN(new_n829));
  OAI211_X1 g0629(.A(new_n829), .B(KEYINPUT37), .C1(new_n825), .C2(new_n826), .ZN(new_n830));
  NAND4_X1  g0630(.A1(new_n824), .A2(new_n828), .A3(KEYINPUT38), .A4(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n819), .A2(new_n831), .ZN(new_n832));
  OAI21_X1  g0632(.A(KEYINPUT95), .B1(new_n786), .B2(new_n798), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n805), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n824), .A2(new_n830), .A3(new_n828), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n835), .A2(new_n818), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n836), .A2(new_n831), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n837), .A2(new_n803), .ZN(new_n838));
  AOI21_X1  g0638(.A(KEYINPUT94), .B1(new_n838), .B2(new_n789), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT94), .ZN(new_n840));
  AOI211_X1 g0640(.A(new_n840), .B(KEYINPUT40), .C1(new_n837), .C2(new_n803), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n834), .B1(new_n839), .B2(new_n841), .ZN(new_n842));
  XNOR2_X1  g0642(.A(new_n788), .B(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(G330), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n837), .A2(KEYINPUT39), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT39), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n364), .A2(new_n808), .ZN(new_n847));
  AND3_X1   g0647(.A1(new_n809), .A2(new_n814), .A3(KEYINPUT37), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n814), .B1(new_n809), .B2(KEYINPUT37), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n847), .B1(new_n850), .B2(new_n813), .ZN(new_n851));
  OAI211_X1 g0651(.A(new_n846), .B(new_n831), .C1(new_n851), .C2(KEYINPUT38), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n845), .A2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n795), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  AOI22_X1  g0655(.A1(new_n794), .A2(new_n389), .B1(new_n417), .B2(new_n796), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(new_n795), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n604), .A2(new_n621), .A3(new_n751), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n858), .B1(new_n859), .B2(new_n750), .ZN(new_n860));
  AOI22_X1  g0660(.A1(new_n860), .A2(new_n837), .B1(new_n355), .B2(new_n618), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n855), .A2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  OAI211_X1 g0663(.A(new_n420), .B(new_n661), .C1(new_n660), .C2(new_n664), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(new_n610), .ZN(new_n865));
  XNOR2_X1  g0665(.A(new_n863), .B(new_n865), .ZN(new_n866));
  XNOR2_X1  g0666(.A(new_n844), .B(new_n866), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n867), .B1(new_n254), .B2(new_n685), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n495), .B1(new_n427), .B2(KEYINPUT35), .ZN(new_n869));
  OAI211_X1 g0669(.A(new_n869), .B(new_n230), .C1(KEYINPUT35), .C2(new_n427), .ZN(new_n870));
  XNOR2_X1  g0670(.A(new_n870), .B(KEYINPUT36), .ZN(new_n871));
  OAI21_X1  g0671(.A(G77), .B1(new_n220), .B2(new_n223), .ZN(new_n872));
  OAI22_X1  g0672(.A1(new_n232), .A2(new_n872), .B1(G50), .B2(new_n223), .ZN(new_n873));
  INV_X1    g0673(.A(G13), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n873), .A2(G1), .A3(new_n874), .ZN(new_n875));
  XNOR2_X1  g0675(.A(new_n875), .B(KEYINPUT90), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n868), .A2(new_n871), .A3(new_n876), .ZN(G367));
  INV_X1    g0677(.A(KEYINPUT98), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n481), .B1(new_n644), .B2(new_n621), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n598), .A2(new_n620), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n580), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n621), .B1(new_n881), .B2(new_n480), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n630), .A2(new_n633), .A3(new_n481), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(KEYINPUT42), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT97), .ZN(new_n886));
  XNOR2_X1  g0686(.A(new_n885), .B(new_n886), .ZN(new_n887));
  OR2_X1    g0687(.A1(new_n883), .A2(KEYINPUT42), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n565), .A2(new_n566), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n620), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n590), .A2(new_n891), .ZN(new_n892));
  OR2_X1    g0692(.A1(new_n603), .A2(new_n891), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n894), .A2(KEYINPUT43), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n878), .B1(new_n889), .B2(new_n896), .ZN(new_n897));
  NAND4_X1  g0697(.A1(new_n887), .A2(KEYINPUT98), .A3(new_n895), .A4(new_n888), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n894), .A2(KEYINPUT43), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n889), .A2(new_n896), .A3(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n897), .A2(new_n898), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n631), .B1(new_n879), .B2(new_n880), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(KEYINPUT99), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  OR2_X1    g0704(.A1(new_n902), .A2(KEYINPUT99), .ZN(new_n905));
  AND2_X1   g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n904), .A2(new_n905), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  XNOR2_X1  g0709(.A(new_n687), .B(KEYINPUT103), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  XNOR2_X1  g0711(.A(new_n630), .B(new_n632), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n912), .B(KEYINPUT101), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n625), .ZN(new_n914));
  AND2_X1   g0714(.A1(new_n914), .A2(KEYINPUT102), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n914), .A2(KEYINPUT102), .ZN(new_n916));
  INV_X1    g0716(.A(new_n631), .ZN(new_n917));
  NOR3_X1   g0717(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(new_n682), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n879), .A2(new_n880), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(new_n634), .ZN(new_n921));
  XOR2_X1   g0721(.A(new_n921), .B(KEYINPUT45), .Z(new_n922));
  NOR2_X1   g0722(.A1(new_n920), .A2(new_n634), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n923), .B(KEYINPUT44), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n919), .A2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(new_n682), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n637), .B(KEYINPUT41), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n911), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n909), .A2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT104), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n932), .B(new_n933), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n315), .B1(new_n722), .B2(G150), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n705), .A2(G77), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n703), .A2(G58), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n730), .A2(G68), .ZN(new_n938));
  NAND4_X1  g0738(.A1(new_n935), .A2(new_n936), .A3(new_n937), .A4(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n716), .A2(G143), .ZN(new_n940));
  INV_X1    g0740(.A(new_n718), .ZN(new_n941));
  OAI221_X1 g0741(.A(new_n940), .B1(new_n202), .B2(new_n712), .C1(new_n941), .C2(new_n766), .ZN(new_n942));
  AOI211_X1 g0742(.A(new_n939), .B(new_n942), .C1(G137), .C2(new_n725), .ZN(new_n943));
  XNOR2_X1  g0743(.A(KEYINPUT106), .B(G317), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n724), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n703), .A2(KEYINPUT46), .A3(G116), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT46), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(new_n702), .B2(new_n495), .ZN(new_n948));
  INV_X1    g0748(.A(new_n521), .ZN(new_n949));
  OAI211_X1 g0749(.A(new_n946), .B(new_n948), .C1(new_n941), .C2(new_n949), .ZN(new_n950));
  XOR2_X1   g0750(.A(new_n950), .B(KEYINPUT105), .Z(new_n951));
  AOI22_X1  g0751(.A1(new_n730), .A2(G107), .B1(new_n705), .B2(G97), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n762), .A2(G283), .ZN(new_n953));
  NAND4_X1  g0753(.A1(new_n951), .A2(new_n315), .A3(new_n952), .A4(new_n953), .ZN(new_n954));
  AOI211_X1 g0754(.A(new_n945), .B(new_n954), .C1(G303), .C2(new_n722), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n716), .A2(G311), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n943), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  XOR2_X1   g0757(.A(new_n957), .B(KEYINPUT47), .Z(new_n958));
  NAND2_X1  g0758(.A1(new_n958), .A2(new_n697), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n892), .A2(new_n743), .A3(new_n893), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n242), .A2(new_n693), .ZN(new_n961));
  OAI211_X1 g0761(.A(new_n961), .B(new_n699), .C1(new_n209), .C2(new_n368), .ZN(new_n962));
  NAND4_X1  g0762(.A1(new_n959), .A2(new_n688), .A3(new_n960), .A4(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n934), .A2(new_n963), .ZN(G387));
  NAND2_X1  g0764(.A1(new_n918), .A2(new_n911), .ZN(new_n965));
  AOI22_X1  g0765(.A1(new_n718), .A2(new_n322), .B1(G68), .B2(new_n762), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT108), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n967), .B1(G97), .B2(new_n705), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n716), .A2(G159), .ZN(new_n969));
  INV_X1    g0769(.A(new_n722), .ZN(new_n970));
  OAI22_X1  g0770(.A1(new_n970), .A2(new_n202), .B1(new_n213), .B2(new_n702), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n368), .A2(new_n729), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n315), .B1(new_n725), .B2(G150), .ZN(new_n974));
  NAND4_X1  g0774(.A1(new_n968), .A2(new_n969), .A3(new_n973), .A4(new_n974), .ZN(new_n975));
  AOI22_X1  g0775(.A1(new_n716), .A2(G322), .B1(G303), .B2(new_n762), .ZN(new_n976));
  OAI221_X1 g0776(.A(new_n976), .B1(new_n707), .B2(new_n941), .C1(new_n970), .C2(new_n944), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(KEYINPUT48), .ZN(new_n978));
  INV_X1    g0778(.A(G283), .ZN(new_n979));
  OAI221_X1 g0779(.A(new_n978), .B1(new_n979), .B2(new_n729), .C1(new_n949), .C2(new_n702), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n980), .B(KEYINPUT49), .Z(new_n981));
  INV_X1    g0781(.A(G326), .ZN(new_n982));
  OAI221_X1 g0782(.A(new_n315), .B1(new_n724), .B2(new_n982), .C1(new_n495), .C2(new_n704), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n975), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(new_n697), .ZN(new_n985));
  OR2_X1    g0785(.A1(new_n630), .A2(new_n744), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n260), .A2(G50), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT107), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n988), .B(KEYINPUT50), .ZN(new_n989));
  INV_X1    g0789(.A(new_n639), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n461), .B1(new_n223), .B2(new_n213), .ZN(new_n991));
  NOR3_X1   g0791(.A1(new_n989), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n990), .A2(new_n209), .A3(new_n271), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n693), .B1(new_n238), .B2(new_n461), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n992), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n209), .A2(G107), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n699), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n985), .A2(new_n688), .A3(new_n986), .A4(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(new_n919), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n637), .B1(new_n918), .B2(new_n682), .ZN(new_n1000));
  OAI211_X1 g0800(.A(new_n965), .B(new_n998), .C1(new_n999), .C2(new_n1000), .ZN(G393));
  XNOR2_X1  g0801(.A(new_n925), .B(new_n631), .ZN(new_n1002));
  OAI211_X1 g0802(.A(new_n928), .B(new_n637), .C1(new_n999), .C2(new_n1002), .ZN(new_n1003));
  OR2_X1    g0803(.A1(new_n1002), .A2(KEYINPUT109), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1002), .A2(KEYINPUT109), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1004), .A2(new_n911), .A3(new_n1005), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(new_n716), .A2(G317), .B1(G311), .B2(new_n722), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(KEYINPUT52), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1008), .B1(G294), .B2(new_n762), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n718), .A2(G303), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n271), .B1(new_n725), .B2(G322), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n702), .A2(new_n979), .ZN(new_n1012));
  AOI211_X1 g0812(.A(new_n734), .B(new_n1012), .C1(G116), .C2(new_n730), .ZN(new_n1013));
  NAND4_X1  g0813(.A1(new_n1009), .A2(new_n1010), .A3(new_n1011), .A4(new_n1013), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n704), .A2(new_n757), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n716), .A2(G150), .B1(G159), .B2(new_n722), .ZN(new_n1016));
  AND2_X1   g0816(.A1(new_n1016), .A2(KEYINPUT51), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n1016), .A2(KEYINPUT51), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(new_n762), .A2(new_n322), .B1(G77), .B2(new_n730), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1019), .B1(new_n941), .B2(new_n202), .ZN(new_n1020));
  NOR3_X1   g0820(.A1(new_n1017), .A2(new_n1018), .A3(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n703), .A2(G68), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n725), .A2(G143), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n1021), .A2(new_n271), .A3(new_n1022), .A4(new_n1023), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1014), .B1(new_n1015), .B2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1025), .A2(new_n697), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n693), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n699), .B1(new_n424), .B2(new_n209), .C1(new_n246), .C2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n879), .A2(new_n698), .A3(new_n880), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n1026), .A2(new_n688), .A3(new_n1028), .A4(new_n1029), .ZN(new_n1030));
  AND3_X1   g0830(.A1(new_n1006), .A2(KEYINPUT110), .A3(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(KEYINPUT110), .B1(new_n1006), .B2(new_n1030), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1003), .B1(new_n1031), .B2(new_n1032), .ZN(G390));
  NAND3_X1  g0833(.A1(new_n845), .A2(new_n852), .A3(new_n777), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(KEYINPUT54), .B(G143), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1035), .B(KEYINPUT115), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n718), .A2(G137), .B1(new_n762), .B2(new_n1036), .ZN(new_n1037));
  XOR2_X1   g0837(.A(new_n1037), .B(KEYINPUT116), .Z(new_n1038));
  AOI21_X1  g0838(.A(new_n315), .B1(new_n730), .B2(G159), .ZN(new_n1039));
  OAI211_X1 g0839(.A(new_n1038), .B(new_n1039), .C1(new_n202), .C2(new_n704), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n722), .A2(G132), .B1(G125), .B2(new_n725), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n716), .ZN(new_n1042));
  INV_X1    g0842(.A(G128), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1041), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n703), .A2(G150), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT53), .ZN(new_n1046));
  NOR3_X1   g0846(.A1(new_n1040), .A2(new_n1044), .A3(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n271), .B1(new_n703), .B2(G87), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n1048), .B1(new_n213), .B2(new_n729), .C1(new_n712), .C2(new_n424), .ZN(new_n1049));
  INV_X1    g0849(.A(G294), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n704), .A2(new_n223), .B1(new_n724), .B2(new_n1050), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT117), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n1052), .B1(new_n1042), .B2(new_n979), .C1(new_n422), .C2(new_n941), .ZN(new_n1053));
  AOI211_X1 g0853(.A(new_n1049), .B(new_n1053), .C1(G116), .C2(new_n722), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n697), .B1(new_n1047), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n779), .A2(new_n260), .ZN(new_n1056));
  AND4_X1   g0856(.A1(new_n688), .A2(new_n1034), .A3(new_n1055), .A4(new_n1056), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n657), .A2(new_n659), .A3(new_n750), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1058), .A2(new_n749), .A3(new_n857), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n854), .B1(new_n819), .B2(new_n831), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n845), .B(new_n852), .C1(new_n860), .C2(new_n854), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n803), .A2(G330), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1066));
  OAI211_X1 g0866(.A(G330), .B(new_n751), .C1(new_n678), .C2(new_n680), .ZN(new_n1067));
  OR2_X1    g0867(.A1(new_n1067), .A2(new_n858), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1061), .A2(new_n1062), .A3(new_n1068), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1066), .A2(KEYINPUT111), .A3(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT111), .ZN(new_n1071));
  AND4_X1   g0871(.A1(new_n1071), .A2(new_n1061), .A3(new_n1068), .A4(new_n1062), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1070), .A2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1057), .B1(new_n1074), .B2(new_n911), .ZN(new_n1075));
  INV_X1    g0875(.A(KEYINPUT118), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1075), .B(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n801), .A2(new_n802), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n753), .A2(G330), .A3(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(new_n858), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1058), .A2(new_n749), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1080), .A2(new_n1068), .A3(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(KEYINPUT113), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n859), .A2(new_n750), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1067), .A2(KEYINPUT112), .A3(new_n858), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1064), .A2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(KEYINPUT112), .B1(new_n1067), .B2(new_n858), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n1083), .B(new_n1084), .C1(new_n1086), .C2(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1067), .A2(new_n858), .ZN(new_n1090));
  INV_X1    g0890(.A(KEYINPUT112), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1092), .A2(new_n1085), .A3(new_n1064), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1083), .B1(new_n1093), .B2(new_n1084), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1082), .B1(new_n1089), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n787), .A2(G330), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n864), .A2(new_n1096), .A3(new_n610), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1095), .A2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1071), .B1(new_n1063), .B2(new_n1065), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1072), .B1(new_n1100), .B2(new_n1069), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n637), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(KEYINPUT114), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1105));
  OAI211_X1 g0905(.A(KEYINPUT114), .B(new_n637), .C1(new_n1099), .C2(new_n1101), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1104), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1077), .A2(new_n1107), .ZN(G378));
  INV_X1    g0908(.A(KEYINPUT120), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1084), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(KEYINPUT113), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1111), .A2(new_n1088), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1097), .B1(new_n1112), .B2(new_n1082), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1074), .A2(new_n1113), .ZN(new_n1114));
  OAI211_X1 g0914(.A(G330), .B(new_n834), .C1(new_n839), .C2(new_n841), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n266), .A2(new_n807), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(new_n295), .B(new_n1116), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1118));
  XNOR2_X1  g0918(.A(new_n1117), .B(new_n1118), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1115), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1115), .A2(new_n1119), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1121), .A2(new_n863), .A3(new_n1122), .ZN(new_n1123));
  AND2_X1   g0923(.A1(new_n1115), .A2(new_n1119), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n862), .B1(new_n1124), .B2(new_n1120), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n1114), .A2(new_n1098), .B1(new_n1123), .B2(new_n1125), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1109), .B1(new_n1126), .B2(KEYINPUT57), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n638), .B1(new_n1126), .B2(KEYINPUT57), .ZN(new_n1128));
  INV_X1    g0928(.A(KEYINPUT57), .ZN(new_n1129));
  AND2_X1   g0929(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1097), .B1(new_n1074), .B2(new_n1113), .ZN(new_n1131));
  OAI211_X1 g0931(.A(KEYINPUT120), .B(new_n1129), .C1(new_n1130), .C2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1127), .A2(new_n1128), .A3(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n691), .B1(new_n1119), .B2(new_n777), .ZN(new_n1134));
  OAI221_X1 g0934(.A(new_n283), .B1(new_n213), .B2(new_n702), .C1(new_n941), .C2(new_n424), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1135), .B1(new_n570), .B2(new_n762), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n704), .A2(new_n220), .ZN(new_n1137));
  AOI211_X1 g0937(.A(new_n271), .B(new_n1137), .C1(new_n716), .C2(G116), .ZN(new_n1138));
  AND3_X1   g0938(.A1(new_n1136), .A2(new_n938), .A3(new_n1138), .ZN(new_n1139));
  OAI221_X1 g0939(.A(new_n1139), .B1(new_n422), .B2(new_n970), .C1(new_n979), .C2(new_n724), .ZN(new_n1140));
  XOR2_X1   g0940(.A(new_n1140), .B(KEYINPUT58), .Z(new_n1141));
  OAI21_X1  g0941(.A(new_n202), .B1(new_n305), .B2(G41), .ZN(new_n1142));
  AOI22_X1  g0942(.A1(new_n716), .A2(G125), .B1(G137), .B2(new_n762), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n718), .A2(G132), .B1(G128), .B2(new_n722), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n730), .A2(G150), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1036), .A2(new_n703), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n1143), .A2(new_n1144), .A3(new_n1145), .A4(new_n1146), .ZN(new_n1147));
  XOR2_X1   g0947(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n1148));
  AOI21_X1  g0948(.A(G41), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(G33), .B1(new_n725), .B2(G124), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n1149), .B(new_n1150), .C1(new_n766), .C2(new_n704), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1142), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n697), .B1(new_n1141), .B2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n779), .A2(new_n202), .ZN(new_n1155));
  AND3_X1   g0955(.A1(new_n1134), .A2(new_n1154), .A3(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1130), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1156), .B1(new_n1157), .B2(new_n911), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1133), .A2(new_n1158), .ZN(G375));
  NAND2_X1  g0959(.A1(new_n858), .A2(new_n777), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n716), .A2(G132), .B1(G150), .B2(new_n762), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n722), .A2(G137), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n718), .A2(new_n1036), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n271), .B1(new_n724), .B2(new_n1043), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n220), .A2(new_n704), .B1(new_n702), .B2(new_n766), .ZN(new_n1165));
  AOI211_X1 g0965(.A(new_n1164), .B(new_n1165), .C1(G50), .C2(new_n730), .ZN(new_n1166));
  NAND4_X1  g0966(.A1(new_n1161), .A2(new_n1162), .A3(new_n1163), .A4(new_n1166), .ZN(new_n1167));
  OAI221_X1 g0967(.A(new_n936), .B1(new_n488), .B2(new_n724), .C1(new_n941), .C2(new_n495), .ZN(new_n1168));
  AOI211_X1 g0968(.A(new_n271), .B(new_n1168), .C1(G294), .C2(new_n716), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n972), .B1(G283), .B2(new_n722), .ZN(new_n1170));
  XOR2_X1   g0970(.A(new_n1170), .B(KEYINPUT121), .Z(new_n1171));
  OAI211_X1 g0971(.A(new_n1169), .B(new_n1171), .C1(new_n422), .C2(new_n712), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n702), .A2(new_n424), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1167), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1174), .A2(new_n697), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n779), .A2(new_n223), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n1160), .A2(new_n688), .A3(new_n1175), .A4(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1082), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(new_n1111), .B2(new_n1088), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1177), .B1(new_n1179), .B2(new_n910), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n930), .B1(new_n1095), .B2(new_n1098), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1181), .B1(new_n1182), .B2(new_n1113), .ZN(G381));
  INV_X1    g0983(.A(G390), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n934), .A2(new_n963), .A3(new_n1184), .ZN(new_n1185));
  NOR3_X1   g0985(.A1(new_n1185), .A2(G396), .A3(G393), .ZN(new_n1186));
  OR2_X1    g0986(.A1(G381), .A2(G384), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  AND3_X1   g0988(.A1(new_n1107), .A2(KEYINPUT122), .A3(new_n1075), .ZN(new_n1189));
  AOI21_X1  g0989(.A(KEYINPUT122), .B1(new_n1107), .B2(new_n1075), .ZN(new_n1190));
  OR2_X1    g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  AND3_X1   g0991(.A1(new_n1191), .A2(new_n1158), .A3(new_n1133), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1186), .A2(new_n1188), .A3(new_n1192), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(new_n1193), .B(KEYINPUT123), .ZN(G407));
  NAND2_X1  g0994(.A1(new_n1192), .A2(new_n619), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(G407), .A2(G213), .A3(new_n1195), .ZN(G409));
  INV_X1    g0996(.A(KEYINPUT126), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1126), .A2(new_n930), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1158), .A2(new_n1198), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1199), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1133), .A2(G378), .A3(new_n1158), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n619), .A2(G213), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1197), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1203), .ZN(new_n1205));
  AOI211_X1 g1005(.A(KEYINPUT126), .B(new_n1205), .C1(new_n1200), .C2(new_n1201), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1179), .A2(KEYINPUT60), .A3(new_n1097), .ZN(new_n1207));
  AND2_X1   g1007(.A1(new_n1207), .A2(new_n637), .ZN(new_n1208));
  AOI21_X1  g1008(.A(KEYINPUT60), .B1(new_n1179), .B2(new_n1097), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n1209), .A2(new_n1113), .ZN(new_n1210));
  AND3_X1   g1010(.A1(new_n1208), .A2(new_n1210), .A3(KEYINPUT124), .ZN(new_n1211));
  AOI21_X1  g1011(.A(KEYINPUT124), .B1(new_n1208), .B2(new_n1210), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1181), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(G384), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  OAI211_X1 g1015(.A(G384), .B(new_n1181), .C1(new_n1211), .C2(new_n1212), .ZN(new_n1216));
  OR2_X1    g1016(.A1(new_n1203), .A2(KEYINPUT125), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1215), .A2(new_n1216), .A3(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1205), .A2(G2897), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1218), .A2(new_n1220), .ZN(new_n1221));
  NAND4_X1  g1021(.A1(new_n1215), .A2(new_n1216), .A3(new_n1219), .A4(new_n1217), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  NOR3_X1   g1023(.A1(new_n1204), .A2(new_n1206), .A3(new_n1223), .ZN(new_n1224));
  OAI21_X1  g1024(.A(KEYINPUT127), .B1(new_n1224), .B2(KEYINPUT61), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1226), .A2(KEYINPUT126), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1223), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1205), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1229), .A2(new_n1197), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1227), .A2(new_n1228), .A3(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT127), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT61), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1231), .A2(new_n1232), .A3(new_n1233), .ZN(new_n1234));
  AND2_X1   g1034(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1229), .A2(new_n1235), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n1236), .A2(KEYINPUT62), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1235), .B1(new_n1204), .B2(new_n1206), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1237), .B1(new_n1238), .B2(KEYINPUT62), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1225), .A2(new_n1234), .A3(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(G387), .A2(G390), .ZN(new_n1241));
  XNOR2_X1  g1041(.A(G393), .B(G396), .ZN(new_n1242));
  AND3_X1   g1042(.A1(new_n1241), .A2(new_n1185), .A3(new_n1242), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1242), .B1(new_n1241), .B2(new_n1185), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1240), .A2(new_n1246), .ZN(new_n1247));
  OAI21_X1  g1047(.A(KEYINPUT63), .B1(new_n1223), .B2(new_n1229), .ZN(new_n1248));
  AOI21_X1  g1048(.A(KEYINPUT61), .B1(new_n1248), .B2(new_n1236), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT63), .ZN(new_n1250));
  OAI211_X1 g1050(.A(new_n1245), .B(new_n1249), .C1(new_n1250), .C2(new_n1238), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1247), .A2(new_n1251), .ZN(G405));
  INV_X1    g1052(.A(new_n1201), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1253), .B1(G375), .B2(new_n1191), .ZN(new_n1254));
  XNOR2_X1  g1054(.A(new_n1254), .B(new_n1235), .ZN(new_n1255));
  XNOR2_X1  g1055(.A(new_n1245), .B(new_n1255), .ZN(G402));
endmodule


