//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 0 0 1 1 1 0 1 1 0 0 0 1 0 0 1 0 0 0 0 0 0 1 0 0 1 0 0 0 1 0 0 1 0 0 0 1 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:09 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n568, new_n569, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n584, new_n585, new_n586, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n627, new_n628, new_n629, new_n632,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1253, new_n1254, new_n1255, new_n1256;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT64), .Z(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  OAI21_X1  g039(.A(G125), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n462), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  OAI21_X1  g042(.A(G137), .B1(new_n463), .B2(new_n464), .ZN(new_n468));
  NAND2_X1  g043(.A1(G101), .A2(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(G2105), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n467), .A2(new_n470), .ZN(G160));
  OR2_X1    g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(G2105), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G136), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n462), .B1(new_n472), .B2(new_n473), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  OR2_X1    g052(.A1(G100), .A2(G2105), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n478), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n475), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G162));
  INV_X1    g056(.A(KEYINPUT65), .ZN(new_n482));
  OAI21_X1  g057(.A(G2104), .B1(new_n462), .B2(G114), .ZN(new_n483));
  NOR2_X1   g058(.A1(G102), .A2(G2105), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n484), .ZN(new_n486));
  INV_X1    g061(.A(G114), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G2105), .ZN(new_n488));
  NAND4_X1  g063(.A1(new_n486), .A2(new_n488), .A3(KEYINPUT65), .A4(G2104), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n485), .A2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(G138), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n491), .A2(G2105), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n492), .B(KEYINPUT66), .C1(new_n464), .C2(new_n463), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n476), .A2(G126), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT66), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n497), .B1(new_n472), .B2(new_n473), .ZN(new_n498));
  NOR3_X1   g073(.A1(new_n494), .A2(new_n491), .A3(G2105), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n490), .A2(new_n495), .A3(new_n496), .A4(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(G164));
  INV_X1    g077(.A(KEYINPUT68), .ZN(new_n503));
  OR2_X1    g078(.A1(KEYINPUT5), .A2(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(KEYINPUT5), .A2(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  XNOR2_X1  g081(.A(KEYINPUT6), .B(G651), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n506), .A2(new_n507), .A3(G88), .ZN(new_n508));
  AND2_X1   g083(.A1(G75), .A2(G543), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n509), .B1(new_n506), .B2(G62), .ZN(new_n510));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n508), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT67), .ZN(new_n513));
  AND2_X1   g088(.A1(G50), .A2(G543), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n513), .B1(new_n507), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n511), .A2(KEYINPUT6), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT6), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G651), .ZN(new_n518));
  AND4_X1   g093(.A1(new_n513), .A2(new_n516), .A3(new_n518), .A4(new_n514), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n515), .A2(new_n519), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n503), .B1(new_n512), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n507), .A2(new_n514), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(KEYINPUT67), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n507), .A2(new_n513), .A3(new_n514), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  AND2_X1   g100(.A1(KEYINPUT5), .A2(G543), .ZN(new_n526));
  NOR2_X1   g101(.A1(KEYINPUT5), .A2(G543), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(G62), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  OAI21_X1  g105(.A(G651), .B1(new_n530), .B2(new_n509), .ZN(new_n531));
  NAND4_X1  g106(.A1(new_n525), .A2(new_n531), .A3(KEYINPUT68), .A4(new_n508), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n521), .A2(new_n532), .ZN(G166));
  NAND3_X1  g108(.A1(new_n506), .A2(G63), .A3(G651), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT69), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n534), .B(new_n535), .ZN(new_n536));
  NAND3_X1  g111(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n537));
  XNOR2_X1  g112(.A(new_n537), .B(KEYINPUT7), .ZN(new_n538));
  OAI211_X1 g113(.A(new_n516), .B(new_n518), .C1(new_n526), .C2(new_n527), .ZN(new_n539));
  INV_X1    g114(.A(G89), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n507), .A2(G543), .ZN(new_n541));
  INV_X1    g116(.A(G51), .ZN(new_n542));
  OAI221_X1 g117(.A(new_n538), .B1(new_n539), .B2(new_n540), .C1(new_n541), .C2(new_n542), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n536), .A2(new_n543), .ZN(G168));
  AOI22_X1  g119(.A1(new_n506), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n545), .A2(new_n511), .ZN(new_n546));
  INV_X1    g121(.A(G52), .ZN(new_n547));
  INV_X1    g122(.A(G90), .ZN(new_n548));
  OAI22_X1  g123(.A1(new_n541), .A2(new_n547), .B1(new_n539), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n546), .A2(new_n549), .ZN(G171));
  INV_X1    g125(.A(G43), .ZN(new_n551));
  INV_X1    g126(.A(G81), .ZN(new_n552));
  OAI22_X1  g127(.A1(new_n541), .A2(new_n551), .B1(new_n539), .B2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT70), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  OAI221_X1 g130(.A(KEYINPUT70), .B1(new_n539), .B2(new_n552), .C1(new_n541), .C2(new_n551), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT71), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n506), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n559));
  OR2_X1    g134(.A1(new_n559), .A2(new_n511), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n557), .A2(new_n558), .A3(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(new_n561), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n558), .B1(new_n557), .B2(new_n560), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G860), .ZN(new_n565));
  XOR2_X1   g140(.A(new_n565), .B(KEYINPUT72), .Z(G153));
  NAND4_X1  g141(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g142(.A1(G1), .A2(G3), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT8), .ZN(new_n569));
  NAND4_X1  g144(.A1(G319), .A2(G483), .A3(G661), .A4(new_n569), .ZN(G188));
  INV_X1    g145(.A(G53), .ZN(new_n571));
  OAI21_X1  g146(.A(KEYINPUT9), .B1(new_n541), .B2(new_n571), .ZN(new_n572));
  AND3_X1   g147(.A1(new_n516), .A2(new_n518), .A3(G543), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT9), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n573), .A2(new_n574), .A3(G53), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n506), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n577));
  OR2_X1    g152(.A1(new_n577), .A2(new_n511), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n506), .A2(new_n507), .A3(G91), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n576), .A2(new_n578), .A3(new_n579), .ZN(G299));
  INV_X1    g155(.A(G171), .ZN(G301));
  INV_X1    g156(.A(G168), .ZN(G286));
  INV_X1    g157(.A(G166), .ZN(G303));
  OAI21_X1  g158(.A(G651), .B1(new_n506), .B2(G74), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n507), .A2(G49), .A3(G543), .ZN(new_n585));
  INV_X1    g160(.A(G87), .ZN(new_n586));
  OAI211_X1 g161(.A(new_n584), .B(new_n585), .C1(new_n586), .C2(new_n539), .ZN(G288));
  INV_X1    g162(.A(G61), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n588), .B1(new_n504), .B2(new_n505), .ZN(new_n589));
  NAND2_X1  g164(.A1(G73), .A2(G543), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(new_n591));
  OAI21_X1  g166(.A(G651), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n506), .A2(new_n507), .A3(G86), .ZN(new_n593));
  NAND4_X1  g168(.A1(new_n516), .A2(new_n518), .A3(G48), .A4(G543), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(G305));
  NAND2_X1  g170(.A1(G72), .A2(G543), .ZN(new_n596));
  INV_X1    g171(.A(G60), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n528), .B2(new_n597), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n511), .B1(new_n598), .B2(KEYINPUT73), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n599), .B1(KEYINPUT73), .B2(new_n598), .ZN(new_n600));
  INV_X1    g175(.A(G47), .ZN(new_n601));
  INV_X1    g176(.A(G85), .ZN(new_n602));
  OAI22_X1  g177(.A1(new_n541), .A2(new_n601), .B1(new_n539), .B2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT74), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n604), .A2(new_n605), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n600), .B1(new_n607), .B2(new_n608), .ZN(G290));
  INV_X1    g184(.A(G868), .ZN(new_n610));
  NOR2_X1   g185(.A1(G301), .A2(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(G92), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n539), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT10), .ZN(new_n614));
  NAND2_X1  g189(.A1(G79), .A2(G543), .ZN(new_n615));
  INV_X1    g190(.A(G66), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n528), .B2(new_n616), .ZN(new_n617));
  AOI22_X1  g192(.A1(new_n617), .A2(G651), .B1(new_n573), .B2(G54), .ZN(new_n618));
  AND2_X1   g193(.A1(new_n614), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n619), .A2(KEYINPUT75), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n614), .A2(new_n618), .ZN(new_n621));
  INV_X1    g196(.A(KEYINPUT75), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n620), .A2(new_n623), .ZN(new_n624));
  AOI21_X1  g199(.A(new_n611), .B1(new_n624), .B2(new_n610), .ZN(G284));
  XOR2_X1   g200(.A(G284), .B(KEYINPUT76), .Z(G321));
  OR3_X1    g201(.A1(G168), .A2(KEYINPUT77), .A3(new_n610), .ZN(new_n627));
  OAI21_X1  g202(.A(KEYINPUT77), .B1(G168), .B2(new_n610), .ZN(new_n628));
  AND3_X1   g203(.A1(new_n576), .A2(new_n578), .A3(new_n579), .ZN(new_n629));
  OAI211_X1 g204(.A(new_n627), .B(new_n628), .C1(G868), .C2(new_n629), .ZN(G297));
  OAI211_X1 g205(.A(new_n627), .B(new_n628), .C1(G868), .C2(new_n629), .ZN(G280));
  XOR2_X1   g206(.A(KEYINPUT78), .B(G559), .Z(new_n632));
  OAI21_X1  g207(.A(new_n624), .B1(G860), .B2(new_n632), .ZN(G148));
  NAND2_X1  g208(.A1(new_n624), .A2(new_n632), .ZN(new_n634));
  INV_X1    g209(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n635), .A2(G868), .ZN(new_n636));
  INV_X1    g211(.A(new_n564), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n636), .B1(G868), .B2(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n638), .B(KEYINPUT11), .Z(G282));
  INV_X1    g214(.A(new_n638), .ZN(G323));
  NAND2_X1  g215(.A1(new_n474), .A2(G2104), .ZN(new_n641));
  XOR2_X1   g216(.A(new_n641), .B(KEYINPUT12), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT79), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(KEYINPUT13), .Z(new_n644));
  INV_X1    g219(.A(G2100), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n644), .A2(new_n645), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n474), .A2(G135), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n476), .A2(G123), .ZN(new_n649));
  NOR2_X1   g224(.A1(G99), .A2(G2105), .ZN(new_n650));
  OAI21_X1  g225(.A(G2104), .B1(new_n462), .B2(G111), .ZN(new_n651));
  OAI211_X1 g226(.A(new_n648), .B(new_n649), .C1(new_n650), .C2(new_n651), .ZN(new_n652));
  INV_X1    g227(.A(G2096), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n646), .A2(new_n647), .A3(new_n654), .ZN(G156));
  XOR2_X1   g230(.A(KEYINPUT15), .B(G2435), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(G2438), .ZN(new_n657));
  XOR2_X1   g232(.A(G2427), .B(G2430), .Z(new_n658));
  OR2_X1    g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(KEYINPUT81), .B(KEYINPUT14), .Z(new_n660));
  NAND2_X1  g235(.A1(new_n657), .A2(new_n658), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n659), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(KEYINPUT80), .B(KEYINPUT16), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(G2443), .B(G2446), .Z(new_n665));
  XNOR2_X1  g240(.A(G2451), .B(G2454), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n664), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1341), .B(G1348), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(KEYINPUT82), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  OAI21_X1  g247(.A(G14), .B1(new_n668), .B2(new_n669), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n672), .A2(new_n673), .ZN(G401));
  XNOR2_X1  g249(.A(G2072), .B(G2078), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT17), .ZN(new_n676));
  XOR2_X1   g251(.A(G2084), .B(G2090), .Z(new_n677));
  XNOR2_X1  g252(.A(G2067), .B(G2678), .ZN(new_n678));
  OAI21_X1  g253(.A(new_n676), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n677), .A2(new_n678), .ZN(new_n680));
  OR3_X1    g255(.A1(new_n677), .A2(new_n675), .A3(new_n678), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n679), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n677), .A2(new_n675), .A3(new_n678), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n683), .B(KEYINPUT18), .Z(new_n684));
  NAND2_X1  g259(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(new_n653), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(G2100), .ZN(G227));
  XOR2_X1   g262(.A(G1971), .B(G1976), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT19), .ZN(new_n689));
  XOR2_X1   g264(.A(G1956), .B(G2474), .Z(new_n690));
  XOR2_X1   g265(.A(G1961), .B(G1966), .Z(new_n691));
  NOR2_X1   g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  AND2_X1   g268(.A1(new_n690), .A2(new_n691), .ZN(new_n694));
  OR2_X1    g269(.A1(new_n694), .A2(new_n692), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n689), .A2(new_n694), .ZN(new_n696));
  XOR2_X1   g271(.A(KEYINPUT83), .B(KEYINPUT20), .Z(new_n697));
  OAI221_X1 g272(.A(new_n693), .B1(new_n695), .B2(new_n689), .C1(new_n696), .C2(new_n697), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n698), .B1(new_n696), .B2(new_n697), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(G1986), .ZN(new_n700));
  XOR2_X1   g275(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  AND2_X1   g277(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n700), .A2(new_n702), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(G1991), .B(G1996), .ZN(new_n706));
  INV_X1    g281(.A(G1981), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  AND2_X1   g283(.A1(new_n705), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n705), .A2(new_n708), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n709), .A2(new_n710), .ZN(G229));
  INV_X1    g286(.A(G16), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(G23), .ZN(new_n713));
  INV_X1    g288(.A(G288), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n713), .B1(new_n714), .B2(new_n712), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT33), .ZN(new_n716));
  XOR2_X1   g291(.A(KEYINPUT86), .B(G1976), .Z(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n712), .A2(G6), .ZN(new_n719));
  INV_X1    g294(.A(G305), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n719), .B1(new_n720), .B2(new_n712), .ZN(new_n721));
  XNOR2_X1  g296(.A(KEYINPUT32), .B(G1981), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT85), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n721), .B(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n718), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(G166), .A2(G16), .ZN(new_n726));
  NOR2_X1   g301(.A1(G16), .A2(G22), .ZN(new_n727));
  INV_X1    g302(.A(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(G1971), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n729), .B(new_n730), .ZN(new_n731));
  OR3_X1    g306(.A1(new_n725), .A2(KEYINPUT34), .A3(new_n731), .ZN(new_n732));
  OAI21_X1  g307(.A(KEYINPUT34), .B1(new_n725), .B2(new_n731), .ZN(new_n733));
  INV_X1    g308(.A(G29), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(G25), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n474), .A2(G131), .ZN(new_n736));
  INV_X1    g311(.A(G119), .ZN(new_n737));
  INV_X1    g312(.A(new_n476), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n736), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(G95), .ZN(new_n740));
  AND3_X1   g315(.A1(new_n740), .A2(new_n462), .A3(KEYINPUT84), .ZN(new_n741));
  AOI21_X1  g316(.A(KEYINPUT84), .B1(new_n740), .B2(new_n462), .ZN(new_n742));
  OAI221_X1 g317(.A(G2104), .B1(G107), .B2(new_n462), .C1(new_n741), .C2(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(new_n743), .ZN(new_n744));
  OR2_X1    g319(.A1(new_n739), .A2(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(new_n745), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n735), .B1(new_n746), .B2(new_n734), .ZN(new_n747));
  XOR2_X1   g322(.A(KEYINPUT35), .B(G1991), .Z(new_n748));
  INV_X1    g323(.A(new_n748), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n747), .B(new_n749), .ZN(new_n750));
  OR2_X1    g325(.A1(G16), .A2(G24), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(G290), .B2(new_n712), .ZN(new_n752));
  INV_X1    g327(.A(G1986), .ZN(new_n753));
  AND2_X1   g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n752), .A2(new_n753), .ZN(new_n755));
  NOR3_X1   g330(.A1(new_n750), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n732), .A2(new_n733), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n757), .A2(KEYINPUT36), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT36), .ZN(new_n759));
  NAND4_X1  g334(.A1(new_n732), .A2(new_n759), .A3(new_n733), .A4(new_n756), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n712), .A2(G20), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT23), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(new_n629), .B2(new_n712), .ZN(new_n764));
  OR2_X1    g339(.A1(new_n764), .A2(KEYINPUT95), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n764), .A2(KEYINPUT95), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g342(.A(G1956), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n734), .A2(G35), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G162), .B2(new_n734), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT29), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n772), .A2(G2090), .ZN(new_n773));
  NAND3_X1  g348(.A1(new_n765), .A2(G1956), .A3(new_n766), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n769), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT96), .ZN(new_n776));
  NOR2_X1   g351(.A1(G168), .A2(new_n712), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(new_n712), .B2(G21), .ZN(new_n778));
  INV_X1    g353(.A(G1966), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  XOR2_X1   g355(.A(KEYINPUT31), .B(G11), .Z(new_n781));
  NOR2_X1   g356(.A1(new_n652), .A2(new_n734), .ZN(new_n782));
  INV_X1    g357(.A(G28), .ZN(new_n783));
  OR2_X1    g358(.A1(new_n783), .A2(KEYINPUT30), .ZN(new_n784));
  AOI21_X1  g359(.A(G29), .B1(new_n783), .B2(KEYINPUT30), .ZN(new_n785));
  AOI211_X1 g360(.A(new_n781), .B(new_n782), .C1(new_n784), .C2(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(G2084), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n734), .B1(KEYINPUT24), .B2(G34), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(KEYINPUT24), .B2(G34), .ZN(new_n789));
  INV_X1    g364(.A(G160), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n789), .B1(new_n790), .B2(G29), .ZN(new_n791));
  OAI211_X1 g366(.A(new_n780), .B(new_n786), .C1(new_n787), .C2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n734), .A2(G33), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n474), .A2(G139), .ZN(new_n794));
  INV_X1    g369(.A(new_n794), .ZN(new_n795));
  OAI21_X1  g370(.A(G127), .B1(new_n463), .B2(new_n464), .ZN(new_n796));
  NAND2_X1  g371(.A1(G115), .A2(G2104), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n462), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT25), .ZN(new_n800));
  NOR3_X1   g375(.A1(new_n795), .A2(new_n798), .A3(new_n800), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n793), .B1(new_n801), .B2(new_n734), .ZN(new_n802));
  XOR2_X1   g377(.A(new_n802), .B(G2072), .Z(new_n803));
  INV_X1    g378(.A(G1961), .ZN(new_n804));
  NOR2_X1   g379(.A1(G171), .A2(new_n712), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(G5), .B2(new_n712), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n803), .B1(new_n804), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(G164), .A2(G29), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(G27), .B2(G29), .ZN(new_n809));
  INV_X1    g384(.A(G2078), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(new_n778), .B2(new_n779), .ZN(new_n812));
  OR3_X1    g387(.A1(new_n792), .A2(new_n807), .A3(new_n812), .ZN(new_n813));
  XOR2_X1   g388(.A(KEYINPUT90), .B(KEYINPUT26), .Z(new_n814));
  NAND3_X1  g389(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n462), .A2(G105), .A3(G2104), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n474), .A2(G141), .ZN(new_n819));
  INV_X1    g394(.A(G129), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n819), .B1(new_n820), .B2(new_n738), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n818), .A2(new_n821), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT91), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n823), .A2(G29), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n734), .A2(G32), .ZN(new_n825));
  XNOR2_X1  g400(.A(KEYINPUT27), .B(G1996), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n824), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT92), .ZN(new_n828));
  NOR2_X1   g403(.A1(G4), .A2(G16), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n829), .B1(new_n624), .B2(G16), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(G1348), .ZN(new_n831));
  NOR3_X1   g406(.A1(new_n813), .A2(new_n828), .A3(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n712), .A2(G19), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n833), .B(KEYINPUT87), .Z(new_n834));
  AOI21_X1  g409(.A(new_n834), .B1(new_n637), .B2(G16), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(G1341), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n734), .A2(G26), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT28), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n476), .A2(G128), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT88), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n839), .B(new_n840), .ZN(new_n841));
  OR2_X1    g416(.A1(G104), .A2(G2105), .ZN(new_n842));
  INV_X1    g417(.A(G2104), .ZN(new_n843));
  INV_X1    g418(.A(G116), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n843), .B1(new_n844), .B2(G2105), .ZN(new_n845));
  AOI22_X1  g420(.A1(new_n474), .A2(G140), .B1(new_n842), .B2(new_n845), .ZN(new_n846));
  AND2_X1   g421(.A1(new_n841), .A2(new_n846), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n838), .B1(new_n847), .B2(new_n734), .ZN(new_n848));
  XNOR2_X1  g423(.A(KEYINPUT89), .B(G2067), .ZN(new_n849));
  INV_X1    g424(.A(new_n849), .ZN(new_n850));
  AND2_X1   g425(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n848), .A2(new_n850), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n809), .A2(new_n810), .ZN(new_n853));
  NOR3_X1   g428(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  OAI21_X1  g429(.A(KEYINPUT94), .B1(new_n772), .B2(G2090), .ZN(new_n855));
  OR3_X1    g430(.A1(new_n772), .A2(KEYINPUT94), .A3(G2090), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n854), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n826), .B1(new_n824), .B2(new_n825), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n806), .A2(new_n804), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n791), .A2(new_n787), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  OR3_X1    g436(.A1(new_n858), .A2(KEYINPUT93), .A3(new_n861), .ZN(new_n862));
  OAI21_X1  g437(.A(KEYINPUT93), .B1(new_n858), .B2(new_n861), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n857), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  AND4_X1   g439(.A1(new_n776), .A2(new_n832), .A3(new_n836), .A4(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT97), .ZN(new_n866));
  AND3_X1   g441(.A1(new_n761), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n866), .B1(new_n761), .B2(new_n865), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n867), .A2(new_n868), .ZN(G311));
  NAND2_X1  g444(.A1(new_n761), .A2(new_n865), .ZN(G150));
  AOI22_X1  g445(.A1(new_n506), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n871), .A2(new_n511), .ZN(new_n872));
  INV_X1    g447(.A(G55), .ZN(new_n873));
  INV_X1    g448(.A(G93), .ZN(new_n874));
  OAI22_X1  g449(.A1(new_n541), .A2(new_n873), .B1(new_n539), .B2(new_n874), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n877), .B1(new_n562), .B2(new_n563), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n557), .A2(new_n560), .A3(new_n876), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(KEYINPUT38), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n624), .A2(G559), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n881), .B(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT39), .ZN(new_n884));
  AOI21_X1  g459(.A(G860), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n885), .B1(new_n884), .B2(new_n883), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n877), .A2(G860), .ZN(new_n887));
  XOR2_X1   g462(.A(new_n887), .B(KEYINPUT37), .Z(new_n888));
  NAND2_X1  g463(.A1(new_n886), .A2(new_n888), .ZN(G145));
  INV_X1    g464(.A(KEYINPUT40), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT101), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n474), .A2(G142), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(KEYINPUT100), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n476), .A2(G130), .ZN(new_n894));
  NOR2_X1   g469(.A1(G106), .A2(G2105), .ZN(new_n895));
  OAI21_X1  g470(.A(G2104), .B1(new_n462), .B2(G118), .ZN(new_n896));
  OAI211_X1 g471(.A(new_n893), .B(new_n894), .C1(new_n895), .C2(new_n896), .ZN(new_n897));
  AND2_X1   g472(.A1(new_n897), .A2(new_n642), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n897), .A2(new_n642), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n745), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  NOR3_X1   g476(.A1(new_n898), .A2(new_n899), .A3(new_n745), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n891), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n902), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n904), .A2(KEYINPUT101), .A3(new_n900), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n822), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n907), .A2(new_n801), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n908), .B1(new_n823), .B2(new_n801), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n501), .A2(KEYINPUT99), .ZN(new_n910));
  AOI22_X1  g485(.A1(G126), .A2(new_n476), .B1(new_n498), .B2(new_n499), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT99), .ZN(new_n912));
  NAND4_X1  g487(.A1(new_n911), .A2(new_n912), .A3(new_n490), .A4(new_n495), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n910), .A2(new_n913), .ZN(new_n914));
  XOR2_X1   g489(.A(new_n847), .B(new_n914), .Z(new_n915));
  OR2_X1    g490(.A1(new_n909), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n909), .A2(new_n915), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n906), .A2(new_n918), .ZN(new_n919));
  NAND4_X1  g494(.A1(new_n916), .A2(new_n903), .A3(new_n905), .A4(new_n917), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  XNOR2_X1  g496(.A(G162), .B(G160), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n922), .B(KEYINPUT98), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n923), .B(new_n652), .ZN(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(G37), .B1(new_n921), .B2(new_n925), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n901), .A2(new_n902), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n916), .A2(new_n917), .A3(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT102), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n916), .A2(new_n927), .A3(KEYINPUT102), .A4(new_n917), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n932), .A2(new_n919), .A3(new_n924), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT103), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n926), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n934), .B1(new_n926), .B2(new_n933), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n890), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n926), .A2(new_n933), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n939), .A2(KEYINPUT103), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n940), .A2(KEYINPUT40), .A3(new_n935), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n938), .A2(new_n941), .ZN(G395));
  INV_X1    g517(.A(KEYINPUT107), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n619), .A2(G299), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n621), .A2(new_n629), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT41), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n944), .A2(KEYINPUT41), .A3(new_n945), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(KEYINPUT104), .ZN(new_n951));
  AOI21_X1  g526(.A(KEYINPUT104), .B1(new_n946), .B2(new_n947), .ZN(new_n952));
  INV_X1    g527(.A(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n635), .A2(new_n880), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n634), .A2(new_n878), .A3(new_n879), .ZN(new_n955));
  AOI22_X1  g530(.A1(new_n951), .A2(new_n953), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  AND3_X1   g531(.A1(new_n954), .A2(new_n955), .A3(new_n946), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(G290), .A2(new_n720), .ZN(new_n959));
  OAI211_X1 g534(.A(G305), .B(new_n600), .C1(new_n607), .C2(new_n608), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(G303), .A2(G288), .ZN(new_n962));
  NAND2_X1  g537(.A1(G166), .A2(new_n714), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n961), .A2(new_n964), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n959), .A2(new_n962), .A3(new_n963), .A4(new_n960), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  XNOR2_X1  g542(.A(KEYINPUT105), .B(KEYINPUT42), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT105), .ZN(new_n970));
  AOI22_X1  g545(.A1(new_n965), .A2(new_n966), .B1(new_n970), .B2(KEYINPUT42), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n943), .B1(new_n958), .B2(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n954), .A2(new_n955), .A3(new_n946), .ZN(new_n975));
  AND2_X1   g550(.A1(new_n954), .A2(new_n955), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n952), .B1(new_n950), .B2(KEYINPUT104), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n975), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  OAI21_X1  g553(.A(KEYINPUT106), .B1(new_n978), .B2(new_n972), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT106), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n958), .A2(new_n980), .A3(new_n973), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n978), .A2(KEYINPUT107), .A3(new_n972), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n974), .A2(new_n979), .A3(new_n981), .A4(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(G868), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(KEYINPUT108), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT108), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n983), .A2(new_n986), .A3(G868), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n877), .A2(new_n610), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n985), .A2(new_n987), .A3(new_n988), .ZN(G295));
  NAND3_X1  g564(.A1(new_n985), .A2(new_n987), .A3(new_n988), .ZN(G331));
  INV_X1    g565(.A(KEYINPUT43), .ZN(new_n991));
  XNOR2_X1  g566(.A(G168), .B(G171), .ZN(new_n992));
  INV_X1    g567(.A(new_n563), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n876), .B1(new_n993), .B2(new_n561), .ZN(new_n994));
  INV_X1    g569(.A(new_n879), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n992), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(new_n946), .ZN(new_n997));
  XNOR2_X1  g572(.A(G168), .B(G301), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n878), .A2(new_n998), .A3(new_n879), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT109), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n878), .A2(new_n998), .A3(KEYINPUT109), .A4(new_n879), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n997), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  AOI22_X1  g578(.A1(new_n996), .A2(new_n999), .B1(new_n948), .B2(new_n949), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n967), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(new_n967), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n996), .A2(new_n946), .A3(new_n999), .ZN(new_n1007));
  AOI22_X1  g582(.A1(new_n1001), .A2(new_n1002), .B1(new_n880), .B2(new_n992), .ZN(new_n1008));
  OAI211_X1 g583(.A(new_n1006), .B(new_n1007), .C1(new_n1008), .C2(new_n977), .ZN(new_n1009));
  INV_X1    g584(.A(G37), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1005), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(KEYINPUT110), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT110), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n1005), .A2(new_n1009), .A3(new_n1013), .A4(new_n1010), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n991), .B1(new_n1012), .B2(new_n1014), .ZN(new_n1015));
  AND2_X1   g590(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1007), .B1(new_n1008), .B2(new_n977), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(new_n967), .ZN(new_n1018));
  AOI21_X1  g593(.A(KEYINPUT43), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g594(.A(KEYINPUT44), .B1(new_n1015), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT44), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n991), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1011), .A2(KEYINPUT43), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1021), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1020), .A2(new_n1024), .ZN(G397));
  NAND3_X1  g600(.A1(new_n521), .A2(new_n532), .A3(G8), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(KEYINPUT55), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT55), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n521), .A2(new_n532), .A3(new_n1028), .A4(G8), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(G1384), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n501), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(KEYINPUT50), .ZN(new_n1033));
  INV_X1    g608(.A(new_n467), .ZN(new_n1034));
  INV_X1    g609(.A(new_n470), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1034), .A2(new_n1035), .A3(G40), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT50), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n501), .A2(new_n1038), .A3(new_n1031), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1033), .A2(new_n1037), .A3(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(G2090), .B1(new_n1040), .B2(KEYINPUT116), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1036), .B1(new_n1032), .B2(KEYINPUT50), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT116), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1042), .A2(new_n1043), .A3(new_n1039), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT45), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1036), .B1(new_n1032), .B2(new_n1045), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1045), .A2(G1384), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n910), .A2(new_n913), .A3(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  AOI22_X1  g624(.A1(new_n1041), .A2(new_n1044), .B1(new_n730), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(G8), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1030), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1027), .A2(G8), .A3(new_n1029), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1049), .A2(new_n730), .ZN(new_n1054));
  INV_X1    g629(.A(G2090), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1042), .A2(new_n1055), .A3(new_n1039), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1053), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(G86), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n594), .B1(new_n539), .B2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g634(.A(G61), .B1(new_n526), .B2(new_n527), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n511), .B1(new_n1060), .B2(new_n590), .ZN(new_n1061));
  OAI21_X1  g636(.A(G1981), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n592), .A2(new_n707), .A3(new_n593), .A4(new_n594), .ZN(new_n1063));
  AND3_X1   g638(.A1(new_n1062), .A2(new_n1063), .A3(KEYINPUT49), .ZN(new_n1064));
  AOI21_X1  g639(.A(KEYINPUT49), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n501), .A2(G160), .A3(G40), .A4(new_n1031), .ZN(new_n1067));
  AND2_X1   g642(.A1(new_n1067), .A2(G8), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n714), .A2(G1976), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1069), .A2(new_n1067), .A3(G8), .ZN(new_n1070));
  AOI22_X1  g645(.A1(new_n1066), .A2(new_n1068), .B1(new_n1070), .B2(KEYINPUT52), .ZN(new_n1071));
  INV_X1    g646(.A(G1976), .ZN(new_n1072));
  AOI21_X1  g647(.A(KEYINPUT52), .B1(G288), .B2(new_n1072), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1069), .A2(new_n1067), .A3(G8), .A4(new_n1073), .ZN(new_n1074));
  AND2_X1   g649(.A1(new_n1074), .A2(KEYINPUT114), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1074), .A2(KEYINPUT114), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1071), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1057), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1052), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(KEYINPUT124), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1046), .A2(new_n810), .A3(new_n1048), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT53), .ZN(new_n1082));
  AOI22_X1  g657(.A1(new_n1081), .A2(new_n1082), .B1(new_n1040), .B2(new_n804), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n910), .A2(new_n1031), .A3(new_n913), .ZN(new_n1084));
  AND2_X1   g659(.A1(new_n1084), .A2(new_n1045), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT123), .ZN(new_n1086));
  NOR3_X1   g661(.A1(new_n1036), .A2(new_n1082), .A3(G2078), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1048), .A2(new_n1087), .ZN(new_n1088));
  NOR3_X1   g663(.A1(new_n1085), .A2(new_n1086), .A3(new_n1088), .ZN(new_n1089));
  AND2_X1   g664(.A1(new_n1048), .A2(new_n1087), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1084), .A2(new_n1045), .ZN(new_n1091));
  AOI21_X1  g666(.A(KEYINPUT123), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  OAI211_X1 g667(.A(G301), .B(new_n1083), .C1(new_n1089), .C2(new_n1092), .ZN(new_n1093));
  AND2_X1   g668(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT122), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n501), .A2(new_n1047), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1082), .A2(G2078), .ZN(new_n1097));
  AND3_X1   g672(.A1(new_n1046), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(G1961), .B1(new_n1042), .B2(new_n1039), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1095), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1040), .A2(new_n804), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1046), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1101), .A2(KEYINPUT122), .A3(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1094), .B1(new_n1100), .B2(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1093), .B1(new_n1104), .B2(G301), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT54), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT124), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1052), .A2(new_n1078), .A3(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(KEYINPUT51), .A2(G8), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1040), .A2(G2084), .ZN(new_n1111));
  AOI21_X1  g686(.A(G1966), .B1(new_n1046), .B2(new_n1096), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(G286), .ZN(new_n1114));
  OAI21_X1  g689(.A(G168), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1110), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1113), .A2(G168), .ZN(new_n1117));
  AOI21_X1  g692(.A(KEYINPUT51), .B1(new_n1117), .B2(G8), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1119));
  AND4_X1   g694(.A1(new_n1080), .A2(new_n1107), .A3(new_n1109), .A4(new_n1119), .ZN(new_n1120));
  OAI211_X1 g695(.A(KEYINPUT126), .B(new_n1083), .C1(new_n1089), .C2(new_n1092), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1121), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1086), .B1(new_n1085), .B2(new_n1088), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1090), .A2(KEYINPUT123), .A3(new_n1091), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(KEYINPUT126), .B1(new_n1125), .B2(new_n1083), .ZN(new_n1126));
  OAI21_X1  g701(.A(G171), .B1(new_n1122), .B2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(G171), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1128));
  NOR3_X1   g703(.A1(new_n1098), .A2(new_n1099), .A3(new_n1095), .ZN(new_n1129));
  AOI21_X1  g704(.A(KEYINPUT122), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1128), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT125), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  OAI211_X1 g708(.A(KEYINPUT125), .B(new_n1128), .C1(new_n1129), .C2(new_n1130), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1127), .A2(new_n1135), .A3(KEYINPUT54), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT127), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  AND3_X1   g713(.A1(new_n1033), .A2(new_n1037), .A3(new_n1039), .ZN(new_n1139));
  XNOR2_X1  g714(.A(KEYINPUT56), .B(G2072), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1140), .ZN(new_n1141));
  OAI22_X1  g716(.A1(new_n1139), .A2(G1956), .B1(new_n1049), .B2(new_n1141), .ZN(new_n1142));
  XNOR2_X1  g717(.A(new_n629), .B(KEYINPUT57), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1145));
  AND2_X1   g720(.A1(new_n620), .A2(new_n623), .ZN(new_n1146));
  INV_X1    g721(.A(G1348), .ZN(new_n1147));
  INV_X1    g722(.A(G2067), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1067), .ZN(new_n1149));
  AOI22_X1  g724(.A1(new_n1040), .A2(new_n1147), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1145), .B1(new_n1146), .B2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1040), .A2(new_n768), .ZN(new_n1152));
  OAI211_X1 g727(.A(new_n1143), .B(new_n1152), .C1(new_n1049), .C2(new_n1141), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1151), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1145), .A2(new_n1153), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT61), .ZN(new_n1156));
  AOI21_X1  g731(.A(KEYINPUT121), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT121), .ZN(new_n1158));
  AOI211_X1 g733(.A(new_n1158), .B(KEYINPUT61), .C1(new_n1145), .C2(new_n1153), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1157), .A2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1150), .A2(KEYINPUT60), .A3(new_n624), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1149), .A2(new_n1148), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1162), .B1(new_n1139), .B2(G1348), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT60), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1146), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1161), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1145), .A2(KEYINPUT61), .A3(new_n1153), .ZN(new_n1168));
  XNOR2_X1  g743(.A(KEYINPUT58), .B(G1341), .ZN(new_n1169));
  OAI22_X1  g744(.A1(new_n1049), .A2(G1996), .B1(new_n1149), .B2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1170), .A2(KEYINPUT119), .A3(new_n564), .ZN(new_n1171));
  XNOR2_X1  g746(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  AND2_X1   g748(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1174));
  OAI211_X1 g749(.A(new_n1167), .B(new_n1168), .C1(new_n1173), .C2(new_n1174), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1154), .B1(new_n1160), .B2(new_n1175), .ZN(new_n1176));
  NAND4_X1  g751(.A1(new_n1127), .A2(new_n1135), .A3(KEYINPUT127), .A4(KEYINPUT54), .ZN(new_n1177));
  NAND4_X1  g752(.A1(new_n1120), .A2(new_n1138), .A3(new_n1176), .A4(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1077), .A2(KEYINPUT115), .ZN(new_n1179));
  XNOR2_X1  g754(.A(new_n1074), .B(KEYINPUT114), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT115), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1180), .A2(new_n1181), .A3(new_n1071), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1179), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1066), .A2(new_n1068), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1184), .A2(new_n1072), .A3(new_n714), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1185), .B1(G1981), .B2(G305), .ZN(new_n1186));
  AOI22_X1  g761(.A1(new_n1183), .A2(new_n1057), .B1(new_n1068), .B2(new_n1186), .ZN(new_n1187));
  XNOR2_X1  g762(.A(KEYINPUT117), .B(KEYINPUT63), .ZN(new_n1188));
  INV_X1    g763(.A(new_n1188), .ZN(new_n1189));
  AOI22_X1  g764(.A1(new_n1139), .A2(new_n1055), .B1(new_n1049), .B2(new_n730), .ZN(new_n1190));
  OAI211_X1 g765(.A(new_n1180), .B(new_n1071), .C1(new_n1190), .C2(new_n1053), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1040), .A2(KEYINPUT116), .ZN(new_n1192));
  AND3_X1   g767(.A1(new_n1192), .A2(new_n1055), .A3(new_n1044), .ZN(new_n1193));
  INV_X1    g768(.A(new_n1054), .ZN(new_n1194));
  OAI21_X1  g769(.A(G8), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1191), .B1(new_n1195), .B2(new_n1030), .ZN(new_n1196));
  OAI211_X1 g771(.A(G8), .B(G168), .C1(new_n1111), .C2(new_n1112), .ZN(new_n1197));
  INV_X1    g772(.A(new_n1197), .ZN(new_n1198));
  AOI21_X1  g773(.A(new_n1189), .B1(new_n1196), .B2(new_n1198), .ZN(new_n1199));
  OAI21_X1  g774(.A(KEYINPUT63), .B1(new_n1190), .B2(new_n1053), .ZN(new_n1200));
  AND3_X1   g775(.A1(new_n1054), .A2(new_n1030), .A3(new_n1056), .ZN(new_n1201));
  NOR3_X1   g776(.A1(new_n1200), .A2(new_n1197), .A3(new_n1201), .ZN(new_n1202));
  AND2_X1   g777(.A1(new_n1202), .A2(new_n1183), .ZN(new_n1203));
  OAI211_X1 g778(.A(KEYINPUT118), .B(new_n1187), .C1(new_n1199), .C2(new_n1203), .ZN(new_n1204));
  INV_X1    g779(.A(KEYINPUT118), .ZN(new_n1205));
  NAND3_X1  g780(.A1(new_n1052), .A2(new_n1078), .A3(new_n1198), .ZN(new_n1206));
  AOI22_X1  g781(.A1(new_n1206), .A2(new_n1188), .B1(new_n1202), .B2(new_n1183), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1183), .A2(new_n1057), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1186), .A2(new_n1068), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  OAI21_X1  g785(.A(new_n1205), .B1(new_n1207), .B2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1204), .A2(new_n1211), .ZN(new_n1212));
  OR2_X1    g787(.A1(new_n1119), .A2(KEYINPUT62), .ZN(new_n1213));
  OR2_X1    g788(.A1(new_n1104), .A2(G301), .ZN(new_n1214));
  AOI21_X1  g789(.A(new_n1214), .B1(new_n1119), .B2(KEYINPUT62), .ZN(new_n1215));
  NAND4_X1  g790(.A1(new_n1213), .A2(new_n1215), .A3(new_n1080), .A4(new_n1109), .ZN(new_n1216));
  NAND3_X1  g791(.A1(new_n1178), .A2(new_n1212), .A3(new_n1216), .ZN(new_n1217));
  NAND3_X1  g792(.A1(new_n1084), .A2(new_n1045), .A3(new_n1037), .ZN(new_n1218));
  OR2_X1    g793(.A1(new_n1218), .A2(KEYINPUT111), .ZN(new_n1219));
  NAND2_X1  g794(.A1(new_n1218), .A2(KEYINPUT111), .ZN(new_n1220));
  AND2_X1   g795(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  XNOR2_X1  g796(.A(new_n847), .B(G2067), .ZN(new_n1222));
  XNOR2_X1  g797(.A(new_n1222), .B(KEYINPUT112), .ZN(new_n1223));
  NAND2_X1  g798(.A1(new_n907), .A2(G1996), .ZN(new_n1224));
  OAI21_X1  g799(.A(new_n1224), .B1(new_n823), .B2(G1996), .ZN(new_n1225));
  OR2_X1    g800(.A1(new_n1223), .A2(new_n1225), .ZN(new_n1226));
  XNOR2_X1  g801(.A(new_n745), .B(new_n749), .ZN(new_n1227));
  OAI21_X1  g802(.A(new_n1221), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1228));
  INV_X1    g803(.A(new_n1221), .ZN(new_n1229));
  XNOR2_X1  g804(.A(G290), .B(new_n753), .ZN(new_n1230));
  OAI21_X1  g805(.A(new_n1228), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  INV_X1    g806(.A(KEYINPUT113), .ZN(new_n1232));
  XNOR2_X1  g807(.A(new_n1231), .B(new_n1232), .ZN(new_n1233));
  NAND2_X1  g808(.A1(new_n1217), .A2(new_n1233), .ZN(new_n1234));
  INV_X1    g809(.A(KEYINPUT46), .ZN(new_n1235));
  OR3_X1    g810(.A1(new_n1229), .A2(new_n1235), .A3(G1996), .ZN(new_n1236));
  OAI21_X1  g811(.A(new_n1221), .B1(new_n1223), .B2(new_n907), .ZN(new_n1237));
  OAI21_X1  g812(.A(new_n1235), .B1(new_n1229), .B2(G1996), .ZN(new_n1238));
  NAND3_X1  g813(.A1(new_n1236), .A2(new_n1237), .A3(new_n1238), .ZN(new_n1239));
  XNOR2_X1  g814(.A(new_n1239), .B(KEYINPUT47), .ZN(new_n1240));
  OR3_X1    g815(.A1(new_n1229), .A2(G1986), .A3(G290), .ZN(new_n1241));
  INV_X1    g816(.A(KEYINPUT48), .ZN(new_n1242));
  OR2_X1    g817(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g818(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1244));
  NAND3_X1  g819(.A1(new_n1243), .A2(new_n1228), .A3(new_n1244), .ZN(new_n1245));
  NAND2_X1  g820(.A1(new_n847), .A2(new_n1148), .ZN(new_n1246));
  NAND2_X1  g821(.A1(new_n746), .A2(new_n748), .ZN(new_n1247));
  OAI21_X1  g822(.A(new_n1246), .B1(new_n1226), .B2(new_n1247), .ZN(new_n1248));
  NAND2_X1  g823(.A1(new_n1248), .A2(new_n1221), .ZN(new_n1249));
  AND3_X1   g824(.A1(new_n1240), .A2(new_n1245), .A3(new_n1249), .ZN(new_n1250));
  NAND2_X1  g825(.A1(new_n1234), .A2(new_n1250), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g826(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1253));
  NOR2_X1   g827(.A1(G227), .A2(new_n460), .ZN(new_n1254));
  OAI221_X1 g828(.A(new_n1254), .B1(new_n672), .B2(new_n673), .C1(new_n709), .C2(new_n710), .ZN(new_n1255));
  INV_X1    g829(.A(new_n939), .ZN(new_n1256));
  NOR3_X1   g830(.A1(new_n1253), .A2(new_n1255), .A3(new_n1256), .ZN(G308));
  OR3_X1    g831(.A1(new_n1253), .A2(new_n1255), .A3(new_n1256), .ZN(G225));
endmodule


