//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 0 0 0 0 1 0 0 0 1 0 0 0 0 1 1 1 0 0 1 0 0 0 1 1 0 1 0 0 0 1 1 0 1 1 1 1 0 0 0 0 1 1 0 0 0 1 0 0 0 0 1 1 1 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:43 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n678, new_n679, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n691,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n746, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n903, new_n904, new_n905,
    new_n906, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980;
  INV_X1    g000(.A(G104), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(KEYINPUT78), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT78), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G104), .ZN(new_n190));
  AOI21_X1  g004(.A(G107), .B1(new_n188), .B2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G107), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n192), .A2(G104), .ZN(new_n193));
  OAI21_X1  g007(.A(G101), .B1(new_n191), .B2(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(KEYINPUT79), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT2), .ZN(new_n196));
  INV_X1    g010(.A(G113), .ZN(new_n197));
  OAI21_X1  g011(.A(KEYINPUT66), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT66), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n199), .A2(KEYINPUT2), .A3(G113), .ZN(new_n200));
  AOI22_X1  g014(.A1(new_n198), .A2(new_n200), .B1(new_n196), .B2(new_n197), .ZN(new_n201));
  XNOR2_X1  g015(.A(G116), .B(G119), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(KEYINPUT5), .ZN(new_n203));
  INV_X1    g017(.A(G116), .ZN(new_n204));
  NOR3_X1   g018(.A1(new_n204), .A2(KEYINPUT5), .A3(G119), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n205), .A2(new_n197), .ZN(new_n206));
  AOI22_X1  g020(.A1(new_n201), .A2(new_n202), .B1(new_n203), .B2(new_n206), .ZN(new_n207));
  XNOR2_X1  g021(.A(KEYINPUT78), .B(G104), .ZN(new_n208));
  OAI21_X1  g022(.A(KEYINPUT3), .B1(new_n208), .B2(G107), .ZN(new_n209));
  NOR3_X1   g023(.A1(new_n187), .A2(KEYINPUT3), .A3(G107), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n210), .B1(new_n208), .B2(G107), .ZN(new_n211));
  INV_X1    g025(.A(G101), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n209), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT79), .ZN(new_n214));
  OAI211_X1 g028(.A(new_n214), .B(G101), .C1(new_n191), .C2(new_n193), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n195), .A2(new_n207), .A3(new_n213), .A4(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT3), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n188), .A2(new_n190), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n217), .B1(new_n218), .B2(new_n192), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n188), .A2(new_n190), .A3(G107), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n217), .A2(new_n192), .A3(G104), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g036(.A(G101), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  AND3_X1   g037(.A1(new_n223), .A2(KEYINPUT4), .A3(new_n213), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n198), .A2(new_n200), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n196), .A2(new_n197), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(new_n202), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n201), .A2(new_n202), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT4), .ZN(new_n232));
  OAI211_X1 g046(.A(new_n232), .B(G101), .C1(new_n219), .C2(new_n222), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n216), .B1(new_n224), .B2(new_n234), .ZN(new_n235));
  XNOR2_X1  g049(.A(G110), .B(G122), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  OAI211_X1 g052(.A(new_n236), .B(new_n216), .C1(new_n224), .C2(new_n234), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n238), .A2(KEYINPUT6), .A3(new_n239), .ZN(new_n240));
  AND2_X1   g054(.A1(KEYINPUT0), .A2(G128), .ZN(new_n241));
  XNOR2_X1  g055(.A(G143), .B(G146), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n241), .B1(new_n242), .B2(KEYINPUT64), .ZN(new_n243));
  INV_X1    g057(.A(G146), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G143), .ZN(new_n245));
  INV_X1    g059(.A(G143), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G146), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  NOR2_X1   g062(.A1(KEYINPUT0), .A2(G128), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n241), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT64), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n248), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n243), .A2(new_n252), .A3(G125), .ZN(new_n253));
  OAI21_X1  g067(.A(KEYINPUT1), .B1(new_n246), .B2(G146), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n246), .A2(G146), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n244), .A2(G143), .ZN(new_n256));
  OAI211_X1 g070(.A(G128), .B(new_n254), .C1(new_n255), .C2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(G128), .ZN(new_n258));
  OAI211_X1 g072(.A(new_n245), .B(new_n247), .C1(KEYINPUT1), .C2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n253), .B1(new_n260), .B2(G125), .ZN(new_n261));
  INV_X1    g075(.A(G953), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G224), .ZN(new_n263));
  XNOR2_X1  g077(.A(new_n263), .B(KEYINPUT83), .ZN(new_n264));
  XNOR2_X1  g078(.A(new_n261), .B(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT6), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n235), .A2(new_n266), .A3(new_n237), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n240), .A2(new_n265), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(KEYINPUT84), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT84), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n240), .A2(new_n270), .A3(new_n265), .A4(new_n267), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(new_n239), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n263), .A2(KEYINPUT7), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(KEYINPUT85), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n261), .A2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(new_n274), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT85), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n276), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n261), .A2(new_n278), .A3(new_n277), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  XOR2_X1   g096(.A(new_n236), .B(KEYINPUT8), .Z(new_n283));
  NAND3_X1  g097(.A1(new_n195), .A2(new_n213), .A3(new_n215), .ZN(new_n284));
  INV_X1    g098(.A(new_n207), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n283), .B1(new_n286), .B2(new_n216), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n282), .A2(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n273), .B1(new_n288), .B2(KEYINPUT86), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT86), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n290), .B1(new_n282), .B2(new_n287), .ZN(new_n291));
  AOI21_X1  g105(.A(G902), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n272), .A2(new_n292), .ZN(new_n293));
  OAI21_X1  g107(.A(G210), .B1(G237), .B2(G902), .ZN(new_n294));
  XOR2_X1   g108(.A(new_n294), .B(KEYINPUT87), .Z(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n293), .A2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(G952), .ZN(new_n298));
  AOI211_X1 g112(.A(G953), .B(new_n298), .C1(G234), .C2(G237), .ZN(new_n299));
  INV_X1    g113(.A(G902), .ZN(new_n300));
  AND2_X1   g114(.A1(KEYINPUT67), .A2(G953), .ZN(new_n301));
  NOR2_X1   g115(.A1(KEYINPUT67), .A2(G953), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  AOI211_X1 g117(.A(new_n300), .B(new_n303), .C1(G234), .C2(G237), .ZN(new_n304));
  XNOR2_X1  g118(.A(KEYINPUT21), .B(G898), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n299), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  OAI21_X1  g121(.A(G214), .B1(G237), .B2(G902), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n272), .A2(new_n292), .A3(new_n295), .ZN(new_n309));
  NAND4_X1  g123(.A1(new_n297), .A2(new_n307), .A3(new_n308), .A4(new_n309), .ZN(new_n310));
  XNOR2_X1  g124(.A(KEYINPUT9), .B(G234), .ZN(new_n311));
  OAI21_X1  g125(.A(G221), .B1(new_n311), .B2(G902), .ZN(new_n312));
  XOR2_X1   g126(.A(KEYINPUT82), .B(G469), .Z(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n303), .A2(G227), .ZN(new_n315));
  XNOR2_X1  g129(.A(new_n315), .B(KEYINPUT77), .ZN(new_n316));
  XNOR2_X1  g130(.A(G110), .B(G140), .ZN(new_n317));
  XNOR2_X1  g131(.A(new_n316), .B(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(G137), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n320), .A2(G134), .ZN(new_n321));
  INV_X1    g135(.A(G134), .ZN(new_n322));
  OAI21_X1  g136(.A(KEYINPUT11), .B1(new_n322), .B2(G137), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT11), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n324), .A2(new_n320), .A3(G134), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n321), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(G131), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  AOI211_X1 g142(.A(G131), .B(new_n321), .C1(new_n323), .C2(new_n325), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  AND2_X1   g144(.A1(new_n257), .A2(new_n259), .ZN(new_n331));
  NAND4_X1  g145(.A1(new_n195), .A2(new_n213), .A3(new_n331), .A4(new_n215), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT80), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT10), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n332), .A2(new_n333), .A3(KEYINPUT10), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n223), .A2(new_n213), .A3(KEYINPUT4), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n339), .A2(new_n243), .A3(new_n252), .A4(new_n233), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n330), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  AND3_X1   g155(.A1(new_n332), .A2(new_n333), .A3(KEYINPUT10), .ZN(new_n342));
  AOI21_X1  g156(.A(KEYINPUT10), .B1(new_n332), .B2(new_n333), .ZN(new_n343));
  OAI211_X1 g157(.A(new_n330), .B(new_n340), .C1(new_n342), .C2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n319), .B1(new_n341), .B2(new_n345), .ZN(new_n346));
  XOR2_X1   g160(.A(KEYINPUT81), .B(KEYINPUT12), .Z(new_n347));
  NAND2_X1  g161(.A1(new_n284), .A2(new_n260), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(new_n332), .ZN(new_n349));
  INV_X1    g163(.A(new_n330), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n347), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NOR2_X1   g165(.A1(KEYINPUT81), .A2(KEYINPUT12), .ZN(new_n352));
  AOI211_X1 g166(.A(new_n330), .B(new_n352), .C1(new_n348), .C2(new_n332), .ZN(new_n353));
  OAI211_X1 g167(.A(new_n344), .B(new_n318), .C1(new_n351), .C2(new_n353), .ZN(new_n354));
  AOI211_X1 g168(.A(G902), .B(new_n314), .C1(new_n346), .C2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(G469), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n344), .B1(new_n351), .B2(new_n353), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(new_n319), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n340), .B1(new_n342), .B2(new_n343), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(new_n350), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n360), .A2(new_n344), .A3(new_n318), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n358), .A2(new_n361), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n356), .B1(new_n362), .B2(new_n300), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n312), .B1(new_n355), .B2(new_n363), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n310), .A2(new_n364), .ZN(new_n365));
  XNOR2_X1  g179(.A(new_n201), .B(new_n228), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n243), .A2(new_n252), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n326), .A2(new_n327), .ZN(new_n368));
  AND2_X1   g182(.A1(new_n323), .A2(new_n325), .ZN(new_n369));
  OAI21_X1  g183(.A(G131), .B1(new_n369), .B2(new_n321), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n367), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  OAI21_X1  g185(.A(KEYINPUT65), .B1(new_n320), .B2(G134), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT65), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n373), .A2(new_n322), .A3(G137), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n320), .A2(G134), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n372), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(G131), .ZN(new_n377));
  AND4_X1   g191(.A1(new_n368), .A2(new_n377), .A3(new_n259), .A4(new_n257), .ZN(new_n378));
  OAI21_X1  g192(.A(KEYINPUT30), .B1(new_n371), .B2(new_n378), .ZN(new_n379));
  OAI211_X1 g193(.A(new_n243), .B(new_n252), .C1(new_n328), .C2(new_n329), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT30), .ZN(new_n381));
  NAND4_X1  g195(.A1(new_n368), .A2(new_n377), .A3(new_n259), .A4(new_n257), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n380), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n366), .B1(new_n379), .B2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(G237), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n303), .A2(G210), .A3(new_n385), .ZN(new_n386));
  XNOR2_X1  g200(.A(new_n386), .B(KEYINPUT27), .ZN(new_n387));
  XOR2_X1   g201(.A(KEYINPUT26), .B(G101), .Z(new_n388));
  XNOR2_X1  g202(.A(new_n387), .B(new_n388), .ZN(new_n389));
  AND3_X1   g203(.A1(new_n380), .A2(new_n366), .A3(new_n382), .ZN(new_n390));
  NOR3_X1   g204(.A1(new_n384), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT31), .ZN(new_n392));
  OAI21_X1  g206(.A(KEYINPUT68), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT69), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n366), .B1(new_n380), .B2(new_n382), .ZN(new_n395));
  OAI211_X1 g209(.A(new_n394), .B(KEYINPUT28), .C1(new_n390), .C2(new_n395), .ZN(new_n396));
  OR2_X1    g210(.A1(new_n390), .A2(KEYINPUT28), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n231), .B1(new_n371), .B2(new_n378), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n380), .A2(new_n366), .A3(new_n382), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n394), .B1(new_n401), .B2(KEYINPUT28), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n389), .B1(new_n398), .B2(new_n402), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n384), .A2(new_n390), .ZN(new_n404));
  INV_X1    g218(.A(new_n389), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n404), .A2(new_n392), .A3(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(new_n383), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n381), .B1(new_n380), .B2(new_n382), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n231), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n409), .A2(new_n405), .A3(new_n400), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT68), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n410), .A2(new_n411), .A3(KEYINPUT31), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n393), .A2(new_n403), .A3(new_n406), .A4(new_n412), .ZN(new_n413));
  NOR2_X1   g227(.A1(G472), .A2(G902), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n413), .A2(KEYINPUT32), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(KEYINPUT71), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n413), .A2(new_n414), .ZN(new_n417));
  XNOR2_X1  g231(.A(KEYINPUT70), .B(KEYINPUT32), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n401), .A2(KEYINPUT28), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(new_n397), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n405), .A2(KEYINPUT29), .ZN(new_n422));
  NOR3_X1   g236(.A1(new_n398), .A2(new_n402), .A3(new_n389), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT29), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n424), .B1(new_n404), .B2(new_n405), .ZN(new_n425));
  OAI221_X1 g239(.A(new_n300), .B1(new_n421), .B2(new_n422), .C1(new_n423), .C2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(G472), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT71), .ZN(new_n428));
  NAND4_X1  g242(.A1(new_n413), .A2(new_n428), .A3(KEYINPUT32), .A4(new_n414), .ZN(new_n429));
  NAND4_X1  g243(.A1(new_n416), .A2(new_n419), .A3(new_n427), .A4(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(G234), .ZN(new_n431));
  OAI21_X1  g245(.A(G217), .B1(new_n431), .B2(G902), .ZN(new_n432));
  OAI21_X1  g246(.A(KEYINPUT23), .B1(new_n258), .B2(G119), .ZN(new_n433));
  INV_X1    g247(.A(G119), .ZN(new_n434));
  OAI211_X1 g248(.A(new_n433), .B(KEYINPUT73), .C1(new_n434), .C2(G128), .ZN(new_n435));
  OAI21_X1  g249(.A(KEYINPUT73), .B1(new_n434), .B2(G128), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n436), .B(KEYINPUT23), .C1(G119), .C2(new_n258), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT72), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n439), .B1(new_n258), .B2(G119), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n434), .A2(KEYINPUT72), .A3(G128), .ZN(new_n441));
  AOI22_X1  g255(.A1(new_n440), .A2(new_n441), .B1(G119), .B2(new_n258), .ZN(new_n442));
  XOR2_X1   g256(.A(KEYINPUT24), .B(G110), .Z(new_n443));
  AOI22_X1  g257(.A1(new_n438), .A2(G110), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT74), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT16), .ZN(new_n446));
  INV_X1    g260(.A(G140), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n446), .A2(new_n447), .A3(G125), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(G125), .ZN(new_n449));
  INV_X1    g263(.A(G125), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(G140), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  OAI211_X1 g266(.A(new_n445), .B(new_n448), .C1(new_n452), .C2(new_n446), .ZN(new_n453));
  XNOR2_X1  g267(.A(G125), .B(G140), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n454), .A2(KEYINPUT74), .A3(KEYINPUT16), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n453), .A2(new_n244), .A3(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n244), .B1(new_n453), .B2(new_n455), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n444), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  OAI22_X1  g273(.A1(new_n438), .A2(G110), .B1(new_n442), .B2(new_n443), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n453), .A2(new_n455), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(G146), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n454), .A2(new_n244), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n460), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n459), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n303), .A2(G221), .A3(G234), .ZN(new_n466));
  XNOR2_X1  g280(.A(KEYINPUT22), .B(G137), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n466), .B(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n465), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n459), .A2(new_n464), .A3(new_n468), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n470), .A2(new_n300), .A3(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT75), .ZN(new_n473));
  AOI21_X1  g287(.A(KEYINPUT76), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT25), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n432), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT76), .ZN(new_n477));
  AND3_X1   g291(.A1(new_n459), .A2(new_n464), .A3(new_n468), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n468), .B1(new_n459), .B2(new_n464), .ZN(new_n479));
  NOR3_X1   g293(.A1(new_n478), .A2(new_n479), .A3(G902), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n477), .B1(new_n480), .B2(KEYINPUT75), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n475), .B1(new_n472), .B2(KEYINPUT76), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n478), .A2(new_n479), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n432), .A2(new_n300), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  AOI22_X1  g300(.A1(new_n476), .A2(new_n483), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT89), .ZN(new_n488));
  OR2_X1    g302(.A1(KEYINPUT67), .A2(G953), .ZN(new_n489));
  NAND2_X1  g303(.A1(KEYINPUT67), .A2(G953), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n489), .A2(G214), .A3(new_n385), .A4(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(new_n246), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n303), .A2(G143), .A3(G214), .A4(new_n385), .ZN(new_n493));
  AND2_X1   g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n488), .B1(new_n494), .B2(new_n327), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n492), .A2(new_n493), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n496), .A2(KEYINPUT89), .A3(G131), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n495), .A2(KEYINPUT17), .A3(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT91), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n457), .A2(new_n458), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT17), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n494), .A2(new_n327), .ZN(new_n503));
  INV_X1    g317(.A(new_n497), .ZN(new_n504));
  AOI21_X1  g318(.A(KEYINPUT89), .B1(new_n496), .B2(G131), .ZN(new_n505));
  OAI211_X1 g319(.A(new_n502), .B(new_n503), .C1(new_n504), .C2(new_n505), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n495), .A2(KEYINPUT91), .A3(KEYINPUT17), .A4(new_n497), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n500), .A2(new_n501), .A3(new_n506), .A4(new_n507), .ZN(new_n508));
  XNOR2_X1  g322(.A(G113), .B(G122), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n509), .B(new_n187), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT18), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n494), .B1(new_n511), .B2(new_n327), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n496), .A2(KEYINPUT18), .A3(G131), .ZN(new_n513));
  AOI21_X1  g327(.A(KEYINPUT88), .B1(new_n454), .B2(new_n244), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n514), .B1(new_n244), .B2(new_n454), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n452), .A2(KEYINPUT88), .A3(G146), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n512), .A2(new_n513), .A3(new_n515), .A4(new_n516), .ZN(new_n517));
  AND3_X1   g331(.A1(new_n508), .A2(new_n510), .A3(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n510), .B1(new_n508), .B2(new_n517), .ZN(new_n519));
  OAI211_X1 g333(.A(KEYINPUT92), .B(new_n300), .C1(new_n518), .C2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(G475), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n508), .A2(new_n517), .ZN(new_n522));
  INV_X1    g336(.A(new_n510), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n508), .A2(new_n510), .A3(new_n517), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(KEYINPUT92), .B1(new_n526), .B2(new_n300), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT20), .ZN(new_n528));
  AOI22_X1  g342(.A1(new_n495), .A2(new_n497), .B1(new_n494), .B2(new_n327), .ZN(new_n529));
  AND2_X1   g343(.A1(KEYINPUT90), .A2(KEYINPUT19), .ZN(new_n530));
  NOR2_X1   g344(.A1(KEYINPUT90), .A2(KEYINPUT19), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n454), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n532), .B1(new_n454), .B2(new_n531), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n462), .B1(G146), .B2(new_n533), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n517), .B1(new_n529), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(new_n523), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n525), .A2(new_n536), .ZN(new_n537));
  NOR2_X1   g351(.A1(G475), .A2(G902), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n528), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  AND3_X1   g353(.A1(new_n537), .A2(new_n528), .A3(new_n538), .ZN(new_n540));
  OAI22_X1  g354(.A1(new_n521), .A2(new_n527), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT97), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT13), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n543), .B1(new_n258), .B2(G143), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n258), .A2(G143), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n246), .A2(KEYINPUT13), .A3(G128), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(G134), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(KEYINPUT94), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT94), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n547), .A2(new_n550), .A3(G134), .ZN(new_n551));
  AND2_X1   g365(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n246), .A2(G128), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n553), .A2(new_n545), .A3(new_n322), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT93), .ZN(new_n555));
  INV_X1    g369(.A(G122), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n555), .B1(new_n556), .B2(G116), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n204), .A2(KEYINPUT93), .A3(G122), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n556), .A2(G116), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n559), .A2(new_n192), .A3(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n192), .B1(new_n559), .B2(new_n560), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n554), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  OAI21_X1  g378(.A(KEYINPUT95), .B1(new_n552), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n553), .A2(new_n545), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(G134), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n562), .B1(new_n554), .B2(new_n567), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n560), .B1(new_n559), .B2(KEYINPUT14), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n559), .A2(KEYINPUT14), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT96), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n559), .A2(KEYINPUT96), .A3(KEYINPUT14), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n569), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n568), .B1(new_n574), .B2(new_n192), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n549), .A2(new_n551), .ZN(new_n576));
  INV_X1    g390(.A(new_n563), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(new_n561), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT95), .ZN(new_n579));
  NAND4_X1  g393(.A1(new_n576), .A2(new_n578), .A3(new_n579), .A4(new_n554), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n565), .A2(new_n575), .A3(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n311), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n582), .A2(G217), .A3(new_n262), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n583), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n565), .A2(new_n575), .A3(new_n580), .A4(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n542), .B1(new_n587), .B2(new_n300), .ZN(new_n588));
  AOI211_X1 g402(.A(KEYINPUT97), .B(G902), .C1(new_n584), .C2(new_n586), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(G478), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n591), .A2(KEYINPUT15), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  OAI211_X1 g407(.A(new_n587), .B(new_n300), .C1(KEYINPUT15), .C2(new_n591), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n541), .A2(new_n595), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n365), .A2(new_n430), .A3(new_n487), .A4(new_n596), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n597), .B(G101), .ZN(G3));
  NAND2_X1  g412(.A1(new_n300), .A2(G478), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n587), .A2(KEYINPUT33), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT33), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n584), .A2(new_n601), .A3(new_n586), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n599), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n603), .B1(new_n590), .B2(new_n591), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n541), .A2(new_n605), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n606), .A2(new_n310), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n413), .A2(new_n300), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT98), .ZN(new_n609));
  INV_X1    g423(.A(G472), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  OAI211_X1 g426(.A(new_n413), .B(new_n300), .C1(new_n609), .C2(new_n610), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n612), .A2(new_n487), .A3(new_n613), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n614), .A2(new_n364), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n607), .A2(new_n615), .ZN(new_n616));
  XOR2_X1   g430(.A(KEYINPUT34), .B(G104), .Z(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(G6));
  OAI21_X1  g432(.A(new_n300), .B1(new_n518), .B2(new_n519), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT92), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n621), .A2(G475), .A3(new_n520), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n537), .A2(new_n538), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(KEYINPUT20), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n537), .A2(new_n528), .A3(new_n538), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n622), .A2(new_n595), .A3(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n310), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(new_n615), .ZN(new_n629));
  XOR2_X1   g443(.A(KEYINPUT35), .B(G107), .Z(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G9));
  NOR2_X1   g445(.A1(new_n469), .A2(KEYINPUT36), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n465), .B(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(new_n486), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n635), .B1(new_n476), .B2(new_n483), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  AND3_X1   g451(.A1(new_n612), .A2(new_n637), .A3(new_n613), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n365), .A2(new_n596), .A3(new_n638), .ZN(new_n639));
  XOR2_X1   g453(.A(KEYINPUT37), .B(G110), .Z(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G12));
  NOR2_X1   g455(.A1(new_n364), .A2(new_n636), .ZN(new_n642));
  AND2_X1   g456(.A1(new_n642), .A2(new_n430), .ZN(new_n643));
  INV_X1    g457(.A(G900), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n304), .A2(KEYINPUT99), .A3(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n299), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  AOI21_X1  g461(.A(KEYINPUT99), .B1(new_n304), .B2(new_n644), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n622), .A2(new_n595), .A3(new_n626), .A4(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n297), .A2(new_n308), .A3(new_n309), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n652), .A2(KEYINPUT100), .A3(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT100), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n656), .B1(new_n651), .B2(new_n653), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n643), .A2(new_n655), .A3(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(KEYINPUT101), .B(G128), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G30));
  XNOR2_X1  g474(.A(KEYINPUT103), .B(KEYINPUT39), .ZN(new_n661));
  XOR2_X1   g475(.A(new_n649), .B(new_n661), .Z(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n364), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(KEYINPUT40), .ZN(new_n665));
  AND3_X1   g479(.A1(new_n541), .A2(new_n595), .A3(new_n308), .ZN(new_n666));
  AND2_X1   g480(.A1(new_n666), .A2(new_n636), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n404), .A2(new_n389), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n300), .B1(new_n405), .B2(new_n401), .ZN(new_n669));
  OAI21_X1  g483(.A(G472), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(KEYINPUT102), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n416), .A2(new_n419), .A3(new_n429), .A4(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n297), .A2(new_n309), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT38), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n665), .A2(new_n667), .A3(new_n672), .A4(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G143), .ZN(G45));
  AOI211_X1 g491(.A(new_n649), .B(new_n604), .C1(new_n622), .C2(new_n626), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n643), .A2(new_n654), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G146), .ZN(G48));
  AND2_X1   g494(.A1(new_n430), .A2(new_n487), .ZN(new_n681));
  INV_X1    g495(.A(new_n354), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n318), .B1(new_n360), .B2(new_n344), .ZN(new_n683));
  OAI211_X1 g497(.A(new_n300), .B(new_n313), .C1(new_n682), .C2(new_n683), .ZN(new_n684));
  AOI21_X1  g498(.A(G902), .B1(new_n346), .B2(new_n354), .ZN(new_n685));
  OAI211_X1 g499(.A(new_n684), .B(new_n312), .C1(new_n685), .C2(new_n356), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n681), .A2(new_n607), .A3(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(KEYINPUT41), .B(G113), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n688), .B(new_n689), .ZN(G15));
  NAND4_X1  g504(.A1(new_n628), .A2(new_n430), .A3(new_n487), .A4(new_n687), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G116), .ZN(G18));
  NOR2_X1   g506(.A1(new_n653), .A2(new_n686), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n636), .A2(new_n306), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n693), .A2(new_n430), .A3(new_n596), .A4(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G119), .ZN(G21));
  AND3_X1   g510(.A1(new_n272), .A2(new_n295), .A3(new_n292), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n295), .B1(new_n272), .B2(new_n292), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(new_n487), .ZN(new_n700));
  XNOR2_X1  g514(.A(KEYINPUT104), .B(G472), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n702), .B1(new_n413), .B2(new_n300), .ZN(new_n703));
  INV_X1    g517(.A(new_n414), .ZN(new_n704));
  AOI22_X1  g518(.A1(new_n392), .A2(new_n391), .B1(new_n421), .B2(new_n389), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n410), .A2(KEYINPUT31), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n704), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  NOR3_X1   g521(.A1(new_n700), .A2(new_n703), .A3(new_n707), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n686), .A2(new_n306), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n666), .A2(new_n699), .A3(new_n708), .A4(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G122), .ZN(G24));
  INV_X1    g525(.A(KEYINPUT105), .ZN(new_n712));
  NOR3_X1   g526(.A1(new_n703), .A2(new_n636), .A3(new_n707), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n713), .A2(new_n699), .A3(new_n308), .A4(new_n687), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n541), .A2(new_n605), .A3(new_n650), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n712), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n693), .A2(new_n678), .A3(KEYINPUT105), .A4(new_n713), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  XOR2_X1   g532(.A(KEYINPUT106), .B(G125), .Z(new_n719));
  XNOR2_X1  g533(.A(new_n718), .B(new_n719), .ZN(G27));
  AOI21_X1  g534(.A(new_n604), .B1(new_n622), .B2(new_n626), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT108), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n358), .A2(G469), .A3(new_n361), .ZN(new_n723));
  NAND2_X1  g537(.A1(G469), .A2(G902), .ZN(new_n724));
  XOR2_X1   g538(.A(new_n724), .B(KEYINPUT107), .Z(new_n725));
  NAND2_X1  g539(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n722), .B1(new_n355), .B2(new_n726), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n684), .A2(KEYINPUT108), .A3(new_n725), .A4(new_n723), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(new_n312), .ZN(new_n730));
  INV_X1    g544(.A(new_n308), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(new_n732), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n733), .B1(new_n297), .B2(new_n309), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n721), .A2(new_n729), .A3(new_n734), .A4(new_n650), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n427), .A2(new_n415), .ZN(new_n736));
  AOI21_X1  g550(.A(KEYINPUT32), .B1(new_n413), .B2(new_n414), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n487), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  OAI21_X1  g552(.A(KEYINPUT42), .B1(new_n735), .B2(new_n738), .ZN(new_n739));
  AND2_X1   g553(.A1(new_n729), .A2(new_n734), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT42), .ZN(new_n741));
  AND4_X1   g555(.A1(new_n741), .A2(new_n541), .A3(new_n605), .A4(new_n650), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n681), .A2(new_n740), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n739), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(new_n327), .ZN(G33));
  NAND4_X1  g559(.A1(new_n430), .A2(new_n729), .A3(new_n734), .A4(new_n487), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n746), .A2(new_n651), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(new_n322), .ZN(G36));
  XNOR2_X1  g562(.A(new_n541), .B(KEYINPUT111), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n749), .A2(KEYINPUT43), .A3(new_n605), .ZN(new_n750));
  INV_X1    g564(.A(new_n541), .ZN(new_n751));
  AOI21_X1  g565(.A(KEYINPUT43), .B1(new_n751), .B2(new_n605), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT110), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  AOI211_X1 g568(.A(KEYINPUT110), .B(KEYINPUT43), .C1(new_n751), .C2(new_n605), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n750), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n636), .B1(new_n612), .B2(new_n613), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT44), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n756), .A2(KEYINPUT44), .A3(new_n757), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT45), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n362), .A2(new_n762), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n358), .A2(KEYINPUT45), .A3(new_n361), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n763), .A2(G469), .A3(new_n764), .ZN(new_n765));
  AND2_X1   g579(.A1(new_n765), .A2(new_n725), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT109), .ZN(new_n767));
  OR3_X1    g581(.A1(new_n766), .A2(new_n767), .A3(KEYINPUT46), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n767), .B1(new_n766), .B2(KEYINPUT46), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n355), .B1(new_n766), .B2(KEYINPUT46), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n768), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(new_n312), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n673), .A2(new_n308), .ZN(new_n773));
  NOR3_X1   g587(.A1(new_n772), .A2(new_n663), .A3(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n760), .A2(new_n761), .A3(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G137), .ZN(G39));
  NOR4_X1   g590(.A1(new_n715), .A2(new_n773), .A3(new_n430), .A4(new_n487), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT113), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n777), .B(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(KEYINPUT112), .B(KEYINPUT47), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n771), .A2(new_n312), .A3(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(new_n780), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n772), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n779), .A2(new_n781), .A3(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G140), .ZN(G42));
  INV_X1    g599(.A(new_n675), .ZN(new_n786));
  INV_X1    g600(.A(new_n672), .ZN(new_n787));
  NOR3_X1   g601(.A1(new_n700), .A2(new_n604), .A3(new_n733), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n684), .B1(new_n685), .B2(new_n356), .ZN(new_n789));
  OR2_X1    g603(.A1(new_n789), .A2(KEYINPUT49), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(KEYINPUT49), .ZN(new_n791));
  AND3_X1   g605(.A1(new_n788), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n786), .A2(new_n787), .A3(new_n749), .A4(new_n792), .ZN(new_n793));
  AND2_X1   g607(.A1(new_n756), .A2(new_n299), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n699), .A2(new_n789), .A3(new_n733), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n794), .A2(new_n713), .A3(new_n795), .ZN(new_n796));
  AND4_X1   g610(.A1(new_n487), .A2(new_n795), .A3(new_n787), .A4(new_n299), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n797), .A2(new_n751), .A3(new_n604), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n699), .A2(new_n731), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n794), .A2(new_n708), .A3(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(new_n789), .ZN(new_n801));
  AOI22_X1  g615(.A1(new_n783), .A2(new_n781), .B1(new_n730), .B2(new_n801), .ZN(new_n802));
  OAI211_X1 g616(.A(new_n796), .B(new_n798), .C1(new_n800), .C2(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT51), .ZN(new_n804));
  NOR3_X1   g618(.A1(new_n675), .A2(new_n308), .A3(new_n686), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n756), .A2(new_n299), .A3(new_n708), .A4(new_n805), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(KEYINPUT50), .ZN(new_n807));
  OR3_X1    g621(.A1(new_n803), .A2(new_n804), .A3(new_n807), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n804), .B1(new_n803), .B2(new_n807), .ZN(new_n809));
  INV_X1    g623(.A(new_n738), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n794), .A2(new_n810), .A3(new_n795), .ZN(new_n811));
  XOR2_X1   g625(.A(KEYINPUT119), .B(KEYINPUT48), .Z(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n794), .A2(new_n693), .A3(new_n708), .ZN(new_n814));
  AOI211_X1 g628(.A(new_n298), .B(G953), .C1(new_n797), .C2(new_n721), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n813), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n811), .A2(new_n812), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n808), .A2(new_n809), .A3(new_n818), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n651), .A2(new_n653), .A3(new_n656), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n642), .A2(new_n430), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  AOI22_X1  g636(.A1(new_n822), .A2(new_n657), .B1(new_n716), .B2(new_n717), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT52), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT116), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n312), .B1(new_n649), .B2(new_n825), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n826), .B1(new_n825), .B2(new_n649), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n729), .A2(new_n636), .A3(new_n827), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n828), .A2(new_n699), .A3(new_n672), .A4(new_n666), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n823), .A2(new_n824), .A3(new_n679), .A4(new_n829), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n688), .A2(new_n691), .A3(new_n695), .A4(new_n710), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT53), .ZN(new_n832));
  NOR3_X1   g646(.A1(new_n831), .A2(new_n744), .A3(new_n832), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n718), .A2(new_n658), .A3(new_n679), .A4(new_n829), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n834), .A2(KEYINPUT52), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n718), .A2(new_n658), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(KEYINPUT52), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n830), .A2(new_n833), .A3(new_n835), .A4(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(new_n310), .ZN(new_n839));
  INV_X1    g653(.A(new_n627), .ZN(new_n840));
  OAI211_X1 g654(.A(new_n615), .B(new_n839), .C1(new_n721), .C2(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n841), .A2(new_n597), .A3(new_n639), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT114), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n841), .A2(new_n597), .A3(KEYINPUT114), .A4(new_n639), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n541), .A2(new_n595), .A3(new_n649), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(new_n799), .ZN(new_n848));
  OAI22_X1  g662(.A1(new_n848), .A2(new_n821), .B1(new_n746), .B2(new_n651), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n740), .A2(new_n678), .A3(new_n713), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT115), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n740), .A2(KEYINPUT115), .A3(new_n678), .A4(new_n713), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n849), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n846), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(KEYINPUT117), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT117), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n846), .A2(new_n857), .A3(new_n854), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n838), .B1(new_n856), .B2(new_n858), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n831), .A2(new_n744), .ZN(new_n860));
  AND3_X1   g674(.A1(new_n846), .A2(new_n860), .A3(new_n854), .ZN(new_n861));
  XNOR2_X1  g675(.A(new_n834), .B(new_n824), .ZN(new_n862));
  AOI21_X1  g676(.A(KEYINPUT53), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n859), .A2(new_n863), .A3(KEYINPUT54), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT54), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n837), .A2(new_n832), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n861), .A2(new_n862), .A3(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n846), .A2(new_n860), .A3(new_n854), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n830), .A2(new_n835), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n832), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n865), .B1(new_n867), .B2(new_n870), .ZN(new_n871));
  OAI21_X1  g685(.A(KEYINPUT118), .B1(new_n864), .B2(new_n871), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n861), .A2(new_n862), .A3(new_n866), .ZN(new_n873));
  OAI21_X1  g687(.A(KEYINPUT54), .B1(new_n873), .B2(new_n863), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT118), .ZN(new_n875));
  AND2_X1   g689(.A1(new_n833), .A2(new_n837), .ZN(new_n876));
  AND3_X1   g690(.A1(new_n846), .A2(new_n857), .A3(new_n854), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n857), .B1(new_n846), .B2(new_n854), .ZN(new_n878));
  OAI211_X1 g692(.A(new_n862), .B(new_n876), .C1(new_n877), .C2(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n879), .A2(new_n865), .A3(new_n870), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n874), .A2(new_n875), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n819), .B1(new_n872), .B2(new_n881), .ZN(new_n882));
  NOR2_X1   g696(.A1(G952), .A2(G953), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n793), .B1(new_n882), .B2(new_n883), .ZN(G75));
  AOI21_X1  g698(.A(new_n300), .B1(new_n879), .B2(new_n870), .ZN(new_n885));
  AOI21_X1  g699(.A(KEYINPUT56), .B1(new_n885), .B2(new_n295), .ZN(new_n886));
  AND2_X1   g700(.A1(new_n240), .A2(new_n267), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n887), .B(new_n265), .ZN(new_n888));
  XOR2_X1   g702(.A(new_n888), .B(KEYINPUT55), .Z(new_n889));
  NOR2_X1   g703(.A1(new_n886), .A2(new_n889), .ZN(new_n890));
  XOR2_X1   g704(.A(KEYINPUT120), .B(KEYINPUT56), .Z(new_n891));
  NAND2_X1  g705(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n892), .B1(new_n885), .B2(new_n295), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n303), .A2(G952), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n890), .A2(new_n893), .A3(new_n894), .ZN(G51));
  XOR2_X1   g709(.A(new_n725), .B(KEYINPUT57), .Z(new_n896));
  AOI21_X1  g710(.A(new_n865), .B1(new_n879), .B2(new_n870), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n896), .B1(new_n864), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n898), .B1(new_n683), .B2(new_n682), .ZN(new_n899));
  INV_X1    g713(.A(new_n765), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n885), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n894), .B1(new_n899), .B2(new_n901), .ZN(G54));
  NAND3_X1  g716(.A1(new_n885), .A2(KEYINPUT58), .A3(G475), .ZN(new_n903));
  INV_X1    g717(.A(new_n537), .ZN(new_n904));
  AND2_X1   g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n903), .A2(new_n904), .ZN(new_n906));
  NOR3_X1   g720(.A1(new_n905), .A2(new_n906), .A3(new_n894), .ZN(G60));
  NAND2_X1  g721(.A1(new_n600), .A2(new_n602), .ZN(new_n908));
  NAND2_X1  g722(.A1(G478), .A2(G902), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n909), .B(KEYINPUT59), .ZN(new_n910));
  OAI211_X1 g724(.A(new_n908), .B(new_n910), .C1(new_n864), .C2(new_n897), .ZN(new_n911));
  INV_X1    g725(.A(new_n894), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(new_n908), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n872), .A2(new_n881), .A3(new_n910), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n913), .B1(new_n914), .B2(new_n915), .ZN(G63));
  NAND2_X1  g730(.A1(G217), .A2(G902), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(KEYINPUT60), .ZN(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n633), .B(KEYINPUT122), .ZN(new_n920));
  OAI211_X1 g734(.A(new_n919), .B(new_n920), .C1(new_n859), .C2(new_n863), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n918), .B1(new_n879), .B2(new_n870), .ZN(new_n922));
  OAI211_X1 g736(.A(new_n921), .B(new_n912), .C1(new_n484), .C2(new_n922), .ZN(new_n923));
  AND3_X1   g737(.A1(new_n923), .A2(KEYINPUT121), .A3(KEYINPUT61), .ZN(new_n924));
  AOI21_X1  g738(.A(KEYINPUT61), .B1(new_n923), .B2(KEYINPUT121), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n924), .A2(new_n925), .ZN(G66));
  INV_X1    g740(.A(G224), .ZN(new_n927));
  OAI21_X1  g741(.A(G953), .B1(new_n305), .B2(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(new_n831), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n846), .A2(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(new_n303), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n928), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(G898), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n887), .B1(new_n934), .B2(new_n932), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n933), .B(new_n935), .Z(G69));
  INV_X1    g750(.A(G227), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n407), .A2(new_n408), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(KEYINPUT123), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n939), .B(new_n533), .ZN(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  OAI221_X1 g755(.A(new_n932), .B1(new_n937), .B2(new_n644), .C1(new_n941), .C2(KEYINPUT125), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n606), .A2(new_n627), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n681), .A2(new_n664), .A3(new_n799), .A4(new_n943), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n944), .B(KEYINPUT124), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n775), .A2(new_n784), .A3(new_n945), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n823), .A2(new_n676), .A3(new_n679), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n947), .B(KEYINPUT62), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n303), .B1(new_n946), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(new_n941), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT126), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n932), .A2(G900), .ZN(new_n952));
  AND2_X1   g766(.A1(new_n823), .A2(new_n679), .ZN(new_n953));
  AND3_X1   g767(.A1(new_n810), .A2(new_n699), .A3(new_n666), .ZN(new_n954));
  AND4_X1   g768(.A1(new_n312), .A2(new_n954), .A3(new_n771), .A4(new_n662), .ZN(new_n955));
  NOR3_X1   g769(.A1(new_n955), .A2(new_n744), .A3(new_n747), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n775), .A2(new_n784), .A3(new_n953), .A4(new_n956), .ZN(new_n957));
  OAI211_X1 g771(.A(new_n940), .B(new_n952), .C1(new_n957), .C2(new_n932), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n950), .A2(new_n951), .A3(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n951), .B1(new_n950), .B2(new_n958), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n942), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(new_n961), .ZN(new_n963));
  INV_X1    g777(.A(new_n942), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n963), .A2(new_n959), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n962), .A2(new_n965), .ZN(G72));
  XNOR2_X1  g780(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n610), .A2(new_n300), .ZN(new_n968));
  XOR2_X1   g782(.A(new_n967), .B(new_n968), .Z(new_n969));
  INV_X1    g783(.A(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT62), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n947), .B(new_n971), .ZN(new_n972));
  NAND4_X1  g786(.A1(new_n972), .A2(new_n775), .A3(new_n784), .A4(new_n945), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n970), .B1(new_n973), .B2(new_n930), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n974), .A2(new_n668), .ZN(new_n975));
  NOR3_X1   g789(.A1(new_n384), .A2(new_n405), .A3(new_n390), .ZN(new_n976));
  NOR3_X1   g790(.A1(new_n668), .A2(new_n976), .A3(new_n969), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n977), .B1(new_n873), .B2(new_n863), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n970), .B1(new_n957), .B2(new_n930), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n894), .B1(new_n979), .B2(new_n976), .ZN(new_n980));
  AND3_X1   g794(.A1(new_n975), .A2(new_n978), .A3(new_n980), .ZN(G57));
endmodule


