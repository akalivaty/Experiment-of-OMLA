//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 1 0 1 1 1 0 0 0 0 0 0 0 1 1 0 1 0 1 0 1 0 1 1 0 1 1 1 0 1 1 0 0 1 1 0 0 0 1 0 1 0 0 1 1 1 0 0 0 1 0 1 0 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:15 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1212, new_n1213,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1269,
    new_n1270, new_n1271, new_n1272, new_n1273;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  NAND2_X1  g0008(.A1(G77), .A2(G244), .ZN(new_n209));
  INV_X1    g0009(.A(G58), .ZN(new_n210));
  INV_X1    g0010(.A(G232), .ZN(new_n211));
  OAI21_X1  g0011(.A(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  AOI21_X1  g0012(.A(new_n212), .B1(G87), .B2(G250), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G107), .A2(G264), .ZN(new_n215));
  AND3_X1   g0015(.A1(new_n213), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  AND2_X1   g0016(.A1(KEYINPUT65), .A2(G68), .ZN(new_n217));
  NOR2_X1   g0017(.A1(KEYINPUT65), .A2(G68), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n219), .A2(G238), .ZN(new_n220));
  INV_X1    g0020(.A(G116), .ZN(new_n221));
  INV_X1    g0021(.A(G270), .ZN(new_n222));
  OAI211_X1 g0022(.A(new_n216), .B(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G20), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  XOR2_X1   g0025(.A(new_n225), .B(KEYINPUT1), .Z(new_n226));
  INV_X1    g0026(.A(new_n201), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n227), .A2(G50), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT64), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  INV_X1    g0030(.A(G20), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n224), .A2(G13), .ZN(new_n233));
  OR2_X1    g0033(.A1(G257), .A2(G264), .ZN(new_n234));
  AND3_X1   g0034(.A1(new_n233), .A2(G250), .A3(new_n234), .ZN(new_n235));
  AOI22_X1  g0035(.A1(new_n229), .A2(new_n232), .B1(KEYINPUT0), .B2(new_n235), .ZN(new_n236));
  OAI211_X1 g0036(.A(new_n226), .B(new_n236), .C1(KEYINPUT0), .C2(new_n235), .ZN(new_n237));
  INV_X1    g0037(.A(new_n237), .ZN(G361));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(new_n211), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT2), .ZN(new_n241));
  INV_X1    g0041(.A(G226), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G250), .B(G257), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT66), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(G264), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(new_n222), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n243), .B(new_n247), .ZN(G358));
  XNOR2_X1  g0048(.A(G50), .B(G68), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(G58), .ZN(new_n250));
  INV_X1    g0050(.A(G77), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(G87), .B(G97), .ZN(new_n253));
  XNOR2_X1  g0053(.A(G107), .B(G116), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n253), .B(new_n254), .ZN(new_n255));
  XOR2_X1   g0055(.A(new_n252), .B(new_n255), .Z(G351));
  NAND2_X1  g0056(.A1(new_n203), .A2(G20), .ZN(new_n257));
  INV_X1    g0057(.A(G150), .ZN(new_n258));
  NOR2_X1   g0058(.A1(G20), .A2(G33), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  XNOR2_X1  g0060(.A(KEYINPUT8), .B(G58), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT68), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n210), .A2(KEYINPUT68), .A3(KEYINPUT8), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n231), .A2(G33), .ZN(new_n266));
  OAI221_X1 g0066(.A(new_n257), .B1(new_n258), .B2(new_n260), .C1(new_n265), .C2(new_n266), .ZN(new_n267));
  NAND3_X1  g0067(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(new_n230), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G13), .ZN(new_n271));
  NOR3_X1   g0071(.A1(new_n271), .A2(new_n231), .A3(G1), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n272), .A2(new_n269), .ZN(new_n273));
  XNOR2_X1  g0073(.A(new_n273), .B(KEYINPUT69), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n231), .A2(G1), .ZN(new_n275));
  XNOR2_X1  g0075(.A(new_n275), .B(KEYINPUT70), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G50), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(KEYINPUT71), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT71), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n276), .A2(new_n279), .A3(G50), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n274), .A2(new_n278), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n272), .A2(new_n202), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n270), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  OR2_X1    g0084(.A1(new_n284), .A2(KEYINPUT9), .ZN(new_n285));
  INV_X1    g0085(.A(G33), .ZN(new_n286));
  INV_X1    g0086(.A(G41), .ZN(new_n287));
  OAI211_X1 g0087(.A(G1), .B(G13), .C1(new_n286), .C2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  AND2_X1   g0089(.A1(KEYINPUT3), .A2(G33), .ZN(new_n290));
  NOR2_X1   g0090(.A1(KEYINPUT3), .A2(G33), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G1698), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(G223), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT3), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(new_n286), .ZN(new_n298));
  NAND2_X1  g0098(.A1(KEYINPUT3), .A2(G33), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(new_n293), .ZN(new_n301));
  INV_X1    g0101(.A(G222), .ZN(new_n302));
  OAI22_X1  g0102(.A1(new_n301), .A2(new_n302), .B1(new_n251), .B2(new_n300), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n289), .B1(new_n296), .B2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G1), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n305), .B1(G41), .B2(G45), .ZN(new_n306));
  INV_X1    g0106(.A(G274), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  AND2_X1   g0109(.A1(new_n288), .A2(new_n306), .ZN(new_n310));
  OR2_X1    g0110(.A1(KEYINPUT67), .A2(G226), .ZN(new_n311));
  NAND2_X1  g0111(.A1(KEYINPUT67), .A2(G226), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n310), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n304), .A2(new_n309), .A3(new_n313), .ZN(new_n314));
  AOI22_X1  g0114(.A1(new_n284), .A2(KEYINPUT9), .B1(G200), .B2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(G190), .ZN(new_n316));
  OR2_X1    g0116(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n285), .A2(new_n315), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(KEYINPUT10), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT10), .ZN(new_n320));
  NAND4_X1  g0120(.A1(new_n285), .A2(new_n315), .A3(new_n320), .A4(new_n317), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  OR2_X1    g0122(.A1(new_n314), .A2(G179), .ZN(new_n323));
  INV_X1    g0123(.A(G169), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n314), .A2(new_n324), .ZN(new_n325));
  AND3_X1   g0125(.A1(new_n323), .A2(new_n283), .A3(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n322), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n300), .A2(G232), .A3(G1698), .ZN(new_n329));
  NAND2_X1  g0129(.A1(G33), .A2(G97), .ZN(new_n330));
  OAI211_X1 g0130(.A(new_n329), .B(new_n330), .C1(new_n301), .C2(new_n242), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n308), .B1(new_n331), .B2(new_n289), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT13), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n310), .A2(G238), .ZN(new_n334));
  AND3_X1   g0134(.A1(new_n332), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n333), .B1(new_n332), .B2(new_n334), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  OAI22_X1  g0137(.A1(new_n337), .A2(new_n324), .B1(KEYINPUT75), .B2(KEYINPUT14), .ZN(new_n338));
  NAND2_X1  g0138(.A1(KEYINPUT75), .A2(KEYINPUT14), .ZN(new_n339));
  NOR2_X1   g0139(.A1(KEYINPUT75), .A2(KEYINPUT14), .ZN(new_n340));
  OAI211_X1 g0140(.A(G169), .B(new_n340), .C1(new_n335), .C2(new_n336), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n337), .A2(G179), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n338), .A2(new_n339), .A3(new_n341), .A4(new_n342), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n276), .A2(G68), .A3(new_n273), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT12), .ZN(new_n345));
  INV_X1    g0145(.A(G68), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n272), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n272), .ZN(new_n348));
  OAI22_X1  g0148(.A1(new_n348), .A2(new_n219), .B1(KEYINPUT74), .B2(KEYINPUT12), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT74), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n350), .A2(new_n345), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n347), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n259), .A2(G50), .ZN(new_n353));
  XNOR2_X1  g0153(.A(new_n353), .B(KEYINPUT73), .ZN(new_n354));
  OAI221_X1 g0154(.A(new_n354), .B1(new_n231), .B2(new_n219), .C1(new_n251), .C2(new_n266), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT11), .ZN(new_n356));
  AND3_X1   g0156(.A1(new_n355), .A2(new_n356), .A3(new_n269), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n356), .B1(new_n355), .B2(new_n269), .ZN(new_n358));
  OAI211_X1 g0158(.A(new_n344), .B(new_n352), .C1(new_n357), .C2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n343), .A2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(new_n359), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n337), .A2(G190), .ZN(new_n362));
  INV_X1    g0162(.A(G200), .ZN(new_n363));
  OAI211_X1 g0163(.A(new_n361), .B(new_n362), .C1(new_n337), .C2(new_n363), .ZN(new_n364));
  OAI22_X1  g0164(.A1(new_n261), .A2(new_n260), .B1(new_n231), .B2(new_n251), .ZN(new_n365));
  XOR2_X1   g0165(.A(new_n365), .B(KEYINPUT72), .Z(new_n366));
  XNOR2_X1  g0166(.A(KEYINPUT15), .B(G87), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n366), .B1(new_n266), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(new_n269), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n272), .A2(new_n251), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n276), .A2(new_n273), .ZN(new_n371));
  OAI211_X1 g0171(.A(new_n369), .B(new_n370), .C1(new_n251), .C2(new_n371), .ZN(new_n372));
  AOI22_X1  g0172(.A1(new_n294), .A2(G238), .B1(G107), .B2(new_n292), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n300), .A2(G232), .A3(new_n293), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(new_n289), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n310), .A2(G244), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n376), .A2(new_n309), .A3(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(new_n378), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n379), .A2(new_n363), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n372), .A2(new_n380), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n381), .B1(new_n316), .B2(new_n378), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n360), .A2(new_n364), .A3(new_n382), .ZN(new_n383));
  AND3_X1   g0183(.A1(new_n276), .A2(new_n264), .A3(new_n263), .ZN(new_n384));
  AOI22_X1  g0184(.A1(new_n274), .A2(new_n384), .B1(new_n272), .B2(new_n265), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n298), .A2(new_n231), .A3(new_n299), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT7), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n298), .A2(KEYINPUT7), .A3(new_n231), .A4(new_n299), .ZN(new_n389));
  AOI21_X1  g0189(.A(KEYINPUT76), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(KEYINPUT7), .B1(new_n292), .B2(new_n231), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT76), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n219), .B1(new_n390), .B2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(G159), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n260), .A2(new_n395), .ZN(new_n396));
  OR2_X1    g0196(.A1(KEYINPUT65), .A2(G68), .ZN(new_n397));
  NAND2_X1  g0197(.A1(KEYINPUT65), .A2(G68), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n397), .A2(G58), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(new_n227), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n396), .B1(new_n400), .B2(G20), .ZN(new_n401));
  AOI21_X1  g0201(.A(KEYINPUT16), .B1(new_n394), .B2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(new_n389), .ZN(new_n403));
  OAI21_X1  g0203(.A(G68), .B1(new_n391), .B2(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n404), .A2(new_n401), .A3(KEYINPUT16), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(new_n269), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n385), .B1(new_n402), .B2(new_n406), .ZN(new_n407));
  OAI211_X1 g0207(.A(G226), .B(G1698), .C1(new_n290), .C2(new_n291), .ZN(new_n408));
  OAI211_X1 g0208(.A(G223), .B(new_n293), .C1(new_n290), .C2(new_n291), .ZN(new_n409));
  INV_X1    g0209(.A(G87), .ZN(new_n410));
  OAI211_X1 g0210(.A(new_n408), .B(new_n409), .C1(new_n286), .C2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(new_n289), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n310), .A2(G232), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n412), .A2(new_n309), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(G169), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n412), .A2(G179), .A3(new_n413), .A4(new_n309), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n415), .A2(KEYINPUT77), .A3(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  AOI21_X1  g0218(.A(KEYINPUT77), .B1(new_n415), .B2(new_n416), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n407), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT18), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  OAI211_X1 g0222(.A(KEYINPUT18), .B(new_n407), .C1(new_n418), .C2(new_n419), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  AND3_X1   g0224(.A1(new_n412), .A2(new_n309), .A3(new_n413), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(G190), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n426), .B(new_n385), .C1(new_n402), .C2(new_n406), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n425), .A2(new_n363), .ZN(new_n428));
  OAI21_X1  g0228(.A(KEYINPUT17), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n274), .A2(new_n384), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n265), .A2(new_n272), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT16), .ZN(new_n433));
  INV_X1    g0233(.A(new_n219), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n392), .B1(new_n391), .B2(new_n403), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n388), .A2(KEYINPUT76), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n434), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n396), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n201), .B1(new_n219), .B2(G58), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n438), .B1(new_n439), .B2(new_n231), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n433), .B1(new_n437), .B2(new_n440), .ZN(new_n441));
  AND2_X1   g0241(.A1(new_n405), .A2(new_n269), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n432), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT17), .ZN(new_n444));
  INV_X1    g0244(.A(new_n428), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n443), .A2(new_n444), .A3(new_n445), .A4(new_n426), .ZN(new_n446));
  AND3_X1   g0246(.A1(new_n429), .A2(KEYINPUT78), .A3(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(KEYINPUT78), .B1(new_n429), .B2(new_n446), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n424), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n378), .A2(new_n324), .ZN(new_n450));
  INV_X1    g0250(.A(G179), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n379), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n372), .A2(new_n450), .A3(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g0254(.A1(new_n328), .A2(new_n383), .A3(new_n449), .A4(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n272), .A2(new_n206), .ZN(new_n456));
  XNOR2_X1  g0256(.A(new_n456), .B(KEYINPUT25), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n273), .B1(G1), .B2(new_n286), .ZN(new_n459));
  AOI21_X1  g0259(.A(G20), .B1(new_n298), .B2(new_n299), .ZN(new_n460));
  NOR2_X1   g0260(.A1(KEYINPUT92), .A2(KEYINPUT22), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(KEYINPUT92), .A2(KEYINPUT22), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n460), .A2(G87), .A3(new_n462), .A4(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n231), .A2(G33), .A3(G116), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n231), .A2(G107), .ZN(new_n466));
  XNOR2_X1  g0266(.A(new_n466), .B(KEYINPUT23), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n231), .B(G87), .C1(new_n290), .C2(new_n291), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(new_n461), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n464), .A2(new_n465), .A3(new_n467), .A4(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT24), .ZN(new_n471));
  XNOR2_X1  g0271(.A(new_n470), .B(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(new_n269), .ZN(new_n473));
  OAI221_X1 g0273(.A(new_n458), .B1(new_n206), .B2(new_n459), .C1(new_n472), .C2(new_n473), .ZN(new_n474));
  OAI211_X1 g0274(.A(G257), .B(G1698), .C1(new_n290), .C2(new_n291), .ZN(new_n475));
  OAI211_X1 g0275(.A(G250), .B(new_n293), .C1(new_n290), .C2(new_n291), .ZN(new_n476));
  NAND2_X1  g0276(.A1(G33), .A2(G294), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n475), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(new_n289), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n305), .B(G45), .C1(new_n287), .C2(KEYINPUT5), .ZN(new_n480));
  AND2_X1   g0280(.A1(new_n287), .A2(KEYINPUT5), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n288), .B(G264), .C1(new_n480), .C2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n479), .A2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT93), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n479), .A2(KEYINPUT93), .A3(new_n482), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(G45), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n488), .A2(G1), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n489), .B(KEYINPUT83), .C1(KEYINPUT5), .C2(new_n287), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n481), .A2(new_n307), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT83), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n480), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n490), .A2(new_n491), .A3(new_n493), .A4(new_n288), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n487), .A2(G179), .A3(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n479), .A2(new_n482), .A3(new_n494), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(G169), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n474), .A2(new_n498), .ZN(new_n499));
  AND2_X1   g0299(.A1(new_n464), .A2(new_n469), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n500), .A2(new_n471), .A3(new_n465), .A4(new_n467), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n470), .A2(KEYINPUT24), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n473), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n459), .A2(new_n206), .ZN(new_n504));
  NOR3_X1   g0304(.A1(new_n503), .A2(new_n504), .A3(new_n457), .ZN(new_n505));
  INV_X1    g0305(.A(new_n494), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n506), .B1(new_n485), .B2(new_n486), .ZN(new_n507));
  OAI22_X1  g0307(.A1(new_n507), .A2(G200), .B1(G190), .B2(new_n496), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n505), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n460), .A2(G68), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT19), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n511), .B1(new_n266), .B2(new_n205), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n231), .B1(new_n330), .B2(new_n511), .ZN(new_n513));
  XNOR2_X1  g0313(.A(new_n513), .B(KEYINPUT87), .ZN(new_n514));
  NOR3_X1   g0314(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n510), .B(new_n512), .C1(new_n514), .C2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(new_n269), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n367), .A2(new_n272), .ZN(new_n518));
  OR2_X1    g0318(.A1(new_n459), .A2(new_n410), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  OAI211_X1 g0320(.A(G244), .B(G1698), .C1(new_n290), .C2(new_n291), .ZN(new_n521));
  OAI211_X1 g0321(.A(G238), .B(new_n293), .C1(new_n290), .C2(new_n291), .ZN(new_n522));
  NAND2_X1  g0322(.A1(G33), .A2(G116), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(KEYINPUT85), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT85), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n521), .A2(new_n522), .A3(new_n526), .A4(new_n523), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n525), .A2(new_n289), .A3(new_n527), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n289), .A2(new_n489), .ZN(new_n529));
  AOI22_X1  g0329(.A1(new_n529), .A2(G250), .B1(G274), .B2(new_n489), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n528), .A2(G190), .A3(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT89), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n528), .A2(KEYINPUT89), .A3(G190), .A4(new_n530), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n520), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n528), .A2(new_n530), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(G200), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n528), .A2(new_n451), .A3(new_n530), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT86), .ZN(new_n540));
  OR2_X1    g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  XNOR2_X1  g0341(.A(new_n367), .B(KEYINPUT88), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n517), .B(new_n518), .C1(new_n459), .C2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n536), .A2(new_n324), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n539), .A2(new_n540), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n541), .A2(new_n543), .A3(new_n544), .A4(new_n545), .ZN(new_n546));
  AND4_X1   g0346(.A1(new_n499), .A2(new_n509), .A3(new_n538), .A4(new_n546), .ZN(new_n547));
  MUX2_X1   g0347(.A(new_n348), .B(new_n459), .S(G97), .Z(new_n548));
  OAI21_X1  g0348(.A(G107), .B1(new_n390), .B2(new_n393), .ZN(new_n549));
  NAND2_X1  g0349(.A1(G97), .A2(G107), .ZN(new_n550));
  AOI21_X1  g0350(.A(KEYINPUT6), .B1(new_n207), .B2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT6), .ZN(new_n552));
  NOR3_X1   g0352(.A1(new_n552), .A2(new_n205), .A3(G107), .ZN(new_n553));
  OAI21_X1  g0353(.A(G20), .B1(new_n551), .B2(new_n553), .ZN(new_n554));
  OR3_X1    g0354(.A1(new_n260), .A2(KEYINPUT79), .A3(new_n251), .ZN(new_n555));
  OAI21_X1  g0355(.A(KEYINPUT79), .B1(new_n260), .B2(new_n251), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT80), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n554), .A2(KEYINPUT80), .A3(new_n555), .A4(new_n556), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n549), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT81), .ZN(new_n562));
  AND3_X1   g0362(.A1(new_n561), .A2(new_n562), .A3(new_n269), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n562), .B1(new_n561), .B2(new_n269), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n548), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT84), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  OAI211_X1 g0367(.A(G244), .B(new_n293), .C1(new_n290), .C2(new_n291), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(KEYINPUT82), .ZN(new_n569));
  OR2_X1    g0369(.A1(new_n569), .A2(KEYINPUT4), .ZN(new_n570));
  NAND2_X1  g0370(.A1(G33), .A2(G283), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n294), .A2(G250), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n569), .A2(KEYINPUT4), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n570), .A2(new_n571), .A3(new_n572), .A4(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n506), .B1(new_n574), .B2(new_n289), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n288), .B(G257), .C1(new_n480), .C2(new_n481), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n575), .A2(G179), .A3(new_n576), .ZN(new_n577));
  AND2_X1   g0377(.A1(new_n575), .A2(new_n576), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n577), .B1(new_n578), .B2(new_n324), .ZN(new_n579));
  OAI211_X1 g0379(.A(KEYINPUT84), .B(new_n548), .C1(new_n563), .C2(new_n564), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n567), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n292), .A2(G303), .ZN(new_n582));
  OAI211_X1 g0382(.A(G257), .B(new_n293), .C1(new_n290), .C2(new_n291), .ZN(new_n583));
  OAI211_X1 g0383(.A(G264), .B(G1698), .C1(new_n290), .C2(new_n291), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT90), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n582), .A2(KEYINPUT90), .A3(new_n583), .A4(new_n584), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n587), .A2(new_n289), .A3(new_n588), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n273), .B(G116), .C1(G1), .C2(new_n286), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n272), .A2(new_n221), .ZN(new_n591));
  AOI22_X1  g0391(.A1(new_n268), .A2(new_n230), .B1(G20), .B2(new_n221), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n571), .B(new_n231), .C1(G33), .C2(new_n205), .ZN(new_n593));
  AOI21_X1  g0393(.A(KEYINPUT20), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  AND3_X1   g0394(.A1(new_n592), .A2(KEYINPUT20), .A3(new_n593), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n590), .B(new_n591), .C1(new_n594), .C2(new_n595), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n288), .B(G270), .C1(new_n480), .C2(new_n481), .ZN(new_n597));
  AND2_X1   g0397(.A1(new_n494), .A2(new_n597), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n589), .A2(new_n596), .A3(G179), .A4(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT91), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n589), .A2(new_n598), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n602), .A2(KEYINPUT21), .A3(G169), .A4(new_n596), .ZN(new_n603));
  AND2_X1   g0403(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n602), .A2(G169), .A3(new_n596), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT21), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  OR2_X1    g0407(.A1(new_n599), .A2(new_n600), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n604), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n602), .A2(new_n316), .ZN(new_n610));
  AOI211_X1 g0410(.A(new_n596), .B(new_n610), .C1(G200), .C2(new_n602), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  OR2_X1    g0412(.A1(new_n563), .A2(new_n564), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n575), .A2(new_n576), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(G200), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n578), .A2(G190), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n613), .A2(new_n548), .A3(new_n615), .A4(new_n616), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n547), .A2(new_n581), .A3(new_n612), .A4(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(new_n618), .ZN(new_n619));
  AND2_X1   g0419(.A1(new_n455), .A2(new_n619), .ZN(G372));
  NAND3_X1  g0420(.A1(new_n543), .A2(new_n544), .A3(new_n539), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n533), .A2(new_n534), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT94), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n537), .A2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n520), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n536), .A2(KEYINPUT94), .A3(G200), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n622), .A2(new_n624), .A3(new_n625), .A4(new_n626), .ZN(new_n627));
  AND3_X1   g0427(.A1(new_n509), .A2(new_n621), .A3(new_n627), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n499), .A2(new_n607), .A3(new_n608), .A4(new_n604), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n581), .A2(new_n628), .A3(new_n617), .A4(new_n629), .ZN(new_n630));
  AND2_X1   g0430(.A1(new_n543), .A2(new_n544), .ZN(new_n631));
  XNOR2_X1  g0431(.A(new_n539), .B(KEYINPUT86), .ZN(new_n632));
  AOI22_X1  g0432(.A1(new_n631), .A2(new_n632), .B1(new_n535), .B2(new_n537), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n633), .A2(new_n567), .A3(new_n579), .A4(new_n580), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(KEYINPUT26), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n579), .A2(new_n565), .A3(new_n627), .A4(new_n621), .ZN(new_n636));
  OR2_X1    g0436(.A1(new_n636), .A2(KEYINPUT26), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n630), .A2(new_n635), .A3(new_n637), .A4(new_n621), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n455), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n454), .A2(new_n364), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n360), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n429), .A2(new_n446), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT78), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n429), .A2(KEYINPUT78), .A3(new_n446), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n641), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n415), .A2(new_n416), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n407), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(new_n421), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n407), .A2(KEYINPUT18), .A3(new_n648), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n647), .A2(new_n652), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n326), .B1(new_n653), .B2(new_n322), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n639), .A2(new_n654), .ZN(G369));
  NOR2_X1   g0455(.A1(new_n271), .A2(G20), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(new_n305), .ZN(new_n657));
  OR2_X1    g0457(.A1(new_n657), .A2(KEYINPUT27), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(KEYINPUT27), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n658), .A2(G213), .A3(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(G343), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n596), .A2(new_n662), .ZN(new_n663));
  MUX2_X1   g0463(.A(new_n609), .B(new_n612), .S(new_n663), .Z(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(G330), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n474), .A2(new_n498), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(new_n662), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n474), .A2(new_n662), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n499), .A2(new_n668), .A3(new_n509), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT95), .ZN(new_n670));
  AND3_X1   g0470(.A1(new_n667), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n670), .B1(new_n667), .B2(new_n669), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n665), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT96), .ZN(new_n675));
  OR2_X1    g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n674), .A2(new_n675), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n662), .ZN(new_n679));
  AND2_X1   g0479(.A1(new_n609), .A2(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n680), .B1(new_n671), .B2(new_n672), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n666), .A2(new_n679), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n678), .A2(new_n684), .ZN(G399));
  INV_X1    g0485(.A(new_n233), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n686), .A2(G41), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n515), .A2(new_n221), .ZN(new_n688));
  NOR3_X1   g0488(.A1(new_n687), .A2(new_n688), .A3(new_n305), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n689), .B1(new_n229), .B2(new_n687), .ZN(new_n690));
  XOR2_X1   g0490(.A(new_n690), .B(KEYINPUT28), .Z(new_n691));
  NAND2_X1  g0491(.A1(new_n638), .A2(new_n679), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT29), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n636), .A2(KEYINPUT26), .ZN(new_n695));
  OAI211_X1 g0495(.A(new_n695), .B(new_n621), .C1(new_n634), .C2(KEYINPUT26), .ZN(new_n696));
  AND4_X1   g0496(.A1(new_n581), .A2(new_n628), .A3(new_n617), .A4(new_n629), .ZN(new_n697));
  OAI211_X1 g0497(.A(KEYINPUT29), .B(new_n679), .C1(new_n696), .C2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n536), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n602), .A2(new_n451), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n578), .A2(new_n487), .A3(new_n699), .A4(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT30), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n699), .B1(new_n575), .B2(new_n576), .ZN(new_n704));
  INV_X1    g0504(.A(new_n507), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n704), .A2(new_n451), .A3(new_n705), .A4(new_n602), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n614), .A2(new_n536), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n707), .A2(KEYINPUT30), .A3(new_n487), .A4(new_n700), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n703), .A2(new_n706), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(new_n662), .ZN(new_n710));
  OAI211_X1 g0510(.A(KEYINPUT31), .B(new_n710), .C1(new_n618), .C2(new_n662), .ZN(new_n711));
  OR2_X1    g0511(.A1(new_n710), .A2(KEYINPUT31), .ZN(new_n712));
  AND2_X1   g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  AOI22_X1  g0513(.A1(new_n694), .A2(new_n698), .B1(new_n713), .B2(G330), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n691), .B1(new_n714), .B2(G1), .ZN(G364));
  AOI21_X1  g0515(.A(new_n230), .B1(G20), .B2(new_n324), .ZN(new_n716));
  NAND2_X1  g0516(.A1(G20), .A2(G179), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT97), .ZN(new_n718));
  XNOR2_X1  g0518(.A(new_n717), .B(new_n718), .ZN(new_n719));
  XNOR2_X1  g0519(.A(new_n719), .B(KEYINPUT98), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n720), .A2(G190), .A3(new_n363), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n720), .A2(new_n316), .A3(new_n363), .ZN(new_n722));
  OAI22_X1  g0522(.A1(new_n210), .A2(new_n721), .B1(new_n722), .B2(new_n251), .ZN(new_n723));
  XOR2_X1   g0523(.A(new_n723), .B(KEYINPUT99), .Z(new_n724));
  NOR2_X1   g0524(.A1(new_n231), .A2(G179), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n725), .A2(new_n316), .A3(G200), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(G107), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n725), .A2(G190), .A3(G200), .ZN(new_n729));
  OAI211_X1 g0529(.A(new_n728), .B(new_n300), .C1(new_n410), .C2(new_n729), .ZN(new_n730));
  XNOR2_X1  g0530(.A(new_n730), .B(KEYINPUT100), .ZN(new_n731));
  NOR3_X1   g0531(.A1(new_n316), .A2(G179), .A3(G200), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n732), .A2(new_n231), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n733), .A2(new_n205), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n719), .A2(G190), .A3(G200), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n734), .B1(new_n736), .B2(G50), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n719), .A2(new_n316), .A3(G200), .ZN(new_n738));
  OAI211_X1 g0538(.A(new_n731), .B(new_n737), .C1(new_n346), .C2(new_n738), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n725), .A2(new_n316), .A3(new_n363), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(G159), .ZN(new_n742));
  XNOR2_X1  g0542(.A(new_n742), .B(KEYINPUT32), .ZN(new_n743));
  NOR3_X1   g0543(.A1(new_n724), .A2(new_n739), .A3(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(G317), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n738), .B1(KEYINPUT33), .B2(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n746), .B1(KEYINPUT33), .B2(new_n745), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n736), .A2(G326), .ZN(new_n748));
  INV_X1    g0548(.A(new_n733), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(G294), .ZN(new_n750));
  INV_X1    g0550(.A(G283), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n292), .B1(new_n726), .B2(new_n751), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n752), .B1(G329), .B2(new_n741), .ZN(new_n753));
  NAND4_X1  g0553(.A1(new_n747), .A2(new_n748), .A3(new_n750), .A4(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(G311), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n722), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(G322), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n721), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(G303), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n729), .A2(new_n759), .ZN(new_n760));
  NOR4_X1   g0560(.A1(new_n754), .A2(new_n756), .A3(new_n758), .A4(new_n760), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n716), .B1(new_n744), .B2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n686), .A2(new_n300), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n229), .A2(new_n488), .ZN(new_n764));
  OAI211_X1 g0564(.A(new_n763), .B(new_n764), .C1(new_n252), .C2(new_n488), .ZN(new_n765));
  NAND3_X1  g0565(.A1(G355), .A2(new_n300), .A3(new_n233), .ZN(new_n766));
  OAI211_X1 g0566(.A(new_n765), .B(new_n766), .C1(G116), .C2(new_n233), .ZN(new_n767));
  NOR2_X1   g0567(.A1(G13), .A2(G33), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(G20), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(new_n716), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n767), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g0572(.A(new_n770), .B(KEYINPUT101), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  OAI211_X1 g0574(.A(new_n762), .B(new_n772), .C1(new_n664), .C2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n687), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n656), .A2(G45), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n776), .A2(G1), .A3(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n775), .A2(new_n779), .ZN(new_n780));
  XOR2_X1   g0580(.A(new_n664), .B(G330), .Z(new_n781));
  OAI21_X1  g0581(.A(new_n780), .B1(new_n781), .B2(new_n779), .ZN(new_n782));
  XOR2_X1   g0582(.A(new_n782), .B(KEYINPUT102), .Z(G396));
  INV_X1    g0583(.A(new_n722), .ZN(new_n784));
  AOI22_X1  g0584(.A1(new_n784), .A2(G159), .B1(G137), .B2(new_n736), .ZN(new_n785));
  INV_X1    g0585(.A(G143), .ZN(new_n786));
  OAI221_X1 g0586(.A(new_n785), .B1(new_n786), .B2(new_n721), .C1(new_n258), .C2(new_n738), .ZN(new_n787));
  XNOR2_X1  g0587(.A(new_n787), .B(KEYINPUT34), .ZN(new_n788));
  OAI22_X1  g0588(.A1(new_n202), .A2(new_n729), .B1(new_n726), .B2(new_n346), .ZN(new_n789));
  AOI211_X1 g0589(.A(new_n292), .B(new_n789), .C1(G58), .C2(new_n749), .ZN(new_n790));
  INV_X1    g0590(.A(G132), .ZN(new_n791));
  OAI211_X1 g0591(.A(new_n788), .B(new_n790), .C1(new_n791), .C2(new_n740), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n300), .B1(new_n741), .B2(G311), .ZN(new_n793));
  OAI221_X1 g0593(.A(new_n793), .B1(new_n751), .B2(new_n738), .C1(new_n722), .C2(new_n221), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n726), .A2(new_n410), .ZN(new_n795));
  INV_X1    g0595(.A(new_n729), .ZN(new_n796));
  AOI211_X1 g0596(.A(new_n795), .B(new_n734), .C1(G107), .C2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(G294), .ZN(new_n798));
  OAI221_X1 g0598(.A(new_n797), .B1(new_n759), .B2(new_n735), .C1(new_n721), .C2(new_n798), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n792), .B1(new_n794), .B2(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n716), .A2(new_n768), .ZN(new_n801));
  AOI22_X1  g0601(.A1(new_n800), .A2(new_n716), .B1(new_n251), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(new_n779), .ZN(new_n803));
  INV_X1    g0603(.A(KEYINPUT103), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n802), .A2(KEYINPUT103), .A3(new_n779), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n454), .A2(new_n679), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n372), .A2(new_n662), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n382), .A2(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n808), .B1(new_n453), .B2(new_n810), .ZN(new_n811));
  OAI211_X1 g0611(.A(new_n805), .B(new_n806), .C1(new_n769), .C2(new_n811), .ZN(new_n812));
  XOR2_X1   g0612(.A(new_n812), .B(KEYINPUT104), .Z(new_n813));
  XNOR2_X1  g0613(.A(new_n692), .B(new_n811), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n713), .A2(G330), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n814), .B(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(new_n778), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n813), .A2(new_n817), .ZN(G384));
  INV_X1    g0618(.A(KEYINPUT40), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n346), .B1(new_n388), .B2(new_n389), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n433), .B1(new_n440), .B2(new_n820), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n821), .A2(new_n269), .A3(new_n405), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n822), .A2(new_n385), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(KEYINPUT107), .ZN(new_n824));
  INV_X1    g0624(.A(new_n660), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT107), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n822), .A2(new_n826), .A3(new_n385), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n824), .A2(new_n825), .A3(new_n827), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n828), .B1(new_n646), .B2(new_n424), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n443), .A2(new_n445), .A3(new_n426), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n407), .A2(new_n825), .ZN(new_n831));
  XOR2_X1   g0631(.A(KEYINPUT109), .B(KEYINPUT37), .Z(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  NAND4_X1  g0633(.A1(new_n420), .A2(new_n830), .A3(new_n831), .A4(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  AND3_X1   g0635(.A1(new_n822), .A2(new_n826), .A3(new_n385), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n826), .B1(new_n822), .B2(new_n385), .ZN(new_n837));
  AND2_X1   g0637(.A1(new_n415), .A2(new_n416), .ZN(new_n838));
  NOR3_X1   g0638(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n427), .A2(new_n428), .ZN(new_n840));
  OAI21_X1  g0640(.A(KEYINPUT108), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n824), .A2(new_n648), .A3(new_n827), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT108), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n842), .A2(new_n843), .A3(new_n830), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n841), .A2(new_n828), .A3(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n835), .B1(new_n845), .B2(KEYINPUT37), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT38), .ZN(new_n847));
  NOR3_X1   g0647(.A1(new_n829), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n844), .A2(new_n828), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n843), .B1(new_n842), .B2(new_n830), .ZN(new_n850));
  OAI21_X1  g0650(.A(KEYINPUT37), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(new_n834), .ZN(new_n852));
  INV_X1    g0652(.A(new_n828), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n449), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g0654(.A(KEYINPUT38), .B1(new_n852), .B2(new_n854), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n848), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n360), .A2(KEYINPUT106), .A3(new_n364), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n359), .A2(new_n662), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  NAND4_X1  g0660(.A1(new_n360), .A2(KEYINPUT106), .A3(new_n364), .A4(new_n858), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND4_X1  g0662(.A1(new_n862), .A2(new_n711), .A3(new_n712), .A4(new_n811), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n819), .B1(new_n856), .B2(new_n863), .ZN(new_n864));
  AND4_X1   g0664(.A1(new_n711), .A2(new_n862), .A3(new_n712), .A4(new_n811), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n830), .A2(new_n649), .A3(new_n831), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT110), .ZN(new_n867));
  AND3_X1   g0667(.A1(new_n866), .A2(new_n867), .A3(new_n832), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n867), .B1(new_n866), .B2(new_n832), .ZN(new_n869));
  NOR3_X1   g0669(.A1(new_n868), .A2(new_n869), .A3(new_n835), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT111), .ZN(new_n871));
  AOI22_X1  g0671(.A1(new_n642), .A2(new_n871), .B1(new_n650), .B2(new_n651), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n429), .A2(KEYINPUT111), .A3(new_n446), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n831), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n847), .B1(new_n870), .B2(new_n874), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n852), .A2(new_n854), .A3(KEYINPUT38), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n819), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n865), .A2(new_n877), .ZN(new_n878));
  AND2_X1   g0678(.A1(new_n864), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n713), .A2(new_n455), .ZN(new_n880));
  XNOR2_X1  g0680(.A(new_n879), .B(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(G330), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n360), .A2(new_n662), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT39), .ZN(new_n884));
  AND3_X1   g0684(.A1(new_n875), .A2(new_n876), .A3(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n847), .B1(new_n829), .B2(new_n846), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n884), .B1(new_n886), .B2(new_n876), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n883), .B1(new_n885), .B2(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n650), .A2(new_n651), .A3(new_n660), .ZN(new_n889));
  AND2_X1   g0689(.A1(new_n860), .A2(new_n861), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n638), .A2(new_n811), .A3(new_n679), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n890), .B1(new_n891), .B2(new_n807), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n886), .A2(new_n876), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n888), .A2(new_n889), .A3(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n694), .A2(new_n455), .A3(new_n698), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(new_n654), .ZN(new_n897));
  XOR2_X1   g0697(.A(new_n895), .B(new_n897), .Z(new_n898));
  XNOR2_X1  g0698(.A(new_n882), .B(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n899), .B1(new_n305), .B2(new_n656), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n551), .A2(new_n553), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT35), .ZN(new_n902));
  AOI211_X1 g0702(.A(new_n231), .B(new_n230), .C1(new_n901), .C2(new_n902), .ZN(new_n903));
  OAI211_X1 g0703(.A(new_n903), .B(G116), .C1(new_n902), .C2(new_n901), .ZN(new_n904));
  XNOR2_X1  g0704(.A(new_n904), .B(KEYINPUT36), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n229), .A2(G77), .A3(new_n399), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n906), .B1(G50), .B2(new_n346), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n907), .A2(G1), .A3(new_n271), .ZN(new_n908));
  XOR2_X1   g0708(.A(new_n908), .B(KEYINPUT105), .Z(new_n909));
  NAND3_X1  g0709(.A1(new_n900), .A2(new_n905), .A3(new_n909), .ZN(G367));
  OAI221_X1 g0710(.A(new_n300), .B1(new_n395), .B2(new_n738), .C1(new_n721), .C2(new_n258), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n727), .A2(G77), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n912), .B1(new_n210), .B2(new_n729), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n913), .B1(G137), .B2(new_n741), .ZN(new_n914));
  OAI221_X1 g0714(.A(new_n914), .B1(new_n346), .B2(new_n733), .C1(new_n786), .C2(new_n735), .ZN(new_n915));
  AOI211_X1 g0715(.A(new_n911), .B(new_n915), .C1(G50), .C2(new_n784), .ZN(new_n916));
  OAI22_X1  g0716(.A1(new_n751), .A2(new_n722), .B1(new_n721), .B2(new_n759), .ZN(new_n917));
  OAI22_X1  g0717(.A1(new_n798), .A2(new_n738), .B1(new_n735), .B2(new_n755), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n300), .B1(new_n741), .B2(G317), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n749), .A2(G107), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n727), .A2(G97), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT46), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n922), .B1(new_n729), .B2(new_n221), .ZN(new_n923));
  NAND4_X1  g0723(.A1(new_n919), .A2(new_n920), .A3(new_n921), .A4(new_n923), .ZN(new_n924));
  NOR3_X1   g0724(.A1(new_n917), .A2(new_n918), .A3(new_n924), .ZN(new_n925));
  NOR3_X1   g0725(.A1(new_n729), .A2(new_n922), .A3(new_n221), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n926), .B(KEYINPUT114), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n916), .B1(new_n925), .B2(new_n927), .ZN(new_n928));
  XOR2_X1   g0728(.A(new_n928), .B(KEYINPUT47), .Z(new_n929));
  AOI21_X1  g0729(.A(new_n778), .B1(new_n929), .B2(new_n716), .ZN(new_n930));
  INV_X1    g0730(.A(new_n763), .ZN(new_n931));
  OAI221_X1 g0731(.A(new_n771), .B1(new_n233), .B2(new_n367), .C1(new_n247), .C2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT112), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n625), .A2(new_n679), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n935), .A2(new_n621), .ZN(new_n936));
  INV_X1    g0736(.A(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n935), .A2(new_n627), .A3(new_n621), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n933), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n939), .B1(new_n933), .B2(new_n937), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  OAI211_X1 g0741(.A(new_n930), .B(new_n932), .C1(new_n774), .C2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n777), .A2(G1), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n565), .A2(new_n662), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n581), .A2(new_n617), .A3(new_n944), .ZN(new_n945));
  OR2_X1    g0745(.A1(new_n945), .A2(KEYINPUT113), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(KEYINPUT113), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  AND2_X1   g0748(.A1(new_n579), .A2(new_n565), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n949), .A2(new_n662), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  AOI21_X1  g0751(.A(KEYINPUT45), .B1(new_n951), .B2(new_n684), .ZN(new_n952));
  AOI22_X1  g0752(.A1(new_n946), .A2(new_n947), .B1(new_n949), .B2(new_n662), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT45), .ZN(new_n954));
  NOR3_X1   g0754(.A1(new_n953), .A2(new_n683), .A3(new_n954), .ZN(new_n955));
  AND3_X1   g0755(.A1(new_n953), .A2(new_n683), .A3(KEYINPUT44), .ZN(new_n956));
  AOI21_X1  g0756(.A(KEYINPUT44), .B1(new_n953), .B2(new_n683), .ZN(new_n957));
  OAI22_X1  g0757(.A1(new_n952), .A2(new_n955), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n674), .B(KEYINPUT96), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT44), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(new_n951), .B2(new_n684), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n953), .A2(new_n683), .A3(KEYINPUT44), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n951), .A2(new_n684), .A3(KEYINPUT45), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n954), .B1(new_n953), .B2(new_n683), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n678), .A2(new_n964), .A3(new_n967), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n680), .B1(new_n664), .B2(G330), .ZN(new_n969));
  XOR2_X1   g0769(.A(new_n969), .B(new_n673), .Z(new_n970));
  NAND4_X1  g0770(.A1(new_n960), .A2(new_n968), .A3(new_n714), .A4(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(new_n714), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n687), .B(KEYINPUT41), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n943), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  OR3_X1    g0774(.A1(new_n953), .A2(KEYINPUT42), .A3(new_n681), .ZN(new_n975));
  OAI21_X1  g0775(.A(KEYINPUT42), .B1(new_n953), .B2(new_n681), .ZN(new_n976));
  INV_X1    g0776(.A(new_n581), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n977), .B1(new_n951), .B2(new_n666), .ZN(new_n978));
  OAI211_X1 g0778(.A(new_n975), .B(new_n976), .C1(new_n662), .C2(new_n978), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n676), .A2(new_n677), .A3(new_n951), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n941), .A2(KEYINPUT43), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n979), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(new_n982), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n980), .B1(new_n979), .B2(new_n981), .ZN(new_n984));
  OAI22_X1  g0784(.A1(new_n983), .A2(new_n984), .B1(KEYINPUT43), .B2(new_n941), .ZN(new_n985));
  INV_X1    g0785(.A(new_n984), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n941), .A2(KEYINPUT43), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n986), .A2(new_n987), .A3(new_n982), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n985), .A2(new_n988), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n942), .B1(new_n974), .B2(new_n989), .ZN(G387));
  INV_X1    g0790(.A(new_n771), .ZN(new_n991));
  OR2_X1    g0791(.A1(new_n243), .A2(new_n488), .ZN(new_n992));
  OR3_X1    g0792(.A1(new_n261), .A2(KEYINPUT50), .A3(G50), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n688), .B1(G68), .B2(G77), .ZN(new_n994));
  OAI21_X1  g0794(.A(KEYINPUT50), .B1(new_n261), .B2(G50), .ZN(new_n995));
  NAND4_X1  g0795(.A1(new_n993), .A2(new_n994), .A3(new_n995), .A4(new_n488), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n996), .A2(new_n763), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(KEYINPUT115), .ZN(new_n998));
  AOI22_X1  g0798(.A1(new_n992), .A2(new_n998), .B1(new_n206), .B2(new_n686), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n688), .A2(new_n233), .A3(new_n300), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n991), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(new_n784), .A2(G303), .B1(G322), .B2(new_n736), .ZN(new_n1002));
  OAI221_X1 g0802(.A(new_n1002), .B1(new_n755), .B2(new_n738), .C1(new_n745), .C2(new_n721), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT48), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n749), .A2(G283), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n796), .A2(G294), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n1004), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT49), .ZN(new_n1008));
  OR2_X1    g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n741), .A2(G326), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n300), .B1(new_n727), .B2(G116), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n1009), .A2(new_n1010), .A3(new_n1011), .A4(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n292), .B1(new_n741), .B2(G150), .ZN(new_n1014));
  OAI211_X1 g0814(.A(new_n1014), .B(new_n921), .C1(new_n251), .C2(new_n729), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n721), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1015), .B1(new_n1016), .B2(G50), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n784), .A2(G68), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n542), .A2(new_n733), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n1019), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n738), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n265), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(G159), .A2(new_n736), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n1017), .A2(new_n1018), .A3(new_n1020), .A4(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1013), .A2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1001), .B1(new_n1025), .B2(new_n716), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n673), .A2(new_n773), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1026), .A2(new_n779), .A3(new_n1027), .ZN(new_n1028));
  XOR2_X1   g0828(.A(new_n1028), .B(KEYINPUT116), .Z(new_n1029));
  NAND2_X1  g0829(.A1(new_n970), .A2(new_n943), .ZN(new_n1030));
  OR2_X1    g0830(.A1(new_n714), .A2(new_n970), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n714), .A2(new_n970), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1031), .A2(new_n687), .A3(new_n1032), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1029), .A2(new_n1030), .A3(new_n1033), .ZN(G393));
  NAND3_X1  g0834(.A1(new_n960), .A2(KEYINPUT117), .A3(new_n968), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT117), .ZN(new_n1036));
  NAND4_X1  g0836(.A1(new_n678), .A2(new_n964), .A3(new_n967), .A4(new_n1036), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1035), .A2(new_n1032), .A3(new_n1037), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1038), .A2(new_n687), .A3(new_n971), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n233), .A2(new_n205), .ZN(new_n1040));
  AOI211_X1 g0840(.A(new_n1040), .B(new_n991), .C1(new_n255), .C2(new_n763), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n1016), .A2(G311), .B1(G317), .B2(new_n736), .ZN(new_n1042));
  OR2_X1    g0842(.A1(new_n1042), .A2(KEYINPUT52), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n728), .B1(new_n751), .B2(new_n729), .C1(new_n221), .C2(new_n733), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1044), .B1(new_n784), .B2(G294), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1042), .A2(KEYINPUT52), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n292), .B1(new_n740), .B2(new_n757), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1047), .B1(new_n1021), .B2(G303), .ZN(new_n1048));
  NAND4_X1  g0848(.A1(new_n1043), .A2(new_n1045), .A3(new_n1046), .A4(new_n1048), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n721), .A2(new_n395), .B1(new_n258), .B2(new_n735), .ZN(new_n1050));
  XOR2_X1   g0850(.A(new_n1050), .B(KEYINPUT51), .Z(new_n1051));
  NOR2_X1   g0851(.A1(new_n722), .A2(new_n261), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n749), .A2(G77), .B1(new_n796), .B2(new_n219), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n1053), .B1(new_n786), .B2(new_n740), .C1(new_n202), .C2(new_n738), .ZN(new_n1054));
  OR4_X1    g0854(.A1(new_n292), .A2(new_n1051), .A3(new_n1052), .A4(new_n1054), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1049), .B1(new_n1055), .B2(new_n795), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1056), .A2(new_n716), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1057), .A2(new_n779), .ZN(new_n1058));
  AOI211_X1 g0858(.A(new_n1041), .B(new_n1058), .C1(new_n953), .C2(new_n770), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1035), .A2(new_n1037), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1059), .B1(new_n1060), .B2(new_n943), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1039), .A2(new_n1061), .ZN(G390));
  OAI21_X1  g0862(.A(KEYINPUT39), .B1(new_n848), .B2(new_n855), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n875), .A2(new_n876), .A3(new_n884), .ZN(new_n1064));
  OAI211_X1 g0864(.A(new_n1063), .B(new_n1064), .C1(new_n892), .C2(new_n883), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n810), .A2(new_n453), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n679), .B(new_n1066), .C1(new_n696), .C2(new_n697), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT118), .ZN(new_n1068));
  AND3_X1   g0868(.A1(new_n1067), .A2(new_n1068), .A3(new_n807), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1068), .B1(new_n1067), .B2(new_n807), .ZN(new_n1070));
  NOR3_X1   g0870(.A1(new_n1069), .A2(new_n1070), .A3(new_n890), .ZN(new_n1071));
  AND2_X1   g0871(.A1(new_n875), .A2(new_n876), .ZN(new_n1072));
  OR2_X1    g0872(.A1(new_n1072), .A2(new_n883), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1065), .B1(new_n1071), .B2(new_n1073), .ZN(new_n1074));
  NAND4_X1  g0874(.A1(new_n711), .A2(G330), .A3(new_n712), .A4(new_n811), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n1075), .A2(new_n890), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1070), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1067), .A2(new_n1068), .A3(new_n807), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1078), .A2(new_n862), .A3(new_n1079), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n1072), .A2(new_n883), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NAND4_X1  g0882(.A1(new_n713), .A2(G330), .A3(new_n811), .A4(new_n862), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1082), .A2(new_n1065), .A3(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1077), .A2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n713), .A2(G330), .A3(new_n455), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n896), .A2(new_n1086), .A3(new_n654), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1075), .A2(new_n890), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n1083), .B(new_n1088), .C1(new_n1069), .C2(new_n1070), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n891), .A2(new_n807), .ZN(new_n1090));
  AND2_X1   g0890(.A1(new_n1075), .A2(new_n890), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1090), .B1(new_n1091), .B2(new_n1076), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1087), .B1(new_n1089), .B2(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1085), .A2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1077), .A2(new_n1084), .A3(new_n1093), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1095), .A2(new_n687), .A3(new_n1096), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1077), .A2(new_n943), .A3(new_n1084), .ZN(new_n1098));
  INV_X1    g0898(.A(KEYINPUT120), .ZN(new_n1099));
  OAI221_X1 g0899(.A(new_n300), .B1(new_n726), .B2(new_n202), .C1(new_n733), .C2(new_n395), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1100), .B1(G128), .B2(new_n736), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n741), .A2(G125), .ZN(new_n1102));
  INV_X1    g0902(.A(G137), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n1101), .B(new_n1102), .C1(new_n1103), .C2(new_n738), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1104), .B1(G132), .B2(new_n1016), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n729), .A2(new_n258), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(new_n1106), .B(KEYINPUT53), .ZN(new_n1107));
  XOR2_X1   g0907(.A(KEYINPUT54), .B(G143), .Z(new_n1108));
  INV_X1    g0908(.A(new_n1108), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n1105), .B(new_n1107), .C1(new_n722), .C2(new_n1109), .ZN(new_n1110));
  XOR2_X1   g0910(.A(new_n1110), .B(KEYINPUT119), .Z(new_n1111));
  NOR2_X1   g0911(.A1(new_n721), .A2(new_n221), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n722), .A2(new_n205), .ZN(new_n1113));
  OAI221_X1 g0913(.A(new_n292), .B1(new_n798), .B2(new_n740), .C1(new_n738), .C2(new_n206), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n749), .A2(G77), .B1(new_n727), .B2(G68), .ZN(new_n1115));
  OAI221_X1 g0915(.A(new_n1115), .B1(new_n410), .B2(new_n729), .C1(new_n751), .C2(new_n735), .ZN(new_n1116));
  NOR4_X1   g0916(.A1(new_n1112), .A2(new_n1113), .A3(new_n1114), .A4(new_n1116), .ZN(new_n1117));
  OR2_X1    g0917(.A1(new_n1111), .A2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n778), .B1(new_n1118), .B2(new_n716), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n801), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1121));
  OAI221_X1 g0921(.A(new_n1119), .B1(new_n1022), .B2(new_n1120), .C1(new_n1121), .C2(new_n769), .ZN(new_n1122));
  AND3_X1   g0922(.A1(new_n1098), .A2(new_n1099), .A3(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1099), .B1(new_n1098), .B2(new_n1122), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1097), .B1(new_n1123), .B2(new_n1124), .ZN(G378));
  AOI22_X1  g0925(.A1(new_n736), .A2(G125), .B1(G150), .B2(new_n749), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1126), .B1(new_n791), .B2(new_n738), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1127), .B1(new_n1016), .B2(G128), .ZN(new_n1128));
  OAI221_X1 g0928(.A(new_n1128), .B1(new_n1103), .B2(new_n722), .C1(new_n729), .C2(new_n1109), .ZN(new_n1129));
  XOR2_X1   g0929(.A(new_n1129), .B(KEYINPUT59), .Z(new_n1130));
  AOI21_X1  g0930(.A(G41), .B1(new_n727), .B2(G159), .ZN(new_n1131));
  AOI21_X1  g0931(.A(G33), .B1(new_n741), .B2(G124), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1130), .A2(new_n1131), .A3(new_n1132), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n202), .B1(new_n290), .B2(G41), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n206), .A2(new_n721), .B1(new_n722), .B2(new_n542), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n749), .A2(G68), .B1(new_n741), .B2(G283), .ZN(new_n1136));
  AOI211_X1 g0936(.A(G41), .B(new_n300), .C1(new_n796), .C2(G77), .ZN(new_n1137));
  OAI221_X1 g0937(.A(new_n1136), .B1(new_n210), .B2(new_n726), .C1(new_n1137), .C2(KEYINPUT121), .ZN(new_n1138));
  OAI22_X1  g0938(.A1(new_n205), .A2(new_n738), .B1(new_n735), .B2(new_n221), .ZN(new_n1139));
  NOR3_X1   g0939(.A1(new_n1135), .A2(new_n1138), .A3(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1137), .A2(KEYINPUT121), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  XNOR2_X1  g0942(.A(new_n1142), .B(KEYINPUT58), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1133), .A2(new_n1134), .A3(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(new_n716), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(new_n1145), .B(KEYINPUT122), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n779), .B1(G50), .B2(new_n1120), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(new_n1147), .B(KEYINPUT123), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT56), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n284), .A2(new_n660), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n328), .A2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1150), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1152), .B1(new_n322), .B2(new_n327), .ZN(new_n1153));
  OAI21_X1  g0953(.A(KEYINPUT55), .B1(new_n1151), .B2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  NOR3_X1   g0955(.A1(new_n1151), .A2(KEYINPUT55), .A3(new_n1153), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1149), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1156), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1158), .A2(KEYINPUT56), .A3(new_n1154), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1157), .A2(new_n1159), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n1146), .B(new_n1148), .C1(new_n1160), .C2(new_n769), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(new_n1161), .B(KEYINPUT124), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n895), .B1(G330), .B2(new_n879), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n864), .A2(G330), .A3(new_n878), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(new_n1121), .A2(new_n883), .B1(new_n893), .B2(new_n892), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1164), .B1(new_n1165), .B2(new_n889), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1160), .B1(new_n1163), .B2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n879), .A2(new_n895), .A3(G330), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1165), .A2(new_n1164), .A3(new_n889), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1160), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1168), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1167), .A2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1162), .B1(new_n1172), .B2(new_n943), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1087), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n1167), .A2(new_n1171), .B1(new_n1096), .B2(new_n1174), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n687), .B1(new_n1175), .B2(KEYINPUT57), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1096), .A2(new_n1174), .ZN(new_n1177));
  AND3_X1   g0977(.A1(new_n1172), .A2(KEYINPUT57), .A3(new_n1177), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1173), .B1(new_n1176), .B2(new_n1178), .ZN(G375));
  INV_X1    g0979(.A(new_n943), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1180), .B1(new_n1089), .B2(new_n1092), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(new_n749), .A2(G50), .B1(new_n796), .B2(G159), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n741), .A2(G128), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1182), .B(new_n1183), .C1(new_n738), .C2(new_n1109), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1184), .B1(G132), .B2(new_n736), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1016), .A2(G137), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n784), .A2(G150), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n292), .B1(new_n727), .B2(G58), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n1185), .A2(new_n1186), .A3(new_n1187), .A4(new_n1188), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(new_n784), .A2(G107), .B1(G294), .B2(new_n736), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1190), .B1(new_n221), .B2(new_n738), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(new_n1191), .B(KEYINPUT125), .ZN(new_n1192));
  OAI221_X1 g0992(.A(new_n292), .B1(new_n740), .B2(new_n759), .C1(new_n205), .C2(new_n729), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(new_n1016), .B2(G283), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1192), .A2(new_n912), .A3(new_n1194), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1189), .B1(new_n1195), .B2(new_n1019), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1196), .A2(new_n716), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1197), .B1(G68), .B2(new_n1120), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1198), .B1(new_n768), .B2(new_n890), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1181), .B1(new_n779), .B2(new_n1199), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1089), .A2(new_n1092), .A3(new_n1087), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1201), .A2(new_n973), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1200), .B1(new_n1202), .B2(new_n1093), .ZN(G381));
  AND2_X1   g1003(.A1(new_n1098), .A2(new_n1122), .ZN(new_n1204));
  AND2_X1   g1004(.A1(new_n1097), .A2(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(G375), .A2(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(G381), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(G393), .A2(G396), .ZN(new_n1209));
  NOR3_X1   g1009(.A1(G387), .A2(G384), .A3(G390), .ZN(new_n1210));
  NAND4_X1  g1010(.A1(new_n1207), .A2(new_n1208), .A3(new_n1209), .A4(new_n1210), .ZN(G407));
  INV_X1    g1011(.A(G213), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1212), .B1(new_n1207), .B2(new_n661), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1213), .A2(G407), .ZN(G409));
  NOR2_X1   g1014(.A1(new_n1212), .A2(G343), .ZN(new_n1215));
  OAI211_X1 g1015(.A(G378), .B(new_n1173), .C1(new_n1176), .C2(new_n1178), .ZN(new_n1216));
  AND2_X1   g1016(.A1(new_n1175), .A2(new_n973), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1162), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1171), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1170), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1218), .B1(new_n1221), .B2(new_n1180), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1205), .B1(new_n1217), .B2(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1215), .B1(new_n1216), .B2(new_n1223), .ZN(new_n1224));
  XNOR2_X1  g1024(.A(KEYINPUT126), .B(KEYINPUT60), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n776), .B1(new_n1201), .B2(new_n1225), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1089), .A2(new_n1092), .A3(KEYINPUT60), .A4(new_n1087), .ZN(new_n1227));
  AND2_X1   g1027(.A1(new_n1227), .A2(KEYINPUT127), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1227), .A2(KEYINPUT127), .ZN(new_n1229));
  OAI211_X1 g1029(.A(new_n1094), .B(new_n1226), .C1(new_n1228), .C2(new_n1229), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1230), .A2(G384), .A3(new_n1200), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(G384), .B1(new_n1230), .B2(new_n1200), .ZN(new_n1233));
  OAI211_X1 g1033(.A(G2897), .B(new_n1215), .C1(new_n1232), .C2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1230), .A2(new_n1200), .ZN(new_n1235));
  INV_X1    g1035(.A(G384), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1215), .A2(G2897), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1237), .A2(new_n1231), .A3(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1234), .A2(new_n1239), .ZN(new_n1240));
  OAI21_X1  g1040(.A(KEYINPUT63), .B1(new_n1224), .B2(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1237), .A2(new_n1231), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1224), .A2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1241), .A2(new_n1244), .ZN(new_n1245));
  XNOR2_X1  g1045(.A(G393), .B(G396), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n973), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1247), .B1(new_n971), .B2(new_n714), .ZN(new_n1248));
  OAI211_X1 g1048(.A(new_n988), .B(new_n985), .C1(new_n1248), .C2(new_n943), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(G390), .A2(new_n1249), .A3(new_n942), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(G390), .B1(new_n942), .B2(new_n1249), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1246), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  XOR2_X1   g1053(.A(G393), .B(G396), .Z(new_n1254));
  NAND3_X1  g1054(.A1(G387), .A2(new_n1061), .A3(new_n1039), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1254), .A2(new_n1250), .A3(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1253), .A2(new_n1256), .ZN(new_n1257));
  AOI211_X1 g1057(.A(new_n1215), .B(new_n1242), .C1(new_n1216), .C2(new_n1223), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1257), .B1(new_n1258), .B2(KEYINPUT63), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT61), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1245), .A2(new_n1259), .A3(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT62), .ZN(new_n1262));
  AND3_X1   g1062(.A1(new_n1224), .A2(new_n1262), .A3(new_n1243), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1260), .B1(new_n1224), .B2(new_n1240), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1262), .B1(new_n1224), .B2(new_n1243), .ZN(new_n1265));
  NOR3_X1   g1065(.A1(new_n1263), .A2(new_n1264), .A3(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1257), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1261), .B1(new_n1266), .B2(new_n1267), .ZN(G405));
  NAND2_X1  g1068(.A1(G375), .A2(new_n1205), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1269), .A2(new_n1216), .A3(new_n1242), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1242), .B1(new_n1269), .B2(new_n1216), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  XNOR2_X1  g1073(.A(new_n1273), .B(new_n1267), .ZN(G402));
endmodule


