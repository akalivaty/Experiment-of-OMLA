

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U551 ( .A(KEYINPUT23), .B(KEYINPUT67), .ZN(n589) );
  AND2_X1 U552 ( .A1(n525), .A2(G2105), .ZN(n891) );
  XNOR2_X1 U553 ( .A(n601), .B(n600), .ZN(n769) );
  OR2_X2 U554 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X2 U555 ( .A(G2104), .B(KEYINPUT65), .ZN(n525) );
  NOR2_X1 U556 ( .A1(n597), .A2(n596), .ZN(n599) );
  XNOR2_X1 U557 ( .A(n727), .B(n604), .ZN(n605) );
  XNOR2_X1 U558 ( .A(n679), .B(n678), .ZN(n703) );
  NAND2_X1 U559 ( .A1(n677), .A2(n676), .ZN(n679) );
  NAND2_X1 U560 ( .A1(n599), .A2(n598), .ZN(n601) );
  XOR2_X1 U561 ( .A(n662), .B(n661), .Z(n518) );
  NOR2_X1 U562 ( .A1(n682), .A2(n681), .ZN(n519) );
  XOR2_X1 U563 ( .A(KEYINPUT92), .B(n716), .Z(n520) );
  OR2_X1 U564 ( .A1(G301), .A2(n663), .ZN(n521) );
  INV_X1 U565 ( .A(KEYINPUT96), .ZN(n610) );
  XNOR2_X1 U566 ( .A(KEYINPUT97), .B(KEYINPUT30), .ZN(n661) );
  INV_X1 U567 ( .A(KEYINPUT29), .ZN(n653) );
  XNOR2_X1 U568 ( .A(n667), .B(KEYINPUT31), .ZN(n668) );
  INV_X1 U569 ( .A(KEYINPUT90), .ZN(n604) );
  INV_X1 U570 ( .A(KEYINPUT32), .ZN(n678) );
  INV_X1 U571 ( .A(KEYINPUT87), .ZN(n602) );
  NOR2_X1 U572 ( .A1(G651), .A2(G543), .ZN(n796) );
  NOR2_X1 U573 ( .A1(G651), .A2(n566), .ZN(n800) );
  NOR2_X1 U574 ( .A1(G2105), .A2(G2104), .ZN(n522) );
  XOR2_X1 U575 ( .A(KEYINPUT17), .B(n522), .Z(n593) );
  BUF_X1 U576 ( .A(n593), .Z(n893) );
  NAND2_X1 U577 ( .A1(G138), .A2(n893), .ZN(n524) );
  NAND2_X1 U578 ( .A1(G126), .A2(n891), .ZN(n523) );
  NAND2_X1 U579 ( .A1(n524), .A2(n523), .ZN(n530) );
  AND2_X1 U580 ( .A1(G2105), .A2(G2104), .ZN(n890) );
  NAND2_X1 U581 ( .A1(G114), .A2(n890), .ZN(n528) );
  NOR2_X2 U582 ( .A1(n525), .A2(G2105), .ZN(n588) );
  INV_X1 U583 ( .A(n588), .ZN(n526) );
  INV_X1 U584 ( .A(n526), .ZN(n894) );
  NAND2_X1 U585 ( .A1(G102), .A2(n894), .ZN(n527) );
  NAND2_X1 U586 ( .A1(n528), .A2(n527), .ZN(n529) );
  NOR2_X1 U587 ( .A1(n530), .A2(n529), .ZN(G164) );
  XOR2_X1 U588 ( .A(KEYINPUT0), .B(G543), .Z(n566) );
  NAND2_X1 U589 ( .A1(n800), .A2(G53), .ZN(n531) );
  XNOR2_X1 U590 ( .A(n531), .B(KEYINPUT70), .ZN(n535) );
  INV_X1 U591 ( .A(G651), .ZN(n537) );
  NOR2_X1 U592 ( .A1(G543), .A2(n537), .ZN(n532) );
  XOR2_X1 U593 ( .A(KEYINPUT1), .B(n532), .Z(n533) );
  XNOR2_X1 U594 ( .A(KEYINPUT68), .B(n533), .ZN(n802) );
  NAND2_X1 U595 ( .A1(G65), .A2(n802), .ZN(n534) );
  NAND2_X1 U596 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U597 ( .A(KEYINPUT71), .B(n536), .ZN(n541) );
  NAND2_X1 U598 ( .A1(G91), .A2(n796), .ZN(n539) );
  NOR2_X1 U599 ( .A1(n566), .A2(n537), .ZN(n797) );
  NAND2_X1 U600 ( .A1(G78), .A2(n797), .ZN(n538) );
  AND2_X1 U601 ( .A1(n539), .A2(n538), .ZN(n540) );
  NAND2_X1 U602 ( .A1(n541), .A2(n540), .ZN(G299) );
  NAND2_X1 U603 ( .A1(n800), .A2(G52), .ZN(n543) );
  NAND2_X1 U604 ( .A1(G64), .A2(n802), .ZN(n542) );
  NAND2_X1 U605 ( .A1(n543), .A2(n542), .ZN(n549) );
  NAND2_X1 U606 ( .A1(G90), .A2(n796), .ZN(n545) );
  NAND2_X1 U607 ( .A1(G77), .A2(n797), .ZN(n544) );
  NAND2_X1 U608 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U609 ( .A(KEYINPUT69), .B(n546), .ZN(n547) );
  XNOR2_X1 U610 ( .A(KEYINPUT9), .B(n547), .ZN(n548) );
  NOR2_X1 U611 ( .A1(n549), .A2(n548), .ZN(G171) );
  INV_X1 U612 ( .A(G171), .ZN(G301) );
  NAND2_X1 U613 ( .A1(n796), .A2(G89), .ZN(n550) );
  XNOR2_X1 U614 ( .A(n550), .B(KEYINPUT4), .ZN(n552) );
  NAND2_X1 U615 ( .A1(G76), .A2(n797), .ZN(n551) );
  NAND2_X1 U616 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U617 ( .A(n553), .B(KEYINPUT5), .ZN(n558) );
  NAND2_X1 U618 ( .A1(n800), .A2(G51), .ZN(n555) );
  NAND2_X1 U619 ( .A1(G63), .A2(n802), .ZN(n554) );
  NAND2_X1 U620 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U621 ( .A(KEYINPUT6), .B(n556), .Z(n557) );
  NAND2_X1 U622 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U623 ( .A(n559), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U624 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U625 ( .A1(G88), .A2(n796), .ZN(n561) );
  NAND2_X1 U626 ( .A1(G75), .A2(n797), .ZN(n560) );
  NAND2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n565) );
  NAND2_X1 U628 ( .A1(n800), .A2(G50), .ZN(n563) );
  NAND2_X1 U629 ( .A1(G62), .A2(n802), .ZN(n562) );
  NAND2_X1 U630 ( .A1(n563), .A2(n562), .ZN(n564) );
  NOR2_X1 U631 ( .A1(n565), .A2(n564), .ZN(G166) );
  INV_X1 U632 ( .A(G166), .ZN(G303) );
  NAND2_X1 U633 ( .A1(n800), .A2(G49), .ZN(n571) );
  NAND2_X1 U634 ( .A1(G87), .A2(n566), .ZN(n568) );
  NAND2_X1 U635 ( .A1(G74), .A2(G651), .ZN(n567) );
  NAND2_X1 U636 ( .A1(n568), .A2(n567), .ZN(n569) );
  NOR2_X1 U637 ( .A1(n802), .A2(n569), .ZN(n570) );
  NAND2_X1 U638 ( .A1(n571), .A2(n570), .ZN(n572) );
  XOR2_X1 U639 ( .A(KEYINPUT81), .B(n572), .Z(G288) );
  NAND2_X1 U640 ( .A1(n797), .A2(G73), .ZN(n574) );
  XNOR2_X1 U641 ( .A(KEYINPUT2), .B(KEYINPUT82), .ZN(n573) );
  XNOR2_X1 U642 ( .A(n574), .B(n573), .ZN(n581) );
  NAND2_X1 U643 ( .A1(n796), .A2(G86), .ZN(n576) );
  NAND2_X1 U644 ( .A1(G61), .A2(n802), .ZN(n575) );
  NAND2_X1 U645 ( .A1(n576), .A2(n575), .ZN(n579) );
  NAND2_X1 U646 ( .A1(G48), .A2(n800), .ZN(n577) );
  XNOR2_X1 U647 ( .A(KEYINPUT83), .B(n577), .ZN(n578) );
  NOR2_X1 U648 ( .A1(n579), .A2(n578), .ZN(n580) );
  NAND2_X1 U649 ( .A1(n581), .A2(n580), .ZN(G305) );
  AND2_X1 U650 ( .A1(G60), .A2(n802), .ZN(n585) );
  NAND2_X1 U651 ( .A1(G85), .A2(n796), .ZN(n583) );
  NAND2_X1 U652 ( .A1(G72), .A2(n797), .ZN(n582) );
  NAND2_X1 U653 ( .A1(n583), .A2(n582), .ZN(n584) );
  NOR2_X1 U654 ( .A1(n585), .A2(n584), .ZN(n587) );
  NAND2_X1 U655 ( .A1(n800), .A2(G47), .ZN(n586) );
  NAND2_X1 U656 ( .A1(n587), .A2(n586), .ZN(G290) );
  NAND2_X1 U657 ( .A1(n588), .A2(G101), .ZN(n592) );
  INV_X1 U658 ( .A(n589), .ZN(n590) );
  XNOR2_X1 U659 ( .A(n590), .B(KEYINPUT66), .ZN(n591) );
  XNOR2_X1 U660 ( .A(n592), .B(n591), .ZN(n597) );
  NAND2_X1 U661 ( .A1(G137), .A2(n593), .ZN(n595) );
  NAND2_X1 U662 ( .A1(G113), .A2(n890), .ZN(n594) );
  NAND2_X1 U663 ( .A1(n595), .A2(n594), .ZN(n596) );
  NAND2_X1 U664 ( .A1(n891), .A2(G125), .ZN(n598) );
  INV_X1 U665 ( .A(KEYINPUT64), .ZN(n600) );
  NAND2_X1 U666 ( .A1(n769), .A2(G40), .ZN(n603) );
  XNOR2_X2 U667 ( .A(n603), .B(n602), .ZN(n727) );
  NOR2_X1 U668 ( .A1(G164), .A2(G1384), .ZN(n728) );
  NAND2_X2 U669 ( .A1(n605), .A2(n728), .ZN(n659) );
  INV_X1 U670 ( .A(n659), .ZN(n606) );
  NAND2_X1 U671 ( .A1(n606), .A2(G1996), .ZN(n607) );
  XNOR2_X1 U672 ( .A(n607), .B(KEYINPUT26), .ZN(n609) );
  BUF_X4 U673 ( .A(n659), .Z(n670) );
  NAND2_X1 U674 ( .A1(G1341), .A2(n670), .ZN(n608) );
  NAND2_X1 U675 ( .A1(n609), .A2(n608), .ZN(n611) );
  XNOR2_X1 U676 ( .A(n611), .B(n610), .ZN(n622) );
  NAND2_X1 U677 ( .A1(G43), .A2(n800), .ZN(n621) );
  NAND2_X1 U678 ( .A1(G56), .A2(n802), .ZN(n612) );
  XNOR2_X1 U679 ( .A(KEYINPUT14), .B(n612), .ZN(n618) );
  NAND2_X1 U680 ( .A1(n796), .A2(G81), .ZN(n613) );
  XNOR2_X1 U681 ( .A(n613), .B(KEYINPUT12), .ZN(n615) );
  NAND2_X1 U682 ( .A1(G68), .A2(n797), .ZN(n614) );
  NAND2_X1 U683 ( .A1(n615), .A2(n614), .ZN(n616) );
  XNOR2_X1 U684 ( .A(KEYINPUT13), .B(n616), .ZN(n617) );
  NAND2_X1 U685 ( .A1(n618), .A2(n617), .ZN(n619) );
  XNOR2_X1 U686 ( .A(KEYINPUT73), .B(n619), .ZN(n620) );
  NAND2_X1 U687 ( .A1(n621), .A2(n620), .ZN(n971) );
  INV_X1 U688 ( .A(n971), .ZN(n773) );
  AND2_X2 U689 ( .A1(n622), .A2(n773), .ZN(n636) );
  NAND2_X1 U690 ( .A1(n796), .A2(G92), .ZN(n624) );
  NAND2_X1 U691 ( .A1(G66), .A2(n802), .ZN(n623) );
  NAND2_X1 U692 ( .A1(n624), .A2(n623), .ZN(n628) );
  NAND2_X1 U693 ( .A1(G79), .A2(n797), .ZN(n626) );
  NAND2_X1 U694 ( .A1(G54), .A2(n800), .ZN(n625) );
  NAND2_X1 U695 ( .A1(n626), .A2(n625), .ZN(n627) );
  NOR2_X1 U696 ( .A1(n628), .A2(n627), .ZN(n630) );
  XNOR2_X1 U697 ( .A(KEYINPUT15), .B(KEYINPUT75), .ZN(n629) );
  XNOR2_X1 U698 ( .A(n630), .B(n629), .ZN(n631) );
  XNOR2_X1 U699 ( .A(KEYINPUT74), .B(n631), .ZN(n956) );
  NAND2_X1 U700 ( .A1(n636), .A2(n956), .ZN(n635) );
  NOR2_X1 U701 ( .A1(G2067), .A2(n670), .ZN(n633) );
  INV_X1 U702 ( .A(n670), .ZN(n655) );
  NOR2_X1 U703 ( .A1(n655), .A2(G1348), .ZN(n632) );
  NOR2_X1 U704 ( .A1(n633), .A2(n632), .ZN(n634) );
  NAND2_X1 U705 ( .A1(n635), .A2(n634), .ZN(n640) );
  INV_X1 U706 ( .A(n636), .ZN(n638) );
  INV_X1 U707 ( .A(n956), .ZN(n637) );
  NAND2_X1 U708 ( .A1(n638), .A2(n637), .ZN(n639) );
  NAND2_X1 U709 ( .A1(n640), .A2(n639), .ZN(n646) );
  INV_X1 U710 ( .A(G299), .ZN(n648) );
  NAND2_X1 U711 ( .A1(n655), .A2(G2072), .ZN(n641) );
  XNOR2_X1 U712 ( .A(KEYINPUT27), .B(n641), .ZN(n644) );
  XOR2_X1 U713 ( .A(G1956), .B(KEYINPUT93), .Z(n988) );
  NAND2_X1 U714 ( .A1(n988), .A2(n670), .ZN(n642) );
  XOR2_X1 U715 ( .A(KEYINPUT94), .B(n642), .Z(n643) );
  NOR2_X1 U716 ( .A1(n644), .A2(n643), .ZN(n647) );
  NAND2_X1 U717 ( .A1(n648), .A2(n647), .ZN(n645) );
  NAND2_X1 U718 ( .A1(n646), .A2(n645), .ZN(n652) );
  NOR2_X1 U719 ( .A1(n648), .A2(n647), .ZN(n650) );
  XNOR2_X1 U720 ( .A(KEYINPUT95), .B(KEYINPUT28), .ZN(n649) );
  XNOR2_X1 U721 ( .A(n650), .B(n649), .ZN(n651) );
  NAND2_X1 U722 ( .A1(n652), .A2(n651), .ZN(n654) );
  XNOR2_X1 U723 ( .A(n654), .B(n653), .ZN(n658) );
  NAND2_X1 U724 ( .A1(G1961), .A2(n670), .ZN(n657) );
  XOR2_X1 U725 ( .A(G2078), .B(KEYINPUT25), .Z(n935) );
  NAND2_X1 U726 ( .A1(n655), .A2(n935), .ZN(n656) );
  NAND2_X1 U727 ( .A1(n657), .A2(n656), .ZN(n663) );
  NAND2_X1 U728 ( .A1(n658), .A2(n521), .ZN(n669) );
  NAND2_X2 U729 ( .A1(G8), .A2(n670), .ZN(n714) );
  NOR2_X1 U730 ( .A1(G1966), .A2(n714), .ZN(n681) );
  NOR2_X1 U731 ( .A1(G2084), .A2(n659), .ZN(n680) );
  NOR2_X1 U732 ( .A1(n681), .A2(n680), .ZN(n660) );
  NAND2_X1 U733 ( .A1(G8), .A2(n660), .ZN(n662) );
  NOR2_X1 U734 ( .A1(G168), .A2(n518), .ZN(n666) );
  NAND2_X1 U735 ( .A1(G301), .A2(n663), .ZN(n664) );
  XOR2_X1 U736 ( .A(KEYINPUT98), .B(n664), .Z(n665) );
  NAND2_X1 U737 ( .A1(n669), .A2(n668), .ZN(n683) );
  NAND2_X1 U738 ( .A1(n683), .A2(G286), .ZN(n677) );
  INV_X1 U739 ( .A(G8), .ZN(n675) );
  NOR2_X1 U740 ( .A1(G1971), .A2(n714), .ZN(n672) );
  NOR2_X1 U741 ( .A1(G2090), .A2(n670), .ZN(n671) );
  NOR2_X1 U742 ( .A1(n672), .A2(n671), .ZN(n673) );
  NAND2_X1 U743 ( .A1(n673), .A2(G303), .ZN(n674) );
  OR2_X1 U744 ( .A1(n675), .A2(n674), .ZN(n676) );
  AND2_X1 U745 ( .A1(G8), .A2(n680), .ZN(n682) );
  NAND2_X1 U746 ( .A1(n683), .A2(n519), .ZN(n702) );
  NOR2_X1 U747 ( .A1(G1976), .A2(G288), .ZN(n965) );
  INV_X1 U748 ( .A(n714), .ZN(n686) );
  NAND2_X1 U749 ( .A1(n965), .A2(n686), .ZN(n684) );
  NAND2_X1 U750 ( .A1(n684), .A2(KEYINPUT33), .ZN(n693) );
  INV_X1 U751 ( .A(n693), .ZN(n689) );
  INV_X1 U752 ( .A(KEYINPUT33), .ZN(n685) );
  NAND2_X1 U753 ( .A1(G1976), .A2(G288), .ZN(n959) );
  AND2_X1 U754 ( .A1(n685), .A2(n959), .ZN(n687) );
  AND2_X1 U755 ( .A1(n687), .A2(n686), .ZN(n688) );
  OR2_X1 U756 ( .A1(n689), .A2(n688), .ZN(n691) );
  AND2_X1 U757 ( .A1(n702), .A2(n691), .ZN(n690) );
  NAND2_X1 U758 ( .A1(n703), .A2(n690), .ZN(n698) );
  INV_X1 U759 ( .A(n691), .ZN(n696) );
  NOR2_X1 U760 ( .A1(G1971), .A2(G303), .ZN(n692) );
  NOR2_X1 U761 ( .A1(n692), .A2(n965), .ZN(n694) );
  AND2_X1 U762 ( .A1(n694), .A2(n693), .ZN(n695) );
  OR2_X1 U763 ( .A1(n696), .A2(n695), .ZN(n697) );
  NAND2_X1 U764 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U765 ( .A(n699), .B(KEYINPUT99), .ZN(n701) );
  XNOR2_X1 U766 ( .A(KEYINPUT100), .B(G1981), .ZN(n700) );
  XNOR2_X1 U767 ( .A(n700), .B(G305), .ZN(n953) );
  NOR2_X1 U768 ( .A1(n701), .A2(n953), .ZN(n710) );
  NAND2_X1 U769 ( .A1(n703), .A2(n702), .ZN(n706) );
  NOR2_X1 U770 ( .A1(G2090), .A2(G303), .ZN(n704) );
  NAND2_X1 U771 ( .A1(G8), .A2(n704), .ZN(n705) );
  NAND2_X1 U772 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U773 ( .A1(n714), .A2(n707), .ZN(n708) );
  XNOR2_X1 U774 ( .A(n708), .B(KEYINPUT101), .ZN(n709) );
  NOR2_X2 U775 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U776 ( .A(n711), .B(KEYINPUT102), .ZN(n717) );
  NOR2_X1 U777 ( .A1(G1981), .A2(G305), .ZN(n712) );
  XNOR2_X1 U778 ( .A(n712), .B(KEYINPUT91), .ZN(n713) );
  XNOR2_X1 U779 ( .A(n713), .B(KEYINPUT24), .ZN(n715) );
  NOR2_X1 U780 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U781 ( .A1(n717), .A2(n520), .ZN(n748) );
  NAND2_X1 U782 ( .A1(G140), .A2(n893), .ZN(n719) );
  NAND2_X1 U783 ( .A1(G104), .A2(n894), .ZN(n718) );
  NAND2_X1 U784 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U785 ( .A(KEYINPUT34), .B(n720), .ZN(n725) );
  NAND2_X1 U786 ( .A1(G128), .A2(n891), .ZN(n722) );
  NAND2_X1 U787 ( .A1(G116), .A2(n890), .ZN(n721) );
  NAND2_X1 U788 ( .A1(n722), .A2(n721), .ZN(n723) );
  XOR2_X1 U789 ( .A(KEYINPUT35), .B(n723), .Z(n724) );
  NOR2_X1 U790 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U791 ( .A(KEYINPUT36), .B(n726), .ZN(n873) );
  XNOR2_X1 U792 ( .A(KEYINPUT37), .B(G2067), .ZN(n762) );
  NOR2_X1 U793 ( .A1(n873), .A2(n762), .ZN(n1005) );
  NOR2_X1 U794 ( .A1(n728), .A2(n727), .ZN(n764) );
  NAND2_X1 U795 ( .A1(n1005), .A2(n764), .ZN(n729) );
  XOR2_X1 U796 ( .A(n729), .B(KEYINPUT88), .Z(n759) );
  NAND2_X1 U797 ( .A1(G105), .A2(n894), .ZN(n730) );
  XOR2_X1 U798 ( .A(KEYINPUT38), .B(n730), .Z(n735) );
  NAND2_X1 U799 ( .A1(G129), .A2(n891), .ZN(n732) );
  NAND2_X1 U800 ( .A1(G117), .A2(n890), .ZN(n731) );
  NAND2_X1 U801 ( .A1(n732), .A2(n731), .ZN(n733) );
  XOR2_X1 U802 ( .A(KEYINPUT89), .B(n733), .Z(n734) );
  NOR2_X1 U803 ( .A1(n735), .A2(n734), .ZN(n737) );
  NAND2_X1 U804 ( .A1(n893), .A2(G141), .ZN(n736) );
  NAND2_X1 U805 ( .A1(n737), .A2(n736), .ZN(n885) );
  AND2_X1 U806 ( .A1(n885), .A2(G1996), .ZN(n745) );
  NAND2_X1 U807 ( .A1(G131), .A2(n893), .ZN(n739) );
  NAND2_X1 U808 ( .A1(G95), .A2(n894), .ZN(n738) );
  NAND2_X1 U809 ( .A1(n739), .A2(n738), .ZN(n743) );
  NAND2_X1 U810 ( .A1(G119), .A2(n891), .ZN(n741) );
  NAND2_X1 U811 ( .A1(G107), .A2(n890), .ZN(n740) );
  NAND2_X1 U812 ( .A1(n741), .A2(n740), .ZN(n742) );
  NOR2_X1 U813 ( .A1(n743), .A2(n742), .ZN(n872) );
  INV_X1 U814 ( .A(G1991), .ZN(n842) );
  NOR2_X1 U815 ( .A1(n872), .A2(n842), .ZN(n744) );
  NOR2_X1 U816 ( .A1(n745), .A2(n744), .ZN(n1007) );
  INV_X1 U817 ( .A(n764), .ZN(n746) );
  NOR2_X1 U818 ( .A1(n1007), .A2(n746), .ZN(n755) );
  NOR2_X1 U819 ( .A1(n759), .A2(n755), .ZN(n747) );
  NAND2_X1 U820 ( .A1(n748), .A2(n747), .ZN(n749) );
  XNOR2_X1 U821 ( .A(n749), .B(KEYINPUT103), .ZN(n751) );
  XNOR2_X1 U822 ( .A(G1986), .B(G290), .ZN(n962) );
  NAND2_X1 U823 ( .A1(n962), .A2(n764), .ZN(n750) );
  NAND2_X1 U824 ( .A1(n751), .A2(n750), .ZN(n767) );
  NOR2_X1 U825 ( .A1(G1996), .A2(n885), .ZN(n1013) );
  NOR2_X1 U826 ( .A1(G1986), .A2(G290), .ZN(n752) );
  AND2_X1 U827 ( .A1(n842), .A2(n872), .ZN(n1009) );
  NOR2_X1 U828 ( .A1(n752), .A2(n1009), .ZN(n753) );
  XNOR2_X1 U829 ( .A(n753), .B(KEYINPUT104), .ZN(n754) );
  NOR2_X1 U830 ( .A1(n755), .A2(n754), .ZN(n756) );
  NOR2_X1 U831 ( .A1(n1013), .A2(n756), .ZN(n757) );
  XOR2_X1 U832 ( .A(KEYINPUT105), .B(n757), .Z(n758) );
  XNOR2_X1 U833 ( .A(n758), .B(KEYINPUT39), .ZN(n761) );
  INV_X1 U834 ( .A(n759), .ZN(n760) );
  NAND2_X1 U835 ( .A1(n761), .A2(n760), .ZN(n763) );
  NAND2_X1 U836 ( .A1(n873), .A2(n762), .ZN(n1010) );
  NAND2_X1 U837 ( .A1(n763), .A2(n1010), .ZN(n765) );
  NAND2_X1 U838 ( .A1(n765), .A2(n764), .ZN(n766) );
  NAND2_X1 U839 ( .A1(n767), .A2(n766), .ZN(n768) );
  XNOR2_X1 U840 ( .A(n768), .B(KEYINPUT40), .ZN(G329) );
  BUF_X1 U841 ( .A(n769), .Z(G160) );
  AND2_X1 U842 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U843 ( .A(G57), .ZN(G237) );
  INV_X1 U844 ( .A(G132), .ZN(G219) );
  INV_X1 U845 ( .A(G82), .ZN(G220) );
  XOR2_X1 U846 ( .A(KEYINPUT11), .B(KEYINPUT72), .Z(n772) );
  NAND2_X1 U847 ( .A1(G7), .A2(G661), .ZN(n770) );
  XOR2_X1 U848 ( .A(n770), .B(KEYINPUT10), .Z(n928) );
  NAND2_X1 U849 ( .A1(G567), .A2(n928), .ZN(n771) );
  XNOR2_X1 U850 ( .A(n772), .B(n771), .ZN(G234) );
  NAND2_X1 U851 ( .A1(n773), .A2(G860), .ZN(G153) );
  NOR2_X1 U852 ( .A1(G868), .A2(n956), .ZN(n774) );
  XOR2_X1 U853 ( .A(KEYINPUT76), .B(n774), .Z(n776) );
  NAND2_X1 U854 ( .A1(G868), .A2(G301), .ZN(n775) );
  NAND2_X1 U855 ( .A1(n776), .A2(n775), .ZN(G284) );
  XNOR2_X1 U856 ( .A(KEYINPUT77), .B(G868), .ZN(n777) );
  NOR2_X1 U857 ( .A1(G286), .A2(n777), .ZN(n779) );
  NOR2_X1 U858 ( .A1(G868), .A2(G299), .ZN(n778) );
  NOR2_X1 U859 ( .A1(n779), .A2(n778), .ZN(G297) );
  INV_X1 U860 ( .A(G860), .ZN(n780) );
  NAND2_X1 U861 ( .A1(n780), .A2(G559), .ZN(n781) );
  NAND2_X1 U862 ( .A1(n781), .A2(n956), .ZN(n782) );
  XNOR2_X1 U863 ( .A(n782), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U864 ( .A1(G868), .A2(n956), .ZN(n783) );
  NOR2_X1 U865 ( .A1(G559), .A2(n783), .ZN(n784) );
  XNOR2_X1 U866 ( .A(n784), .B(KEYINPUT78), .ZN(n786) );
  NOR2_X1 U867 ( .A1(n971), .A2(G868), .ZN(n785) );
  NOR2_X1 U868 ( .A1(n786), .A2(n785), .ZN(G282) );
  NAND2_X1 U869 ( .A1(G111), .A2(n890), .ZN(n788) );
  NAND2_X1 U870 ( .A1(G99), .A2(n894), .ZN(n787) );
  NAND2_X1 U871 ( .A1(n788), .A2(n787), .ZN(n789) );
  XNOR2_X1 U872 ( .A(n789), .B(KEYINPUT79), .ZN(n791) );
  NAND2_X1 U873 ( .A1(G135), .A2(n893), .ZN(n790) );
  NAND2_X1 U874 ( .A1(n791), .A2(n790), .ZN(n794) );
  NAND2_X1 U875 ( .A1(n891), .A2(G123), .ZN(n792) );
  XOR2_X1 U876 ( .A(KEYINPUT18), .B(n792), .Z(n793) );
  NOR2_X1 U877 ( .A1(n794), .A2(n793), .ZN(n1004) );
  XNOR2_X1 U878 ( .A(G2096), .B(n1004), .ZN(n795) );
  INV_X1 U879 ( .A(G2100), .ZN(n859) );
  NAND2_X1 U880 ( .A1(n795), .A2(n859), .ZN(G156) );
  NAND2_X1 U881 ( .A1(G93), .A2(n796), .ZN(n799) );
  NAND2_X1 U882 ( .A1(G80), .A2(n797), .ZN(n798) );
  NAND2_X1 U883 ( .A1(n799), .A2(n798), .ZN(n806) );
  NAND2_X1 U884 ( .A1(G55), .A2(n800), .ZN(n801) );
  XNOR2_X1 U885 ( .A(n801), .B(KEYINPUT80), .ZN(n804) );
  NAND2_X1 U886 ( .A1(G67), .A2(n802), .ZN(n803) );
  NAND2_X1 U887 ( .A1(n804), .A2(n803), .ZN(n805) );
  NOR2_X1 U888 ( .A1(n806), .A2(n805), .ZN(n810) );
  NAND2_X1 U889 ( .A1(G559), .A2(n956), .ZN(n818) );
  XNOR2_X1 U890 ( .A(n971), .B(n818), .ZN(n807) );
  NOR2_X1 U891 ( .A1(G860), .A2(n807), .ZN(n808) );
  XNOR2_X1 U892 ( .A(n810), .B(n808), .ZN(G145) );
  NOR2_X1 U893 ( .A1(G868), .A2(n810), .ZN(n809) );
  XNOR2_X1 U894 ( .A(n809), .B(KEYINPUT85), .ZN(n821) );
  XOR2_X1 U895 ( .A(KEYINPUT19), .B(KEYINPUT84), .Z(n812) );
  XOR2_X1 U896 ( .A(G303), .B(n810), .Z(n811) );
  XNOR2_X1 U897 ( .A(n812), .B(n811), .ZN(n815) );
  XOR2_X1 U898 ( .A(n971), .B(G305), .Z(n813) );
  XNOR2_X1 U899 ( .A(n813), .B(G288), .ZN(n814) );
  XNOR2_X1 U900 ( .A(n815), .B(n814), .ZN(n817) );
  XOR2_X1 U901 ( .A(G290), .B(G299), .Z(n816) );
  XNOR2_X1 U902 ( .A(n817), .B(n816), .ZN(n907) );
  XNOR2_X1 U903 ( .A(n907), .B(n818), .ZN(n819) );
  NAND2_X1 U904 ( .A1(G868), .A2(n819), .ZN(n820) );
  NAND2_X1 U905 ( .A1(n821), .A2(n820), .ZN(G295) );
  NAND2_X1 U906 ( .A1(G2078), .A2(G2084), .ZN(n822) );
  XOR2_X1 U907 ( .A(KEYINPUT20), .B(n822), .Z(n823) );
  NAND2_X1 U908 ( .A1(G2090), .A2(n823), .ZN(n824) );
  XNOR2_X1 U909 ( .A(KEYINPUT21), .B(n824), .ZN(n825) );
  NAND2_X1 U910 ( .A1(n825), .A2(G2072), .ZN(n826) );
  XNOR2_X1 U911 ( .A(KEYINPUT86), .B(n826), .ZN(G158) );
  XNOR2_X1 U912 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U913 ( .A1(G220), .A2(G219), .ZN(n827) );
  XOR2_X1 U914 ( .A(KEYINPUT22), .B(n827), .Z(n828) );
  NOR2_X1 U915 ( .A1(G218), .A2(n828), .ZN(n829) );
  NAND2_X1 U916 ( .A1(G96), .A2(n829), .ZN(n839) );
  NAND2_X1 U917 ( .A1(n839), .A2(G2106), .ZN(n833) );
  NAND2_X1 U918 ( .A1(G69), .A2(G120), .ZN(n830) );
  NOR2_X1 U919 ( .A1(G237), .A2(n830), .ZN(n831) );
  NAND2_X1 U920 ( .A1(G108), .A2(n831), .ZN(n840) );
  NAND2_X1 U921 ( .A1(n840), .A2(G567), .ZN(n832) );
  NAND2_X1 U922 ( .A1(n833), .A2(n832), .ZN(n841) );
  NAND2_X1 U923 ( .A1(G661), .A2(G483), .ZN(n834) );
  NOR2_X1 U924 ( .A1(n841), .A2(n834), .ZN(n836) );
  NAND2_X1 U925 ( .A1(n836), .A2(G36), .ZN(G176) );
  NAND2_X1 U926 ( .A1(G2106), .A2(n928), .ZN(G217) );
  AND2_X1 U927 ( .A1(G15), .A2(G2), .ZN(n835) );
  NAND2_X1 U928 ( .A1(G661), .A2(n835), .ZN(G259) );
  NAND2_X1 U929 ( .A1(G1), .A2(G3), .ZN(n837) );
  NAND2_X1 U930 ( .A1(n837), .A2(n836), .ZN(n838) );
  XNOR2_X1 U931 ( .A(n838), .B(KEYINPUT108), .ZN(G188) );
  XNOR2_X1 U932 ( .A(G96), .B(KEYINPUT109), .ZN(G221) );
  NOR2_X1 U933 ( .A1(n840), .A2(n839), .ZN(G325) );
  XOR2_X1 U934 ( .A(KEYINPUT110), .B(G325), .Z(G261) );
  INV_X1 U936 ( .A(G120), .ZN(G236) );
  INV_X1 U937 ( .A(G69), .ZN(G235) );
  INV_X1 U938 ( .A(n841), .ZN(G319) );
  XOR2_X1 U939 ( .A(G2474), .B(G1981), .Z(n844) );
  XOR2_X1 U940 ( .A(G1996), .B(n842), .Z(n843) );
  XNOR2_X1 U941 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U942 ( .A(n845), .B(KEYINPUT112), .Z(n847) );
  XNOR2_X1 U943 ( .A(G1976), .B(G1956), .ZN(n846) );
  XNOR2_X1 U944 ( .A(n847), .B(n846), .ZN(n851) );
  XOR2_X1 U945 ( .A(G1961), .B(G1966), .Z(n849) );
  XNOR2_X1 U946 ( .A(G1986), .B(G1971), .ZN(n848) );
  XNOR2_X1 U947 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U948 ( .A(n851), .B(n850), .Z(n853) );
  XNOR2_X1 U949 ( .A(KEYINPUT113), .B(KEYINPUT41), .ZN(n852) );
  XNOR2_X1 U950 ( .A(n853), .B(n852), .ZN(G229) );
  XOR2_X1 U951 ( .A(KEYINPUT42), .B(G2090), .Z(n855) );
  XNOR2_X1 U952 ( .A(G2067), .B(G2078), .ZN(n854) );
  XNOR2_X1 U953 ( .A(n855), .B(n854), .ZN(n856) );
  XOR2_X1 U954 ( .A(n856), .B(G2096), .Z(n858) );
  XNOR2_X1 U955 ( .A(G2072), .B(G2084), .ZN(n857) );
  XNOR2_X1 U956 ( .A(n858), .B(n857), .ZN(n863) );
  XOR2_X1 U957 ( .A(KEYINPUT43), .B(KEYINPUT111), .Z(n861) );
  XOR2_X1 U958 ( .A(G2678), .B(n859), .Z(n860) );
  XNOR2_X1 U959 ( .A(n861), .B(n860), .ZN(n862) );
  XOR2_X1 U960 ( .A(n863), .B(n862), .Z(G227) );
  NAND2_X1 U961 ( .A1(n893), .A2(G136), .ZN(n870) );
  NAND2_X1 U962 ( .A1(G112), .A2(n890), .ZN(n865) );
  NAND2_X1 U963 ( .A1(G100), .A2(n894), .ZN(n864) );
  NAND2_X1 U964 ( .A1(n865), .A2(n864), .ZN(n868) );
  NAND2_X1 U965 ( .A1(n891), .A2(G124), .ZN(n866) );
  XOR2_X1 U966 ( .A(KEYINPUT44), .B(n866), .Z(n867) );
  NOR2_X1 U967 ( .A1(n868), .A2(n867), .ZN(n869) );
  NAND2_X1 U968 ( .A1(n870), .A2(n869), .ZN(n871) );
  XOR2_X1 U969 ( .A(KEYINPUT114), .B(n871), .Z(G162) );
  XNOR2_X1 U970 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n875) );
  XNOR2_X1 U971 ( .A(n873), .B(n872), .ZN(n874) );
  XNOR2_X1 U972 ( .A(n875), .B(n874), .ZN(n884) );
  NAND2_X1 U973 ( .A1(G139), .A2(n893), .ZN(n877) );
  NAND2_X1 U974 ( .A1(G103), .A2(n894), .ZN(n876) );
  NAND2_X1 U975 ( .A1(n877), .A2(n876), .ZN(n878) );
  XOR2_X1 U976 ( .A(KEYINPUT117), .B(n878), .Z(n883) );
  NAND2_X1 U977 ( .A1(G127), .A2(n891), .ZN(n880) );
  NAND2_X1 U978 ( .A1(G115), .A2(n890), .ZN(n879) );
  NAND2_X1 U979 ( .A1(n880), .A2(n879), .ZN(n881) );
  XOR2_X1 U980 ( .A(KEYINPUT47), .B(n881), .Z(n882) );
  NOR2_X1 U981 ( .A1(n883), .A2(n882), .ZN(n1019) );
  XOR2_X1 U982 ( .A(n884), .B(n1019), .Z(n887) );
  XOR2_X1 U983 ( .A(G164), .B(n885), .Z(n886) );
  XNOR2_X1 U984 ( .A(n887), .B(n886), .ZN(n888) );
  XNOR2_X1 U985 ( .A(n888), .B(G160), .ZN(n889) );
  XNOR2_X1 U986 ( .A(n889), .B(G162), .ZN(n905) );
  NAND2_X1 U987 ( .A1(G118), .A2(n890), .ZN(n902) );
  NAND2_X1 U988 ( .A1(n891), .A2(G130), .ZN(n892) );
  XNOR2_X1 U989 ( .A(KEYINPUT115), .B(n892), .ZN(n900) );
  NAND2_X1 U990 ( .A1(G142), .A2(n893), .ZN(n896) );
  NAND2_X1 U991 ( .A1(G106), .A2(n894), .ZN(n895) );
  NAND2_X1 U992 ( .A1(n896), .A2(n895), .ZN(n897) );
  XOR2_X1 U993 ( .A(KEYINPUT116), .B(n897), .Z(n898) );
  XNOR2_X1 U994 ( .A(KEYINPUT45), .B(n898), .ZN(n899) );
  NOR2_X1 U995 ( .A1(n900), .A2(n899), .ZN(n901) );
  NAND2_X1 U996 ( .A1(n902), .A2(n901), .ZN(n903) );
  XNOR2_X1 U997 ( .A(n903), .B(n1004), .ZN(n904) );
  XNOR2_X1 U998 ( .A(n905), .B(n904), .ZN(n906) );
  NOR2_X1 U999 ( .A1(G37), .A2(n906), .ZN(G395) );
  XOR2_X1 U1000 ( .A(n956), .B(G286), .Z(n908) );
  XNOR2_X1 U1001 ( .A(n908), .B(n907), .ZN(n909) );
  XOR2_X1 U1002 ( .A(n909), .B(G301), .Z(n910) );
  NOR2_X1 U1003 ( .A1(G37), .A2(n910), .ZN(G397) );
  XNOR2_X1 U1004 ( .A(G2451), .B(G2427), .ZN(n920) );
  XOR2_X1 U1005 ( .A(G2430), .B(G2443), .Z(n912) );
  XNOR2_X1 U1006 ( .A(KEYINPUT107), .B(G2435), .ZN(n911) );
  XNOR2_X1 U1007 ( .A(n912), .B(n911), .ZN(n916) );
  XOR2_X1 U1008 ( .A(G2438), .B(G2454), .Z(n914) );
  XNOR2_X1 U1009 ( .A(G1348), .B(G1341), .ZN(n913) );
  XNOR2_X1 U1010 ( .A(n914), .B(n913), .ZN(n915) );
  XOR2_X1 U1011 ( .A(n916), .B(n915), .Z(n918) );
  XNOR2_X1 U1012 ( .A(G2446), .B(KEYINPUT106), .ZN(n917) );
  XNOR2_X1 U1013 ( .A(n918), .B(n917), .ZN(n919) );
  XNOR2_X1 U1014 ( .A(n920), .B(n919), .ZN(n921) );
  NAND2_X1 U1015 ( .A1(n921), .A2(G14), .ZN(n927) );
  NAND2_X1 U1016 ( .A1(G319), .A2(n927), .ZN(n924) );
  NOR2_X1 U1017 ( .A1(G229), .A2(G227), .ZN(n922) );
  XNOR2_X1 U1018 ( .A(KEYINPUT49), .B(n922), .ZN(n923) );
  NOR2_X1 U1019 ( .A1(n924), .A2(n923), .ZN(n926) );
  NOR2_X1 U1020 ( .A1(G395), .A2(G397), .ZN(n925) );
  NAND2_X1 U1021 ( .A1(n926), .A2(n925), .ZN(G225) );
  INV_X1 U1022 ( .A(G225), .ZN(G308) );
  INV_X1 U1023 ( .A(G108), .ZN(G238) );
  INV_X1 U1024 ( .A(n927), .ZN(G401) );
  INV_X1 U1025 ( .A(n928), .ZN(G223) );
  XOR2_X1 U1026 ( .A(G29), .B(KEYINPUT122), .Z(n949) );
  XOR2_X1 U1027 ( .A(G2067), .B(G26), .Z(n930) );
  XOR2_X1 U1028 ( .A(G1996), .B(G32), .Z(n929) );
  NAND2_X1 U1029 ( .A1(n930), .A2(n929), .ZN(n932) );
  XNOR2_X1 U1030 ( .A(G33), .B(G2072), .ZN(n931) );
  NOR2_X1 U1031 ( .A1(n932), .A2(n931), .ZN(n940) );
  XOR2_X1 U1032 ( .A(G1991), .B(G25), .Z(n933) );
  NAND2_X1 U1033 ( .A1(n933), .A2(G28), .ZN(n934) );
  XNOR2_X1 U1034 ( .A(n934), .B(KEYINPUT120), .ZN(n938) );
  XOR2_X1 U1035 ( .A(n935), .B(G27), .Z(n936) );
  XNOR2_X1 U1036 ( .A(KEYINPUT121), .B(n936), .ZN(n937) );
  NOR2_X1 U1037 ( .A1(n938), .A2(n937), .ZN(n939) );
  NAND2_X1 U1038 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1039 ( .A(n941), .B(KEYINPUT53), .ZN(n944) );
  XOR2_X1 U1040 ( .A(G2084), .B(KEYINPUT54), .Z(n942) );
  XNOR2_X1 U1041 ( .A(G34), .B(n942), .ZN(n943) );
  NAND2_X1 U1042 ( .A1(n944), .A2(n943), .ZN(n946) );
  XNOR2_X1 U1043 ( .A(G35), .B(G2090), .ZN(n945) );
  NOR2_X1 U1044 ( .A1(n946), .A2(n945), .ZN(n947) );
  INV_X1 U1045 ( .A(KEYINPUT55), .ZN(n1027) );
  XOR2_X1 U1046 ( .A(n947), .B(n1027), .Z(n948) );
  NAND2_X1 U1047 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1048 ( .A1(n950), .A2(G11), .ZN(n951) );
  XNOR2_X1 U1049 ( .A(n951), .B(KEYINPUT123), .ZN(n1034) );
  INV_X1 U1050 ( .A(G16), .ZN(n1001) );
  XOR2_X1 U1051 ( .A(n1001), .B(KEYINPUT56), .Z(n977) );
  XOR2_X1 U1052 ( .A(G1966), .B(G168), .Z(n952) );
  NOR2_X1 U1053 ( .A1(n953), .A2(n952), .ZN(n954) );
  XOR2_X1 U1054 ( .A(KEYINPUT57), .B(n954), .Z(n975) );
  XOR2_X1 U1055 ( .A(G303), .B(G1971), .Z(n955) );
  XNOR2_X1 U1056 ( .A(n955), .B(KEYINPUT125), .ZN(n958) );
  XOR2_X1 U1057 ( .A(G1348), .B(n956), .Z(n957) );
  NOR2_X1 U1058 ( .A1(n958), .A2(n957), .ZN(n964) );
  XOR2_X1 U1059 ( .A(G1961), .B(G301), .Z(n960) );
  NAND2_X1 U1060 ( .A1(n960), .A2(n959), .ZN(n961) );
  NOR2_X1 U1061 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1062 ( .A1(n964), .A2(n963), .ZN(n969) );
  XOR2_X1 U1063 ( .A(n965), .B(KEYINPUT124), .Z(n967) );
  XOR2_X1 U1064 ( .A(G1956), .B(G299), .Z(n966) );
  NAND2_X1 U1065 ( .A1(n967), .A2(n966), .ZN(n968) );
  NOR2_X1 U1066 ( .A1(n969), .A2(n968), .ZN(n970) );
  XOR2_X1 U1067 ( .A(KEYINPUT126), .B(n970), .Z(n973) );
  XNOR2_X1 U1068 ( .A(n971), .B(G1341), .ZN(n972) );
  NOR2_X1 U1069 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1070 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1071 ( .A1(n977), .A2(n976), .ZN(n1003) );
  XOR2_X1 U1072 ( .A(G1976), .B(G23), .Z(n979) );
  XOR2_X1 U1073 ( .A(G1971), .B(G22), .Z(n978) );
  NAND2_X1 U1074 ( .A1(n979), .A2(n978), .ZN(n981) );
  XNOR2_X1 U1075 ( .A(G24), .B(G1986), .ZN(n980) );
  NOR2_X1 U1076 ( .A1(n981), .A2(n980), .ZN(n982) );
  XOR2_X1 U1077 ( .A(KEYINPUT58), .B(n982), .Z(n998) );
  XOR2_X1 U1078 ( .A(G1961), .B(G5), .Z(n993) );
  XNOR2_X1 U1079 ( .A(G1348), .B(KEYINPUT59), .ZN(n983) );
  XNOR2_X1 U1080 ( .A(n983), .B(G4), .ZN(n987) );
  XNOR2_X1 U1081 ( .A(G1981), .B(G6), .ZN(n985) );
  XNOR2_X1 U1082 ( .A(G1341), .B(G19), .ZN(n984) );
  NOR2_X1 U1083 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1084 ( .A1(n987), .A2(n986), .ZN(n990) );
  XNOR2_X1 U1085 ( .A(G20), .B(n988), .ZN(n989) );
  NOR2_X1 U1086 ( .A1(n990), .A2(n989), .ZN(n991) );
  XNOR2_X1 U1087 ( .A(KEYINPUT60), .B(n991), .ZN(n992) );
  NAND2_X1 U1088 ( .A1(n993), .A2(n992), .ZN(n995) );
  XNOR2_X1 U1089 ( .A(G21), .B(G1966), .ZN(n994) );
  NOR2_X1 U1090 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1091 ( .A(KEYINPUT127), .B(n996), .ZN(n997) );
  NOR2_X1 U1092 ( .A1(n998), .A2(n997), .ZN(n999) );
  XNOR2_X1 U1093 ( .A(KEYINPUT61), .B(n999), .ZN(n1000) );
  NAND2_X1 U1094 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1095 ( .A1(n1003), .A2(n1002), .ZN(n1032) );
  NOR2_X1 U1096 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1097 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NOR2_X1 U1098 ( .A1(n1009), .A2(n1008), .ZN(n1018) );
  XNOR2_X1 U1099 ( .A(G2084), .B(G160), .ZN(n1011) );
  NAND2_X1 U1100 ( .A1(n1011), .A2(n1010), .ZN(n1016) );
  XOR2_X1 U1101 ( .A(G2090), .B(G162), .Z(n1012) );
  NOR2_X1 U1102 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1103 ( .A(n1014), .B(KEYINPUT51), .ZN(n1015) );
  NOR2_X1 U1104 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1105 ( .A1(n1018), .A2(n1017), .ZN(n1025) );
  XOR2_X1 U1106 ( .A(G2072), .B(n1019), .Z(n1021) );
  XOR2_X1 U1107 ( .A(G164), .B(G2078), .Z(n1020) );
  NOR2_X1 U1108 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XOR2_X1 U1109 ( .A(KEYINPUT50), .B(n1022), .Z(n1023) );
  XNOR2_X1 U1110 ( .A(KEYINPUT118), .B(n1023), .ZN(n1024) );
  NOR2_X1 U1111 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XNOR2_X1 U1112 ( .A(n1026), .B(KEYINPUT52), .ZN(n1028) );
  NAND2_X1 U1113 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NAND2_X1 U1114 ( .A1(G29), .A2(n1029), .ZN(n1030) );
  XNOR2_X1 U1115 ( .A(KEYINPUT119), .B(n1030), .ZN(n1031) );
  NOR2_X1 U1116 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  NAND2_X1 U1117 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  XNOR2_X1 U1118 ( .A(KEYINPUT62), .B(n1035), .ZN(G150) );
  INV_X1 U1119 ( .A(G150), .ZN(G311) );
endmodule

