//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 1 0 0 0 1 1 0 0 1 0 0 1 0 1 1 0 0 1 0 0 1 1 0 0 0 1 0 1 0 0 1 0 0 1 0 0 1 1 1 1 1 0 1 1 1 1 0 0 1 1 0 1 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:43 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n446, new_n448, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n570, new_n571, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n636, new_n638, new_n639, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n845, new_n846, new_n847, new_n848, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n939, new_n940, new_n941, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1186, new_n1187, new_n1188;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT64), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT65), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT66), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  NAND2_X1  g020(.A1(G94), .A2(G452), .ZN(new_n446));
  XNOR2_X1  g021(.A(new_n446), .B(KEYINPUT67), .ZN(G173));
  XNOR2_X1  g022(.A(KEYINPUT68), .B(KEYINPUT1), .ZN(new_n448));
  AND2_X1   g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n448), .B(new_n449), .ZN(G223));
  NAND2_X1  g025(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n449), .A2(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  XOR2_X1   g032(.A(G325), .B(KEYINPUT69), .Z(G261));
  AND2_X1   g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  INV_X1    g034(.A(KEYINPUT70), .ZN(new_n460));
  OR2_X1    g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  AOI22_X1  g036(.A1(new_n459), .A2(new_n460), .B1(G567), .B2(new_n456), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  OR2_X1    g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(G2105), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  AOI22_X1  g044(.A1(new_n467), .A2(G137), .B1(G101), .B2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G125), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n471), .B1(new_n465), .B2(new_n466), .ZN(new_n472));
  AND2_X1   g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  OAI21_X1  g048(.A(G2105), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  AND2_X1   g049(.A1(new_n470), .A2(new_n474), .ZN(G160));
  NAND2_X1  g050(.A1(new_n467), .A2(G136), .ZN(new_n476));
  XOR2_X1   g051(.A(new_n476), .B(KEYINPUT71), .Z(new_n477));
  AND2_X1   g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  NOR2_X1   g053(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(G2105), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NOR2_X1   g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n483), .B(KEYINPUT72), .ZN(new_n484));
  INV_X1    g059(.A(G112), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n468), .B1(new_n485), .B2(G2105), .ZN(new_n486));
  AOI22_X1  g061(.A1(G124), .A2(new_n482), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  AND2_X1   g062(.A1(new_n477), .A2(new_n487), .ZN(G162));
  XNOR2_X1  g063(.A(KEYINPUT3), .B(G2104), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n489), .A2(G126), .A3(G2105), .ZN(new_n490));
  OR2_X1    g065(.A1(G102), .A2(G2105), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n491), .B(G2104), .C1(G114), .C2(new_n481), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  OAI211_X1 g068(.A(G138), .B(new_n481), .C1(new_n478), .C2(new_n479), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT73), .ZN(new_n495));
  OR2_X1    g070(.A1(new_n495), .A2(KEYINPUT4), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n489), .A2(G138), .A3(new_n496), .A4(new_n481), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n495), .A2(KEYINPUT4), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n493), .B1(new_n500), .B2(new_n501), .ZN(G164));
  NAND2_X1  g077(.A1(KEYINPUT74), .A2(KEYINPUT5), .ZN(new_n503));
  INV_X1    g078(.A(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g080(.A1(KEYINPUT74), .A2(KEYINPUT5), .A3(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n507), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n508));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  OR2_X1    g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n504), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G50), .ZN(new_n514));
  INV_X1    g089(.A(G88), .ZN(new_n515));
  AND3_X1   g090(.A1(KEYINPUT74), .A2(KEYINPUT5), .A3(G543), .ZN(new_n516));
  AOI21_X1  g091(.A(G543), .B1(KEYINPUT74), .B2(KEYINPUT5), .ZN(new_n517));
  AND2_X1   g092(.A1(KEYINPUT6), .A2(G651), .ZN(new_n518));
  NOR2_X1   g093(.A1(KEYINPUT6), .A2(G651), .ZN(new_n519));
  OAI22_X1  g094(.A1(new_n516), .A2(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n514), .B1(new_n515), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n510), .A2(new_n521), .ZN(G166));
  INV_X1    g097(.A(KEYINPUT77), .ZN(new_n523));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(KEYINPUT7), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT7), .ZN(new_n526));
  NAND4_X1  g101(.A1(new_n526), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(G89), .ZN(new_n529));
  OAI211_X1 g104(.A(KEYINPUT76), .B(new_n528), .C1(new_n520), .C2(new_n529), .ZN(new_n530));
  XOR2_X1   g105(.A(KEYINPUT75), .B(G51), .Z(new_n531));
  AND2_X1   g106(.A1(G63), .A2(G651), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n513), .A2(new_n531), .B1(new_n507), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n530), .A2(new_n533), .ZN(new_n534));
  XNOR2_X1  g109(.A(KEYINPUT6), .B(G651), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n507), .A2(G89), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g111(.A(KEYINPUT76), .B1(new_n536), .B2(new_n528), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n523), .B1(new_n534), .B2(new_n537), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n528), .B1(new_n520), .B2(new_n529), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT76), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND4_X1  g116(.A1(new_n541), .A2(KEYINPUT77), .A3(new_n530), .A4(new_n533), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n538), .A2(new_n542), .ZN(G168));
  INV_X1    g118(.A(G64), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n544), .B1(new_n505), .B2(new_n506), .ZN(new_n545));
  NAND2_X1  g120(.A1(G77), .A2(G543), .ZN(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(new_n547));
  OAI21_X1  g122(.A(KEYINPUT78), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(KEYINPUT78), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n516), .A2(new_n517), .ZN(new_n550));
  OAI211_X1 g125(.A(new_n549), .B(new_n546), .C1(new_n550), .C2(new_n544), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n548), .A2(new_n551), .A3(G651), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n505), .A2(new_n506), .B1(new_n511), .B2(new_n512), .ZN(new_n553));
  AOI22_X1  g128(.A1(new_n553), .A2(G90), .B1(new_n513), .B2(G52), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n552), .A2(new_n554), .ZN(G301));
  INV_X1    g130(.A(G301), .ZN(G171));
  INV_X1    g131(.A(G56), .ZN(new_n557));
  AOI21_X1  g132(.A(new_n557), .B1(new_n505), .B2(new_n506), .ZN(new_n558));
  NAND2_X1  g133(.A1(G68), .A2(G543), .ZN(new_n559));
  INV_X1    g134(.A(new_n559), .ZN(new_n560));
  OAI21_X1  g135(.A(KEYINPUT79), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT79), .ZN(new_n562));
  OAI211_X1 g137(.A(new_n562), .B(new_n559), .C1(new_n550), .C2(new_n557), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n561), .A2(new_n563), .A3(G651), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n553), .A2(G81), .B1(new_n513), .B2(G43), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G860), .ZN(G153));
  NAND4_X1  g143(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g144(.A1(G1), .A2(G3), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT8), .ZN(new_n571));
  NAND4_X1  g146(.A1(G319), .A2(G483), .A3(G661), .A4(new_n571), .ZN(G188));
  NAND2_X1  g147(.A1(G78), .A2(G543), .ZN(new_n573));
  INV_X1    g148(.A(G65), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n573), .B1(new_n550), .B2(new_n574), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n575), .A2(G651), .B1(new_n553), .B2(G91), .ZN(new_n576));
  AND2_X1   g151(.A1(KEYINPUT80), .A2(G53), .ZN(new_n577));
  OAI211_X1 g152(.A(G543), .B(new_n577), .C1(new_n518), .C2(new_n519), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n578), .A2(KEYINPUT9), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT9), .ZN(new_n580));
  NAND4_X1  g155(.A1(new_n535), .A2(new_n580), .A3(G543), .A4(new_n577), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n579), .A2(new_n581), .A3(KEYINPUT81), .ZN(new_n582));
  INV_X1    g157(.A(new_n582), .ZN(new_n583));
  AOI21_X1  g158(.A(KEYINPUT81), .B1(new_n579), .B2(new_n581), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n576), .B1(new_n583), .B2(new_n584), .ZN(G299));
  INV_X1    g160(.A(G168), .ZN(G286));
  INV_X1    g161(.A(G166), .ZN(G303));
  AOI22_X1  g162(.A1(new_n553), .A2(G87), .B1(new_n513), .B2(G49), .ZN(new_n588));
  OAI21_X1  g163(.A(G651), .B1(new_n507), .B2(G74), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n588), .A2(new_n589), .ZN(G288));
  AOI22_X1  g165(.A1(new_n507), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n591), .A2(new_n509), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n513), .A2(G48), .ZN(new_n593));
  INV_X1    g168(.A(G86), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n594), .B2(new_n520), .ZN(new_n595));
  OR2_X1    g170(.A1(new_n592), .A2(new_n595), .ZN(G305));
  AOI22_X1  g171(.A1(new_n507), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n597), .A2(new_n509), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n513), .A2(G47), .ZN(new_n599));
  INV_X1    g174(.A(G85), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n600), .B2(new_n520), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(new_n602), .ZN(G290));
  NAND2_X1  g178(.A1(G301), .A2(G868), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT82), .ZN(new_n605));
  OAI21_X1  g180(.A(G66), .B1(new_n516), .B2(new_n517), .ZN(new_n606));
  NAND2_X1  g181(.A1(G79), .A2(G543), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n509), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  OAI211_X1 g183(.A(G54), .B(G543), .C1(new_n518), .C2(new_n519), .ZN(new_n609));
  INV_X1    g184(.A(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n605), .B1(new_n608), .B2(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(G66), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n612), .B1(new_n505), .B2(new_n506), .ZN(new_n613));
  INV_X1    g188(.A(new_n607), .ZN(new_n614));
  OAI21_X1  g189(.A(G651), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n615), .A2(KEYINPUT82), .A3(new_n609), .ZN(new_n616));
  INV_X1    g191(.A(KEYINPUT10), .ZN(new_n617));
  INV_X1    g192(.A(G92), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n520), .B2(new_n618), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n553), .A2(KEYINPUT10), .A3(G92), .ZN(new_n620));
  AOI22_X1  g195(.A1(new_n611), .A2(new_n616), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n604), .B1(new_n621), .B2(G868), .ZN(G284));
  OAI21_X1  g197(.A(new_n604), .B1(new_n621), .B2(G868), .ZN(G321));
  NAND2_X1  g198(.A1(new_n553), .A2(G91), .ZN(new_n624));
  AOI22_X1  g199(.A1(new_n507), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n624), .B1(new_n625), .B2(new_n509), .ZN(new_n626));
  INV_X1    g201(.A(KEYINPUT81), .ZN(new_n627));
  AOI21_X1  g202(.A(new_n580), .B1(new_n513), .B2(new_n577), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n578), .A2(KEYINPUT9), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n627), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n626), .B1(new_n630), .B2(new_n582), .ZN(new_n631));
  OAI21_X1  g206(.A(KEYINPUT83), .B1(new_n631), .B2(G868), .ZN(new_n632));
  NAND2_X1  g207(.A1(G286), .A2(G868), .ZN(new_n633));
  MUX2_X1   g208(.A(KEYINPUT83), .B(new_n632), .S(new_n633), .Z(G297));
  MUX2_X1   g209(.A(KEYINPUT83), .B(new_n632), .S(new_n633), .Z(G280));
  INV_X1    g210(.A(G559), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n621), .B1(new_n636), .B2(G860), .ZN(G148));
  NAND2_X1  g212(.A1(new_n621), .A2(new_n636), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n638), .A2(G868), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n639), .B1(G868), .B2(new_n567), .ZN(G323));
  XNOR2_X1  g215(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g216(.A1(new_n489), .A2(new_n469), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT12), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2100), .ZN(new_n644));
  XOR2_X1   g219(.A(KEYINPUT84), .B(KEYINPUT13), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n467), .A2(G135), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n647), .B(KEYINPUT85), .Z(new_n648));
  NAND2_X1  g223(.A1(new_n482), .A2(G123), .ZN(new_n649));
  NOR2_X1   g224(.A1(new_n481), .A2(G111), .ZN(new_n650));
  OAI21_X1  g225(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n651));
  OAI211_X1 g226(.A(new_n648), .B(new_n649), .C1(new_n650), .C2(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(KEYINPUT86), .Z(new_n653));
  AND2_X1   g228(.A1(new_n653), .A2(G2096), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n653), .A2(G2096), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n646), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n656), .B(KEYINPUT87), .Z(G156));
  XNOR2_X1  g232(.A(G2427), .B(G2438), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(G2430), .ZN(new_n659));
  XNOR2_X1  g234(.A(KEYINPUT15), .B(G2435), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n659), .A2(new_n660), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n661), .A2(new_n662), .A3(KEYINPUT14), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1341), .B(G1348), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2443), .B(G2446), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n663), .B(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G2451), .B(G2454), .Z(new_n668));
  XNOR2_X1  g243(.A(KEYINPUT88), .B(KEYINPUT16), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  OR2_X1    g245(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n667), .A2(new_n670), .ZN(new_n672));
  AND3_X1   g247(.A1(new_n671), .A2(G14), .A3(new_n672), .ZN(G401));
  XOR2_X1   g248(.A(G2084), .B(G2090), .Z(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G2067), .B(G2678), .ZN(new_n676));
  XNOR2_X1  g251(.A(G2072), .B(G2078), .ZN(new_n677));
  OAI21_X1  g252(.A(new_n675), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(KEYINPUT17), .ZN(new_n679));
  AOI21_X1  g254(.A(new_n678), .B1(new_n679), .B2(new_n676), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT89), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n674), .A2(new_n676), .A3(new_n677), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT18), .ZN(new_n683));
  NOR3_X1   g258(.A1(new_n679), .A2(new_n676), .A3(new_n675), .ZN(new_n684));
  NOR3_X1   g259(.A1(new_n681), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G2096), .B(G2100), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(G227));
  XOR2_X1   g262(.A(G1971), .B(G1976), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT19), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1956), .B(G2474), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1961), .B(G1966), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT20), .ZN(new_n694));
  AND2_X1   g269(.A1(new_n690), .A2(new_n691), .ZN(new_n695));
  NOR3_X1   g270(.A1(new_n689), .A2(new_n692), .A3(new_n695), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(new_n689), .B2(new_n695), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n694), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XOR2_X1   g275(.A(G1991), .B(G1996), .Z(new_n701));
  XOR2_X1   g276(.A(new_n701), .B(KEYINPUT90), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n700), .B(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(G1981), .B(G1986), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(G229));
  NOR2_X1   g280(.A1(G6), .A2(G16), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n592), .A2(new_n595), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n706), .B1(new_n707), .B2(G16), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT32), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(G1981), .ZN(new_n710));
  INV_X1    g285(.A(G16), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(G22), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(G166), .B2(new_n711), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(G1971), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n714), .A2(KEYINPUT94), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n714), .A2(KEYINPUT94), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n711), .A2(G23), .ZN(new_n717));
  INV_X1    g292(.A(G288), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n717), .B1(new_n718), .B2(new_n711), .ZN(new_n719));
  XNOR2_X1  g294(.A(KEYINPUT33), .B(G1976), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n716), .A2(new_n721), .ZN(new_n722));
  NOR3_X1   g297(.A1(new_n710), .A2(new_n715), .A3(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(KEYINPUT34), .ZN(new_n724));
  OR2_X1    g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n723), .A2(new_n724), .ZN(new_n726));
  INV_X1    g301(.A(G29), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(G25), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n467), .A2(G131), .ZN(new_n729));
  INV_X1    g304(.A(G119), .ZN(new_n730));
  INV_X1    g305(.A(new_n482), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n729), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(G95), .ZN(new_n733));
  AND3_X1   g308(.A1(new_n733), .A2(new_n481), .A3(KEYINPUT91), .ZN(new_n734));
  AOI21_X1  g309(.A(KEYINPUT91), .B1(new_n733), .B2(new_n481), .ZN(new_n735));
  OAI221_X1 g310(.A(G2104), .B1(G107), .B2(new_n481), .C1(new_n734), .C2(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(new_n736), .ZN(new_n737));
  OR2_X1    g312(.A1(new_n732), .A2(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(new_n738), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n728), .B1(new_n739), .B2(new_n727), .ZN(new_n740));
  XOR2_X1   g315(.A(KEYINPUT35), .B(G1991), .Z(new_n741));
  XOR2_X1   g316(.A(new_n741), .B(KEYINPUT92), .Z(new_n742));
  XNOR2_X1  g317(.A(new_n740), .B(new_n742), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n711), .B1(G290), .B2(KEYINPUT93), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(KEYINPUT93), .B2(G290), .ZN(new_n745));
  INV_X1    g320(.A(G24), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n745), .B1(G16), .B2(new_n746), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n743), .B1(new_n747), .B2(G1986), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(G1986), .B2(new_n747), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n725), .A2(new_n726), .A3(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(KEYINPUT95), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n751), .A2(KEYINPUT36), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n750), .B(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n653), .A2(G29), .ZN(new_n754));
  NAND2_X1  g329(.A1(G115), .A2(G2104), .ZN(new_n755));
  INV_X1    g330(.A(G127), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n755), .B1(new_n480), .B2(new_n756), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n481), .B1(new_n757), .B2(KEYINPUT98), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(KEYINPUT98), .B2(new_n757), .ZN(new_n759));
  INV_X1    g334(.A(KEYINPUT25), .ZN(new_n760));
  NAND2_X1  g335(.A1(G103), .A2(G2104), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n760), .B1(new_n761), .B2(G2105), .ZN(new_n762));
  NAND4_X1  g337(.A1(new_n481), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n763));
  AOI22_X1  g338(.A1(new_n467), .A2(G139), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  AND2_X1   g339(.A1(new_n759), .A2(new_n764), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n765), .A2(new_n727), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(new_n727), .B2(G33), .ZN(new_n767));
  INV_X1    g342(.A(G2072), .ZN(new_n768));
  AOI22_X1  g343(.A1(new_n754), .A2(KEYINPUT100), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n711), .A2(G20), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT23), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(new_n631), .B2(new_n711), .ZN(new_n772));
  INV_X1    g347(.A(G1956), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  OAI211_X1 g349(.A(new_n769), .B(new_n774), .C1(new_n768), .C2(new_n767), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n727), .A2(G35), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(G162), .B2(new_n727), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(KEYINPUT29), .Z(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(G2090), .Z(new_n779));
  INV_X1    g354(.A(KEYINPUT30), .ZN(new_n780));
  AND2_X1   g355(.A1(new_n780), .A2(G28), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n727), .B1(new_n780), .B2(G28), .ZN(new_n782));
  AND2_X1   g357(.A1(KEYINPUT31), .A2(G11), .ZN(new_n783));
  NOR2_X1   g358(.A1(KEYINPUT31), .A2(G11), .ZN(new_n784));
  OAI22_X1  g359(.A1(new_n781), .A2(new_n782), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(G34), .ZN(new_n786));
  AOI21_X1  g361(.A(G29), .B1(new_n786), .B2(KEYINPUT24), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(KEYINPUT24), .B2(new_n786), .ZN(new_n788));
  INV_X1    g363(.A(G160), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n788), .B1(new_n789), .B2(new_n727), .ZN(new_n790));
  INV_X1    g365(.A(G2084), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n785), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  OAI221_X1 g367(.A(new_n792), .B1(new_n791), .B2(new_n790), .C1(new_n754), .C2(KEYINPUT100), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n482), .A2(G129), .ZN(new_n794));
  AOI22_X1  g369(.A1(new_n467), .A2(G141), .B1(G105), .B2(new_n469), .ZN(new_n795));
  NAND3_X1  g370(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(KEYINPUT26), .Z(new_n797));
  NAND3_X1  g372(.A1(new_n794), .A2(new_n795), .A3(new_n797), .ZN(new_n798));
  MUX2_X1   g373(.A(G32), .B(new_n798), .S(G29), .Z(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT27), .ZN(new_n800));
  INV_X1    g375(.A(G1996), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n800), .B(new_n801), .ZN(new_n802));
  NOR4_X1   g377(.A1(new_n775), .A2(new_n779), .A3(new_n793), .A4(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n711), .A2(G5), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(G171), .B2(new_n711), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT101), .ZN(new_n806));
  INV_X1    g381(.A(G1961), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n467), .A2(G140), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT96), .ZN(new_n811));
  OAI21_X1  g386(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n812));
  INV_X1    g387(.A(G116), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n812), .B1(new_n813), .B2(G2105), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n814), .B1(new_n482), .B2(G128), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n811), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n816), .A2(G29), .ZN(new_n817));
  XOR2_X1   g392(.A(new_n817), .B(KEYINPUT97), .Z(new_n818));
  NAND2_X1  g393(.A1(new_n727), .A2(G26), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT28), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(G2067), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n727), .A2(G27), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n824), .B1(G164), .B2(new_n727), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(G2078), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n826), .B(KEYINPUT102), .Z(new_n827));
  NAND2_X1  g402(.A1(new_n711), .A2(G19), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n828), .B1(new_n567), .B2(new_n711), .ZN(new_n829));
  XOR2_X1   g404(.A(new_n829), .B(G1341), .Z(new_n830));
  AND3_X1   g405(.A1(new_n823), .A2(new_n827), .A3(new_n830), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n803), .A2(new_n809), .A3(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n711), .A2(G4), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n833), .B1(new_n621), .B2(new_n711), .ZN(new_n834));
  INV_X1    g409(.A(G1348), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n834), .B(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n711), .A2(G21), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n837), .B1(G168), .B2(new_n711), .ZN(new_n838));
  XOR2_X1   g413(.A(KEYINPUT99), .B(G1966), .Z(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  OR2_X1    g415(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n838), .A2(new_n840), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n836), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  NOR3_X1   g418(.A1(new_n753), .A2(new_n832), .A3(new_n843), .ZN(G311));
  AND3_X1   g419(.A1(new_n803), .A2(new_n809), .A3(new_n831), .ZN(new_n845));
  INV_X1    g420(.A(new_n843), .ZN(new_n846));
  AND3_X1   g421(.A1(new_n750), .A2(new_n751), .A3(KEYINPUT36), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n750), .B1(new_n751), .B2(KEYINPUT36), .ZN(new_n848));
  OAI211_X1 g423(.A(new_n845), .B(new_n846), .C1(new_n847), .C2(new_n848), .ZN(G150));
  NAND2_X1  g424(.A1(new_n621), .A2(G559), .ZN(new_n850));
  XOR2_X1   g425(.A(KEYINPUT103), .B(KEYINPUT38), .Z(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT104), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n850), .B(new_n852), .ZN(new_n853));
  OAI21_X1  g428(.A(G67), .B1(new_n516), .B2(new_n517), .ZN(new_n854));
  NAND2_X1  g429(.A1(G80), .A2(G543), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n509), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  AOI22_X1  g432(.A1(new_n553), .A2(G93), .B1(new_n513), .B2(G55), .ZN(new_n858));
  AOI22_X1  g433(.A1(new_n564), .A2(new_n565), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n535), .A2(G55), .A3(G543), .ZN(new_n861));
  INV_X1    g436(.A(G93), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n861), .B1(new_n862), .B2(new_n520), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n863), .A2(new_n856), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n864), .A2(new_n564), .A3(new_n565), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n860), .A2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n853), .B(new_n866), .ZN(new_n867));
  OR2_X1    g442(.A1(new_n867), .A2(KEYINPUT39), .ZN(new_n868));
  INV_X1    g443(.A(G860), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n867), .A2(KEYINPUT39), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n868), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n864), .A2(new_n869), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(KEYINPUT37), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n871), .A2(new_n873), .ZN(G145));
  XNOR2_X1  g449(.A(new_n653), .B(new_n789), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(G162), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n816), .B(new_n798), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(new_n738), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n765), .A2(KEYINPUT106), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT105), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n879), .B(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n881), .A2(G164), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n879), .B(KEYINPUT105), .ZN(new_n883));
  INV_X1    g458(.A(G164), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n882), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n482), .A2(G130), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n467), .A2(G142), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n481), .A2(G118), .ZN(new_n889));
  OAI21_X1  g464(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n890));
  OAI211_X1 g465(.A(new_n887), .B(new_n888), .C1(new_n889), .C2(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(new_n643), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n886), .A2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n892), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n882), .A2(new_n885), .A3(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n878), .B1(new_n893), .B2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n893), .A2(new_n878), .A3(new_n895), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n876), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(G37), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n897), .A2(new_n876), .A3(new_n898), .ZN(new_n902));
  NAND4_X1  g477(.A1(new_n900), .A2(KEYINPUT40), .A3(new_n901), .A4(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT40), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n902), .A2(new_n901), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n904), .B1(new_n905), .B2(new_n899), .ZN(new_n906));
  AND2_X1   g481(.A1(new_n903), .A2(new_n906), .ZN(G395));
  XNOR2_X1  g482(.A(new_n866), .B(new_n638), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n620), .A2(new_n619), .ZN(new_n909));
  NOR3_X1   g484(.A1(new_n608), .A2(new_n605), .A3(new_n610), .ZN(new_n910));
  AOI21_X1  g485(.A(KEYINPUT82), .B1(new_n615), .B2(new_n609), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n909), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(new_n631), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n621), .A2(G299), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n908), .A2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT107), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n917), .B1(new_n621), .B2(G299), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n912), .A2(KEYINPUT107), .A3(new_n631), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n918), .A2(new_n919), .A3(new_n914), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT41), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n921), .B1(new_n621), .B2(G299), .ZN(new_n922));
  AOI22_X1  g497(.A1(new_n920), .A2(new_n921), .B1(new_n913), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n916), .B1(new_n923), .B2(new_n908), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT108), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n925), .A2(KEYINPUT42), .ZN(new_n926));
  OR2_X1    g501(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n718), .B(G166), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n707), .B(new_n602), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n928), .B(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n930), .B1(new_n925), .B2(KEYINPUT42), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n924), .A2(new_n926), .ZN(new_n932));
  AND3_X1   g507(.A1(new_n927), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n931), .B1(new_n927), .B2(new_n932), .ZN(new_n934));
  OAI21_X1  g509(.A(G868), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n864), .A2(G868), .ZN(new_n936));
  INV_X1    g511(.A(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n935), .A2(new_n937), .ZN(G295));
  NAND2_X1  g513(.A1(G295), .A2(KEYINPUT109), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT109), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n935), .A2(new_n940), .A3(new_n937), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n939), .A2(new_n941), .ZN(G331));
  INV_X1    g517(.A(KEYINPUT44), .ZN(new_n943));
  AND3_X1   g518(.A1(new_n538), .A2(new_n542), .A3(G301), .ZN(new_n944));
  AOI21_X1  g519(.A(G301), .B1(new_n538), .B2(new_n542), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n866), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(G168), .A2(G171), .ZN(new_n947));
  AND3_X1   g522(.A1(new_n864), .A2(new_n564), .A3(new_n565), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n948), .A2(new_n859), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n538), .A2(new_n542), .A3(G301), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n947), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n946), .A2(new_n951), .A3(new_n915), .ZN(new_n952));
  AND2_X1   g527(.A1(new_n946), .A2(new_n951), .ZN(new_n953));
  OAI211_X1 g528(.A(new_n930), .B(new_n952), .C1(new_n953), .C2(new_n923), .ZN(new_n954));
  AND2_X1   g529(.A1(new_n954), .A2(new_n901), .ZN(new_n955));
  INV_X1    g530(.A(new_n930), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT111), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n946), .A2(new_n951), .A3(new_n957), .A4(new_n915), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n952), .A2(KEYINPUT111), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n912), .A2(new_n631), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n621), .A2(G299), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n921), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n918), .A2(new_n922), .A3(new_n919), .ZN(new_n963));
  AOI22_X1  g538(.A1(new_n951), .A2(new_n946), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  OAI211_X1 g539(.A(new_n956), .B(new_n958), .C1(new_n959), .C2(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(KEYINPUT112), .B1(new_n955), .B2(new_n965), .ZN(new_n966));
  AND4_X1   g541(.A1(KEYINPUT112), .A2(new_n965), .A3(new_n901), .A4(new_n954), .ZN(new_n967));
  OAI21_X1  g542(.A(KEYINPUT43), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT43), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n920), .A2(new_n921), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n922), .A2(new_n913), .ZN(new_n971));
  AOI22_X1  g546(.A1(new_n970), .A2(new_n971), .B1(new_n951), .B2(new_n946), .ZN(new_n972));
  INV_X1    g547(.A(new_n952), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n956), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n974), .A2(KEYINPUT110), .A3(new_n901), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(new_n954), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n952), .B1(new_n953), .B2(new_n923), .ZN(new_n977));
  AOI21_X1  g552(.A(G37), .B1(new_n977), .B2(new_n956), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n978), .A2(KEYINPUT110), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n969), .B1(new_n976), .B2(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n943), .B1(new_n968), .B2(new_n980), .ZN(new_n981));
  OAI21_X1  g556(.A(KEYINPUT43), .B1(new_n976), .B2(new_n979), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n965), .A2(new_n901), .A3(new_n954), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n983), .A2(KEYINPUT43), .ZN(new_n984));
  INV_X1    g559(.A(new_n984), .ZN(new_n985));
  AOI21_X1  g560(.A(KEYINPUT44), .B1(new_n982), .B2(new_n985), .ZN(new_n986));
  OAI21_X1  g561(.A(KEYINPUT113), .B1(new_n981), .B2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT112), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n983), .A2(new_n988), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n955), .A2(KEYINPUT112), .A3(new_n965), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n969), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  OR2_X1    g566(.A1(new_n978), .A2(KEYINPUT110), .ZN(new_n992));
  INV_X1    g567(.A(new_n954), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n993), .B1(new_n978), .B2(KEYINPUT110), .ZN(new_n994));
  AOI21_X1  g569(.A(KEYINPUT43), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  OAI21_X1  g570(.A(KEYINPUT44), .B1(new_n991), .B2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT113), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n969), .B1(new_n992), .B2(new_n994), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n943), .B1(new_n998), .B2(new_n984), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n996), .A2(new_n997), .A3(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n987), .A2(new_n1000), .ZN(G397));
  XOR2_X1   g576(.A(KEYINPUT114), .B(G1384), .Z(new_n1002));
  NAND2_X1  g577(.A1(new_n884), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT45), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n470), .A2(new_n474), .A3(G40), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  XOR2_X1   g582(.A(new_n1007), .B(KEYINPUT115), .Z(new_n1008));
  NAND2_X1  g583(.A1(new_n816), .A2(G2067), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n811), .A2(new_n822), .A3(new_n815), .ZN(new_n1010));
  AND2_X1   g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  XNOR2_X1  g586(.A(new_n798), .B(new_n801), .ZN(new_n1012));
  AND2_X1   g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n739), .A2(new_n741), .ZN(new_n1014));
  OR2_X1    g589(.A1(new_n739), .A2(new_n741), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1013), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(G1986), .ZN(new_n1017));
  XNOR2_X1  g592(.A(new_n602), .B(new_n1017), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1008), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(G1384), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1006), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n884), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  AND2_X1   g597(.A1(new_n1022), .A2(G8), .ZN(new_n1023));
  NAND2_X1  g598(.A1(G305), .A2(G1981), .ZN(new_n1024));
  INV_X1    g599(.A(G1981), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n707), .A2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT49), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1024), .A2(KEYINPUT49), .A3(new_n1026), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1029), .A2(new_n1023), .A3(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(G1976), .ZN(new_n1032));
  AND3_X1   g607(.A1(new_n1031), .A2(new_n1032), .A3(new_n718), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1026), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1023), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n718), .A2(G1976), .ZN(new_n1036));
  AOI21_X1  g611(.A(KEYINPUT52), .B1(G288), .B2(new_n1032), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1023), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1022), .A2(G8), .A3(new_n1036), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(KEYINPUT52), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1031), .A2(new_n1038), .A3(new_n1040), .ZN(new_n1041));
  AND2_X1   g616(.A1(new_n1041), .A2(KEYINPUT116), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1041), .A2(KEYINPUT116), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g619(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT50), .ZN(new_n1046));
  AOI22_X1  g621(.A1(new_n498), .A2(new_n499), .B1(new_n495), .B2(KEYINPUT4), .ZN(new_n1047));
  OAI211_X1 g622(.A(new_n1046), .B(new_n1020), .C1(new_n1047), .C2(new_n493), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1045), .A2(new_n1021), .A3(new_n1048), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1049), .A2(G2090), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1020), .B1(new_n1047), .B2(new_n493), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1006), .B1(new_n1051), .B2(new_n1004), .ZN(new_n1052));
  OAI211_X1 g627(.A(KEYINPUT45), .B(new_n1002), .C1(new_n1047), .C2(new_n493), .ZN(new_n1053));
  AOI21_X1  g628(.A(G1971), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(G8), .B1(new_n1050), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(G303), .A2(G8), .ZN(new_n1056));
  XNOR2_X1  g631(.A(new_n1056), .B(KEYINPUT55), .ZN(new_n1057));
  OR2_X1    g632(.A1(new_n1055), .A2(new_n1057), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1035), .B1(new_n1044), .B2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1055), .A2(new_n1057), .ZN(new_n1060));
  AND2_X1   g635(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1004), .B1(G164), .B2(G1384), .ZN(new_n1062));
  OAI211_X1 g637(.A(KEYINPUT45), .B(new_n1020), .C1(new_n1047), .C2(new_n493), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1062), .A2(new_n1021), .A3(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(new_n839), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1045), .A2(new_n1021), .A3(new_n791), .A4(new_n1048), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1067), .A2(G8), .A3(G168), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT63), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  OAI211_X1 g645(.A(new_n1061), .B(new_n1070), .C1(new_n1042), .C2(new_n1043), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1041), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1058), .A2(new_n1072), .A3(new_n1060), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1069), .B1(new_n1073), .B2(new_n1068), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1059), .B1(new_n1071), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1049), .A2(new_n773), .ZN(new_n1076));
  AOI21_X1  g651(.A(KEYINPUT57), .B1(new_n579), .B2(new_n581), .ZN(new_n1077));
  AOI22_X1  g652(.A1(G299), .A2(KEYINPUT57), .B1(new_n1077), .B2(new_n576), .ZN(new_n1078));
  XNOR2_X1  g653(.A(KEYINPUT56), .B(G2072), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1052), .A2(new_n1053), .A3(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1076), .A2(new_n1078), .A3(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(KEYINPUT117), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT117), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1076), .A2(new_n1083), .A3(new_n1078), .A4(new_n1080), .ZN(new_n1084));
  AND2_X1   g659(.A1(new_n1082), .A2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1078), .B1(new_n1076), .B2(new_n1080), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1049), .A2(new_n835), .ZN(new_n1087));
  NOR4_X1   g662(.A1(G164), .A2(new_n1006), .A3(G1384), .A4(G2067), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1088), .ZN(new_n1089));
  AOI21_X1  g664(.A(KEYINPUT118), .B1(new_n1087), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT118), .ZN(new_n1091));
  AOI211_X1 g666(.A(new_n1091), .B(new_n1088), .C1(new_n1049), .C2(new_n835), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(new_n621), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1086), .B1(new_n1094), .B2(KEYINPUT119), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT119), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1093), .A2(new_n1096), .A3(new_n621), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1085), .B1(new_n1095), .B2(new_n1097), .ZN(new_n1098));
  OAI21_X1  g673(.A(KEYINPUT60), .B1(new_n1090), .B2(new_n1092), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(KEYINPUT121), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT121), .ZN(new_n1101));
  OAI211_X1 g676(.A(new_n1101), .B(KEYINPUT60), .C1(new_n1090), .C2(new_n1092), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1090), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1092), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT60), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1103), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1106));
  AOI22_X1  g681(.A1(new_n1100), .A2(new_n1102), .B1(new_n1106), .B2(new_n621), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1052), .A2(new_n801), .A3(new_n1053), .ZN(new_n1108));
  XOR2_X1   g683(.A(KEYINPUT58), .B(G1341), .Z(new_n1109));
  NAND2_X1  g684(.A1(new_n1022), .A2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n566), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1111));
  XNOR2_X1  g686(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1112), .ZN(new_n1113));
  XNOR2_X1  g688(.A(new_n1111), .B(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1086), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1115), .A2(KEYINPUT61), .A3(new_n1081), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1086), .B1(new_n1082), .B2(new_n1084), .ZN(new_n1117));
  OAI211_X1 g692(.A(new_n1114), .B(new_n1116), .C1(new_n1117), .C2(KEYINPUT61), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1107), .A2(new_n1118), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1100), .A2(new_n621), .A3(new_n1106), .A4(new_n1102), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1098), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(G2078), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1052), .A2(new_n1122), .A3(new_n1053), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT53), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1049), .A2(new_n807), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1122), .A2(KEYINPUT53), .ZN(new_n1127));
  OAI211_X1 g702(.A(new_n1125), .B(new_n1126), .C1(new_n1064), .C2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g703(.A(KEYINPUT54), .B1(new_n1128), .B2(G171), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1053), .ZN(new_n1130));
  NOR3_X1   g705(.A1(new_n1130), .A2(new_n1006), .A3(new_n1127), .ZN(new_n1131));
  AOI22_X1  g706(.A1(new_n1124), .A2(new_n1123), .B1(new_n1131), .B2(new_n1005), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT124), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1126), .A2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1049), .A2(KEYINPUT124), .A3(new_n807), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1132), .A2(new_n1134), .A3(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1129), .B1(G171), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1128), .A2(G171), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1132), .A2(G301), .A3(new_n1134), .A4(new_n1135), .ZN(new_n1139));
  AOI21_X1  g714(.A(KEYINPUT54), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  NOR3_X1   g715(.A1(new_n1137), .A2(new_n1073), .A3(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT123), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1065), .A2(G168), .A3(new_n1066), .ZN(new_n1143));
  OAI21_X1  g718(.A(G8), .B1(KEYINPUT122), .B2(KEYINPUT51), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(KEYINPUT122), .A2(KEYINPUT51), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1143), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1067), .A2(G8), .A3(G286), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1146), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1142), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1143), .A2(new_n1145), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1146), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1154), .A2(KEYINPUT123), .A3(new_n1148), .A4(new_n1147), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1151), .A2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1141), .A2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1075), .B1(new_n1121), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT62), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1151), .A2(new_n1159), .A3(new_n1155), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n1073), .A2(new_n1138), .ZN(new_n1161));
  AND3_X1   g736(.A1(new_n1160), .A2(KEYINPUT125), .A3(new_n1161), .ZN(new_n1162));
  AOI21_X1  g737(.A(KEYINPUT125), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1159), .B1(new_n1151), .B2(new_n1155), .ZN(new_n1164));
  NOR3_X1   g739(.A1(new_n1162), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1019), .B1(new_n1158), .B2(new_n1165), .ZN(new_n1166));
  XOR2_X1   g741(.A(new_n1014), .B(KEYINPUT126), .Z(new_n1167));
  INV_X1    g742(.A(new_n1013), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1010), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1169), .A2(new_n1008), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1008), .A2(new_n1017), .A3(new_n602), .ZN(new_n1171));
  XOR2_X1   g746(.A(new_n1171), .B(KEYINPUT48), .Z(new_n1172));
  NAND2_X1  g747(.A1(new_n1008), .A2(new_n1016), .ZN(new_n1173));
  XNOR2_X1  g748(.A(new_n1173), .B(KEYINPUT127), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1170), .B1(new_n1172), .B2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1008), .A2(new_n801), .ZN(new_n1176));
  XNOR2_X1  g751(.A(new_n1176), .B(KEYINPUT46), .ZN(new_n1177));
  INV_X1    g752(.A(new_n1011), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1008), .B1(new_n798), .B2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1177), .A2(new_n1179), .ZN(new_n1180));
  OR2_X1    g755(.A1(new_n1180), .A2(KEYINPUT47), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1180), .A2(KEYINPUT47), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1175), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1166), .A2(new_n1183), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g759(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(new_n1186));
  NOR4_X1   g760(.A1(G229), .A2(new_n463), .A3(G401), .A4(G227), .ZN(new_n1187));
  NAND2_X1  g761(.A1(new_n982), .A2(new_n985), .ZN(new_n1188));
  AND3_X1   g762(.A1(new_n1186), .A2(new_n1187), .A3(new_n1188), .ZN(G308));
  NAND3_X1  g763(.A1(new_n1186), .A2(new_n1188), .A3(new_n1187), .ZN(G225));
endmodule


