

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U551 ( .A1(n655), .A2(n596), .ZN(n598) );
  XNOR2_X1 U552 ( .A(KEYINPUT99), .B(KEYINPUT31), .ZN(n650) );
  XNOR2_X1 U553 ( .A(n651), .B(n650), .ZN(n652) );
  INV_X1 U554 ( .A(n989), .ZN(n674) );
  AND2_X1 U555 ( .A1(n676), .A2(n675), .ZN(n677) );
  NAND2_X1 U556 ( .A1(n582), .A2(n725), .ZN(n655) );
  NOR2_X1 U557 ( .A1(G164), .A2(G1384), .ZN(n725) );
  NOR2_X1 U558 ( .A1(G651), .A2(n557), .ZN(n771) );
  INV_X1 U559 ( .A(KEYINPUT85), .ZN(n522) );
  INV_X1 U560 ( .A(G2105), .ZN(n519) );
  AND2_X1 U561 ( .A1(n519), .A2(G2104), .ZN(n883) );
  NAND2_X1 U562 ( .A1(G102), .A2(n883), .ZN(n518) );
  NOR2_X1 U563 ( .A1(G2104), .A2(G2105), .ZN(n516) );
  XOR2_X2 U564 ( .A(KEYINPUT17), .B(n516), .Z(n881) );
  NAND2_X1 U565 ( .A1(G138), .A2(n881), .ZN(n517) );
  NAND2_X1 U566 ( .A1(n518), .A2(n517), .ZN(n525) );
  NOR2_X2 U567 ( .A1(G2104), .A2(n519), .ZN(n877) );
  NAND2_X1 U568 ( .A1(G126), .A2(n877), .ZN(n521) );
  AND2_X1 U569 ( .A1(G2104), .A2(G2105), .ZN(n876) );
  NAND2_X1 U570 ( .A1(G114), .A2(n876), .ZN(n520) );
  NAND2_X1 U571 ( .A1(n521), .A2(n520), .ZN(n523) );
  XNOR2_X1 U572 ( .A(n523), .B(n522), .ZN(n524) );
  NOR2_X1 U573 ( .A1(n525), .A2(n524), .ZN(G164) );
  XNOR2_X1 U574 ( .A(G651), .B(KEYINPUT67), .ZN(n530) );
  NOR2_X1 U575 ( .A1(G543), .A2(n530), .ZN(n526) );
  XOR2_X1 U576 ( .A(KEYINPUT1), .B(n526), .Z(n770) );
  NAND2_X1 U577 ( .A1(G64), .A2(n770), .ZN(n528) );
  XOR2_X1 U578 ( .A(KEYINPUT0), .B(G543), .Z(n557) );
  NAND2_X1 U579 ( .A1(G52), .A2(n771), .ZN(n527) );
  NAND2_X1 U580 ( .A1(n528), .A2(n527), .ZN(n535) );
  NOR2_X1 U581 ( .A1(G651), .A2(G543), .ZN(n529) );
  XOR2_X1 U582 ( .A(KEYINPUT65), .B(n529), .Z(n774) );
  NAND2_X1 U583 ( .A1(G90), .A2(n774), .ZN(n532) );
  NOR2_X1 U584 ( .A1(n557), .A2(n530), .ZN(n775) );
  NAND2_X1 U585 ( .A1(G77), .A2(n775), .ZN(n531) );
  NAND2_X1 U586 ( .A1(n532), .A2(n531), .ZN(n533) );
  XOR2_X1 U587 ( .A(KEYINPUT9), .B(n533), .Z(n534) );
  NOR2_X1 U588 ( .A1(n535), .A2(n534), .ZN(G171) );
  INV_X1 U589 ( .A(G171), .ZN(G301) );
  NAND2_X1 U590 ( .A1(n771), .A2(G51), .ZN(n536) );
  XNOR2_X1 U591 ( .A(n536), .B(KEYINPUT74), .ZN(n538) );
  NAND2_X1 U592 ( .A1(G63), .A2(n770), .ZN(n537) );
  NAND2_X1 U593 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U594 ( .A(KEYINPUT6), .B(n539), .ZN(n545) );
  NAND2_X1 U595 ( .A1(n774), .A2(G89), .ZN(n540) );
  XNOR2_X1 U596 ( .A(n540), .B(KEYINPUT4), .ZN(n542) );
  NAND2_X1 U597 ( .A1(G76), .A2(n775), .ZN(n541) );
  NAND2_X1 U598 ( .A1(n542), .A2(n541), .ZN(n543) );
  XOR2_X1 U599 ( .A(n543), .B(KEYINPUT5), .Z(n544) );
  NOR2_X1 U600 ( .A1(n545), .A2(n544), .ZN(n546) );
  XOR2_X1 U601 ( .A(KEYINPUT75), .B(n546), .Z(n547) );
  XOR2_X1 U602 ( .A(KEYINPUT7), .B(n547), .Z(G168) );
  XOR2_X1 U603 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U604 ( .A1(G88), .A2(n774), .ZN(n549) );
  NAND2_X1 U605 ( .A1(G75), .A2(n775), .ZN(n548) );
  NAND2_X1 U606 ( .A1(n549), .A2(n548), .ZN(n553) );
  NAND2_X1 U607 ( .A1(G62), .A2(n770), .ZN(n551) );
  NAND2_X1 U608 ( .A1(G50), .A2(n771), .ZN(n550) );
  NAND2_X1 U609 ( .A1(n551), .A2(n550), .ZN(n552) );
  NOR2_X1 U610 ( .A1(n553), .A2(n552), .ZN(G166) );
  XOR2_X1 U611 ( .A(KEYINPUT86), .B(G166), .Z(G303) );
  NAND2_X1 U612 ( .A1(G49), .A2(n771), .ZN(n555) );
  NAND2_X1 U613 ( .A1(G74), .A2(G651), .ZN(n554) );
  NAND2_X1 U614 ( .A1(n555), .A2(n554), .ZN(n556) );
  NOR2_X1 U615 ( .A1(n770), .A2(n556), .ZN(n560) );
  NAND2_X1 U616 ( .A1(G87), .A2(n557), .ZN(n558) );
  XOR2_X1 U617 ( .A(KEYINPUT79), .B(n558), .Z(n559) );
  NAND2_X1 U618 ( .A1(n560), .A2(n559), .ZN(G288) );
  NAND2_X1 U619 ( .A1(G86), .A2(n774), .ZN(n562) );
  NAND2_X1 U620 ( .A1(G61), .A2(n770), .ZN(n561) );
  NAND2_X1 U621 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U622 ( .A(KEYINPUT80), .B(n563), .ZN(n566) );
  NAND2_X1 U623 ( .A1(n775), .A2(G73), .ZN(n564) );
  XOR2_X1 U624 ( .A(KEYINPUT2), .B(n564), .Z(n565) );
  NOR2_X1 U625 ( .A1(n566), .A2(n565), .ZN(n568) );
  NAND2_X1 U626 ( .A1(n771), .A2(G48), .ZN(n567) );
  NAND2_X1 U627 ( .A1(n568), .A2(n567), .ZN(G305) );
  AND2_X1 U628 ( .A1(n775), .A2(G72), .ZN(n572) );
  NAND2_X1 U629 ( .A1(G85), .A2(n774), .ZN(n570) );
  NAND2_X1 U630 ( .A1(G47), .A2(n771), .ZN(n569) );
  NAND2_X1 U631 ( .A1(n570), .A2(n569), .ZN(n571) );
  NOR2_X1 U632 ( .A1(n572), .A2(n571), .ZN(n574) );
  NAND2_X1 U633 ( .A1(n770), .A2(G60), .ZN(n573) );
  NAND2_X1 U634 ( .A1(n574), .A2(n573), .ZN(G290) );
  NAND2_X1 U635 ( .A1(G113), .A2(n876), .ZN(n576) );
  NAND2_X1 U636 ( .A1(G125), .A2(n877), .ZN(n575) );
  AND2_X1 U637 ( .A1(n576), .A2(n575), .ZN(n745) );
  AND2_X1 U638 ( .A1(n745), .A2(G40), .ZN(n581) );
  NAND2_X1 U639 ( .A1(G137), .A2(n881), .ZN(n577) );
  XNOR2_X1 U640 ( .A(n577), .B(KEYINPUT66), .ZN(n580) );
  NAND2_X1 U641 ( .A1(G101), .A2(n883), .ZN(n578) );
  XOR2_X1 U642 ( .A(KEYINPUT23), .B(n578), .Z(n579) );
  AND2_X1 U643 ( .A1(n580), .A2(n579), .ZN(n744) );
  NAND2_X1 U644 ( .A1(n581), .A2(n744), .ZN(n724) );
  INV_X1 U645 ( .A(n724), .ZN(n582) );
  NAND2_X1 U646 ( .A1(G1961), .A2(n655), .ZN(n584) );
  INV_X1 U647 ( .A(n655), .ZN(n602) );
  XOR2_X1 U648 ( .A(G2078), .B(KEYINPUT25), .Z(n909) );
  NAND2_X1 U649 ( .A1(n602), .A2(n909), .ZN(n583) );
  NAND2_X1 U650 ( .A1(n584), .A2(n583), .ZN(n639) );
  OR2_X1 U651 ( .A1(G301), .A2(n639), .ZN(n638) );
  NAND2_X1 U652 ( .A1(G2072), .A2(n602), .ZN(n585) );
  XNOR2_X1 U653 ( .A(n585), .B(KEYINPUT27), .ZN(n586) );
  XNOR2_X1 U654 ( .A(KEYINPUT94), .B(n586), .ZN(n588) );
  AND2_X1 U655 ( .A1(n655), .A2(G1956), .ZN(n587) );
  NOR2_X1 U656 ( .A1(n588), .A2(n587), .ZN(n631) );
  NAND2_X1 U657 ( .A1(G65), .A2(n770), .ZN(n590) );
  NAND2_X1 U658 ( .A1(G53), .A2(n771), .ZN(n589) );
  NAND2_X1 U659 ( .A1(n590), .A2(n589), .ZN(n594) );
  NAND2_X1 U660 ( .A1(G91), .A2(n774), .ZN(n592) );
  NAND2_X1 U661 ( .A1(G78), .A2(n775), .ZN(n591) );
  NAND2_X1 U662 ( .A1(n592), .A2(n591), .ZN(n593) );
  NOR2_X1 U663 ( .A1(n594), .A2(n593), .ZN(n988) );
  NOR2_X1 U664 ( .A1(n631), .A2(n988), .ZN(n595) );
  XOR2_X1 U665 ( .A(n595), .B(KEYINPUT28), .Z(n635) );
  INV_X1 U666 ( .A(G1996), .ZN(n596) );
  XOR2_X1 U667 ( .A(KEYINPUT64), .B(KEYINPUT26), .Z(n597) );
  XNOR2_X1 U668 ( .A(n598), .B(n597), .ZN(n600) );
  NAND2_X1 U669 ( .A1(n655), .A2(G1341), .ZN(n599) );
  NAND2_X1 U670 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U671 ( .A(n601), .B(KEYINPUT95), .ZN(n613) );
  NAND2_X1 U672 ( .A1(G1348), .A2(n655), .ZN(n604) );
  NAND2_X1 U673 ( .A1(G2067), .A2(n602), .ZN(n603) );
  NAND2_X1 U674 ( .A1(n604), .A2(n603), .ZN(n627) );
  NAND2_X1 U675 ( .A1(G66), .A2(n770), .ZN(n606) );
  NAND2_X1 U676 ( .A1(G54), .A2(n771), .ZN(n605) );
  NAND2_X1 U677 ( .A1(n606), .A2(n605), .ZN(n610) );
  NAND2_X1 U678 ( .A1(G92), .A2(n774), .ZN(n608) );
  NAND2_X1 U679 ( .A1(G79), .A2(n775), .ZN(n607) );
  NAND2_X1 U680 ( .A1(n608), .A2(n607), .ZN(n609) );
  NOR2_X1 U681 ( .A1(n610), .A2(n609), .ZN(n611) );
  XNOR2_X1 U682 ( .A(n611), .B(KEYINPUT15), .ZN(n999) );
  NAND2_X1 U683 ( .A1(n627), .A2(n999), .ZN(n612) );
  NAND2_X1 U684 ( .A1(n613), .A2(n612), .ZN(n626) );
  NAND2_X1 U685 ( .A1(n774), .A2(G81), .ZN(n614) );
  XNOR2_X1 U686 ( .A(n614), .B(KEYINPUT12), .ZN(n616) );
  NAND2_X1 U687 ( .A1(G68), .A2(n775), .ZN(n615) );
  NAND2_X1 U688 ( .A1(n616), .A2(n615), .ZN(n617) );
  XNOR2_X1 U689 ( .A(KEYINPUT13), .B(n617), .ZN(n624) );
  XOR2_X1 U690 ( .A(KEYINPUT14), .B(KEYINPUT70), .Z(n619) );
  NAND2_X1 U691 ( .A1(G56), .A2(n770), .ZN(n618) );
  XNOR2_X1 U692 ( .A(n619), .B(n618), .ZN(n622) );
  NAND2_X1 U693 ( .A1(G43), .A2(n771), .ZN(n620) );
  XNOR2_X1 U694 ( .A(KEYINPUT71), .B(n620), .ZN(n621) );
  NOR2_X1 U695 ( .A1(n622), .A2(n621), .ZN(n623) );
  NAND2_X1 U696 ( .A1(n624), .A2(n623), .ZN(n625) );
  XNOR2_X1 U697 ( .A(KEYINPUT72), .B(n625), .ZN(n997) );
  NOR2_X1 U698 ( .A1(n626), .A2(n997), .ZN(n629) );
  NOR2_X1 U699 ( .A1(n627), .A2(n999), .ZN(n628) );
  NOR2_X1 U700 ( .A1(n629), .A2(n628), .ZN(n630) );
  XNOR2_X1 U701 ( .A(n630), .B(KEYINPUT96), .ZN(n633) );
  NAND2_X1 U702 ( .A1(n631), .A2(n988), .ZN(n632) );
  NAND2_X1 U703 ( .A1(n633), .A2(n632), .ZN(n634) );
  NAND2_X1 U704 ( .A1(n635), .A2(n634), .ZN(n636) );
  XOR2_X1 U705 ( .A(KEYINPUT29), .B(n636), .Z(n637) );
  NAND2_X1 U706 ( .A1(n638), .A2(n637), .ZN(n653) );
  NAND2_X1 U707 ( .A1(G301), .A2(n639), .ZN(n640) );
  XOR2_X1 U708 ( .A(KEYINPUT98), .B(n640), .Z(n649) );
  XOR2_X1 U709 ( .A(KEYINPUT30), .B(KEYINPUT97), .Z(n646) );
  INV_X1 U710 ( .A(KEYINPUT93), .ZN(n642) );
  NAND2_X1 U711 ( .A1(G8), .A2(n655), .ZN(n693) );
  NOR2_X1 U712 ( .A1(G1966), .A2(n693), .ZN(n641) );
  XNOR2_X1 U713 ( .A(n642), .B(n641), .ZN(n667) );
  NOR2_X1 U714 ( .A1(n655), .A2(G2084), .ZN(n643) );
  XNOR2_X1 U715 ( .A(n643), .B(KEYINPUT92), .ZN(n664) );
  NOR2_X1 U716 ( .A1(n667), .A2(n664), .ZN(n644) );
  NAND2_X1 U717 ( .A1(n644), .A2(G8), .ZN(n645) );
  XNOR2_X1 U718 ( .A(n646), .B(n645), .ZN(n647) );
  NOR2_X1 U719 ( .A1(G168), .A2(n647), .ZN(n648) );
  NOR2_X1 U720 ( .A1(n649), .A2(n648), .ZN(n651) );
  NAND2_X1 U721 ( .A1(n653), .A2(n652), .ZN(n665) );
  AND2_X1 U722 ( .A1(G286), .A2(G8), .ZN(n654) );
  NAND2_X1 U723 ( .A1(n665), .A2(n654), .ZN(n662) );
  INV_X1 U724 ( .A(G8), .ZN(n660) );
  NOR2_X1 U725 ( .A1(G1971), .A2(n693), .ZN(n657) );
  NOR2_X1 U726 ( .A1(G2090), .A2(n655), .ZN(n656) );
  NOR2_X1 U727 ( .A1(n657), .A2(n656), .ZN(n658) );
  NAND2_X1 U728 ( .A1(G303), .A2(n658), .ZN(n659) );
  OR2_X1 U729 ( .A1(n660), .A2(n659), .ZN(n661) );
  AND2_X1 U730 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U731 ( .A(n663), .B(KEYINPUT32), .ZN(n671) );
  NAND2_X1 U732 ( .A1(n664), .A2(G8), .ZN(n669) );
  INV_X1 U733 ( .A(n665), .ZN(n666) );
  NOR2_X1 U734 ( .A1(n667), .A2(n666), .ZN(n668) );
  NAND2_X1 U735 ( .A1(n669), .A2(n668), .ZN(n670) );
  NAND2_X1 U736 ( .A1(n671), .A2(n670), .ZN(n691) );
  NOR2_X1 U737 ( .A1(G1976), .A2(G288), .ZN(n680) );
  NOR2_X1 U738 ( .A1(G303), .A2(G1971), .ZN(n672) );
  NOR2_X1 U739 ( .A1(n680), .A2(n672), .ZN(n996) );
  XNOR2_X1 U740 ( .A(KEYINPUT100), .B(n996), .ZN(n673) );
  NAND2_X1 U741 ( .A1(n691), .A2(n673), .ZN(n676) );
  NAND2_X1 U742 ( .A1(G1976), .A2(G288), .ZN(n989) );
  NOR2_X1 U743 ( .A1(n693), .A2(n674), .ZN(n675) );
  NOR2_X1 U744 ( .A1(KEYINPUT33), .A2(n677), .ZN(n679) );
  XOR2_X1 U745 ( .A(G1981), .B(G305), .Z(n985) );
  INV_X1 U746 ( .A(n985), .ZN(n678) );
  NOR2_X1 U747 ( .A1(n679), .A2(n678), .ZN(n683) );
  NAND2_X1 U748 ( .A1(n680), .A2(KEYINPUT33), .ZN(n681) );
  OR2_X1 U749 ( .A1(n693), .A2(n681), .ZN(n682) );
  NAND2_X1 U750 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X1 U751 ( .A(n684), .B(KEYINPUT101), .ZN(n688) );
  NOR2_X1 U752 ( .A1(G1981), .A2(G305), .ZN(n685) );
  XOR2_X1 U753 ( .A(n685), .B(KEYINPUT24), .Z(n686) );
  NOR2_X1 U754 ( .A1(n693), .A2(n686), .ZN(n687) );
  NOR2_X1 U755 ( .A1(n688), .A2(n687), .ZN(n695) );
  NOR2_X1 U756 ( .A1(G2090), .A2(G303), .ZN(n689) );
  NAND2_X1 U757 ( .A1(G8), .A2(n689), .ZN(n690) );
  NAND2_X1 U758 ( .A1(n691), .A2(n690), .ZN(n692) );
  NAND2_X1 U759 ( .A1(n693), .A2(n692), .ZN(n694) );
  NAND2_X1 U760 ( .A1(n695), .A2(n694), .ZN(n728) );
  NAND2_X1 U761 ( .A1(G104), .A2(n883), .ZN(n697) );
  NAND2_X1 U762 ( .A1(G140), .A2(n881), .ZN(n696) );
  NAND2_X1 U763 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U764 ( .A(KEYINPUT34), .B(n698), .ZN(n703) );
  NAND2_X1 U765 ( .A1(G116), .A2(n876), .ZN(n700) );
  NAND2_X1 U766 ( .A1(G128), .A2(n877), .ZN(n699) );
  NAND2_X1 U767 ( .A1(n700), .A2(n699), .ZN(n701) );
  XOR2_X1 U768 ( .A(KEYINPUT35), .B(n701), .Z(n702) );
  NOR2_X1 U769 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U770 ( .A(KEYINPUT36), .B(n704), .ZN(n873) );
  XOR2_X1 U771 ( .A(G2067), .B(KEYINPUT37), .Z(n705) );
  XNOR2_X1 U772 ( .A(KEYINPUT87), .B(n705), .ZN(n737) );
  NOR2_X1 U773 ( .A1(n873), .A2(n737), .ZN(n734) );
  XOR2_X1 U774 ( .A(KEYINPUT89), .B(G1991), .Z(n913) );
  NAND2_X1 U775 ( .A1(G107), .A2(n876), .ZN(n707) );
  NAND2_X1 U776 ( .A1(G95), .A2(n883), .ZN(n706) );
  NAND2_X1 U777 ( .A1(n707), .A2(n706), .ZN(n710) );
  NAND2_X1 U778 ( .A1(n881), .A2(G131), .ZN(n708) );
  XOR2_X1 U779 ( .A(KEYINPUT88), .B(n708), .Z(n709) );
  NOR2_X1 U780 ( .A1(n710), .A2(n709), .ZN(n712) );
  NAND2_X1 U781 ( .A1(n877), .A2(G119), .ZN(n711) );
  NAND2_X1 U782 ( .A1(n712), .A2(n711), .ZN(n892) );
  NAND2_X1 U783 ( .A1(n913), .A2(n892), .ZN(n713) );
  XNOR2_X1 U784 ( .A(n713), .B(KEYINPUT90), .ZN(n723) );
  NAND2_X1 U785 ( .A1(G117), .A2(n876), .ZN(n715) );
  NAND2_X1 U786 ( .A1(G129), .A2(n877), .ZN(n714) );
  NAND2_X1 U787 ( .A1(n715), .A2(n714), .ZN(n719) );
  NAND2_X1 U788 ( .A1(G105), .A2(n883), .ZN(n716) );
  XNOR2_X1 U789 ( .A(n716), .B(KEYINPUT38), .ZN(n717) );
  XNOR2_X1 U790 ( .A(n717), .B(KEYINPUT91), .ZN(n718) );
  NOR2_X1 U791 ( .A1(n719), .A2(n718), .ZN(n721) );
  NAND2_X1 U792 ( .A1(n881), .A2(G141), .ZN(n720) );
  NAND2_X1 U793 ( .A1(n721), .A2(n720), .ZN(n894) );
  NAND2_X1 U794 ( .A1(G1996), .A2(n894), .ZN(n722) );
  NAND2_X1 U795 ( .A1(n723), .A2(n722), .ZN(n731) );
  NOR2_X1 U796 ( .A1(n734), .A2(n731), .ZN(n972) );
  XOR2_X1 U797 ( .A(G1986), .B(G290), .Z(n992) );
  NAND2_X1 U798 ( .A1(n972), .A2(n992), .ZN(n726) );
  NOR2_X1 U799 ( .A1(n725), .A2(n724), .ZN(n739) );
  NAND2_X1 U800 ( .A1(n726), .A2(n739), .ZN(n727) );
  NAND2_X1 U801 ( .A1(n728), .A2(n727), .ZN(n742) );
  NOR2_X1 U802 ( .A1(G1996), .A2(n894), .ZN(n966) );
  NOR2_X1 U803 ( .A1(n913), .A2(n892), .ZN(n962) );
  NOR2_X1 U804 ( .A1(G1986), .A2(G290), .ZN(n729) );
  NOR2_X1 U805 ( .A1(n962), .A2(n729), .ZN(n730) );
  NOR2_X1 U806 ( .A1(n731), .A2(n730), .ZN(n732) );
  NOR2_X1 U807 ( .A1(n966), .A2(n732), .ZN(n733) );
  XNOR2_X1 U808 ( .A(KEYINPUT39), .B(n733), .ZN(n736) );
  INV_X1 U809 ( .A(n734), .ZN(n735) );
  NAND2_X1 U810 ( .A1(n736), .A2(n735), .ZN(n738) );
  NAND2_X1 U811 ( .A1(n873), .A2(n737), .ZN(n963) );
  NAND2_X1 U812 ( .A1(n738), .A2(n963), .ZN(n740) );
  NAND2_X1 U813 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U814 ( .A1(n742), .A2(n741), .ZN(n743) );
  XNOR2_X1 U815 ( .A(n743), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U816 ( .A1(n745), .A2(n744), .ZN(G160) );
  NAND2_X1 U817 ( .A1(G123), .A2(n877), .ZN(n746) );
  XNOR2_X1 U818 ( .A(n746), .B(KEYINPUT18), .ZN(n753) );
  NAND2_X1 U819 ( .A1(G111), .A2(n876), .ZN(n748) );
  NAND2_X1 U820 ( .A1(G135), .A2(n881), .ZN(n747) );
  NAND2_X1 U821 ( .A1(n748), .A2(n747), .ZN(n751) );
  NAND2_X1 U822 ( .A1(n883), .A2(G99), .ZN(n749) );
  XOR2_X1 U823 ( .A(KEYINPUT76), .B(n749), .Z(n750) );
  NOR2_X1 U824 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U825 ( .A1(n753), .A2(n752), .ZN(n959) );
  XNOR2_X1 U826 ( .A(G2096), .B(n959), .ZN(n754) );
  OR2_X1 U827 ( .A1(G2100), .A2(n754), .ZN(G156) );
  INV_X1 U828 ( .A(G132), .ZN(G219) );
  INV_X1 U829 ( .A(G82), .ZN(G220) );
  INV_X1 U830 ( .A(G120), .ZN(G236) );
  INV_X1 U831 ( .A(G69), .ZN(G235) );
  INV_X1 U832 ( .A(G108), .ZN(G238) );
  NAND2_X1 U833 ( .A1(G94), .A2(G452), .ZN(n755) );
  XOR2_X1 U834 ( .A(KEYINPUT68), .B(n755), .Z(G173) );
  NAND2_X1 U835 ( .A1(G7), .A2(G661), .ZN(n756) );
  XNOR2_X1 U836 ( .A(n756), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U837 ( .A(G223), .ZN(n823) );
  NAND2_X1 U838 ( .A1(n823), .A2(G567), .ZN(n757) );
  XOR2_X1 U839 ( .A(KEYINPUT11), .B(n757), .Z(G234) );
  XOR2_X1 U840 ( .A(G860), .B(KEYINPUT73), .Z(n764) );
  INV_X1 U841 ( .A(n997), .ZN(n758) );
  NAND2_X1 U842 ( .A1(n764), .A2(n758), .ZN(G153) );
  NAND2_X1 U843 ( .A1(G868), .A2(G301), .ZN(n760) );
  INV_X1 U844 ( .A(G868), .ZN(n794) );
  NAND2_X1 U845 ( .A1(n999), .A2(n794), .ZN(n759) );
  NAND2_X1 U846 ( .A1(n760), .A2(n759), .ZN(G284) );
  XNOR2_X1 U847 ( .A(n988), .B(KEYINPUT69), .ZN(G299) );
  NAND2_X1 U848 ( .A1(G286), .A2(G868), .ZN(n762) );
  NAND2_X1 U849 ( .A1(n794), .A2(G299), .ZN(n761) );
  NAND2_X1 U850 ( .A1(n762), .A2(n761), .ZN(G297) );
  INV_X1 U851 ( .A(G559), .ZN(n763) );
  NOR2_X1 U852 ( .A1(n764), .A2(n763), .ZN(n765) );
  NOR2_X1 U853 ( .A1(n999), .A2(n765), .ZN(n766) );
  XOR2_X1 U854 ( .A(KEYINPUT16), .B(n766), .Z(G148) );
  NOR2_X1 U855 ( .A1(n997), .A2(G868), .ZN(n769) );
  INV_X1 U856 ( .A(n999), .ZN(n899) );
  NAND2_X1 U857 ( .A1(G868), .A2(n899), .ZN(n767) );
  NOR2_X1 U858 ( .A1(G559), .A2(n767), .ZN(n768) );
  NOR2_X1 U859 ( .A1(n769), .A2(n768), .ZN(G282) );
  NAND2_X1 U860 ( .A1(G67), .A2(n770), .ZN(n773) );
  NAND2_X1 U861 ( .A1(G55), .A2(n771), .ZN(n772) );
  NAND2_X1 U862 ( .A1(n773), .A2(n772), .ZN(n779) );
  NAND2_X1 U863 ( .A1(G93), .A2(n774), .ZN(n777) );
  NAND2_X1 U864 ( .A1(G80), .A2(n775), .ZN(n776) );
  NAND2_X1 U865 ( .A1(n777), .A2(n776), .ZN(n778) );
  OR2_X1 U866 ( .A1(n779), .A2(n778), .ZN(n793) );
  NAND2_X1 U867 ( .A1(G559), .A2(n899), .ZN(n780) );
  XOR2_X1 U868 ( .A(KEYINPUT77), .B(n780), .Z(n791) );
  XNOR2_X1 U869 ( .A(n997), .B(n791), .ZN(n781) );
  NOR2_X1 U870 ( .A1(G860), .A2(n781), .ZN(n782) );
  XOR2_X1 U871 ( .A(n793), .B(n782), .Z(n783) );
  XNOR2_X1 U872 ( .A(n783), .B(KEYINPUT78), .ZN(G145) );
  XNOR2_X1 U873 ( .A(n997), .B(G305), .ZN(n790) );
  XNOR2_X1 U874 ( .A(KEYINPUT81), .B(KEYINPUT19), .ZN(n784) );
  XOR2_X1 U875 ( .A(n784), .B(n793), .Z(n787) );
  XNOR2_X1 U876 ( .A(G166), .B(G290), .ZN(n785) );
  XNOR2_X1 U877 ( .A(n785), .B(G299), .ZN(n786) );
  XNOR2_X1 U878 ( .A(n787), .B(n786), .ZN(n788) );
  XNOR2_X1 U879 ( .A(n788), .B(G288), .ZN(n789) );
  XNOR2_X1 U880 ( .A(n790), .B(n789), .ZN(n898) );
  XNOR2_X1 U881 ( .A(n791), .B(n898), .ZN(n792) );
  NAND2_X1 U882 ( .A1(n792), .A2(G868), .ZN(n796) );
  NAND2_X1 U883 ( .A1(n794), .A2(n793), .ZN(n795) );
  NAND2_X1 U884 ( .A1(n796), .A2(n795), .ZN(G295) );
  NAND2_X1 U885 ( .A1(G2078), .A2(G2084), .ZN(n797) );
  XOR2_X1 U886 ( .A(KEYINPUT20), .B(n797), .Z(n798) );
  NAND2_X1 U887 ( .A1(G2090), .A2(n798), .ZN(n799) );
  XNOR2_X1 U888 ( .A(KEYINPUT21), .B(n799), .ZN(n800) );
  NAND2_X1 U889 ( .A1(n800), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U890 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U891 ( .A1(G483), .A2(G661), .ZN(n810) );
  NOR2_X1 U892 ( .A1(G235), .A2(G236), .ZN(n801) );
  XNOR2_X1 U893 ( .A(n801), .B(KEYINPUT83), .ZN(n802) );
  NOR2_X1 U894 ( .A1(G238), .A2(n802), .ZN(n803) );
  NAND2_X1 U895 ( .A1(G57), .A2(n803), .ZN(n830) );
  NAND2_X1 U896 ( .A1(n830), .A2(G567), .ZN(n809) );
  NOR2_X1 U897 ( .A1(G220), .A2(G219), .ZN(n804) );
  XOR2_X1 U898 ( .A(KEYINPUT22), .B(n804), .Z(n805) );
  NOR2_X1 U899 ( .A1(G218), .A2(n805), .ZN(n806) );
  NAND2_X1 U900 ( .A1(G96), .A2(n806), .ZN(n829) );
  NAND2_X1 U901 ( .A1(G2106), .A2(n829), .ZN(n807) );
  XNOR2_X1 U902 ( .A(KEYINPUT82), .B(n807), .ZN(n808) );
  NAND2_X1 U903 ( .A1(n809), .A2(n808), .ZN(n831) );
  NOR2_X1 U904 ( .A1(n810), .A2(n831), .ZN(n811) );
  XNOR2_X1 U905 ( .A(n811), .B(KEYINPUT84), .ZN(n828) );
  NAND2_X1 U906 ( .A1(G36), .A2(n828), .ZN(G176) );
  XNOR2_X1 U907 ( .A(G2443), .B(G2435), .ZN(n821) );
  XOR2_X1 U908 ( .A(G2454), .B(G2430), .Z(n813) );
  XNOR2_X1 U909 ( .A(G2446), .B(KEYINPUT103), .ZN(n812) );
  XNOR2_X1 U910 ( .A(n813), .B(n812), .ZN(n817) );
  XOR2_X1 U911 ( .A(G2451), .B(G2427), .Z(n815) );
  XNOR2_X1 U912 ( .A(G1348), .B(G1341), .ZN(n814) );
  XNOR2_X1 U913 ( .A(n815), .B(n814), .ZN(n816) );
  XOR2_X1 U914 ( .A(n817), .B(n816), .Z(n819) );
  XNOR2_X1 U915 ( .A(G2438), .B(KEYINPUT102), .ZN(n818) );
  XNOR2_X1 U916 ( .A(n819), .B(n818), .ZN(n820) );
  XNOR2_X1 U917 ( .A(n821), .B(n820), .ZN(n822) );
  NAND2_X1 U918 ( .A1(n822), .A2(G14), .ZN(n903) );
  XOR2_X1 U919 ( .A(KEYINPUT104), .B(n903), .Z(G401) );
  NAND2_X1 U920 ( .A1(G2106), .A2(n823), .ZN(G217) );
  NAND2_X1 U921 ( .A1(G15), .A2(G2), .ZN(n825) );
  INV_X1 U922 ( .A(G661), .ZN(n824) );
  NOR2_X1 U923 ( .A1(n825), .A2(n824), .ZN(n826) );
  XNOR2_X1 U924 ( .A(n826), .B(KEYINPUT105), .ZN(G259) );
  NAND2_X1 U925 ( .A1(G3), .A2(G1), .ZN(n827) );
  NAND2_X1 U926 ( .A1(n828), .A2(n827), .ZN(G188) );
  XOR2_X1 U927 ( .A(G96), .B(KEYINPUT106), .Z(G221) );
  NOR2_X1 U929 ( .A1(n830), .A2(n829), .ZN(G325) );
  INV_X1 U930 ( .A(G325), .ZN(G261) );
  INV_X1 U931 ( .A(n831), .ZN(G319) );
  XOR2_X1 U932 ( .A(KEYINPUT107), .B(G2090), .Z(n833) );
  XNOR2_X1 U933 ( .A(G2067), .B(G2084), .ZN(n832) );
  XNOR2_X1 U934 ( .A(n833), .B(n832), .ZN(n834) );
  XOR2_X1 U935 ( .A(n834), .B(G2100), .Z(n836) );
  XNOR2_X1 U936 ( .A(G2078), .B(G2072), .ZN(n835) );
  XNOR2_X1 U937 ( .A(n836), .B(n835), .ZN(n840) );
  XOR2_X1 U938 ( .A(G2096), .B(KEYINPUT43), .Z(n838) );
  XNOR2_X1 U939 ( .A(G2678), .B(KEYINPUT42), .ZN(n837) );
  XNOR2_X1 U940 ( .A(n838), .B(n837), .ZN(n839) );
  XOR2_X1 U941 ( .A(n840), .B(n839), .Z(G227) );
  XOR2_X1 U942 ( .A(KEYINPUT109), .B(G1956), .Z(n842) );
  XNOR2_X1 U943 ( .A(G1996), .B(G1991), .ZN(n841) );
  XNOR2_X1 U944 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U945 ( .A(n843), .B(KEYINPUT41), .Z(n845) );
  XNOR2_X1 U946 ( .A(G1966), .B(G1971), .ZN(n844) );
  XNOR2_X1 U947 ( .A(n845), .B(n844), .ZN(n849) );
  XOR2_X1 U948 ( .A(G1976), .B(G1981), .Z(n847) );
  XNOR2_X1 U949 ( .A(G1986), .B(G1961), .ZN(n846) );
  XNOR2_X1 U950 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U951 ( .A(n849), .B(n848), .Z(n851) );
  XNOR2_X1 U952 ( .A(KEYINPUT108), .B(G2474), .ZN(n850) );
  XNOR2_X1 U953 ( .A(n851), .B(n850), .ZN(G229) );
  NAND2_X1 U954 ( .A1(G124), .A2(n877), .ZN(n852) );
  XNOR2_X1 U955 ( .A(n852), .B(KEYINPUT44), .ZN(n853) );
  XNOR2_X1 U956 ( .A(n853), .B(KEYINPUT110), .ZN(n855) );
  NAND2_X1 U957 ( .A1(G100), .A2(n883), .ZN(n854) );
  NAND2_X1 U958 ( .A1(n855), .A2(n854), .ZN(n859) );
  NAND2_X1 U959 ( .A1(G112), .A2(n876), .ZN(n857) );
  NAND2_X1 U960 ( .A1(G136), .A2(n881), .ZN(n856) );
  NAND2_X1 U961 ( .A1(n857), .A2(n856), .ZN(n858) );
  NOR2_X1 U962 ( .A1(n859), .A2(n858), .ZN(n860) );
  XOR2_X1 U963 ( .A(KEYINPUT111), .B(n860), .Z(G162) );
  XNOR2_X1 U964 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n862) );
  XNOR2_X1 U965 ( .A(n959), .B(KEYINPUT114), .ZN(n861) );
  XNOR2_X1 U966 ( .A(n862), .B(n861), .ZN(n863) );
  XNOR2_X1 U967 ( .A(G162), .B(n863), .ZN(n875) );
  NAND2_X1 U968 ( .A1(G103), .A2(n883), .ZN(n865) );
  NAND2_X1 U969 ( .A1(G139), .A2(n881), .ZN(n864) );
  NAND2_X1 U970 ( .A1(n865), .A2(n864), .ZN(n871) );
  NAND2_X1 U971 ( .A1(n876), .A2(G115), .ZN(n866) );
  XOR2_X1 U972 ( .A(KEYINPUT115), .B(n866), .Z(n868) );
  NAND2_X1 U973 ( .A1(n877), .A2(G127), .ZN(n867) );
  NAND2_X1 U974 ( .A1(n868), .A2(n867), .ZN(n869) );
  XOR2_X1 U975 ( .A(KEYINPUT47), .B(n869), .Z(n870) );
  NOR2_X1 U976 ( .A1(n871), .A2(n870), .ZN(n872) );
  XOR2_X1 U977 ( .A(KEYINPUT116), .B(n872), .Z(n973) );
  XNOR2_X1 U978 ( .A(n873), .B(n973), .ZN(n874) );
  XNOR2_X1 U979 ( .A(n875), .B(n874), .ZN(n890) );
  NAND2_X1 U980 ( .A1(G118), .A2(n876), .ZN(n879) );
  NAND2_X1 U981 ( .A1(G130), .A2(n877), .ZN(n878) );
  NAND2_X1 U982 ( .A1(n879), .A2(n878), .ZN(n880) );
  XNOR2_X1 U983 ( .A(KEYINPUT112), .B(n880), .ZN(n888) );
  NAND2_X1 U984 ( .A1(n881), .A2(G142), .ZN(n882) );
  XOR2_X1 U985 ( .A(KEYINPUT113), .B(n882), .Z(n885) );
  NAND2_X1 U986 ( .A1(n883), .A2(G106), .ZN(n884) );
  NAND2_X1 U987 ( .A1(n885), .A2(n884), .ZN(n886) );
  XOR2_X1 U988 ( .A(n886), .B(KEYINPUT45), .Z(n887) );
  NOR2_X1 U989 ( .A1(n888), .A2(n887), .ZN(n889) );
  XOR2_X1 U990 ( .A(n890), .B(n889), .Z(n896) );
  XOR2_X1 U991 ( .A(G164), .B(G160), .Z(n891) );
  XNOR2_X1 U992 ( .A(n892), .B(n891), .ZN(n893) );
  XNOR2_X1 U993 ( .A(n894), .B(n893), .ZN(n895) );
  XNOR2_X1 U994 ( .A(n896), .B(n895), .ZN(n897) );
  NOR2_X1 U995 ( .A1(G37), .A2(n897), .ZN(G395) );
  XOR2_X1 U996 ( .A(n898), .B(G286), .Z(n901) );
  XNOR2_X1 U997 ( .A(G171), .B(n899), .ZN(n900) );
  XNOR2_X1 U998 ( .A(n901), .B(n900), .ZN(n902) );
  NOR2_X1 U999 ( .A1(G37), .A2(n902), .ZN(G397) );
  NAND2_X1 U1000 ( .A1(G319), .A2(n903), .ZN(n906) );
  NOR2_X1 U1001 ( .A1(G227), .A2(G229), .ZN(n904) );
  XNOR2_X1 U1002 ( .A(KEYINPUT49), .B(n904), .ZN(n905) );
  NOR2_X1 U1003 ( .A1(n906), .A2(n905), .ZN(n908) );
  NOR2_X1 U1004 ( .A1(G395), .A2(G397), .ZN(n907) );
  NAND2_X1 U1005 ( .A1(n908), .A2(n907), .ZN(G225) );
  INV_X1 U1006 ( .A(G225), .ZN(G308) );
  INV_X1 U1007 ( .A(G57), .ZN(G237) );
  XOR2_X1 U1008 ( .A(n909), .B(G27), .Z(n912) );
  XOR2_X1 U1009 ( .A(G33), .B(KEYINPUT120), .Z(n910) );
  XNOR2_X1 U1010 ( .A(G2072), .B(n910), .ZN(n911) );
  NAND2_X1 U1011 ( .A1(n912), .A2(n911), .ZN(n921) );
  XOR2_X1 U1012 ( .A(n913), .B(G25), .Z(n914) );
  NAND2_X1 U1013 ( .A1(G28), .A2(n914), .ZN(n915) );
  XNOR2_X1 U1014 ( .A(n915), .B(KEYINPUT119), .ZN(n919) );
  XNOR2_X1 U1015 ( .A(G2067), .B(G26), .ZN(n917) );
  XNOR2_X1 U1016 ( .A(G32), .B(G1996), .ZN(n916) );
  NOR2_X1 U1017 ( .A1(n917), .A2(n916), .ZN(n918) );
  NAND2_X1 U1018 ( .A1(n919), .A2(n918), .ZN(n920) );
  NOR2_X1 U1019 ( .A1(n921), .A2(n920), .ZN(n922) );
  XOR2_X1 U1020 ( .A(KEYINPUT53), .B(n922), .Z(n926) );
  XNOR2_X1 U1021 ( .A(KEYINPUT54), .B(KEYINPUT121), .ZN(n923) );
  XNOR2_X1 U1022 ( .A(n923), .B(G34), .ZN(n924) );
  XNOR2_X1 U1023 ( .A(G2084), .B(n924), .ZN(n925) );
  NAND2_X1 U1024 ( .A1(n926), .A2(n925), .ZN(n928) );
  XNOR2_X1 U1025 ( .A(G35), .B(G2090), .ZN(n927) );
  NOR2_X1 U1026 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1027 ( .A(KEYINPUT55), .B(n929), .ZN(n931) );
  INV_X1 U1028 ( .A(G29), .ZN(n930) );
  NAND2_X1 U1029 ( .A1(n931), .A2(n930), .ZN(n932) );
  NAND2_X1 U1030 ( .A1(n932), .A2(G11), .ZN(n933) );
  XNOR2_X1 U1031 ( .A(n933), .B(KEYINPUT122), .ZN(n958) );
  XNOR2_X1 U1032 ( .A(G21), .B(G1966), .ZN(n934) );
  XNOR2_X1 U1033 ( .A(n934), .B(KEYINPUT127), .ZN(n954) );
  XOR2_X1 U1034 ( .A(G1961), .B(G5), .Z(n945) );
  XNOR2_X1 U1035 ( .A(G1348), .B(KEYINPUT59), .ZN(n935) );
  XNOR2_X1 U1036 ( .A(n935), .B(G4), .ZN(n939) );
  XNOR2_X1 U1037 ( .A(G1956), .B(G20), .ZN(n937) );
  XNOR2_X1 U1038 ( .A(G6), .B(G1981), .ZN(n936) );
  NOR2_X1 U1039 ( .A1(n937), .A2(n936), .ZN(n938) );
  NAND2_X1 U1040 ( .A1(n939), .A2(n938), .ZN(n942) );
  XNOR2_X1 U1041 ( .A(G19), .B(G1341), .ZN(n940) );
  XNOR2_X1 U1042 ( .A(KEYINPUT126), .B(n940), .ZN(n941) );
  NOR2_X1 U1043 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1044 ( .A(KEYINPUT60), .B(n943), .ZN(n944) );
  NAND2_X1 U1045 ( .A1(n945), .A2(n944), .ZN(n952) );
  XNOR2_X1 U1046 ( .A(G1971), .B(G22), .ZN(n947) );
  XNOR2_X1 U1047 ( .A(G23), .B(G1976), .ZN(n946) );
  NOR2_X1 U1048 ( .A1(n947), .A2(n946), .ZN(n949) );
  XOR2_X1 U1049 ( .A(G1986), .B(G24), .Z(n948) );
  NAND2_X1 U1050 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1051 ( .A(KEYINPUT58), .B(n950), .ZN(n951) );
  NOR2_X1 U1052 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1053 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1054 ( .A(KEYINPUT61), .B(n955), .ZN(n956) );
  NOR2_X1 U1055 ( .A1(n956), .A2(G16), .ZN(n957) );
  NOR2_X1 U1056 ( .A1(n958), .A2(n957), .ZN(n984) );
  XNOR2_X1 U1057 ( .A(G160), .B(G2084), .ZN(n960) );
  NAND2_X1 U1058 ( .A1(n960), .A2(n959), .ZN(n961) );
  NOR2_X1 U1059 ( .A1(n962), .A2(n961), .ZN(n964) );
  NAND2_X1 U1060 ( .A1(n964), .A2(n963), .ZN(n970) );
  XNOR2_X1 U1061 ( .A(G2090), .B(G162), .ZN(n965) );
  XNOR2_X1 U1062 ( .A(n965), .B(KEYINPUT117), .ZN(n967) );
  NOR2_X1 U1063 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1064 ( .A(KEYINPUT51), .B(n968), .ZN(n969) );
  NOR2_X1 U1065 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1066 ( .A1(n972), .A2(n971), .ZN(n978) );
  XOR2_X1 U1067 ( .A(G164), .B(G2078), .Z(n975) );
  XNOR2_X1 U1068 ( .A(G2072), .B(n973), .ZN(n974) );
  NOR2_X1 U1069 ( .A1(n975), .A2(n974), .ZN(n976) );
  XOR2_X1 U1070 ( .A(KEYINPUT50), .B(n976), .Z(n977) );
  NOR2_X1 U1071 ( .A1(n978), .A2(n977), .ZN(n979) );
  XOR2_X1 U1072 ( .A(KEYINPUT52), .B(n979), .Z(n980) );
  NOR2_X1 U1073 ( .A1(KEYINPUT55), .A2(n980), .ZN(n981) );
  XOR2_X1 U1074 ( .A(KEYINPUT118), .B(n981), .Z(n982) );
  NAND2_X1 U1075 ( .A1(G29), .A2(n982), .ZN(n983) );
  NAND2_X1 U1076 ( .A1(n984), .A2(n983), .ZN(n1013) );
  XOR2_X1 U1077 ( .A(G16), .B(KEYINPUT56), .Z(n1011) );
  XNOR2_X1 U1078 ( .A(G1966), .B(G168), .ZN(n986) );
  NAND2_X1 U1079 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1080 ( .A(n987), .B(KEYINPUT57), .ZN(n1008) );
  XNOR2_X1 U1081 ( .A(n988), .B(G1956), .ZN(n990) );
  NAND2_X1 U1082 ( .A1(n990), .A2(n989), .ZN(n994) );
  NAND2_X1 U1083 ( .A1(G303), .A2(G1971), .ZN(n991) );
  NAND2_X1 U1084 ( .A1(n992), .A2(n991), .ZN(n993) );
  NOR2_X1 U1085 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1086 ( .A1(n996), .A2(n995), .ZN(n1006) );
  XOR2_X1 U1087 ( .A(n997), .B(G1341), .Z(n1004) );
  XNOR2_X1 U1088 ( .A(G171), .B(G1961), .ZN(n998) );
  XNOR2_X1 U1089 ( .A(n998), .B(KEYINPUT123), .ZN(n1001) );
  XNOR2_X1 U1090 ( .A(G1348), .B(n999), .ZN(n1000) );
  NOR2_X1 U1091 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1092 ( .A(KEYINPUT124), .B(n1002), .ZN(n1003) );
  NAND2_X1 U1093 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NOR2_X1 U1094 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1095 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1096 ( .A(n1009), .B(KEYINPUT125), .ZN(n1010) );
  NOR2_X1 U1097 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NOR2_X1 U1098 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1099 ( .A(n1014), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1100 ( .A(G311), .ZN(G150) );
endmodule

