//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 1 0 1 0 1 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 0 1 0 0 0 0 1 1 0 0 0 1 1 1 0 1 0 0 0 1 0 1 0 0 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:32 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n716, new_n717, new_n718, new_n719, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n750, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n912,
    new_n913, new_n915, new_n916, new_n917, new_n918, new_n919, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973;
  INV_X1    g000(.A(KEYINPUT10), .ZN(new_n187));
  INV_X1    g001(.A(G101), .ZN(new_n188));
  INV_X1    g002(.A(G104), .ZN(new_n189));
  AND2_X1   g003(.A1(KEYINPUT79), .A2(G107), .ZN(new_n190));
  NOR2_X1   g004(.A1(KEYINPUT79), .A2(G107), .ZN(new_n191));
  OAI21_X1  g005(.A(new_n189), .B1(new_n190), .B2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G107), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G104), .ZN(new_n194));
  AOI211_X1 g008(.A(KEYINPUT80), .B(new_n188), .C1(new_n192), .C2(new_n194), .ZN(new_n195));
  AOI21_X1  g009(.A(new_n188), .B1(new_n192), .B2(new_n194), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT80), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT79), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(new_n193), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT3), .ZN(new_n201));
  NAND2_X1  g015(.A1(KEYINPUT79), .A2(G107), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n200), .A2(new_n201), .A3(G104), .A4(new_n202), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n201), .B1(new_n193), .B2(G104), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(new_n194), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n203), .A2(new_n205), .A3(new_n188), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n195), .B1(new_n198), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G128), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n208), .A2(KEYINPUT1), .ZN(new_n209));
  INV_X1    g023(.A(G143), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G146), .ZN(new_n211));
  INV_X1    g025(.A(G146), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G143), .ZN(new_n213));
  AND3_X1   g027(.A1(new_n209), .A2(new_n211), .A3(new_n213), .ZN(new_n214));
  AND2_X1   g028(.A1(new_n211), .A2(new_n213), .ZN(new_n215));
  INV_X1    g029(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n213), .A2(KEYINPUT1), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G128), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n214), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n187), .B1(new_n207), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n201), .A2(G104), .ZN(new_n221));
  NOR3_X1   g035(.A1(new_n221), .A2(new_n190), .A3(new_n191), .ZN(new_n222));
  AOI21_X1  g036(.A(KEYINPUT3), .B1(new_n189), .B2(G107), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n189), .A2(G107), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g039(.A(G101), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n226), .A2(KEYINPUT4), .A3(new_n206), .ZN(new_n227));
  OAI21_X1  g041(.A(KEYINPUT64), .B1(new_n210), .B2(G146), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT64), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n229), .A2(new_n212), .A3(G143), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n228), .A2(new_n230), .A3(new_n211), .ZN(new_n231));
  AND2_X1   g045(.A1(KEYINPUT0), .A2(G128), .ZN(new_n232));
  NOR2_X1   g046(.A1(KEYINPUT0), .A2(G128), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  AOI22_X1  g048(.A1(new_n231), .A2(new_n234), .B1(new_n215), .B2(new_n232), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT4), .ZN(new_n236));
  OAI211_X1 g050(.A(new_n236), .B(G101), .C1(new_n222), .C2(new_n225), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n227), .A2(new_n235), .A3(new_n237), .ZN(new_n238));
  AOI21_X1  g052(.A(G104), .B1(new_n200), .B2(new_n202), .ZN(new_n239));
  OAI21_X1  g053(.A(G101), .B1(new_n239), .B2(new_n224), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n240), .A2(new_n206), .A3(KEYINPUT80), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n196), .A2(new_n197), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n214), .B1(new_n218), .B2(new_n231), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n244), .A2(new_n187), .ZN(new_n245));
  AND3_X1   g059(.A1(new_n243), .A2(KEYINPUT81), .A3(new_n245), .ZN(new_n246));
  AOI21_X1  g060(.A(KEYINPUT81), .B1(new_n243), .B2(new_n245), .ZN(new_n247));
  OAI211_X1 g061(.A(new_n220), .B(new_n238), .C1(new_n246), .C2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT11), .ZN(new_n249));
  INV_X1    g063(.A(G134), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n249), .B1(new_n250), .B2(G137), .ZN(new_n251));
  INV_X1    g065(.A(G137), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n252), .A2(KEYINPUT11), .A3(G134), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n250), .A2(G137), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n251), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  XNOR2_X1  g070(.A(KEYINPUT65), .B(G131), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT66), .ZN(new_n259));
  AND2_X1   g073(.A1(new_n255), .A2(new_n259), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n251), .A2(new_n253), .A3(KEYINPUT66), .A4(new_n254), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G131), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n258), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  XOR2_X1   g077(.A(new_n263), .B(KEYINPUT82), .Z(new_n264));
  NOR2_X1   g078(.A1(new_n248), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT84), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n219), .B1(new_n241), .B2(new_n242), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n238), .B1(new_n267), .B2(KEYINPUT10), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT81), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n218), .A2(new_n231), .ZN(new_n270));
  INV_X1    g084(.A(new_n214), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(KEYINPUT10), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n269), .B1(new_n207), .B2(new_n273), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n243), .A2(KEYINPUT81), .A3(new_n245), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n268), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(new_n263), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n266), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n248), .A2(KEYINPUT84), .A3(new_n263), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n265), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  OR2_X1    g094(.A1(KEYINPUT70), .A2(G953), .ZN(new_n281));
  NAND2_X1  g095(.A1(KEYINPUT70), .A2(G953), .ZN(new_n282));
  AND2_X1   g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(G227), .ZN(new_n284));
  XOR2_X1   g098(.A(G110), .B(G140), .Z(new_n285));
  XNOR2_X1  g099(.A(new_n284), .B(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  OAI21_X1  g101(.A(KEYINPUT86), .B1(new_n280), .B2(new_n287), .ZN(new_n288));
  OR2_X1    g102(.A1(new_n248), .A2(new_n264), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n274), .A2(new_n275), .ZN(new_n290));
  INV_X1    g104(.A(new_n268), .ZN(new_n291));
  AOI211_X1 g105(.A(new_n266), .B(new_n277), .C1(new_n290), .C2(new_n291), .ZN(new_n292));
  AOI21_X1  g106(.A(KEYINPUT84), .B1(new_n248), .B2(new_n263), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n289), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT86), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n294), .A2(new_n295), .A3(new_n286), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n243), .A2(new_n272), .ZN(new_n297));
  OAI211_X1 g111(.A(KEYINPUT12), .B(new_n263), .C1(new_n297), .C2(new_n267), .ZN(new_n298));
  OR2_X1    g112(.A1(new_n298), .A2(KEYINPUT83), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(KEYINPUT83), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n297), .A2(new_n267), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n301), .A2(new_n277), .ZN(new_n302));
  OAI211_X1 g116(.A(new_n299), .B(new_n300), .C1(KEYINPUT12), .C2(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n303), .A2(new_n289), .A3(new_n287), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n288), .A2(new_n296), .A3(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(G902), .ZN(new_n306));
  XOR2_X1   g120(.A(KEYINPUT85), .B(G469), .Z(new_n307));
  NAND3_X1  g121(.A1(new_n305), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n287), .B1(new_n303), .B2(new_n289), .ZN(new_n309));
  AOI211_X1 g123(.A(new_n286), .B(new_n265), .C1(new_n278), .C2(new_n279), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n306), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(G469), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n308), .A2(new_n312), .ZN(new_n313));
  XNOR2_X1  g127(.A(KEYINPUT9), .B(G234), .ZN(new_n314));
  OAI21_X1  g128(.A(G221), .B1(new_n314), .B2(G902), .ZN(new_n315));
  OAI21_X1  g129(.A(G214), .B1(G237), .B2(G902), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  OAI21_X1  g131(.A(G210), .B1(G237), .B2(G902), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT67), .ZN(new_n320));
  AND2_X1   g134(.A1(KEYINPUT69), .A2(G116), .ZN(new_n321));
  NOR2_X1   g135(.A1(KEYINPUT69), .A2(G116), .ZN(new_n322));
  INV_X1    g136(.A(G119), .ZN(new_n323));
  NOR3_X1   g137(.A1(new_n321), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT68), .ZN(new_n325));
  INV_X1    g139(.A(G116), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n325), .B1(new_n326), .B2(G119), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n323), .A2(KEYINPUT68), .A3(G116), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n320), .B1(new_n324), .B2(new_n329), .ZN(new_n330));
  XNOR2_X1  g144(.A(KEYINPUT2), .B(G113), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  OAI211_X1 g147(.A(new_n320), .B(new_n331), .C1(new_n324), .C2(new_n329), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n335), .A2(new_n237), .A3(new_n227), .ZN(new_n336));
  NOR3_X1   g150(.A1(new_n324), .A2(new_n329), .A3(new_n331), .ZN(new_n337));
  INV_X1    g151(.A(new_n324), .ZN(new_n338));
  INV_X1    g152(.A(new_n329), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n338), .A2(new_n339), .A3(KEYINPUT5), .ZN(new_n340));
  NOR3_X1   g154(.A1(new_n326), .A2(KEYINPUT5), .A3(G119), .ZN(new_n341));
  INV_X1    g155(.A(G113), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n337), .B1(new_n340), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n243), .A2(new_n344), .ZN(new_n345));
  XNOR2_X1  g159(.A(G110), .B(G122), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n336), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(KEYINPUT6), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n336), .A2(new_n345), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT87), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n346), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n348), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n349), .A2(KEYINPUT6), .A3(new_n351), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  XNOR2_X1  g169(.A(KEYINPUT77), .B(G125), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n235), .A2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT88), .ZN(new_n359));
  AOI22_X1  g173(.A1(new_n358), .A2(new_n359), .B1(new_n357), .B2(new_n244), .ZN(new_n360));
  OAI21_X1  g174(.A(KEYINPUT88), .B1(new_n235), .B2(new_n357), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(G224), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n363), .A2(G953), .ZN(new_n364));
  XNOR2_X1  g178(.A(new_n362), .B(new_n364), .ZN(new_n365));
  AND2_X1   g179(.A1(new_n355), .A2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT7), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n364), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n360), .A2(new_n361), .A3(new_n368), .ZN(new_n369));
  XNOR2_X1  g183(.A(new_n369), .B(KEYINPUT89), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n362), .B1(new_n367), .B2(new_n364), .ZN(new_n371));
  XNOR2_X1  g185(.A(new_n346), .B(KEYINPUT8), .ZN(new_n372));
  INV_X1    g186(.A(new_n345), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n243), .A2(new_n344), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n372), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n371), .A2(new_n375), .A3(new_n347), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n306), .B1(new_n370), .B2(new_n376), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n319), .B1(new_n366), .B2(new_n377), .ZN(new_n378));
  OR2_X1    g192(.A1(new_n370), .A2(new_n376), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n355), .A2(new_n365), .ZN(new_n380));
  NAND4_X1  g194(.A1(new_n379), .A2(new_n306), .A3(new_n380), .A4(new_n318), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n317), .B1(new_n378), .B2(new_n381), .ZN(new_n382));
  AND3_X1   g196(.A1(new_n313), .A2(new_n315), .A3(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(G237), .ZN(new_n384));
  OR2_X1    g198(.A1(KEYINPUT90), .A2(G143), .ZN(new_n385));
  NAND4_X1  g199(.A1(new_n283), .A2(G214), .A3(new_n384), .A4(new_n385), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n281), .A2(G214), .A3(new_n384), .A4(new_n282), .ZN(new_n387));
  XNOR2_X1  g201(.A(KEYINPUT90), .B(G143), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(new_n257), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT17), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n386), .A2(new_n389), .A3(new_n257), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n392), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT16), .ZN(new_n396));
  INV_X1    g210(.A(G140), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n356), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  NOR2_X1   g212(.A1(G125), .A2(G140), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n399), .B1(new_n356), .B2(G140), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n398), .B1(new_n400), .B2(new_n396), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(new_n212), .ZN(new_n402));
  OAI211_X1 g216(.A(G146), .B(new_n398), .C1(new_n400), .C2(new_n396), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n390), .A2(KEYINPUT17), .A3(new_n391), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n395), .A2(new_n402), .A3(new_n403), .A4(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(KEYINPUT18), .A2(G131), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  OAI21_X1  g221(.A(KEYINPUT91), .B1(new_n390), .B2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT91), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n386), .A2(new_n409), .A3(new_n406), .A4(new_n389), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  XNOR2_X1  g225(.A(G125), .B(G140), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(new_n212), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n400), .A2(G146), .ZN(new_n414));
  AOI22_X1  g228(.A1(new_n390), .A2(new_n407), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n411), .A2(new_n415), .ZN(new_n416));
  XNOR2_X1  g230(.A(G113), .B(G122), .ZN(new_n417));
  XNOR2_X1  g231(.A(KEYINPUT93), .B(G104), .ZN(new_n418));
  XOR2_X1   g232(.A(new_n417), .B(new_n418), .Z(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n405), .A2(new_n416), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(KEYINPUT94), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT94), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n405), .A2(new_n416), .A3(new_n423), .A4(new_n420), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n405), .A2(new_n416), .ZN(new_n425));
  AOI22_X1  g239(.A1(new_n422), .A2(new_n424), .B1(new_n419), .B2(new_n425), .ZN(new_n426));
  OAI21_X1  g240(.A(KEYINPUT95), .B1(new_n426), .B2(G902), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n425), .A2(new_n419), .ZN(new_n428));
  AND3_X1   g242(.A1(new_n404), .A2(new_n402), .A3(new_n403), .ZN(new_n429));
  AOI22_X1  g243(.A1(new_n429), .A2(new_n395), .B1(new_n411), .B2(new_n415), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n423), .B1(new_n430), .B2(new_n420), .ZN(new_n431));
  INV_X1    g245(.A(new_n424), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n428), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT95), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n433), .A2(new_n434), .A3(new_n306), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n427), .A2(new_n435), .A3(G475), .ZN(new_n436));
  MUX2_X1   g250(.A(new_n412), .B(new_n400), .S(KEYINPUT19), .Z(new_n437));
  INV_X1    g251(.A(KEYINPUT92), .ZN(new_n438));
  OR3_X1    g252(.A1(new_n437), .A2(new_n438), .A3(G146), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n392), .A2(new_n394), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n438), .B1(new_n437), .B2(G146), .ZN(new_n441));
  NAND4_X1  g255(.A1(new_n439), .A2(new_n440), .A3(new_n403), .A4(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(new_n416), .ZN(new_n443));
  AOI22_X1  g257(.A1(new_n422), .A2(new_n424), .B1(new_n419), .B2(new_n443), .ZN(new_n444));
  NOR2_X1   g258(.A1(G475), .A2(G902), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(KEYINPUT20), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n443), .A2(new_n419), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n448), .B1(new_n431), .B2(new_n432), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT20), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n449), .A2(new_n450), .A3(new_n445), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n447), .A2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(G953), .ZN(new_n453));
  AND2_X1   g267(.A1(new_n453), .A2(G952), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n455), .B1(G234), .B2(G237), .ZN(new_n456));
  AOI211_X1 g270(.A(new_n306), .B(new_n283), .C1(G234), .C2(G237), .ZN(new_n457));
  XNOR2_X1  g271(.A(KEYINPUT21), .B(G898), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n456), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  XNOR2_X1  g274(.A(KEYINPUT74), .B(G217), .ZN(new_n461));
  NOR3_X1   g275(.A1(new_n461), .A2(new_n314), .A3(G953), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n326), .A2(G122), .ZN(new_n464));
  XNOR2_X1  g278(.A(new_n464), .B(KEYINPUT96), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n321), .A2(new_n322), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(G122), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n190), .A2(new_n191), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n465), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(KEYINPUT99), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n208), .A2(G143), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT98), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n471), .B(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n210), .A2(G128), .ZN(new_n474));
  AOI21_X1  g288(.A(G134), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n473), .A2(G134), .A3(new_n474), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT99), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n465), .A2(new_n467), .A3(new_n478), .A4(new_n468), .ZN(new_n479));
  NAND4_X1  g293(.A1(new_n470), .A2(new_n476), .A3(new_n477), .A4(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n467), .A2(KEYINPUT14), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT14), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n466), .A2(new_n482), .A3(G122), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n481), .A2(new_n465), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(G107), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT100), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n484), .A2(KEYINPUT100), .A3(G107), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n480), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  OAI21_X1  g303(.A(G134), .B1(KEYINPUT97), .B2(KEYINPUT13), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n490), .B1(KEYINPUT97), .B2(KEYINPUT13), .ZN(new_n491));
  INV_X1    g305(.A(new_n477), .ZN(new_n492));
  OAI211_X1 g306(.A(new_n473), .B(new_n491), .C1(new_n492), .C2(new_n475), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n473), .A2(new_n491), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n476), .A2(new_n477), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n465), .A2(new_n467), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n496), .B1(new_n191), .B2(new_n190), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(new_n469), .ZN(new_n498));
  AND3_X1   g312(.A1(new_n493), .A2(new_n495), .A3(new_n498), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n463), .B1(new_n489), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n493), .A2(new_n498), .A3(new_n495), .ZN(new_n501));
  AND2_X1   g315(.A1(new_n487), .A2(new_n488), .ZN(new_n502));
  OAI211_X1 g316(.A(new_n501), .B(new_n462), .C1(new_n502), .C2(new_n480), .ZN(new_n503));
  AOI21_X1  g317(.A(G902), .B1(new_n500), .B2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(G478), .ZN(new_n505));
  OR2_X1    g319(.A1(KEYINPUT101), .A2(KEYINPUT15), .ZN(new_n506));
  NAND2_X1  g320(.A1(KEYINPUT101), .A2(KEYINPUT15), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n505), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n504), .B(new_n508), .ZN(new_n509));
  NAND4_X1  g323(.A1(new_n436), .A2(new_n452), .A3(new_n460), .A4(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT102), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n510), .B(new_n511), .ZN(new_n512));
  AND2_X1   g326(.A1(new_n383), .A2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT30), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n263), .A2(new_n235), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n252), .A2(G134), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(new_n254), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(G131), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n518), .B1(new_n391), .B2(new_n255), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(new_n272), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n514), .B1(new_n515), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n231), .A2(new_n234), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n215), .A2(new_n232), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n255), .A2(new_n259), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n526), .A2(G131), .A3(new_n261), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n525), .B1(new_n527), .B2(new_n258), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n244), .A2(new_n519), .ZN(new_n529));
  NOR3_X1   g343(.A1(new_n528), .A2(KEYINPUT30), .A3(new_n529), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n335), .B1(new_n522), .B2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT31), .ZN(new_n532));
  AND2_X1   g346(.A1(new_n333), .A2(new_n334), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n515), .A2(new_n533), .A3(new_n521), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n283), .A2(G210), .A3(new_n384), .ZN(new_n535));
  OR2_X1    g349(.A1(new_n535), .A2(KEYINPUT27), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(KEYINPUT27), .ZN(new_n537));
  XNOR2_X1  g351(.A(KEYINPUT26), .B(G101), .ZN(new_n538));
  AND3_X1   g352(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n538), .B1(new_n536), .B2(new_n537), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND4_X1  g355(.A1(new_n531), .A2(new_n532), .A3(new_n534), .A4(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT71), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NOR3_X1   g358(.A1(new_n528), .A2(new_n335), .A3(new_n529), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n515), .A2(new_n514), .A3(new_n521), .ZN(new_n546));
  OAI21_X1  g360(.A(KEYINPUT30), .B1(new_n528), .B2(new_n529), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n545), .B1(new_n548), .B2(new_n335), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n549), .A2(KEYINPUT71), .A3(new_n532), .A4(new_n541), .ZN(new_n550));
  AOI22_X1  g364(.A1(new_n263), .A2(new_n235), .B1(new_n272), .B2(new_n520), .ZN(new_n551));
  AOI21_X1  g365(.A(KEYINPUT28), .B1(new_n551), .B2(new_n533), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n335), .B1(new_n528), .B2(new_n529), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n534), .A2(new_n553), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n552), .B1(new_n554), .B2(KEYINPUT28), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n532), .B1(new_n555), .B2(new_n541), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n549), .A2(new_n541), .ZN(new_n557));
  AOI22_X1  g371(.A1(new_n544), .A2(new_n550), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NOR2_X1   g372(.A1(G472), .A2(G902), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  OAI21_X1  g374(.A(KEYINPUT32), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n544), .A2(new_n550), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n556), .A2(new_n557), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT32), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n564), .A2(new_n565), .A3(new_n559), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT73), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n533), .B1(new_n515), .B2(new_n521), .ZN(new_n568));
  OAI21_X1  g382(.A(KEYINPUT28), .B1(new_n568), .B2(new_n545), .ZN(new_n569));
  INV_X1    g383(.A(new_n552), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT29), .ZN(new_n571));
  NOR3_X1   g385(.A1(new_n539), .A2(new_n540), .A3(new_n571), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n569), .A2(KEYINPUT72), .A3(new_n570), .A4(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(new_n306), .ZN(new_n574));
  AOI21_X1  g388(.A(KEYINPUT72), .B1(new_n555), .B2(new_n572), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n567), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n569), .A2(new_n570), .A3(new_n572), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT72), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND4_X1  g393(.A1(new_n579), .A2(KEYINPUT73), .A3(new_n306), .A4(new_n573), .ZN(new_n580));
  INV_X1    g394(.A(new_n541), .ZN(new_n581));
  AND2_X1   g395(.A1(new_n549), .A2(new_n581), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n555), .A2(new_n581), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n571), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n576), .A2(new_n580), .A3(new_n584), .ZN(new_n585));
  AOI22_X1  g399(.A1(new_n561), .A2(new_n566), .B1(G472), .B2(new_n585), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n461), .B1(G234), .B2(new_n306), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT25), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n208), .A2(G119), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n323), .A2(G128), .ZN(new_n591));
  AND2_X1   g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  XOR2_X1   g406(.A(KEYINPUT24), .B(G110), .Z(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  OR2_X1    g408(.A1(new_n594), .A2(KEYINPUT75), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(KEYINPUT75), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT76), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n590), .A2(new_n597), .ZN(new_n598));
  OR2_X1    g412(.A1(new_n598), .A2(KEYINPUT23), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(KEYINPUT23), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n599), .A2(new_n591), .A3(new_n600), .ZN(new_n601));
  AOI22_X1  g415(.A1(new_n595), .A2(new_n596), .B1(new_n601), .B2(G110), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n402), .A2(new_n403), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  OAI22_X1  g418(.A1(new_n601), .A2(G110), .B1(new_n592), .B2(new_n593), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n605), .A2(new_n413), .A3(new_n403), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n283), .A2(G221), .A3(G234), .ZN(new_n608));
  XNOR2_X1  g422(.A(KEYINPUT22), .B(G137), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n608), .B(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n607), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n604), .A2(new_n606), .A3(new_n610), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n589), .B1(new_n614), .B2(G902), .ZN(new_n615));
  NAND4_X1  g429(.A1(new_n612), .A2(KEYINPUT25), .A3(new_n306), .A4(new_n613), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n588), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NOR3_X1   g431(.A1(new_n614), .A2(G902), .A3(new_n587), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  OAI21_X1  g434(.A(KEYINPUT78), .B1(new_n586), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n585), .A2(G472), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n565), .B1(new_n564), .B2(new_n559), .ZN(new_n623));
  NOR3_X1   g437(.A1(new_n558), .A2(KEYINPUT32), .A3(new_n560), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n622), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT78), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n625), .A2(new_n626), .A3(new_n619), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n621), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n513), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(G101), .ZN(G3));
  OAI21_X1  g444(.A(G472), .B1(new_n558), .B2(G902), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n564), .A2(new_n559), .ZN(new_n632));
  AND3_X1   g446(.A1(new_n631), .A2(new_n632), .A3(new_n619), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n313), .A2(new_n315), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(KEYINPUT103), .ZN(new_n635));
  INV_X1    g449(.A(new_n315), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n636), .B1(new_n308), .B2(new_n312), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT103), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n637), .A2(new_n638), .A3(new_n633), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n436), .A2(new_n452), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n500), .A2(new_n503), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n500), .A2(KEYINPUT104), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n641), .A2(new_n642), .A3(KEYINPUT33), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT33), .ZN(new_n644));
  OAI211_X1 g458(.A(new_n500), .B(new_n503), .C1(KEYINPUT104), .C2(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n643), .A2(G478), .A3(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n504), .A2(new_n505), .ZN(new_n647));
  NAND2_X1  g461(.A1(G478), .A2(G902), .ZN(new_n648));
  AND3_X1   g462(.A1(new_n646), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n640), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n382), .A2(new_n460), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n635), .A2(new_n639), .A3(new_n652), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT34), .B(G104), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G6));
  INV_X1    g469(.A(new_n640), .ZN(new_n656));
  AOI211_X1 g470(.A(new_n459), .B(new_n317), .C1(new_n378), .C2(new_n381), .ZN(new_n657));
  XOR2_X1   g471(.A(new_n504), .B(new_n508), .Z(new_n658));
  NAND4_X1  g472(.A1(new_n656), .A2(new_n657), .A3(KEYINPUT105), .A4(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT105), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n436), .A2(new_n658), .A3(new_n452), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n660), .B1(new_n651), .B2(new_n661), .ZN(new_n662));
  AND2_X1   g476(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n663), .A2(new_n635), .A3(new_n639), .ZN(new_n664));
  XOR2_X1   g478(.A(KEYINPUT35), .B(G107), .Z(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G9));
  NAND2_X1  g480(.A1(new_n631), .A2(new_n632), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n587), .A2(G902), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n611), .A2(KEYINPUT36), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n607), .B(new_n669), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n617), .B1(new_n668), .B2(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n667), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n513), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(KEYINPUT106), .ZN(new_n674));
  XNOR2_X1  g488(.A(KEYINPUT37), .B(G110), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G12));
  NAND2_X1  g490(.A1(new_n561), .A2(new_n566), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n671), .B1(new_n677), .B2(new_n622), .ZN(new_n678));
  INV_X1    g492(.A(G900), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n456), .B1(new_n457), .B2(new_n679), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n661), .A2(new_n680), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n637), .A2(new_n678), .A3(new_n382), .A4(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G128), .ZN(G30));
  XNOR2_X1  g497(.A(new_n680), .B(KEYINPUT39), .ZN(new_n684));
  AOI211_X1 g498(.A(new_n636), .B(new_n684), .C1(new_n308), .C2(new_n312), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(KEYINPUT40), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT107), .ZN(new_n687));
  OR2_X1    g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n686), .A2(new_n687), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n671), .A2(new_n658), .ZN(new_n690));
  NOR3_X1   g504(.A1(new_n656), .A2(new_n690), .A3(new_n317), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n549), .A2(new_n581), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n306), .B1(new_n554), .B2(new_n541), .ZN(new_n693));
  OAI21_X1  g507(.A(G472), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n677), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n378), .A2(new_n381), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(KEYINPUT38), .ZN(new_n697));
  AND3_X1   g511(.A1(new_n691), .A2(new_n695), .A3(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n688), .A2(new_n689), .A3(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G143), .ZN(G45));
  INV_X1    g514(.A(new_n680), .ZN(new_n701));
  AND3_X1   g515(.A1(new_n640), .A2(new_n649), .A3(new_n701), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n637), .A2(new_n702), .A3(new_n678), .A4(new_n382), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G146), .ZN(G48));
  NAND2_X1  g518(.A1(new_n305), .A2(new_n306), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(G469), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n706), .A2(new_n315), .A3(new_n308), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n620), .B1(new_n677), .B2(new_n622), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(new_n652), .ZN(new_n711));
  XNOR2_X1  g525(.A(KEYINPUT41), .B(G113), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n711), .B(new_n712), .ZN(G15));
  NAND2_X1  g527(.A1(new_n710), .A2(new_n663), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G116), .ZN(G18));
  XNOR2_X1  g529(.A(new_n510), .B(KEYINPUT102), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n706), .A2(new_n315), .A3(new_n308), .A4(new_n382), .ZN(new_n717));
  INV_X1    g531(.A(new_n678), .ZN(new_n718));
  NOR3_X1   g532(.A1(new_n716), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(new_n323), .ZN(G21));
  INV_X1    g534(.A(new_n707), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n619), .A2(KEYINPUT108), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT108), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n723), .B1(new_n617), .B2(new_n618), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n725), .A2(new_n632), .A3(new_n631), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n640), .A2(new_n382), .A3(new_n460), .A4(new_n658), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n721), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G122), .ZN(G24));
  INV_X1    g544(.A(new_n717), .ZN(new_n731));
  OAI21_X1  g545(.A(KEYINPUT109), .B1(new_n667), .B2(new_n671), .ZN(new_n732));
  INV_X1    g546(.A(new_n617), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n670), .A2(new_n668), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT109), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n735), .A2(new_n631), .A3(new_n736), .A4(new_n632), .ZN(new_n737));
  AND2_X1   g551(.A1(new_n732), .A2(new_n737), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n731), .A2(new_n702), .A3(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G125), .ZN(G27));
  INV_X1    g554(.A(new_n702), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n741), .A2(KEYINPUT42), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n378), .A2(new_n381), .A3(new_n315), .A4(new_n316), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n743), .B1(new_n308), .B2(new_n312), .ZN(new_n744));
  AND2_X1   g558(.A1(new_n744), .A2(new_n708), .ZN(new_n745));
  AOI22_X1  g559(.A1(new_n677), .A2(new_n622), .B1(new_n722), .B2(new_n724), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n744), .A2(new_n746), .A3(new_n702), .ZN(new_n747));
  AOI22_X1  g561(.A1(new_n742), .A2(new_n745), .B1(new_n747), .B2(KEYINPUT42), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G131), .ZN(G33));
  NAND3_X1  g563(.A1(new_n744), .A2(new_n708), .A3(new_n681), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G134), .ZN(G36));
  AND2_X1   g565(.A1(G469), .A2(G902), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n309), .A2(new_n310), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(KEYINPUT45), .ZN(new_n754));
  XOR2_X1   g568(.A(new_n754), .B(KEYINPUT110), .Z(new_n755));
  OAI21_X1  g569(.A(G469), .B1(new_n753), .B2(KEYINPUT45), .ZN(new_n756));
  INV_X1    g570(.A(new_n756), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n752), .B1(new_n755), .B2(new_n757), .ZN(new_n758));
  AND2_X1   g572(.A1(new_n758), .A2(KEYINPUT46), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n308), .B1(new_n758), .B2(KEYINPUT46), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n315), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  OR3_X1    g575(.A1(new_n761), .A2(KEYINPUT111), .A3(new_n684), .ZN(new_n762));
  OAI21_X1  g576(.A(KEYINPUT111), .B1(new_n761), .B2(new_n684), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n378), .A2(new_n316), .A3(new_n381), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(KEYINPUT112), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n656), .A2(new_n649), .ZN(new_n766));
  XOR2_X1   g580(.A(new_n766), .B(KEYINPUT43), .Z(new_n767));
  NAND3_X1  g581(.A1(new_n767), .A2(new_n667), .A3(new_n735), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(KEYINPUT44), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n762), .A2(new_n763), .A3(new_n765), .A4(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G137), .ZN(G39));
  INV_X1    g585(.A(KEYINPUT47), .ZN(new_n772));
  OR2_X1    g586(.A1(new_n761), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n761), .A2(new_n772), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NOR3_X1   g589(.A1(new_n741), .A2(new_n619), .A3(new_n764), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n775), .A2(new_n586), .A3(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G140), .ZN(G42));
  INV_X1    g592(.A(new_n456), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n726), .A2(new_n779), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n767), .A2(new_n780), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n707), .A2(new_n316), .A3(new_n697), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  XOR2_X1   g597(.A(new_n783), .B(KEYINPUT50), .Z(new_n784));
  AND2_X1   g598(.A1(new_n706), .A2(new_n308), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n743), .A2(new_n779), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n767), .A2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n677), .A2(new_n619), .A3(new_n694), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n787), .A2(new_n791), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n640), .A2(new_n649), .ZN(new_n793));
  AOI22_X1  g607(.A1(new_n790), .A2(new_n738), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n784), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n781), .A2(new_n765), .ZN(new_n796));
  INV_X1    g610(.A(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n785), .A2(new_n636), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n773), .A2(new_n774), .A3(new_n798), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n795), .B1(new_n797), .B2(new_n799), .ZN(new_n800));
  OAI21_X1  g614(.A(KEYINPUT117), .B1(new_n800), .B2(KEYINPUT51), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT117), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT51), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n799), .A2(new_n797), .ZN(new_n804));
  OAI211_X1 g618(.A(new_n802), .B(new_n803), .C1(new_n804), .C2(new_n795), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n801), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n790), .A2(new_n746), .ZN(new_n807));
  XOR2_X1   g621(.A(KEYINPUT119), .B(KEYINPUT48), .Z(new_n808));
  XNOR2_X1  g622(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NOR3_X1   g623(.A1(new_n787), .A2(new_n650), .A3(new_n791), .ZN(new_n810));
  AOI211_X1 g624(.A(new_n455), .B(new_n810), .C1(new_n781), .C2(new_n731), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(KEYINPUT120), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n796), .B1(new_n799), .B2(KEYINPUT118), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n814), .B1(KEYINPUT118), .B2(new_n799), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n795), .A2(new_n803), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n813), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n806), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n702), .A2(new_n732), .A3(new_n737), .ZN(new_n819));
  OAI211_X1 g633(.A(new_n703), .B(new_n682), .C1(new_n717), .C2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n640), .A2(new_n382), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n821), .A2(new_n680), .A3(new_n690), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n822), .A2(new_n637), .A3(new_n695), .ZN(new_n823));
  INV_X1    g637(.A(new_n823), .ZN(new_n824));
  OAI21_X1  g638(.A(KEYINPUT52), .B1(new_n820), .B2(new_n824), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n703), .A2(new_n682), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT52), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n826), .A2(new_n827), .A3(new_n739), .A4(new_n823), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n825), .A2(new_n828), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n744), .A2(new_n702), .A3(new_n732), .A4(new_n737), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n378), .A2(new_n381), .A3(new_n316), .A4(new_n701), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n640), .A2(new_n831), .A3(new_n658), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n637), .A2(new_n678), .A3(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n830), .A2(new_n750), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n834), .A2(KEYINPUT113), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT113), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n830), .A2(new_n750), .A3(new_n833), .A4(new_n836), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  OAI211_X1 g652(.A(new_n512), .B(new_n383), .C1(new_n628), .C2(new_n672), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n651), .A2(new_n661), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n635), .A2(new_n639), .A3(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n839), .A2(new_n653), .A3(new_n841), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n829), .A2(new_n838), .A3(new_n842), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n716), .A2(new_n718), .ZN(new_n844));
  AOI22_X1  g658(.A1(new_n731), .A2(new_n844), .B1(new_n710), .B2(new_n663), .ZN(new_n845));
  AOI22_X1  g659(.A1(new_n710), .A2(new_n652), .B1(new_n721), .B2(new_n728), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n845), .A2(new_n748), .A3(KEYINPUT53), .A4(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n843), .A2(new_n848), .ZN(new_n849));
  OR2_X1    g663(.A1(new_n849), .A2(KEYINPUT114), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n845), .A2(new_n846), .ZN(new_n851));
  INV_X1    g665(.A(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n843), .A2(new_n748), .A3(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT53), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n849), .A2(KEYINPUT114), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n850), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n857), .A2(KEYINPUT54), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT54), .ZN(new_n859));
  AND3_X1   g673(.A1(new_n839), .A2(new_n653), .A3(new_n841), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT115), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n835), .A2(new_n837), .ZN(new_n862));
  AND3_X1   g676(.A1(new_n860), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n861), .B1(new_n860), .B2(new_n862), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n829), .A2(new_n847), .ZN(new_n866));
  AOI21_X1  g680(.A(KEYINPUT116), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  OAI21_X1  g681(.A(KEYINPUT115), .B1(new_n838), .B2(new_n842), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n860), .A2(new_n861), .A3(new_n862), .ZN(new_n869));
  AND4_X1   g683(.A1(KEYINPUT116), .A2(new_n866), .A3(new_n868), .A4(new_n869), .ZN(new_n870));
  OAI211_X1 g684(.A(new_n855), .B(new_n859), .C1(new_n867), .C2(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n858), .A2(new_n871), .ZN(new_n872));
  OAI22_X1  g686(.A1(new_n818), .A2(new_n872), .B1(G952), .B2(G953), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT49), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n785), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n725), .A2(new_n315), .A3(new_n316), .ZN(new_n876));
  NOR4_X1   g690(.A1(new_n697), .A2(new_n876), .A3(new_n766), .A4(new_n695), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n785), .A2(new_n874), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n873), .B1(new_n875), .B2(new_n879), .ZN(G75));
  NOR2_X1   g694(.A1(new_n283), .A2(G952), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n881), .B(KEYINPUT122), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n855), .B1(new_n867), .B2(new_n870), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n883), .A2(G210), .A3(G902), .ZN(new_n884));
  INV_X1    g698(.A(new_n884), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n355), .B(new_n365), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n886), .B(KEYINPUT55), .ZN(new_n887));
  OR2_X1    g701(.A1(new_n887), .A2(KEYINPUT56), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n882), .B1(new_n885), .B2(new_n888), .ZN(new_n889));
  AOI21_X1  g703(.A(KEYINPUT56), .B1(new_n884), .B2(KEYINPUT121), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n890), .B1(KEYINPUT121), .B2(new_n884), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n889), .B1(new_n891), .B2(new_n887), .ZN(G51));
  INV_X1    g706(.A(new_n881), .ZN(new_n893));
  INV_X1    g707(.A(new_n305), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n883), .A2(KEYINPUT54), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n895), .A2(new_n871), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n752), .B(KEYINPUT57), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n894), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  AND2_X1   g712(.A1(new_n755), .A2(new_n757), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n883), .A2(G902), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(KEYINPUT123), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT123), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n883), .A2(new_n902), .A3(G902), .A4(new_n899), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n893), .B1(new_n898), .B2(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT124), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  OAI211_X1 g721(.A(KEYINPUT124), .B(new_n893), .C1(new_n898), .C2(new_n904), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(G54));
  INV_X1    g723(.A(new_n883), .ZN(new_n910));
  NAND2_X1  g724(.A1(KEYINPUT58), .A2(G475), .ZN(new_n911));
  NOR3_X1   g725(.A1(new_n910), .A2(new_n306), .A3(new_n911), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n893), .B1(new_n912), .B2(new_n449), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n913), .B1(new_n449), .B2(new_n912), .ZN(G60));
  NAND2_X1  g728(.A1(new_n643), .A2(new_n645), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n648), .B(KEYINPUT59), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n896), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(new_n882), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n915), .B1(new_n872), .B2(new_n916), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n918), .A2(new_n919), .ZN(G63));
  NAND2_X1  g734(.A1(G217), .A2(G902), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(KEYINPUT60), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n910), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(new_n670), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n614), .B1(new_n910), .B2(new_n922), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n924), .A2(new_n882), .A3(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT61), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n926), .B(new_n927), .ZN(G66));
  NAND2_X1  g742(.A1(new_n852), .A2(new_n860), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n929), .A2(new_n283), .ZN(new_n930));
  OAI21_X1  g744(.A(G953), .B1(new_n458), .B2(new_n363), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  OAI211_X1 g746(.A(new_n353), .B(new_n354), .C1(G898), .C2(new_n283), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n932), .B(new_n933), .ZN(G69));
  INV_X1    g748(.A(new_n820), .ZN(new_n935));
  AND3_X1   g749(.A1(new_n935), .A2(new_n748), .A3(new_n750), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n762), .A2(new_n763), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n821), .A2(new_n509), .ZN(new_n938));
  AOI22_X1  g752(.A1(new_n769), .A2(new_n765), .B1(new_n938), .B2(new_n746), .ZN(new_n939));
  OAI211_X1 g753(.A(new_n777), .B(new_n936), .C1(new_n937), .C2(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(new_n283), .ZN(new_n941));
  OR2_X1    g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n548), .B(new_n437), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n943), .B1(G900), .B2(new_n941), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n764), .B1(new_n650), .B2(new_n661), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n628), .A2(new_n685), .A3(new_n946), .ZN(new_n947));
  AND2_X1   g761(.A1(new_n777), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n699), .A2(new_n935), .ZN(new_n949));
  OR2_X1    g763(.A1(new_n949), .A2(KEYINPUT62), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(KEYINPUT62), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n948), .A2(new_n770), .A3(new_n950), .A4(new_n951), .ZN(new_n952));
  AND2_X1   g766(.A1(new_n952), .A2(new_n283), .ZN(new_n953));
  INV_X1    g767(.A(new_n943), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n945), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(G227), .ZN(new_n956));
  OAI221_X1 g770(.A(new_n941), .B1(new_n956), .B2(new_n679), .C1(new_n943), .C2(KEYINPUT125), .ZN(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n955), .A2(new_n958), .ZN(new_n959));
  OAI211_X1 g773(.A(new_n945), .B(new_n957), .C1(new_n953), .C2(new_n954), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n959), .A2(new_n960), .ZN(G72));
  NAND2_X1  g775(.A1(G472), .A2(G902), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n962), .B(KEYINPUT63), .Z(new_n963));
  OAI21_X1  g777(.A(new_n963), .B1(new_n952), .B2(new_n929), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(new_n692), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n963), .B1(new_n940), .B2(new_n929), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT126), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  OAI211_X1 g782(.A(KEYINPUT126), .B(new_n963), .C1(new_n940), .C2(new_n929), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n968), .A2(new_n582), .A3(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(new_n582), .ZN(new_n971));
  INV_X1    g785(.A(new_n692), .ZN(new_n972));
  NAND4_X1  g786(.A1(new_n857), .A2(new_n971), .A3(new_n972), .A4(new_n963), .ZN(new_n973));
  AND4_X1   g787(.A1(new_n893), .A2(new_n965), .A3(new_n970), .A4(new_n973), .ZN(G57));
endmodule


