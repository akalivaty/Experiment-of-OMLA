//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 0 0 0 1 1 0 0 0 1 0 0 1 0 1 0 0 0 1 0 1 0 0 0 0 1 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 1 0 0 0 0 1 1 1 0 0 0 0 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:39 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n733, new_n734,
    new_n735, new_n737, new_n738, new_n739, new_n741, new_n742, new_n743,
    new_n744, new_n746, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n847, new_n848, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n934, new_n936, new_n937, new_n938, new_n939, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n967, new_n968, new_n969, new_n970, new_n972, new_n973;
  INV_X1    g000(.A(KEYINPUT3), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT74), .ZN(new_n203));
  AND2_X1   g002(.A1(G211gat), .A2(G218gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(G211gat), .A2(G218gat), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n203), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(G211gat), .ZN(new_n207));
  INV_X1    g006(.A(G218gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(G211gat), .A2(G218gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n209), .A2(KEYINPUT74), .A3(new_n210), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n206), .A2(new_n211), .A3(KEYINPUT73), .ZN(new_n212));
  INV_X1    g011(.A(G197gat), .ZN(new_n213));
  INV_X1    g012(.A(G204gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(G197gat), .A2(G204gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT22), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n210), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  XNOR2_X1  g019(.A(new_n212), .B(new_n220), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n202), .B1(new_n221), .B2(KEYINPUT29), .ZN(new_n222));
  INV_X1    g021(.A(G148gat), .ZN(new_n223));
  OAI21_X1  g022(.A(KEYINPUT78), .B1(new_n223), .B2(G141gat), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT78), .ZN(new_n225));
  INV_X1    g024(.A(G141gat), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n225), .A2(new_n226), .A3(G148gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n223), .A2(G141gat), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n224), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(G155gat), .ZN(new_n230));
  INV_X1    g029(.A(G162gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(G155gat), .A2(G162gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(KEYINPUT2), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(KEYINPUT79), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT79), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n233), .A2(new_n237), .A3(KEYINPUT2), .ZN(new_n238));
  NAND4_X1  g037(.A1(new_n229), .A2(new_n234), .A3(new_n236), .A4(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(G141gat), .B(G148gat), .ZN(new_n240));
  XNOR2_X1  g039(.A(KEYINPUT77), .B(KEYINPUT2), .ZN(new_n241));
  OAI211_X1 g040(.A(new_n233), .B(new_n232), .C1(new_n240), .C2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n239), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n222), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT29), .ZN(new_n245));
  XNOR2_X1  g044(.A(KEYINPUT80), .B(KEYINPUT3), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n245), .B1(new_n243), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(new_n221), .ZN(new_n248));
  NAND4_X1  g047(.A1(new_n244), .A2(G228gat), .A3(G233gat), .A4(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n206), .A2(new_n211), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(new_n220), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n206), .A2(new_n211), .A3(new_n219), .A4(new_n217), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n251), .A2(new_n245), .A3(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n246), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT85), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n255), .A2(new_n256), .A3(new_n243), .ZN(new_n257));
  AOI21_X1  g056(.A(KEYINPUT29), .B1(new_n250), .B2(new_n220), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n246), .B1(new_n258), .B2(new_n252), .ZN(new_n259));
  AND2_X1   g058(.A1(new_n239), .A2(new_n242), .ZN(new_n260));
  OAI21_X1  g059(.A(KEYINPUT85), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n257), .A2(new_n261), .A3(new_n248), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT86), .ZN(new_n263));
  NAND2_X1  g062(.A1(G228gat), .A2(G233gat), .ZN(new_n264));
  AND3_X1   g063(.A1(new_n262), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n263), .B1(new_n262), .B2(new_n264), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n249), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(KEYINPUT31), .B(G50gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(G78gat), .B(G106gat), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n270), .B(G22gat), .ZN(new_n271));
  INV_X1    g070(.A(new_n268), .ZN(new_n272));
  OAI211_X1 g071(.A(new_n272), .B(new_n249), .C1(new_n265), .C2(new_n266), .ZN(new_n273));
  AND3_X1   g072(.A1(new_n269), .A2(new_n271), .A3(new_n273), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n271), .B1(new_n269), .B2(new_n273), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(G57gat), .B(G85gat), .ZN(new_n277));
  XNOR2_X1  g076(.A(KEYINPUT83), .B(KEYINPUT0), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n277), .B(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(G1gat), .B(G29gat), .ZN(new_n280));
  XOR2_X1   g079(.A(new_n279), .B(new_n280), .Z(new_n281));
  INV_X1    g080(.A(G113gat), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n282), .A2(G120gat), .ZN(new_n283));
  INV_X1    g082(.A(G120gat), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n284), .A2(G113gat), .ZN(new_n285));
  OAI21_X1  g084(.A(KEYINPUT69), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(G127gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(G134gat), .ZN(new_n288));
  INV_X1    g087(.A(G134gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(G127gat), .ZN(new_n290));
  AND2_X1   g089(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n284), .A2(G113gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n282), .A2(G120gat), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT69), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n292), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(KEYINPUT70), .B(KEYINPUT1), .ZN(new_n296));
  NAND4_X1  g095(.A1(new_n286), .A2(new_n291), .A3(new_n295), .A4(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT68), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n288), .A2(new_n290), .A3(new_n298), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n287), .A2(KEYINPUT68), .A3(G134gat), .ZN(new_n300));
  XNOR2_X1  g099(.A(G113gat), .B(G120gat), .ZN(new_n301));
  OAI211_X1 g100(.A(new_n299), .B(new_n300), .C1(KEYINPUT1), .C2(new_n301), .ZN(new_n302));
  AND2_X1   g101(.A1(new_n297), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT81), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n303), .A2(new_n260), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n297), .A2(new_n302), .ZN(new_n306));
  OAI21_X1  g105(.A(KEYINPUT81), .B1(new_n306), .B2(new_n243), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n243), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n305), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(G225gat), .A2(G233gat), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT82), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT4), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n305), .A2(new_n315), .A3(new_n307), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n202), .B1(new_n239), .B2(new_n242), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  OAI211_X1 g117(.A(new_n318), .B(new_n306), .C1(new_n243), .C2(new_n246), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n303), .A2(new_n260), .A3(KEYINPUT4), .ZN(new_n320));
  NAND4_X1  g119(.A1(new_n316), .A2(new_n310), .A3(new_n319), .A4(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n309), .A2(KEYINPUT82), .A3(new_n311), .ZN(new_n322));
  NAND4_X1  g121(.A1(new_n314), .A2(KEYINPUT5), .A3(new_n321), .A4(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT87), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n306), .B1(new_n243), .B2(new_n246), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n325), .A2(new_n317), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n305), .A2(new_n307), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n326), .B1(new_n327), .B2(KEYINPUT4), .ZN(new_n328));
  AOI21_X1  g127(.A(KEYINPUT4), .B1(new_n303), .B2(new_n260), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n311), .A2(KEYINPUT5), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n328), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  AND3_X1   g131(.A1(new_n323), .A2(new_n324), .A3(new_n332), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n324), .B1(new_n323), .B2(new_n332), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  AOI21_X1  g134(.A(KEYINPUT39), .B1(new_n328), .B2(new_n330), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n315), .B1(new_n305), .B2(new_n307), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT39), .ZN(new_n338));
  NOR4_X1   g137(.A1(new_n337), .A2(new_n326), .A3(new_n338), .A4(new_n329), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n311), .B1(new_n336), .B2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(new_n281), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n309), .A2(KEYINPUT39), .A3(new_n310), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n340), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(KEYINPUT40), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT40), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n340), .A2(new_n345), .A3(new_n341), .A4(new_n342), .ZN(new_n346));
  AOI22_X1  g145(.A1(new_n281), .A2(new_n335), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT30), .ZN(new_n348));
  NAND2_X1  g147(.A1(G226gat), .A2(G233gat), .ZN(new_n349));
  XNOR2_X1  g148(.A(new_n349), .B(KEYINPUT75), .ZN(new_n350));
  NAND2_X1  g149(.A1(G169gat), .A2(G176gat), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT24), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n352), .A2(G183gat), .A3(G190gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(G183gat), .A2(G190gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(KEYINPUT24), .ZN(new_n355));
  NOR2_X1   g154(.A1(G183gat), .A2(G190gat), .ZN(new_n356));
  OAI211_X1 g155(.A(new_n351), .B(new_n353), .C1(new_n355), .C2(new_n356), .ZN(new_n357));
  NOR2_X1   g156(.A1(G169gat), .A2(G176gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(KEYINPUT23), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT23), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n360), .B1(G169gat), .B2(G176gat), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  OAI21_X1  g161(.A(KEYINPUT65), .B1(new_n357), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(KEYINPUT25), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT25), .ZN(new_n365));
  OAI211_X1 g164(.A(KEYINPUT65), .B(new_n365), .C1(new_n357), .C2(new_n362), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT26), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n351), .A2(new_n368), .ZN(new_n369));
  MUX2_X1   g168(.A(new_n369), .B(new_n368), .S(new_n358), .Z(new_n370));
  INV_X1    g169(.A(KEYINPUT28), .ZN(new_n371));
  NOR2_X1   g170(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n373), .A2(KEYINPUT67), .A3(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT67), .ZN(new_n376));
  AND2_X1   g175(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n376), .B1(new_n377), .B2(new_n372), .ZN(new_n378));
  AOI211_X1 g177(.A(new_n371), .B(G190gat), .C1(new_n375), .C2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(G190gat), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n380), .B1(new_n377), .B2(new_n372), .ZN(new_n381));
  XNOR2_X1  g180(.A(KEYINPUT66), .B(KEYINPUT28), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n381), .A2(new_n354), .A3(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n370), .B1(new_n379), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n367), .A2(new_n385), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n350), .B1(new_n386), .B2(new_n245), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n375), .A2(new_n378), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n388), .A2(KEYINPUT28), .A3(new_n380), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(new_n383), .ZN(new_n390));
  AOI22_X1  g189(.A1(new_n390), .A2(new_n370), .B1(new_n364), .B2(new_n366), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n391), .A2(new_n349), .ZN(new_n392));
  INV_X1    g191(.A(new_n221), .ZN(new_n393));
  NOR3_X1   g192(.A1(new_n387), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  AOI21_X1  g193(.A(KEYINPUT29), .B1(new_n367), .B2(new_n385), .ZN(new_n395));
  INV_X1    g194(.A(new_n349), .ZN(new_n396));
  OAI21_X1  g195(.A(KEYINPUT76), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n386), .A2(new_n350), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT76), .ZN(new_n399));
  OAI211_X1 g198(.A(new_n399), .B(new_n349), .C1(new_n391), .C2(KEYINPUT29), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n397), .A2(new_n398), .A3(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n394), .B1(new_n393), .B2(new_n401), .ZN(new_n402));
  XNOR2_X1  g201(.A(G8gat), .B(G36gat), .ZN(new_n403));
  XNOR2_X1  g202(.A(G64gat), .B(G92gat), .ZN(new_n404));
  XNOR2_X1  g203(.A(new_n403), .B(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n348), .B1(new_n402), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n401), .A2(new_n393), .ZN(new_n407));
  INV_X1    g206(.A(new_n394), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n405), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n406), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n409), .A2(new_n348), .A3(new_n410), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n276), .B1(new_n347), .B2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT88), .ZN(new_n417));
  NOR3_X1   g216(.A1(new_n333), .A2(new_n334), .A3(new_n341), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n323), .A2(new_n341), .A3(new_n332), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT6), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n417), .B1(new_n418), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n323), .A2(new_n332), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n423), .A2(KEYINPUT6), .A3(new_n281), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT89), .ZN(new_n425));
  XNOR2_X1  g224(.A(new_n424), .B(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n423), .A2(KEYINPUT87), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n323), .A2(new_n324), .A3(new_n332), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n427), .A2(new_n281), .A3(new_n428), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n429), .A2(KEYINPUT88), .A3(new_n420), .A4(new_n419), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n422), .A2(new_n426), .A3(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n407), .A2(KEYINPUT37), .A3(new_n408), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n432), .A2(KEYINPUT90), .A3(new_n405), .ZN(new_n433));
  OR2_X1    g232(.A1(new_n402), .A2(KEYINPUT37), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g234(.A(KEYINPUT90), .B1(new_n432), .B2(new_n405), .ZN(new_n436));
  OAI21_X1  g235(.A(KEYINPUT38), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n393), .B1(new_n387), .B2(new_n392), .ZN(new_n438));
  OAI211_X1 g237(.A(KEYINPUT37), .B(new_n438), .C1(new_n401), .C2(new_n393), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(new_n405), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n440), .A2(KEYINPUT38), .ZN(new_n441));
  AOI22_X1  g240(.A1(new_n441), .A2(new_n434), .B1(new_n409), .B2(new_n410), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n437), .A2(new_n442), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n416), .B1(new_n431), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n386), .A2(new_n306), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n391), .A2(new_n303), .ZN(new_n446));
  NAND2_X1  g245(.A1(G227gat), .A2(G233gat), .ZN(new_n447));
  XNOR2_X1  g246(.A(new_n447), .B(KEYINPUT64), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n445), .A2(new_n446), .A3(new_n449), .ZN(new_n450));
  XNOR2_X1  g249(.A(new_n450), .B(KEYINPUT34), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  XNOR2_X1  g251(.A(G15gat), .B(G43gat), .ZN(new_n453));
  INV_X1    g252(.A(G71gat), .ZN(new_n454));
  XNOR2_X1  g253(.A(new_n453), .B(new_n454), .ZN(new_n455));
  XNOR2_X1  g254(.A(new_n455), .B(G99gat), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n449), .B1(new_n445), .B2(new_n446), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n456), .B1(new_n457), .B2(KEYINPUT33), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT32), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  NOR2_X1   g259(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n462));
  AOI221_X4 g261(.A(new_n459), .B1(KEYINPUT33), .B2(new_n456), .C1(new_n462), .C2(new_n448), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n452), .B1(new_n461), .B2(new_n463), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n386), .A2(new_n306), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n303), .B1(new_n367), .B2(new_n385), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n448), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(KEYINPUT32), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT33), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n468), .A2(new_n470), .A3(new_n456), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n458), .A2(new_n460), .ZN(new_n472));
  AOI21_X1  g271(.A(KEYINPUT71), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  OAI22_X1  g272(.A1(new_n464), .A2(KEYINPUT71), .B1(new_n473), .B2(new_n452), .ZN(new_n474));
  AND3_X1   g273(.A1(new_n471), .A2(new_n472), .A3(new_n451), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n451), .B1(new_n471), .B2(new_n472), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  XOR2_X1   g276(.A(KEYINPUT72), .B(KEYINPUT36), .Z(new_n478));
  AOI22_X1  g277(.A1(new_n474), .A2(KEYINPUT36), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  AND3_X1   g278(.A1(new_n419), .A2(KEYINPUT84), .A3(new_n420), .ZN(new_n480));
  AOI21_X1  g279(.A(KEYINPUT84), .B1(new_n419), .B2(new_n420), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n341), .B1(new_n323), .B2(new_n332), .ZN(new_n482));
  NOR3_X1   g281(.A1(new_n480), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(new_n424), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n414), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n479), .B1(new_n485), .B2(new_n276), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n444), .A2(new_n486), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n276), .A2(new_n477), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n431), .A2(new_n414), .A3(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT35), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(new_n485), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n474), .B1(new_n274), .B2(new_n275), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT91), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(new_n276), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n496), .A2(KEYINPUT91), .A3(new_n474), .ZN(new_n497));
  NAND4_X1  g296(.A1(new_n492), .A2(new_n495), .A3(new_n497), .A4(KEYINPUT35), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n487), .A2(new_n491), .A3(new_n498), .ZN(new_n499));
  XNOR2_X1  g298(.A(G15gat), .B(G22gat), .ZN(new_n500));
  INV_X1    g299(.A(G1gat), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(KEYINPUT16), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n503), .B1(G1gat), .B2(new_n500), .ZN(new_n504));
  XOR2_X1   g303(.A(new_n504), .B(G8gat), .Z(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(KEYINPUT96), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n504), .B(G8gat), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT96), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT21), .ZN(new_n511));
  XNOR2_X1  g310(.A(G71gat), .B(G78gat), .ZN(new_n512));
  INV_X1    g311(.A(G57gat), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(G64gat), .ZN(new_n514));
  INV_X1    g313(.A(G64gat), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(G57gat), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n512), .B1(KEYINPUT9), .B2(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n518), .B(KEYINPUT97), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT98), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n516), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n515), .A2(KEYINPUT98), .A3(G57gat), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n521), .A2(new_n514), .A3(new_n522), .ZN(new_n523));
  AND2_X1   g322(.A1(G71gat), .A2(G78gat), .ZN(new_n524));
  OAI211_X1 g323(.A(new_n523), .B(new_n512), .C1(KEYINPUT9), .C2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n519), .A2(new_n525), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n510), .B1(new_n511), .B2(new_n526), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n527), .B(G183gat), .ZN(new_n528));
  INV_X1    g327(.A(new_n526), .ZN(new_n529));
  XNOR2_X1  g328(.A(KEYINPUT99), .B(KEYINPUT21), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  OR2_X1    g330(.A1(new_n527), .A2(G183gat), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n527), .A2(G183gat), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n529), .A2(new_n530), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n531), .A2(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(G127gat), .B(G155gat), .ZN(new_n537));
  XOR2_X1   g336(.A(new_n537), .B(KEYINPUT20), .Z(new_n538));
  NAND2_X1  g337(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(new_n538), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n531), .A2(new_n535), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  XNOR2_X1  g341(.A(KEYINPUT100), .B(KEYINPUT19), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n543), .B(G211gat), .ZN(new_n544));
  AND2_X1   g343(.A1(G231gat), .A2(G233gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n544), .B(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n542), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n539), .A2(new_n546), .A3(new_n541), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(G190gat), .B(G218gat), .ZN(new_n552));
  XOR2_X1   g351(.A(G43gat), .B(G50gat), .Z(new_n553));
  INV_X1    g352(.A(KEYINPUT15), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT95), .ZN(new_n556));
  NAND2_X1  g355(.A1(G29gat), .A2(G36gat), .ZN(new_n557));
  XOR2_X1   g356(.A(new_n557), .B(KEYINPUT93), .Z(new_n558));
  AOI21_X1  g357(.A(new_n555), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  OR2_X1    g358(.A1(new_n558), .A2(new_n556), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n553), .A2(new_n554), .ZN(new_n561));
  OR3_X1    g360(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n562));
  OR2_X1    g361(.A1(new_n562), .A2(KEYINPUT94), .ZN(new_n563));
  OAI21_X1  g362(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n562), .A2(KEYINPUT94), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  NAND4_X1  g365(.A1(new_n559), .A2(new_n560), .A3(new_n561), .A4(new_n566), .ZN(new_n567));
  AND2_X1   g366(.A1(new_n562), .A2(new_n564), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n555), .B1(new_n558), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT17), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n570), .B(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(G85gat), .A2(G92gat), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n573), .A2(KEYINPUT101), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT101), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n575), .A2(G85gat), .A3(G92gat), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n574), .A2(new_n576), .A3(KEYINPUT7), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT102), .ZN(new_n578));
  OAI211_X1 g377(.A(new_n577), .B(new_n578), .C1(KEYINPUT7), .C2(new_n573), .ZN(new_n579));
  NAND2_X1  g378(.A1(G99gat), .A2(G106gat), .ZN(new_n580));
  INV_X1    g379(.A(G85gat), .ZN(new_n581));
  INV_X1    g380(.A(G92gat), .ZN(new_n582));
  AOI22_X1  g381(.A1(KEYINPUT8), .A2(new_n580), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  OAI211_X1 g382(.A(new_n579), .B(new_n583), .C1(new_n578), .C2(new_n577), .ZN(new_n584));
  XOR2_X1   g383(.A(G99gat), .B(G106gat), .Z(new_n585));
  OR2_X1    g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n584), .A2(new_n585), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n586), .A2(KEYINPUT103), .A3(new_n587), .ZN(new_n588));
  OR3_X1    g387(.A1(new_n584), .A2(KEYINPUT103), .A3(new_n585), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n572), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n570), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n552), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n570), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(new_n571), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n570), .A2(KEYINPUT17), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n600), .A2(new_n589), .A3(new_n588), .ZN(new_n601));
  AND4_X1   g400(.A1(new_n595), .A2(new_n601), .A3(new_n592), .A4(new_n552), .ZN(new_n602));
  OAI21_X1  g401(.A(KEYINPUT104), .B1(new_n596), .B2(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n594), .A2(new_n595), .A3(new_n552), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n601), .A2(new_n595), .A3(new_n592), .ZN(new_n605));
  INV_X1    g404(.A(new_n552), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT104), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n604), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(G134gat), .B(G162gat), .ZN(new_n610));
  AOI21_X1  g409(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n610), .B(new_n611), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n603), .A2(new_n609), .A3(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n612), .ZN(new_n614));
  OAI211_X1 g413(.A(KEYINPUT104), .B(new_n614), .C1(new_n596), .C2(new_n602), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n551), .A2(new_n617), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n507), .B1(new_n598), .B2(new_n599), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n506), .A2(new_n509), .A3(new_n570), .ZN(new_n621));
  NAND2_X1  g420(.A1(G229gat), .A2(G233gat), .ZN(new_n622));
  NAND4_X1  g421(.A1(new_n620), .A2(KEYINPUT18), .A3(new_n621), .A4(new_n622), .ZN(new_n623));
  OAI211_X1 g422(.A(new_n621), .B(new_n622), .C1(new_n572), .C2(new_n507), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT18), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n510), .A2(new_n597), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n627), .A2(new_n621), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n622), .B(KEYINPUT13), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n623), .A2(new_n626), .A3(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(G169gat), .B(G197gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(KEYINPUT92), .B(KEYINPUT11), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(G113gat), .B(G141gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n638), .B(KEYINPUT12), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n633), .A2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n639), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n632), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(G230gat), .ZN(new_n645));
  INV_X1    g444(.A(G233gat), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n585), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n584), .B(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n649), .A2(new_n529), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(KEYINPUT105), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT10), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n588), .A2(new_n526), .A3(new_n589), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT105), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n649), .A2(new_n529), .A3(new_n654), .ZN(new_n655));
  NAND4_X1  g454(.A1(new_n651), .A2(new_n652), .A3(new_n653), .A4(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n590), .A2(KEYINPUT10), .A3(new_n529), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n647), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n647), .ZN(new_n659));
  AND2_X1   g458(.A1(new_n653), .A2(new_n655), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n659), .B1(new_n660), .B2(new_n651), .ZN(new_n661));
  OAI21_X1  g460(.A(KEYINPUT106), .B1(new_n658), .B2(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(G120gat), .B(G148gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(G176gat), .B(G204gat), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n663), .B(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n662), .A2(new_n666), .ZN(new_n667));
  OAI211_X1 g466(.A(KEYINPUT106), .B(new_n665), .C1(new_n658), .C2(new_n661), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n644), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n499), .A2(new_n618), .A3(new_n670), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(KEYINPUT107), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n483), .A2(new_n484), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(new_n501), .ZN(G1324gat));
  INV_X1    g475(.A(KEYINPUT108), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n677), .A2(KEYINPUT42), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n672), .A2(new_n414), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n679), .B1(new_n677), .B2(KEYINPUT42), .ZN(new_n680));
  XNOR2_X1  g479(.A(KEYINPUT16), .B(G8gat), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n678), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  OAI21_X1  g481(.A(G8gat), .B1(new_n672), .B2(new_n414), .ZN(new_n683));
  INV_X1    g482(.A(new_n681), .ZN(new_n684));
  NAND4_X1  g483(.A1(new_n679), .A2(new_n677), .A3(KEYINPUT42), .A4(new_n684), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n682), .A2(new_n683), .A3(new_n685), .ZN(G1325gat));
  NOR2_X1   g485(.A1(new_n672), .A2(new_n477), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n687), .A2(G15gat), .ZN(new_n688));
  INV_X1    g487(.A(new_n479), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n672), .A2(new_n689), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n688), .B1(G15gat), .B2(new_n690), .ZN(G1326gat));
  NOR2_X1   g490(.A1(new_n672), .A2(new_n496), .ZN(new_n692));
  XOR2_X1   g491(.A(KEYINPUT43), .B(G22gat), .Z(new_n693));
  XNOR2_X1  g492(.A(new_n692), .B(new_n693), .ZN(G1327gat));
  AOI22_X1  g493(.A1(new_n444), .A2(new_n486), .B1(new_n489), .B2(new_n490), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n616), .B1(new_n695), .B2(new_n498), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n551), .A2(new_n670), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(G29gat), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n700), .A2(new_n701), .A3(new_n673), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(KEYINPUT45), .ZN(new_n703));
  AND3_X1   g502(.A1(new_n613), .A2(new_n615), .A3(KEYINPUT109), .ZN(new_n704));
  AOI21_X1  g503(.A(KEYINPUT109), .B1(new_n613), .B2(new_n615), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT44), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n499), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n709), .B1(new_n696), .B2(new_n708), .ZN(new_n710));
  AND2_X1   g509(.A1(new_n710), .A2(new_n698), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(new_n673), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n703), .B1(new_n713), .B2(new_n701), .ZN(G1328gat));
  NOR3_X1   g513(.A1(new_n699), .A2(G36gat), .A3(new_n414), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT46), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  XOR2_X1   g516(.A(new_n717), .B(KEYINPUT110), .Z(new_n718));
  NAND2_X1  g517(.A1(new_n711), .A2(new_n415), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(G36gat), .ZN(new_n720));
  OAI211_X1 g519(.A(new_n718), .B(new_n720), .C1(new_n716), .C2(new_n715), .ZN(G1329gat));
  NAND3_X1  g520(.A1(new_n711), .A2(G43gat), .A3(new_n479), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n699), .A2(new_n477), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n722), .B1(G43gat), .B2(new_n723), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n724), .B(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g524(.A1(new_n711), .A2(new_n276), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(G50gat), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT48), .ZN(new_n728));
  OR3_X1    g527(.A1(new_n699), .A2(G50gat), .A3(new_n496), .ZN(new_n729));
  AND3_X1   g528(.A1(new_n727), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n728), .B1(new_n727), .B2(new_n729), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n730), .A2(new_n731), .ZN(G1331gat));
  AND3_X1   g531(.A1(new_n499), .A2(new_n618), .A3(new_n644), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(new_n669), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n734), .A2(new_n674), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(new_n513), .ZN(G1332gat));
  NAND3_X1  g535(.A1(new_n733), .A2(new_n669), .A3(new_n415), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n737), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n738));
  XOR2_X1   g537(.A(KEYINPUT49), .B(G64gat), .Z(new_n739));
  OAI21_X1  g538(.A(new_n738), .B1(new_n737), .B2(new_n739), .ZN(G1333gat));
  OAI21_X1  g539(.A(new_n454), .B1(new_n734), .B2(new_n477), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n689), .A2(new_n454), .ZN(new_n742));
  INV_X1    g541(.A(new_n742), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n741), .B1(new_n734), .B2(new_n743), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g544(.A1(new_n734), .A2(new_n496), .ZN(new_n746));
  XOR2_X1   g545(.A(new_n746), .B(G78gat), .Z(G1335gat));
  INV_X1    g546(.A(new_n669), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n550), .A2(new_n643), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n499), .A2(new_n617), .A3(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT51), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND4_X1  g551(.A1(new_n499), .A2(KEYINPUT51), .A3(new_n617), .A4(new_n749), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n748), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  AOI21_X1  g553(.A(G85gat), .B1(new_n754), .B2(new_n673), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n708), .B1(new_n499), .B2(new_n617), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n708), .B1(new_n704), .B2(new_n705), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n757), .B1(new_n695), .B2(new_n498), .ZN(new_n758));
  OAI211_X1 g557(.A(new_n669), .B(new_n749), .C1(new_n756), .C2(new_n758), .ZN(new_n759));
  NOR3_X1   g558(.A1(new_n759), .A2(new_n581), .A3(new_n674), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n755), .A2(new_n760), .ZN(G1336gat));
  OR3_X1    g560(.A1(new_n759), .A2(KEYINPUT112), .A3(new_n414), .ZN(new_n762));
  OAI21_X1  g561(.A(KEYINPUT112), .B1(new_n759), .B2(new_n414), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n762), .A2(G92gat), .A3(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT52), .ZN(new_n765));
  INV_X1    g564(.A(new_n754), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n415), .A2(new_n582), .ZN(new_n767));
  OAI211_X1 g566(.A(new_n764), .B(new_n765), .C1(new_n766), .C2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT111), .ZN(new_n769));
  AOI21_X1  g568(.A(KEYINPUT51), .B1(new_n696), .B2(new_n749), .ZN(new_n770));
  INV_X1    g569(.A(new_n753), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n769), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n769), .B1(new_n750), .B2(new_n751), .ZN(new_n773));
  INV_X1    g572(.A(new_n773), .ZN(new_n774));
  AOI211_X1 g573(.A(new_n748), .B(new_n767), .C1(new_n772), .C2(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(new_n759), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n582), .B1(new_n776), .B2(new_n415), .ZN(new_n777));
  OAI21_X1  g576(.A(KEYINPUT52), .B1(new_n775), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n768), .A2(new_n778), .ZN(G1337gat));
  OAI21_X1  g578(.A(G99gat), .B1(new_n759), .B2(new_n689), .ZN(new_n780));
  OR2_X1    g579(.A1(new_n477), .A2(G99gat), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n780), .B1(new_n766), .B2(new_n781), .ZN(G1338gat));
  INV_X1    g581(.A(KEYINPUT114), .ZN(new_n783));
  OAI21_X1  g582(.A(G106gat), .B1(new_n759), .B2(new_n496), .ZN(new_n784));
  NOR3_X1   g583(.A1(new_n748), .A2(new_n496), .A3(G106gat), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n785), .B1(new_n770), .B2(new_n771), .ZN(new_n786));
  XNOR2_X1  g585(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n784), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n774), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n710), .A2(new_n669), .A3(new_n276), .A4(new_n749), .ZN(new_n790));
  AOI22_X1  g589(.A1(new_n789), .A2(new_n785), .B1(G106gat), .B2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT53), .ZN(new_n792));
  OAI211_X1 g591(.A(new_n783), .B(new_n788), .C1(new_n791), .C2(new_n792), .ZN(new_n793));
  AOI21_X1  g592(.A(KEYINPUT111), .B1(new_n752), .B2(new_n753), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n785), .B1(new_n794), .B2(new_n773), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n792), .B1(new_n795), .B2(new_n784), .ZN(new_n796));
  AND3_X1   g595(.A1(new_n784), .A2(new_n786), .A3(new_n787), .ZN(new_n797));
  OAI21_X1  g596(.A(KEYINPUT114), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n793), .A2(new_n798), .ZN(G1339gat));
  INV_X1    g598(.A(KEYINPUT55), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n656), .A2(new_n657), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(new_n659), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n656), .A2(new_n647), .A3(new_n657), .ZN(new_n803));
  AND3_X1   g602(.A1(new_n802), .A2(KEYINPUT54), .A3(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT54), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n666), .B1(new_n658), .B2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(new_n806), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n800), .B1(new_n804), .B2(new_n807), .ZN(new_n808));
  OR3_X1    g607(.A1(new_n658), .A2(new_n661), .A3(new_n665), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n802), .A2(KEYINPUT54), .A3(new_n803), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n810), .A2(KEYINPUT55), .A3(new_n806), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n808), .A2(new_n643), .A3(new_n809), .A4(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(new_n622), .ZN(new_n813));
  INV_X1    g612(.A(new_n621), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n813), .B1(new_n619), .B2(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT115), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n627), .A2(new_n621), .A3(new_n629), .ZN(new_n818));
  OAI211_X1 g617(.A(KEYINPUT115), .B(new_n813), .C1(new_n619), .C2(new_n814), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n817), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  AOI22_X1  g619(.A1(new_n633), .A2(new_n639), .B1(new_n820), .B2(new_n638), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(new_n669), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT116), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n821), .A2(new_n669), .A3(KEYINPUT116), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n812), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(new_n706), .ZN(new_n827));
  AND2_X1   g626(.A1(new_n811), .A2(new_n809), .ZN(new_n828));
  AND2_X1   g627(.A1(new_n828), .A2(new_n808), .ZN(new_n829));
  OAI211_X1 g628(.A(new_n829), .B(new_n821), .C1(new_n704), .C2(new_n705), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n550), .B1(new_n827), .B2(new_n830), .ZN(new_n831));
  NOR4_X1   g630(.A1(new_n551), .A2(new_n643), .A3(new_n669), .A4(new_n617), .ZN(new_n832));
  OR2_X1    g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n833), .A2(new_n673), .A3(new_n414), .A4(new_n488), .ZN(new_n834));
  NOR3_X1   g633(.A1(new_n834), .A2(new_n282), .A3(new_n644), .ZN(new_n835));
  AND2_X1   g634(.A1(new_n497), .A2(new_n495), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n833), .A2(new_n673), .A3(new_n414), .A4(new_n836), .ZN(new_n837));
  OR2_X1    g636(.A1(new_n837), .A2(new_n644), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n835), .B1(new_n282), .B2(new_n838), .ZN(G1340gat));
  OR3_X1    g638(.A1(new_n834), .A2(new_n284), .A3(new_n748), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n284), .B1(new_n837), .B2(new_n748), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(KEYINPUT117), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT117), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n840), .A2(new_n844), .A3(new_n841), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n843), .A2(new_n845), .ZN(G1341gat));
  OAI21_X1  g645(.A(G127gat), .B1(new_n834), .B2(new_n551), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n550), .A2(new_n287), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n847), .B1(new_n837), .B2(new_n848), .ZN(G1342gat));
  OAI21_X1  g648(.A(G134gat), .B1(new_n834), .B2(new_n616), .ZN(new_n850));
  NOR3_X1   g649(.A1(new_n616), .A2(G134gat), .A3(new_n415), .ZN(new_n851));
  NAND4_X1  g650(.A1(new_n833), .A2(new_n673), .A3(new_n836), .A4(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT56), .ZN(new_n853));
  AND2_X1   g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n852), .A2(new_n853), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n850), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT118), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  OAI211_X1 g657(.A(KEYINPUT118), .B(new_n850), .C1(new_n854), .C2(new_n855), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(G1343gat));
  NOR2_X1   g659(.A1(new_n674), .A2(new_n479), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(new_n414), .ZN(new_n862));
  INV_X1    g661(.A(new_n862), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n833), .A2(new_n276), .A3(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(new_n864), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n865), .A2(new_n226), .A3(new_n643), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT57), .ZN(new_n867));
  OAI211_X1 g666(.A(new_n867), .B(new_n276), .C1(new_n831), .C2(new_n832), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n828), .A2(new_n808), .A3(new_n821), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n706), .A2(new_n869), .ZN(new_n870));
  OAI21_X1  g669(.A(KEYINPUT119), .B1(new_n804), .B2(new_n807), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT119), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n810), .A2(new_n872), .A3(new_n806), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n871), .A2(new_n800), .A3(new_n873), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n874), .A2(new_n828), .A3(new_n643), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n617), .B1(new_n875), .B2(new_n822), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n551), .B1(new_n870), .B2(new_n876), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n618), .A2(new_n644), .A3(new_n748), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n496), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  OAI211_X1 g678(.A(new_n868), .B(new_n863), .C1(new_n879), .C2(new_n867), .ZN(new_n880));
  OAI21_X1  g679(.A(G141gat), .B1(new_n880), .B2(new_n644), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n866), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(KEYINPUT58), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT58), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n866), .A2(new_n881), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n883), .A2(new_n885), .ZN(G1344gat));
  NAND3_X1  g685(.A1(new_n865), .A2(new_n223), .A3(new_n669), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT120), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND4_X1  g688(.A1(new_n865), .A2(KEYINPUT120), .A3(new_n223), .A4(new_n669), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT59), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n276), .B1(new_n831), .B2(new_n832), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(KEYINPUT57), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n869), .A2(new_n616), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n551), .B1(new_n876), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(new_n878), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n496), .A2(KEYINPUT57), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  XNOR2_X1  g698(.A(new_n862), .B(KEYINPUT121), .ZN(new_n900));
  NAND4_X1  g699(.A1(new_n894), .A2(new_n669), .A3(new_n899), .A4(new_n900), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT122), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n223), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  AOI22_X1  g702(.A1(new_n893), .A2(KEYINPUT57), .B1(new_n897), .B2(new_n898), .ZN(new_n904));
  NAND4_X1  g703(.A1(new_n904), .A2(KEYINPUT122), .A3(new_n669), .A4(new_n900), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n892), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  OAI211_X1 g705(.A(new_n892), .B(G148gat), .C1(new_n880), .C2(new_n748), .ZN(new_n907));
  INV_X1    g706(.A(new_n907), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n891), .B1(new_n906), .B2(new_n908), .ZN(G1345gat));
  NAND2_X1  g708(.A1(new_n550), .A2(G155gat), .ZN(new_n910));
  XOR2_X1   g709(.A(new_n910), .B(KEYINPUT124), .Z(new_n911));
  NOR2_X1   g710(.A1(new_n880), .A2(new_n911), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n864), .A2(new_n551), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT123), .ZN(new_n914));
  XNOR2_X1  g713(.A(new_n913), .B(new_n914), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n912), .B1(new_n915), .B2(new_n230), .ZN(G1346gat));
  OAI21_X1  g715(.A(G162gat), .B1(new_n880), .B2(new_n706), .ZN(new_n917));
  INV_X1    g716(.A(new_n893), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n616), .A2(new_n415), .ZN(new_n919));
  NAND4_X1  g718(.A1(new_n918), .A2(new_n231), .A3(new_n919), .A4(new_n861), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n917), .A2(new_n920), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT125), .ZN(new_n922));
  XNOR2_X1  g721(.A(new_n921), .B(new_n922), .ZN(G1347gat));
  NOR2_X1   g722(.A1(new_n673), .A2(new_n414), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n833), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(new_n488), .ZN(new_n926));
  OAI21_X1  g725(.A(G169gat), .B1(new_n926), .B2(new_n644), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n925), .A2(new_n836), .ZN(new_n928));
  OR2_X1    g727(.A1(new_n644), .A2(G169gat), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n927), .B1(new_n928), .B2(new_n929), .ZN(G1348gat));
  INV_X1    g729(.A(G176gat), .ZN(new_n931));
  NOR3_X1   g730(.A1(new_n926), .A2(new_n931), .A3(new_n748), .ZN(new_n932));
  INV_X1    g731(.A(new_n928), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n933), .A2(new_n669), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n932), .B1(new_n931), .B2(new_n934), .ZN(G1349gat));
  NAND4_X1  g734(.A1(new_n833), .A2(new_n550), .A3(new_n488), .A4(new_n924), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n936), .A2(G183gat), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n550), .A2(new_n388), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n937), .B1(new_n928), .B2(new_n938), .ZN(new_n939));
  XNOR2_X1  g738(.A(new_n939), .B(KEYINPUT60), .ZN(G1350gat));
  NAND4_X1  g739(.A1(new_n833), .A2(new_n617), .A3(new_n488), .A4(new_n924), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(G190gat), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n942), .A2(KEYINPUT126), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT126), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n941), .A2(new_n944), .A3(G190gat), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n943), .A2(KEYINPUT61), .A3(new_n945), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n933), .A2(new_n380), .A3(new_n707), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT61), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n942), .A2(KEYINPUT126), .A3(new_n948), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n946), .A2(new_n947), .A3(new_n949), .ZN(G1351gat));
  NAND2_X1  g749(.A1(new_n924), .A2(new_n689), .ZN(new_n951));
  INV_X1    g750(.A(new_n951), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n918), .A2(new_n952), .ZN(new_n953));
  INV_X1    g752(.A(new_n953), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n954), .A2(new_n213), .A3(new_n643), .ZN(new_n955));
  INV_X1    g754(.A(new_n904), .ZN(new_n956));
  NOR3_X1   g755(.A1(new_n956), .A2(new_n644), .A3(new_n951), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n955), .B1(new_n957), .B2(new_n213), .ZN(G1352gat));
  NAND3_X1  g757(.A1(new_n918), .A2(new_n214), .A3(new_n952), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT127), .ZN(new_n960));
  OAI22_X1  g759(.A1(new_n959), .A2(new_n748), .B1(new_n960), .B2(KEYINPUT62), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT62), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n961), .B1(KEYINPUT127), .B2(new_n962), .ZN(new_n963));
  OAI211_X1 g762(.A(new_n960), .B(KEYINPUT62), .C1(new_n959), .C2(new_n748), .ZN(new_n964));
  NOR3_X1   g763(.A1(new_n956), .A2(new_n748), .A3(new_n951), .ZN(new_n965));
  OAI211_X1 g764(.A(new_n963), .B(new_n964), .C1(new_n214), .C2(new_n965), .ZN(G1353gat));
  NAND3_X1  g765(.A1(new_n954), .A2(new_n207), .A3(new_n550), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n904), .A2(new_n550), .A3(new_n952), .ZN(new_n968));
  AND3_X1   g767(.A1(new_n968), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n969));
  AOI21_X1  g768(.A(KEYINPUT63), .B1(new_n968), .B2(G211gat), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n967), .B1(new_n969), .B2(new_n970), .ZN(G1354gat));
  NAND3_X1  g770(.A1(new_n954), .A2(new_n208), .A3(new_n707), .ZN(new_n972));
  NOR3_X1   g771(.A1(new_n956), .A2(new_n616), .A3(new_n951), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n972), .B1(new_n973), .B2(new_n208), .ZN(G1355gat));
endmodule


