//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 1 0 1 1 1 0 1 0 0 1 0 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 0 1 1 1 1 0 0 1 0 0 0 1 1 0 0 1 1 0 1 1 0 1 1 1 0 0 1 1 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:11 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n713, new_n714, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n729, new_n730, new_n731, new_n732, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n773,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n797, new_n798, new_n799, new_n800, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n928, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000;
  INV_X1    g000(.A(KEYINPUT79), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT25), .ZN(new_n188));
  INV_X1    g002(.A(G902), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT77), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT24), .B(G110), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G128), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G119), .ZN(new_n194));
  INV_X1    g008(.A(G119), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G128), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT75), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n194), .A2(new_n196), .A3(KEYINPUT75), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n192), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT23), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n202), .B1(new_n195), .B2(G128), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n193), .A2(KEYINPUT23), .A3(G119), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n203), .A2(new_n196), .A3(new_n204), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n205), .A2(G110), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n190), .B1(new_n201), .B2(new_n206), .ZN(new_n207));
  OR2_X1    g021(.A1(new_n205), .A2(G110), .ZN(new_n208));
  AND3_X1   g022(.A1(new_n194), .A2(new_n196), .A3(KEYINPUT75), .ZN(new_n209));
  AOI21_X1  g023(.A(KEYINPUT75), .B1(new_n194), .B2(new_n196), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n191), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n208), .A2(new_n211), .A3(KEYINPUT77), .ZN(new_n212));
  INV_X1    g026(.A(G140), .ZN(new_n213));
  INV_X1    g027(.A(G125), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(KEYINPUT76), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT76), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G125), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n213), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  NOR2_X1   g032(.A1(G125), .A2(G140), .ZN(new_n219));
  OAI21_X1  g033(.A(KEYINPUT16), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n215), .A2(new_n217), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT16), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n221), .A2(new_n222), .A3(new_n213), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n220), .A2(G146), .A3(new_n223), .ZN(new_n224));
  XNOR2_X1  g038(.A(G125), .B(G140), .ZN(new_n225));
  INV_X1    g039(.A(G146), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n207), .A2(new_n212), .A3(new_n224), .A4(new_n227), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n209), .A2(new_n210), .ZN(new_n229));
  AOI22_X1  g043(.A1(new_n229), .A2(new_n192), .B1(G110), .B2(new_n205), .ZN(new_n230));
  AND3_X1   g044(.A1(new_n220), .A2(G146), .A3(new_n223), .ZN(new_n231));
  AOI21_X1  g045(.A(G146), .B1(new_n220), .B2(new_n223), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n230), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n228), .A2(new_n233), .A3(KEYINPUT78), .ZN(new_n234));
  XNOR2_X1  g048(.A(KEYINPUT22), .B(G137), .ZN(new_n235));
  INV_X1    g049(.A(G221), .ZN(new_n236));
  INV_X1    g050(.A(G234), .ZN(new_n237));
  NOR3_X1   g051(.A1(new_n236), .A2(new_n237), .A3(G953), .ZN(new_n238));
  XOR2_X1   g052(.A(new_n235), .B(new_n238), .Z(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n234), .A2(new_n240), .ZN(new_n241));
  AOI21_X1  g055(.A(KEYINPUT78), .B1(new_n228), .B2(new_n233), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n228), .A2(new_n233), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT78), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n244), .A2(new_n245), .A3(new_n239), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  OAI211_X1 g061(.A(new_n188), .B(new_n189), .C1(new_n243), .C2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(G217), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n249), .B1(G234), .B2(new_n189), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n244), .A2(new_n245), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n252), .A2(new_n240), .A3(new_n234), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(new_n246), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n188), .B1(new_n254), .B2(new_n189), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n187), .B1(new_n251), .B2(new_n255), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n189), .B1(new_n243), .B2(new_n247), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(KEYINPUT25), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n258), .A2(KEYINPUT79), .A3(new_n248), .A4(new_n250), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n250), .A2(G902), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n254), .A2(new_n260), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n256), .A2(new_n259), .A3(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(G237), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(KEYINPUT71), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT71), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(G237), .ZN(new_n266));
  AOI21_X1  g080(.A(G953), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G210), .ZN(new_n268));
  XOR2_X1   g082(.A(new_n268), .B(KEYINPUT27), .Z(new_n269));
  XNOR2_X1  g083(.A(KEYINPUT26), .B(G101), .ZN(new_n270));
  XNOR2_X1  g084(.A(new_n269), .B(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  XNOR2_X1  g086(.A(KEYINPUT72), .B(KEYINPUT28), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n226), .A2(G143), .ZN(new_n274));
  INV_X1    g088(.A(G143), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(G146), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT0), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n278), .A2(new_n193), .ZN(new_n279));
  OR2_X1    g093(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  NOR2_X1   g094(.A1(KEYINPUT0), .A2(G128), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n277), .B1(new_n281), .B2(new_n279), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT11), .ZN(new_n284));
  INV_X1    g098(.A(G134), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n284), .B1(new_n285), .B2(G137), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT64), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  OAI211_X1 g102(.A(KEYINPUT64), .B(new_n284), .C1(new_n285), .C2(G137), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(G131), .ZN(new_n291));
  INV_X1    g105(.A(G137), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n292), .A2(KEYINPUT11), .A3(G134), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n285), .A2(G137), .ZN(new_n294));
  AND2_X1   g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND4_X1  g109(.A1(new_n290), .A2(KEYINPUT65), .A3(new_n291), .A4(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n293), .A2(new_n294), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n298), .B1(new_n288), .B2(new_n289), .ZN(new_n299));
  AOI21_X1  g113(.A(KEYINPUT65), .B1(new_n299), .B2(new_n291), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(KEYINPUT66), .B1(new_n299), .B2(new_n291), .ZN(new_n302));
  INV_X1    g116(.A(new_n289), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n292), .A2(G134), .ZN(new_n304));
  AOI21_X1  g118(.A(KEYINPUT64), .B1(new_n304), .B2(new_n284), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n295), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT66), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n306), .A2(new_n307), .A3(G131), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n302), .A2(new_n308), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n283), .B1(new_n301), .B2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT70), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n291), .B1(new_n304), .B2(new_n294), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n301), .A2(new_n312), .ZN(new_n313));
  AND2_X1   g127(.A1(new_n274), .A2(new_n276), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n193), .B1(new_n274), .B2(KEYINPUT1), .ZN(new_n315));
  XNOR2_X1  g129(.A(new_n314), .B(new_n315), .ZN(new_n316));
  AOI22_X1  g130(.A1(new_n310), .A2(new_n311), .B1(new_n313), .B2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT69), .ZN(new_n318));
  INV_X1    g132(.A(G116), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n319), .A2(G119), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n195), .A2(G116), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n318), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  XOR2_X1   g136(.A(KEYINPUT2), .B(G113), .Z(new_n323));
  XNOR2_X1  g137(.A(new_n322), .B(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  OAI211_X1 g139(.A(new_n295), .B(new_n291), .C1(new_n303), .C2(new_n305), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT65), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(new_n296), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n329), .A2(new_n302), .A3(new_n308), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n330), .A2(KEYINPUT70), .A3(new_n283), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n317), .A2(new_n325), .A3(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT67), .ZN(new_n334));
  INV_X1    g148(.A(new_n312), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n334), .B1(new_n329), .B2(new_n335), .ZN(new_n336));
  AOI211_X1 g150(.A(KEYINPUT67), .B(new_n312), .C1(new_n328), .C2(new_n296), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n316), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n325), .B1(new_n338), .B2(new_n310), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n273), .B1(new_n333), .B2(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n329), .A2(new_n335), .A3(new_n316), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n310), .A2(new_n325), .A3(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT28), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n272), .B1(new_n340), .B2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n310), .A2(new_n311), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n347), .A2(KEYINPUT30), .A3(new_n331), .A4(new_n341), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n338), .A2(new_n310), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT30), .ZN(new_n350));
  AOI22_X1  g164(.A1(new_n348), .A2(KEYINPUT68), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT68), .ZN(new_n352));
  AOI211_X1 g166(.A(new_n352), .B(KEYINPUT30), .C1(new_n338), .C2(new_n310), .ZN(new_n353));
  NOR3_X1   g167(.A1(new_n351), .A2(new_n325), .A3(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT31), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n332), .A2(new_n272), .ZN(new_n356));
  NOR3_X1   g170(.A1(new_n354), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n348), .A2(KEYINPUT68), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n349), .A2(new_n350), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(new_n353), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n360), .A2(new_n324), .A3(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(new_n356), .ZN(new_n363));
  AOI21_X1  g177(.A(KEYINPUT31), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n346), .B1(new_n357), .B2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(G472), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n365), .A2(new_n366), .A3(new_n189), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(KEYINPUT32), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n355), .B1(new_n354), .B2(new_n356), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n362), .A2(KEYINPUT31), .A3(new_n363), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  AOI21_X1  g185(.A(G902), .B1(new_n371), .B2(new_n346), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT32), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n372), .A2(new_n373), .A3(new_n366), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n368), .A2(new_n374), .ZN(new_n375));
  NOR3_X1   g189(.A1(new_n354), .A2(new_n272), .A3(new_n333), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT29), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n325), .B1(new_n317), .B2(new_n331), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n332), .B1(new_n379), .B2(KEYINPUT73), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT73), .ZN(new_n381));
  NAND4_X1  g195(.A1(new_n317), .A2(new_n381), .A3(new_n325), .A4(new_n331), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n343), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  XOR2_X1   g197(.A(new_n344), .B(KEYINPUT74), .Z(new_n384));
  NOR2_X1   g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n385), .A2(new_n377), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n340), .A2(new_n344), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n272), .B1(new_n387), .B2(KEYINPUT29), .ZN(new_n388));
  OAI211_X1 g202(.A(new_n189), .B(new_n378), .C1(new_n386), .C2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(G472), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n262), .B1(new_n375), .B2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT4), .ZN(new_n392));
  INV_X1    g206(.A(G104), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(KEYINPUT81), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT81), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(G104), .ZN(new_n396));
  AOI21_X1  g210(.A(G107), .B1(new_n394), .B2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT3), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(G107), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n398), .A2(new_n400), .A3(G104), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n394), .A2(new_n396), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n401), .B1(new_n402), .B2(new_n400), .ZN(new_n403));
  OAI211_X1 g217(.A(new_n392), .B(G101), .C1(new_n399), .C2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(new_n283), .ZN(new_n405));
  OAI21_X1  g219(.A(G101), .B1(new_n399), .B2(new_n403), .ZN(new_n406));
  XNOR2_X1  g220(.A(KEYINPUT81), .B(G104), .ZN(new_n407));
  OAI21_X1  g221(.A(KEYINPUT3), .B1(new_n407), .B2(G107), .ZN(new_n408));
  INV_X1    g222(.A(G101), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n407), .A2(G107), .ZN(new_n410));
  NAND4_X1  g224(.A1(new_n408), .A2(new_n409), .A3(new_n410), .A4(new_n401), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n406), .A2(new_n411), .A3(KEYINPUT4), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(KEYINPUT82), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT82), .ZN(new_n414));
  NAND4_X1  g228(.A1(new_n406), .A2(new_n411), .A3(new_n414), .A4(KEYINPUT4), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n405), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT83), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n400), .A2(G104), .ZN(new_n419));
  OAI211_X1 g233(.A(new_n418), .B(G101), .C1(new_n397), .C2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n419), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n422), .B1(new_n407), .B2(G107), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n418), .B1(new_n423), .B2(G101), .ZN(new_n424));
  OAI211_X1 g238(.A(new_n316), .B(new_n411), .C1(new_n421), .C2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT10), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  OAI21_X1  g241(.A(G101), .B1(new_n397), .B2(new_n419), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(KEYINPUT83), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(new_n420), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n430), .A2(KEYINPUT10), .A3(new_n316), .A4(new_n411), .ZN(new_n431));
  AND2_X1   g245(.A1(new_n427), .A2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(new_n330), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n417), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n427), .A2(new_n431), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n330), .B1(new_n416), .B2(new_n435), .ZN(new_n436));
  XNOR2_X1  g250(.A(G110), .B(G140), .ZN(new_n437));
  INV_X1    g251(.A(G953), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(G227), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n437), .B(new_n439), .ZN(new_n440));
  AND3_X1   g254(.A1(new_n434), .A2(new_n436), .A3(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(new_n425), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n316), .B1(new_n430), .B2(new_n411), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n330), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT12), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  OAI211_X1 g260(.A(KEYINPUT12), .B(new_n330), .C1(new_n442), .C2(new_n443), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n440), .B1(new_n448), .B2(new_n434), .ZN(new_n449));
  OAI21_X1  g263(.A(KEYINPUT84), .B1(new_n441), .B2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT84), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n434), .A2(new_n436), .A3(new_n440), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n416), .A2(new_n435), .ZN(new_n453));
  AOI22_X1  g267(.A1(new_n433), .A2(new_n453), .B1(new_n446), .B2(new_n447), .ZN(new_n454));
  OAI211_X1 g268(.A(new_n451), .B(new_n452), .C1(new_n454), .C2(new_n440), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n450), .A2(G469), .A3(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(G469), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n457), .A2(new_n189), .ZN(new_n458));
  INV_X1    g272(.A(new_n440), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n433), .B1(new_n417), .B2(new_n432), .ZN(new_n460));
  NOR3_X1   g274(.A1(new_n416), .A2(new_n435), .A3(new_n330), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n459), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n448), .A2(new_n434), .A3(new_n440), .ZN(new_n463));
  AOI21_X1  g277(.A(G902), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n458), .B1(new_n464), .B2(new_n457), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n456), .A2(new_n465), .ZN(new_n466));
  XOR2_X1   g280(.A(KEYINPUT9), .B(G234), .Z(new_n467));
  XNOR2_X1  g281(.A(new_n467), .B(KEYINPUT80), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n236), .B1(new_n468), .B2(new_n189), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  XOR2_X1   g284(.A(KEYINPUT91), .B(G475), .Z(new_n471));
  XNOR2_X1  g285(.A(G113), .B(G122), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n472), .B(new_n393), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n267), .A2(G214), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(new_n275), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n267), .A2(G143), .A3(G214), .ZN(new_n476));
  NAND2_X1  g290(.A1(KEYINPUT18), .A2(G131), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n475), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(new_n219), .ZN(new_n479));
  INV_X1    g293(.A(new_n221), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n479), .B1(new_n480), .B2(new_n213), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n227), .B1(new_n481), .B2(new_n226), .ZN(new_n482));
  AND3_X1   g296(.A1(new_n267), .A2(G143), .A3(G214), .ZN(new_n483));
  AOI21_X1  g297(.A(G143), .B1(new_n267), .B2(G214), .ZN(new_n484));
  OAI21_X1  g298(.A(G131), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT18), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n478), .B(new_n482), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n475), .A2(new_n291), .A3(new_n476), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT17), .ZN(new_n489));
  AND3_X1   g303(.A1(new_n485), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  OAI211_X1 g304(.A(KEYINPUT17), .B(G131), .C1(new_n483), .C2(new_n484), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n220), .A2(new_n223), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(new_n226), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n491), .A2(new_n493), .A3(new_n224), .ZN(new_n494));
  OAI211_X1 g308(.A(new_n473), .B(new_n487), .C1(new_n490), .C2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n485), .A2(new_n488), .A3(new_n489), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n231), .A2(new_n232), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n497), .A2(new_n498), .A3(new_n491), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n473), .B1(new_n499), .B2(new_n487), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n189), .B1(new_n496), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(KEYINPUT92), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT92), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n503), .B(new_n189), .C1(new_n496), .C2(new_n500), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n471), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT20), .ZN(new_n506));
  AND2_X1   g320(.A1(new_n485), .A2(new_n488), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n225), .A2(KEYINPUT19), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n508), .B1(new_n481), .B2(KEYINPUT19), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n224), .B1(new_n509), .B2(G146), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n487), .B1(new_n507), .B2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(new_n473), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(new_n495), .ZN(new_n514));
  NOR2_X1   g328(.A1(G475), .A2(G902), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n506), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(new_n515), .ZN(new_n517));
  AOI211_X1 g331(.A(KEYINPUT20), .B(new_n517), .C1(new_n513), .C2(new_n495), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT95), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n520), .B1(new_n193), .B2(G143), .ZN(new_n521));
  NOR3_X1   g335(.A1(new_n275), .A2(KEYINPUT95), .A3(G128), .ZN(new_n522));
  OR2_X1    g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n275), .A2(G128), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT13), .ZN(new_n525));
  OAI211_X1 g339(.A(new_n523), .B(new_n524), .C1(new_n525), .C2(new_n285), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n524), .B1(new_n521), .B2(new_n522), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n521), .A2(new_n522), .ZN(new_n528));
  OAI211_X1 g342(.A(new_n527), .B(G134), .C1(new_n528), .C2(KEYINPUT13), .ZN(new_n529));
  INV_X1    g343(.A(G122), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(KEYINPUT93), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT93), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(G122), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(G116), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT94), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n536), .B1(new_n530), .B2(G116), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n319), .A2(KEYINPUT94), .A3(G122), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n535), .A2(new_n400), .A3(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n400), .B1(new_n535), .B2(new_n539), .ZN(new_n542));
  OAI211_X1 g356(.A(new_n526), .B(new_n529), .C1(new_n541), .C2(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n468), .A2(G217), .A3(new_n438), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n539), .A2(KEYINPUT14), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT96), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n546), .A2(new_n547), .A3(new_n535), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT14), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n537), .A2(new_n549), .A3(new_n538), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT97), .ZN(new_n551));
  OR2_X1    g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n549), .B1(new_n537), .B2(new_n538), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n319), .B1(new_n531), .B2(new_n533), .ZN(new_n554));
  OAI21_X1  g368(.A(KEYINPUT96), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n550), .A2(new_n551), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n548), .A2(new_n552), .A3(new_n555), .A4(new_n556), .ZN(new_n557));
  AND2_X1   g371(.A1(new_n557), .A2(G107), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n523), .A2(G134), .A3(new_n524), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n527), .A2(new_n285), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n559), .A2(new_n540), .A3(new_n560), .ZN(new_n561));
  OAI211_X1 g375(.A(new_n543), .B(new_n545), .C1(new_n558), .C2(new_n561), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n561), .B1(new_n557), .B2(G107), .ZN(new_n563));
  INV_X1    g377(.A(new_n543), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n544), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(new_n189), .ZN(new_n567));
  INV_X1    g381(.A(G478), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n568), .A2(KEYINPUT15), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  OAI211_X1 g384(.A(new_n566), .B(new_n189), .C1(KEYINPUT15), .C2(new_n568), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AND2_X1   g386(.A1(new_n438), .A2(G952), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n573), .B1(new_n237), .B2(new_n263), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  AOI211_X1 g389(.A(new_n189), .B(new_n438), .C1(G234), .C2(G237), .ZN(new_n576));
  XNOR2_X1  g390(.A(KEYINPUT21), .B(G898), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n575), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NOR4_X1   g392(.A1(new_n505), .A2(new_n519), .A3(new_n572), .A4(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n466), .A2(new_n470), .A3(new_n579), .ZN(new_n580));
  OAI21_X1  g394(.A(G214), .B1(G237), .B2(G902), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n413), .A2(new_n415), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n404), .A2(new_n324), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n320), .A2(new_n321), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(KEYINPUT5), .ZN(new_n587));
  INV_X1    g401(.A(G113), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT5), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n588), .B1(new_n320), .B2(new_n589), .ZN(new_n590));
  AOI22_X1  g404(.A1(new_n587), .A2(new_n590), .B1(new_n323), .B2(new_n586), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n430), .A2(new_n411), .A3(new_n591), .ZN(new_n592));
  XNOR2_X1  g406(.A(G110), .B(G122), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n585), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n593), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n583), .B1(new_n413), .B2(new_n415), .ZN(new_n596));
  INV_X1    g410(.A(new_n592), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n595), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n594), .A2(KEYINPUT6), .A3(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT85), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n594), .A2(new_n598), .A3(KEYINPUT85), .A4(KEYINPUT6), .ZN(new_n602));
  OR2_X1    g416(.A1(new_n598), .A2(KEYINPUT6), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n315), .B(new_n277), .ZN(new_n604));
  AND3_X1   g418(.A1(new_n604), .A2(KEYINPUT88), .A3(new_n480), .ZN(new_n605));
  AOI21_X1  g419(.A(KEYINPUT88), .B1(new_n604), .B2(new_n480), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT86), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n609), .B1(new_n283), .B2(new_n480), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n280), .A2(KEYINPUT86), .A3(new_n282), .A4(new_n221), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n610), .A2(KEYINPUT87), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n610), .A2(new_n611), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT87), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n608), .A2(new_n612), .A3(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(G224), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n617), .A2(G953), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n616), .B(new_n618), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n601), .A2(new_n602), .A3(new_n603), .A4(new_n619), .ZN(new_n620));
  OAI21_X1  g434(.A(G210), .B1(G237), .B2(G902), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT7), .ZN(new_n622));
  OAI22_X1  g436(.A1(new_n607), .A2(new_n613), .B1(new_n622), .B2(new_n618), .ZN(new_n623));
  OR2_X1    g437(.A1(new_n618), .A2(KEYINPUT90), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n618), .A2(KEYINPUT90), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n622), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n608), .A2(new_n612), .A3(new_n615), .A4(new_n626), .ZN(new_n627));
  AND3_X1   g441(.A1(new_n594), .A2(new_n623), .A3(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n593), .B(KEYINPUT8), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n591), .B1(new_n430), .B2(new_n411), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n629), .B1(new_n597), .B2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT89), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(new_n633));
  AOI21_X1  g447(.A(G902), .B1(new_n628), .B2(new_n633), .ZN(new_n634));
  AND3_X1   g448(.A1(new_n620), .A2(new_n621), .A3(new_n634), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n621), .B1(new_n620), .B2(new_n634), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n581), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n580), .A2(new_n637), .ZN(new_n638));
  AND2_X1   g452(.A1(new_n391), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g453(.A(KEYINPUT98), .B(G101), .Z(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G3));
  AOI21_X1  g455(.A(new_n345), .B1(new_n369), .B2(new_n370), .ZN(new_n642));
  OAI21_X1  g456(.A(G472), .B1(new_n642), .B2(G902), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(new_n367), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n469), .B1(new_n456), .B2(new_n465), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  NOR3_X1   g460(.A1(new_n644), .A2(new_n262), .A3(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n578), .ZN(new_n648));
  OAI211_X1 g462(.A(new_n581), .B(new_n648), .C1(new_n635), .C2(new_n636), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n567), .A2(G478), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT33), .ZN(new_n651));
  AND3_X1   g465(.A1(new_n562), .A2(new_n565), .A3(new_n651), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n651), .B1(new_n562), .B2(new_n565), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n189), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n650), .B1(new_n654), .B2(G478), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n655), .B1(new_n505), .B2(new_n519), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n649), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n647), .A2(new_n657), .ZN(new_n658));
  XOR2_X1   g472(.A(KEYINPUT34), .B(G104), .Z(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G6));
  NOR2_X1   g474(.A1(new_n505), .A2(new_n519), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(new_n572), .ZN(new_n663));
  NOR3_X1   g477(.A1(new_n649), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n647), .A2(new_n664), .ZN(new_n665));
  XOR2_X1   g479(.A(KEYINPUT35), .B(G107), .Z(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(G9));
  NOR2_X1   g481(.A1(new_n240), .A2(KEYINPUT36), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n244), .B(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(new_n260), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n256), .A2(new_n259), .A3(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT99), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n256), .A2(new_n259), .A3(KEYINPUT99), .A4(new_n670), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n638), .A2(new_n367), .A3(new_n643), .A4(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(KEYINPUT100), .ZN(new_n677));
  XNOR2_X1  g491(.A(KEYINPUT37), .B(G110), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n677), .B(new_n678), .ZN(G12));
  AOI21_X1  g493(.A(new_n373), .B1(new_n372), .B2(new_n366), .ZN(new_n680));
  NOR4_X1   g494(.A1(new_n642), .A2(KEYINPUT32), .A3(G472), .A4(G902), .ZN(new_n681));
  OAI21_X1  g495(.A(new_n390), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(new_n675), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n683), .A2(new_n637), .ZN(new_n684));
  AND2_X1   g498(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  NOR3_X1   g499(.A1(new_n505), .A2(new_n663), .A3(new_n519), .ZN(new_n686));
  INV_X1    g500(.A(G900), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n576), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(new_n574), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n645), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n685), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G128), .ZN(G30));
  INV_X1    g509(.A(new_n636), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n620), .A2(new_n621), .A3(new_n634), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  XOR2_X1   g512(.A(KEYINPUT101), .B(KEYINPUT38), .Z(new_n699));
  XNOR2_X1  g513(.A(new_n698), .B(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(new_n581), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n662), .A2(new_n572), .ZN(new_n702));
  NOR4_X1   g516(.A1(new_n700), .A2(new_n701), .A3(new_n675), .A4(new_n702), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n272), .B1(new_n380), .B2(new_n382), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n704), .B1(new_n362), .B2(new_n363), .ZN(new_n705));
  OAI21_X1  g519(.A(G472), .B1(new_n705), .B2(G902), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n375), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n689), .B(KEYINPUT39), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n645), .A2(new_n708), .ZN(new_n709));
  XOR2_X1   g523(.A(new_n709), .B(KEYINPUT40), .Z(new_n710));
  NAND3_X1  g524(.A1(new_n703), .A2(new_n707), .A3(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G143), .ZN(G45));
  INV_X1    g526(.A(new_n656), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(new_n689), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n646), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n685), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G146), .ZN(G48));
  INV_X1    g531(.A(new_n262), .ZN(new_n718));
  OR2_X1    g532(.A1(new_n464), .A2(new_n457), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n464), .A2(new_n457), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n721), .A2(new_n469), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n682), .A2(new_n718), .A3(new_n657), .A4(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(KEYINPUT102), .ZN(new_n724));
  XOR2_X1   g538(.A(KEYINPUT41), .B(G113), .Z(new_n725));
  XNOR2_X1  g539(.A(new_n724), .B(new_n725), .ZN(G15));
  NAND4_X1  g540(.A1(new_n682), .A2(new_n718), .A3(new_n664), .A4(new_n722), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G116), .ZN(G18));
  NOR3_X1   g542(.A1(new_n721), .A2(new_n469), .A3(new_n578), .ZN(new_n729));
  AND3_X1   g543(.A1(new_n729), .A2(new_n661), .A3(new_n663), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n682), .A2(new_n684), .A3(new_n730), .ZN(new_n731));
  XOR2_X1   g545(.A(KEYINPUT103), .B(G119), .Z(new_n732));
  XNOR2_X1  g546(.A(new_n731), .B(new_n732), .ZN(G21));
  AOI21_X1  g547(.A(new_n701), .B1(new_n696), .B2(new_n697), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n734), .A2(KEYINPUT105), .A3(new_n662), .A4(new_n572), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT105), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n736), .B1(new_n637), .B2(new_n702), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n271), .B1(new_n383), .B2(new_n384), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n739), .B1(new_n357), .B2(new_n364), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n366), .A2(new_n189), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(KEYINPUT104), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  AND3_X1   g557(.A1(new_n643), .A2(new_n718), .A3(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n738), .A2(new_n729), .A3(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G122), .ZN(G24));
  NAND3_X1  g560(.A1(new_n643), .A2(new_n675), .A3(new_n743), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT106), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n643), .A2(new_n675), .A3(new_n743), .A4(KEYINPUT106), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(new_n714), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n752), .A2(new_n734), .A3(new_n722), .ZN(new_n753));
  INV_X1    g567(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n751), .A2(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT107), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n751), .A2(KEYINPUT107), .A3(new_n754), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G125), .ZN(G27));
  NAND3_X1  g574(.A1(new_n696), .A2(new_n581), .A3(new_n697), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n761), .A2(new_n469), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n441), .A2(new_n449), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n763), .A2(G469), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n465), .A2(new_n764), .ZN(new_n765));
  AND2_X1   g579(.A1(new_n762), .A2(new_n765), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n682), .A2(new_n718), .A3(new_n766), .A4(new_n752), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT42), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n391), .A2(KEYINPUT42), .A3(new_n752), .A4(new_n766), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G131), .ZN(G33));
  NAND3_X1  g586(.A1(new_n391), .A2(new_n691), .A3(new_n766), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G134), .ZN(G36));
  INV_X1    g588(.A(new_n655), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n662), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(KEYINPUT43), .ZN(new_n777));
  AND2_X1   g591(.A1(new_n777), .A2(new_n675), .ZN(new_n778));
  AOI21_X1  g592(.A(KEYINPUT44), .B1(new_n778), .B2(new_n644), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n779), .A2(new_n761), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n778), .A2(KEYINPUT44), .A3(new_n644), .ZN(new_n781));
  AND2_X1   g595(.A1(new_n450), .A2(new_n455), .ZN(new_n782));
  OR2_X1    g596(.A1(new_n782), .A2(KEYINPUT45), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n763), .A2(KEYINPUT45), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT108), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n763), .A2(KEYINPUT108), .A3(KEYINPUT45), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n457), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n458), .B1(new_n783), .B2(new_n788), .ZN(new_n789));
  OR2_X1    g603(.A1(new_n789), .A2(KEYINPUT46), .ZN(new_n790));
  AOI22_X1  g604(.A1(new_n789), .A2(KEYINPUT46), .B1(new_n457), .B2(new_n464), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n469), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n780), .A2(new_n708), .A3(new_n781), .A4(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(KEYINPUT110), .ZN(new_n794));
  XNOR2_X1  g608(.A(KEYINPUT109), .B(G137), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n794), .B(new_n795), .ZN(G39));
  NOR4_X1   g610(.A1(new_n682), .A2(new_n718), .A3(new_n714), .A4(new_n761), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n792), .A2(KEYINPUT47), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n792), .A2(KEYINPUT47), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n797), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(G140), .ZN(G42));
  NOR2_X1   g615(.A1(G952), .A2(G953), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(KEYINPUT118), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n769), .A2(new_n770), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n656), .A2(KEYINPUT112), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT112), .ZN(new_n806));
  OAI211_X1 g620(.A(new_n655), .B(new_n806), .C1(new_n505), .C2(new_n519), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n686), .B1(new_n805), .B2(new_n807), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n808), .A2(new_n649), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n645), .A2(new_n718), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n809), .A2(new_n367), .A3(new_n643), .A4(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(new_n676), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n812), .B1(new_n391), .B2(new_n638), .ZN(new_n813));
  AND3_X1   g627(.A1(new_n762), .A2(new_n752), .A3(new_n765), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n661), .A2(new_n663), .A3(new_n689), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(KEYINPUT113), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT113), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n661), .A2(new_n817), .A3(new_n663), .A4(new_n689), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n816), .A2(new_n645), .A3(new_n818), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n683), .A2(new_n819), .A3(new_n761), .ZN(new_n820));
  AOI22_X1  g634(.A1(new_n751), .A2(new_n814), .B1(new_n682), .B2(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n813), .A2(new_n821), .A3(new_n773), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n723), .A2(new_n727), .A3(new_n731), .A4(new_n745), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n804), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(new_n671), .ZN(new_n825));
  AND3_X1   g639(.A1(new_n765), .A2(new_n470), .A3(new_n689), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n707), .A2(new_n825), .A3(new_n738), .A4(new_n826), .ZN(new_n827));
  OAI211_X1 g641(.A(new_n682), .B(new_n684), .C1(new_n693), .C2(new_n715), .ZN(new_n828));
  AOI21_X1  g642(.A(KEYINPUT107), .B1(new_n751), .B2(new_n754), .ZN(new_n829));
  AOI211_X1 g643(.A(new_n756), .B(new_n753), .C1(new_n749), .C2(new_n750), .ZN(new_n830));
  OAI211_X1 g644(.A(new_n827), .B(new_n828), .C1(new_n829), .C2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT52), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n831), .A2(new_n832), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n824), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(KEYINPUT53), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n759), .A2(KEYINPUT52), .A3(new_n827), .A4(new_n828), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n831), .A2(new_n832), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT114), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n837), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  OR3_X1    g654(.A1(new_n831), .A2(new_n839), .A3(new_n832), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT53), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n840), .A2(new_n841), .A3(new_n842), .A4(new_n824), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n836), .A2(new_n843), .A3(KEYINPUT54), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n835), .A2(new_n842), .ZN(new_n845));
  AND4_X1   g659(.A1(new_n723), .A2(new_n727), .A3(new_n731), .A4(new_n745), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n846), .A2(new_n771), .A3(KEYINPUT53), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT115), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n822), .A2(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n813), .A2(new_n821), .A3(KEYINPUT115), .A4(new_n773), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n847), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n851), .A2(new_n840), .A3(new_n841), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT54), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n845), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n844), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n734), .A2(new_n722), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n777), .A2(new_n575), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n857), .A2(new_n744), .ZN(new_n858));
  INV_X1    g672(.A(new_n721), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n762), .A2(new_n718), .A3(new_n575), .A4(new_n859), .ZN(new_n860));
  OR2_X1    g674(.A1(new_n707), .A2(new_n860), .ZN(new_n861));
  OAI221_X1 g675(.A(new_n573), .B1(new_n856), .B2(new_n858), .C1(new_n861), .C2(new_n656), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n700), .A2(new_n701), .A3(new_n722), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n858), .A2(new_n863), .ZN(new_n864));
  XNOR2_X1  g678(.A(new_n864), .B(KEYINPUT50), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n751), .A2(new_n859), .A3(new_n857), .A4(new_n762), .ZN(new_n866));
  OR3_X1    g680(.A1(new_n861), .A2(new_n662), .A3(new_n655), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT51), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n798), .A2(new_n799), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n859), .A2(new_n469), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n858), .A2(new_n761), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n870), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n862), .B1(new_n869), .B2(new_n875), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n391), .A2(new_n859), .A3(new_n762), .A4(new_n857), .ZN(new_n877));
  OAI21_X1  g691(.A(KEYINPUT48), .B1(new_n877), .B2(KEYINPUT117), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(KEYINPUT117), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n878), .B(new_n879), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n872), .B(KEYINPUT116), .ZN(new_n881));
  AOI211_X1 g695(.A(new_n761), .B(new_n858), .C1(new_n871), .C2(new_n881), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n870), .B1(new_n882), .B2(new_n868), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n876), .A2(new_n880), .A3(new_n883), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n803), .B1(new_n855), .B2(new_n884), .ZN(new_n885));
  AND4_X1   g699(.A1(new_n718), .A2(new_n776), .A3(new_n581), .A4(new_n470), .ZN(new_n886));
  AND2_X1   g700(.A1(new_n886), .A2(KEYINPUT111), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n886), .A2(KEYINPUT111), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n721), .B(KEYINPUT49), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n887), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n890), .A2(new_n700), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n885), .B1(new_n707), .B2(new_n891), .ZN(G75));
  NAND3_X1  g706(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n893), .B(new_n619), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n894), .B(KEYINPUT55), .ZN(new_n895));
  AND3_X1   g709(.A1(new_n851), .A2(new_n841), .A3(new_n840), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n837), .A2(new_n838), .ZN(new_n897));
  AOI21_X1  g711(.A(KEYINPUT53), .B1(new_n897), .B2(new_n824), .ZN(new_n898));
  OAI211_X1 g712(.A(G210), .B(G902), .C1(new_n896), .C2(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT119), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n189), .B1(new_n845), .B2(new_n852), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n902), .A2(KEYINPUT119), .A3(G210), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT56), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n895), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n438), .A2(G952), .ZN(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n895), .A2(new_n905), .ZN(new_n909));
  AOI211_X1 g723(.A(KEYINPUT120), .B(new_n909), .C1(new_n902), .C2(G210), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT120), .ZN(new_n911));
  INV_X1    g725(.A(new_n909), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n911), .B1(new_n899), .B2(new_n912), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n908), .B1(new_n910), .B2(new_n913), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n906), .A2(new_n914), .ZN(G51));
  NAND2_X1  g729(.A1(new_n462), .A2(new_n463), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n845), .A2(new_n852), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(KEYINPUT54), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n918), .A2(new_n854), .ZN(new_n919));
  INV_X1    g733(.A(new_n919), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n458), .B(KEYINPUT57), .Z(new_n921));
  OAI21_X1  g735(.A(new_n916), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n902), .A2(new_n783), .A3(new_n788), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n907), .B1(new_n922), .B2(new_n923), .ZN(G54));
  NAND3_X1  g738(.A1(new_n902), .A2(KEYINPUT58), .A3(G475), .ZN(new_n925));
  INV_X1    g739(.A(new_n514), .ZN(new_n926));
  AND2_X1   g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n925), .A2(new_n926), .ZN(new_n928));
  NOR3_X1   g742(.A1(new_n927), .A2(new_n928), .A3(new_n907), .ZN(G60));
  NAND2_X1  g743(.A1(G478), .A2(G902), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n930), .B(KEYINPUT59), .Z(new_n931));
  AOI21_X1  g745(.A(new_n931), .B1(new_n844), .B2(new_n854), .ZN(new_n932));
  INV_X1    g746(.A(new_n932), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n652), .A2(new_n653), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n933), .A2(KEYINPUT121), .A3(new_n934), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n934), .A2(new_n931), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n907), .B1(new_n919), .B2(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT121), .ZN(new_n938));
  INV_X1    g752(.A(new_n934), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n938), .B1(new_n932), .B2(new_n939), .ZN(new_n940));
  AND3_X1   g754(.A1(new_n935), .A2(new_n937), .A3(new_n940), .ZN(G63));
  XNOR2_X1  g755(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n249), .A2(new_n189), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n942), .B(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n917), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n945), .A2(new_n246), .A3(new_n253), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n917), .A2(new_n669), .A3(new_n944), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n946), .A2(new_n908), .A3(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT61), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n946), .A2(KEYINPUT61), .A3(new_n908), .A4(new_n947), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n951), .ZN(G66));
  NOR3_X1   g766(.A1(new_n577), .A2(new_n617), .A3(new_n438), .ZN(new_n953));
  NOR3_X1   g767(.A1(new_n823), .A2(new_n639), .A3(new_n812), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n953), .B1(new_n954), .B2(new_n438), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n893), .B1(G898), .B2(new_n438), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n956), .B(KEYINPUT123), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n955), .B(new_n957), .ZN(G69));
  AOI21_X1  g772(.A(new_n438), .B1(G227), .B2(G900), .ZN(new_n959));
  NAND4_X1  g773(.A1(new_n792), .A2(new_n391), .A3(new_n708), .A4(new_n738), .ZN(new_n960));
  AND2_X1   g774(.A1(new_n960), .A2(new_n773), .ZN(new_n961));
  AND4_X1   g775(.A1(new_n771), .A2(new_n793), .A3(new_n800), .A4(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n759), .A2(new_n828), .ZN(new_n963));
  INV_X1    g777(.A(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(G953), .B1(new_n962), .B2(new_n964), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n438), .A2(G900), .ZN(new_n966));
  NOR3_X1   g780(.A1(new_n965), .A2(KEYINPUT125), .A3(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n351), .A2(new_n353), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n969), .B(KEYINPUT124), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n970), .B(new_n509), .Z(new_n971));
  INV_X1    g785(.A(new_n971), .ZN(new_n972));
  OAI21_X1  g786(.A(KEYINPUT125), .B1(new_n965), .B2(new_n966), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n968), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  NOR3_X1   g788(.A1(new_n709), .A2(new_n808), .A3(new_n761), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n391), .A2(new_n975), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n800), .A2(new_n793), .A3(new_n976), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n964), .A2(KEYINPUT62), .A3(new_n711), .ZN(new_n978));
  INV_X1    g792(.A(KEYINPUT62), .ZN(new_n979));
  INV_X1    g793(.A(new_n711), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n979), .B1(new_n963), .B2(new_n980), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n977), .B1(new_n978), .B2(new_n981), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n971), .B1(new_n982), .B2(G953), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n959), .B1(new_n974), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n973), .A2(new_n972), .ZN(new_n985));
  OAI211_X1 g799(.A(new_n983), .B(new_n959), .C1(new_n985), .C2(new_n967), .ZN(new_n986));
  INV_X1    g800(.A(new_n986), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n984), .A2(new_n987), .ZN(G72));
  AOI21_X1  g802(.A(new_n271), .B1(new_n362), .B2(new_n332), .ZN(new_n989));
  AND2_X1   g803(.A1(new_n982), .A2(new_n989), .ZN(new_n990));
  AND3_X1   g804(.A1(new_n962), .A2(new_n376), .A3(new_n964), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n954), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  OR2_X1    g806(.A1(new_n376), .A2(new_n989), .ZN(new_n993));
  XNOR2_X1  g807(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n366), .A2(new_n189), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n994), .B(new_n995), .ZN(new_n996));
  NOR2_X1   g810(.A1(new_n993), .A2(new_n996), .ZN(new_n997));
  XOR2_X1   g811(.A(new_n997), .B(KEYINPUT127), .Z(new_n998));
  NAND3_X1  g812(.A1(new_n836), .A2(new_n843), .A3(new_n998), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n907), .B1(new_n993), .B2(new_n996), .ZN(new_n1000));
  AND3_X1   g814(.A1(new_n992), .A2(new_n999), .A3(new_n1000), .ZN(G57));
endmodule


