//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 1 1 0 0 0 1 1 0 1 1 0 0 0 1 1 0 1 1 1 0 0 1 1 1 1 1 1 0 0 1 0 1 1 1 0 0 0 0 1 0 0 0 1 1 0 1 0 0 1 1 1 0 1 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:49 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n734, new_n735, new_n736, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n766, new_n767, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n783, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n975, new_n976, new_n977, new_n978,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT86), .ZN(new_n188));
  INV_X1    g002(.A(G104), .ZN(new_n189));
  OR3_X1    g003(.A1(new_n189), .A2(KEYINPUT80), .A3(G107), .ZN(new_n190));
  OAI21_X1  g004(.A(KEYINPUT80), .B1(new_n189), .B2(G107), .ZN(new_n191));
  INV_X1    g005(.A(G107), .ZN(new_n192));
  OAI211_X1 g006(.A(new_n190), .B(new_n191), .C1(G104), .C2(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G101), .ZN(new_n194));
  XNOR2_X1  g008(.A(G116), .B(G119), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(KEYINPUT5), .ZN(new_n196));
  INV_X1    g010(.A(G116), .ZN(new_n197));
  NOR3_X1   g011(.A1(new_n197), .A2(KEYINPUT5), .A3(G119), .ZN(new_n198));
  INV_X1    g012(.A(G113), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  XNOR2_X1  g014(.A(KEYINPUT2), .B(G113), .ZN(new_n201));
  INV_X1    g015(.A(new_n201), .ZN(new_n202));
  AOI22_X1  g016(.A1(new_n196), .A2(new_n200), .B1(new_n202), .B2(new_n195), .ZN(new_n203));
  INV_X1    g017(.A(G101), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT77), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT3), .ZN(new_n206));
  AOI22_X1  g020(.A1(new_n205), .A2(new_n206), .B1(new_n189), .B2(G107), .ZN(new_n207));
  NAND2_X1  g021(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n208));
  NOR3_X1   g022(.A1(new_n208), .A2(new_n189), .A3(G107), .ZN(new_n209));
  AOI22_X1  g023(.A1(new_n192), .A2(G104), .B1(KEYINPUT77), .B2(KEYINPUT3), .ZN(new_n210));
  OAI211_X1 g024(.A(new_n204), .B(new_n207), .C1(new_n209), .C2(new_n210), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n211), .A2(KEYINPUT78), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT78), .ZN(new_n213));
  OAI22_X1  g027(.A1(new_n192), .A2(G104), .B1(KEYINPUT77), .B2(KEYINPUT3), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n208), .B1(new_n189), .B2(G107), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n192), .A2(KEYINPUT77), .A3(KEYINPUT3), .A4(G104), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n213), .B1(new_n217), .B2(new_n204), .ZN(new_n218));
  OAI211_X1 g032(.A(new_n194), .B(new_n203), .C1(new_n212), .C2(new_n218), .ZN(new_n219));
  XNOR2_X1  g033(.A(G110), .B(G122), .ZN(new_n220));
  OAI21_X1  g034(.A(KEYINPUT4), .B1(new_n217), .B2(new_n204), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n217), .A2(new_n213), .A3(new_n204), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n211), .A2(KEYINPUT78), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n221), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  XOR2_X1   g038(.A(new_n195), .B(new_n201), .Z(new_n225));
  OAI21_X1  g039(.A(new_n207), .B1(new_n209), .B2(new_n210), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT4), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n226), .A2(new_n227), .A3(G101), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n225), .A2(new_n228), .ZN(new_n229));
  OAI211_X1 g043(.A(new_n219), .B(new_n220), .C1(new_n224), .C2(new_n229), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n227), .B1(new_n226), .B2(G101), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n231), .B1(new_n212), .B2(new_n218), .ZN(new_n232));
  NOR3_X1   g046(.A1(new_n217), .A2(KEYINPUT4), .A3(new_n204), .ZN(new_n233));
  XNOR2_X1  g047(.A(new_n195), .B(new_n201), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  AOI22_X1  g049(.A1(new_n223), .A2(new_n222), .B1(G101), .B2(new_n193), .ZN(new_n236));
  AOI22_X1  g050(.A1(new_n232), .A2(new_n235), .B1(new_n236), .B2(new_n203), .ZN(new_n237));
  XNOR2_X1  g051(.A(new_n220), .B(KEYINPUT83), .ZN(new_n238));
  OAI211_X1 g052(.A(new_n230), .B(KEYINPUT6), .C1(new_n237), .C2(new_n238), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n219), .B1(new_n224), .B2(new_n229), .ZN(new_n240));
  INV_X1    g054(.A(new_n238), .ZN(new_n241));
  XNOR2_X1  g055(.A(KEYINPUT84), .B(KEYINPUT6), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n240), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  XNOR2_X1  g057(.A(KEYINPUT0), .B(G128), .ZN(new_n244));
  INV_X1    g058(.A(G146), .ZN(new_n245));
  OAI21_X1  g059(.A(KEYINPUT64), .B1(new_n245), .B2(G143), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(G143), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n245), .A2(KEYINPUT64), .A3(G143), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n244), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(G143), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G146), .ZN(new_n252));
  AND2_X1   g066(.A1(KEYINPUT0), .A2(G128), .ZN(new_n253));
  AND3_X1   g067(.A1(new_n247), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  OAI21_X1  g068(.A(G125), .B1(new_n250), .B2(new_n254), .ZN(new_n255));
  AND2_X1   g069(.A1(new_n247), .A2(new_n252), .ZN(new_n256));
  INV_X1    g070(.A(G128), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n257), .A2(KEYINPUT1), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(G125), .ZN(new_n260));
  AND3_X1   g074(.A1(new_n245), .A2(KEYINPUT64), .A3(G143), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n261), .B1(new_n247), .B2(new_n246), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n257), .B1(new_n247), .B2(KEYINPUT1), .ZN(new_n263));
  OAI211_X1 g077(.A(new_n259), .B(new_n260), .C1(new_n262), .C2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n255), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(G224), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n266), .A2(G953), .ZN(new_n267));
  XNOR2_X1  g081(.A(new_n265), .B(new_n267), .ZN(new_n268));
  AND3_X1   g082(.A1(new_n239), .A2(new_n243), .A3(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(G902), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT7), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n267), .A2(new_n271), .ZN(new_n272));
  AND3_X1   g086(.A1(new_n255), .A2(new_n264), .A3(new_n272), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n272), .B1(new_n255), .B2(new_n264), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n230), .A2(new_n275), .ZN(new_n276));
  XNOR2_X1  g090(.A(KEYINPUT85), .B(KEYINPUT8), .ZN(new_n277));
  XNOR2_X1  g091(.A(new_n220), .B(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n223), .A2(new_n222), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(new_n194), .ZN(new_n281));
  INV_X1    g095(.A(new_n203), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n279), .B1(new_n283), .B2(new_n219), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n270), .B1(new_n276), .B2(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n188), .B1(new_n269), .B2(new_n285), .ZN(new_n286));
  OAI21_X1  g100(.A(G210), .B1(G237), .B2(G902), .ZN(new_n287));
  INV_X1    g101(.A(new_n287), .ZN(new_n288));
  AND2_X1   g102(.A1(new_n230), .A2(new_n275), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n283), .A2(new_n219), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(new_n278), .ZN(new_n291));
  AOI21_X1  g105(.A(G902), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n239), .A2(new_n243), .A3(new_n268), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n292), .A2(new_n293), .A3(KEYINPUT86), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n286), .A2(new_n288), .A3(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n292), .A2(new_n293), .A3(new_n287), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n251), .A2(G128), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n257), .A2(G143), .ZN(new_n299));
  AND2_X1   g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(G134), .ZN(new_n301));
  XNOR2_X1  g115(.A(new_n300), .B(new_n301), .ZN(new_n302));
  OR2_X1    g116(.A1(KEYINPUT88), .A2(G122), .ZN(new_n303));
  NAND2_X1  g117(.A1(KEYINPUT88), .A2(G122), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n197), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n197), .A2(G122), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  NOR3_X1   g121(.A1(new_n305), .A2(G107), .A3(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  XNOR2_X1  g123(.A(new_n306), .B(KEYINPUT14), .ZN(new_n310));
  OAI21_X1  g124(.A(G107), .B1(new_n310), .B2(new_n305), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n302), .A2(new_n309), .A3(new_n311), .ZN(new_n312));
  XNOR2_X1  g126(.A(KEYINPUT9), .B(G234), .ZN(new_n313));
  INV_X1    g127(.A(G217), .ZN(new_n314));
  NOR3_X1   g128(.A1(new_n313), .A2(new_n314), .A3(G953), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT92), .ZN(new_n316));
  XNOR2_X1  g130(.A(KEYINPUT89), .B(KEYINPUT13), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n316), .B1(new_n317), .B2(new_n298), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT13), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(KEYINPUT89), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT89), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(KEYINPUT13), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(new_n298), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n323), .A2(KEYINPUT92), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n318), .A2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT90), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n327), .B1(new_n323), .B2(new_n324), .ZN(new_n328));
  NAND4_X1  g142(.A1(new_n298), .A2(new_n320), .A3(new_n322), .A4(KEYINPUT90), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n328), .A2(new_n299), .A3(new_n329), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n326), .B1(new_n330), .B2(KEYINPUT91), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT91), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n328), .A2(new_n332), .A3(new_n299), .A4(new_n329), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n301), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n300), .A2(new_n301), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n303), .A2(new_n304), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(G116), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n192), .B1(new_n337), .B2(new_n306), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n335), .B1(new_n338), .B2(new_n308), .ZN(new_n339));
  OAI211_X1 g153(.A(new_n312), .B(new_n315), .C1(new_n334), .C2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(new_n315), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n329), .A2(new_n299), .ZN(new_n342));
  AOI21_X1  g156(.A(KEYINPUT90), .B1(new_n317), .B2(new_n298), .ZN(new_n343));
  OAI21_X1  g157(.A(KEYINPUT91), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NOR3_X1   g158(.A1(new_n317), .A2(new_n316), .A3(new_n298), .ZN(new_n345));
  AOI21_X1  g159(.A(KEYINPUT92), .B1(new_n323), .B2(new_n324), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n344), .A2(new_n333), .A3(new_n347), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n339), .B1(new_n348), .B2(G134), .ZN(new_n349));
  INV_X1    g163(.A(new_n312), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n341), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n340), .A2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(G478), .ZN(new_n353));
  OAI21_X1  g167(.A(KEYINPUT93), .B1(new_n353), .B2(KEYINPUT15), .ZN(new_n354));
  OR3_X1    g168(.A1(new_n353), .A2(KEYINPUT93), .A3(KEYINPUT15), .ZN(new_n355));
  NAND4_X1  g169(.A1(new_n352), .A2(new_n270), .A3(new_n354), .A4(new_n355), .ZN(new_n356));
  AOI21_X1  g170(.A(G902), .B1(new_n340), .B2(new_n351), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n356), .B1(new_n357), .B2(new_n354), .ZN(new_n358));
  INV_X1    g172(.A(G952), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n359), .A2(G953), .ZN(new_n360));
  INV_X1    g174(.A(G234), .ZN(new_n361));
  INV_X1    g175(.A(G237), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n360), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  AND2_X1   g178(.A1(KEYINPUT67), .A2(G953), .ZN(new_n365));
  NOR2_X1   g179(.A1(KEYINPUT67), .A2(G953), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  AOI211_X1 g181(.A(new_n270), .B(new_n367), .C1(G234), .C2(G237), .ZN(new_n368));
  XNOR2_X1  g182(.A(KEYINPUT21), .B(G898), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n364), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  OR2_X1    g185(.A1(KEYINPUT67), .A2(G953), .ZN(new_n372));
  NAND2_X1  g186(.A1(KEYINPUT67), .A2(G953), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n372), .A2(G214), .A3(new_n362), .A4(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(new_n251), .ZN(new_n375));
  NAND4_X1  g189(.A1(new_n367), .A2(G143), .A3(G214), .A4(new_n362), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(KEYINPUT18), .A2(G131), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(G140), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(G125), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n260), .A2(G140), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(KEYINPUT74), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT74), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n382), .A2(new_n383), .A3(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n385), .A2(new_n245), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n384), .A2(G146), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n375), .A2(new_n376), .A3(new_n378), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n380), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(G131), .ZN(new_n393));
  AND3_X1   g207(.A1(new_n375), .A2(new_n376), .A3(new_n393), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n393), .B1(new_n375), .B2(new_n376), .ZN(new_n395));
  NOR3_X1   g209(.A1(new_n394), .A2(new_n395), .A3(KEYINPUT17), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n377), .A2(KEYINPUT17), .A3(G131), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n382), .A2(new_n383), .A3(KEYINPUT16), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT16), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n399), .A2(new_n381), .A3(G125), .ZN(new_n400));
  AND3_X1   g214(.A1(new_n398), .A2(G146), .A3(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(G146), .B1(new_n398), .B2(new_n400), .ZN(new_n402));
  OAI21_X1  g216(.A(KEYINPUT87), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n398), .A2(new_n400), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(new_n245), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT87), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n398), .A2(new_n400), .A3(G146), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n405), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n397), .A2(new_n403), .A3(new_n408), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n392), .B1(new_n396), .B2(new_n409), .ZN(new_n410));
  XNOR2_X1  g224(.A(G113), .B(G122), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n411), .B(new_n189), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n410), .A2(new_n413), .ZN(new_n414));
  OAI211_X1 g228(.A(new_n412), .B(new_n392), .C1(new_n396), .C2(new_n409), .ZN(new_n415));
  AOI21_X1  g229(.A(G902), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(G475), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT20), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT19), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n385), .A2(new_n419), .A3(new_n387), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n384), .A2(KEYINPUT19), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n420), .A2(new_n245), .A3(new_n421), .ZN(new_n422));
  OAI211_X1 g236(.A(new_n422), .B(new_n407), .C1(new_n394), .C2(new_n395), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(new_n392), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(new_n413), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(new_n415), .ZN(new_n426));
  NOR2_X1   g240(.A1(G475), .A2(G902), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n418), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n427), .ZN(new_n429));
  AOI211_X1 g243(.A(KEYINPUT20), .B(new_n429), .C1(new_n425), .C2(new_n415), .ZN(new_n430));
  OAI221_X1 g244(.A(new_n371), .B1(new_n416), .B2(new_n417), .C1(new_n428), .C2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  AND4_X1   g246(.A1(new_n187), .A2(new_n297), .A3(new_n358), .A4(new_n432), .ZN(new_n433));
  OAI21_X1  g247(.A(G221), .B1(new_n313), .B2(G902), .ZN(new_n434));
  XNOR2_X1  g248(.A(new_n434), .B(KEYINPUT76), .ZN(new_n435));
  INV_X1    g249(.A(G469), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n367), .A2(G227), .ZN(new_n437));
  XOR2_X1   g251(.A(G110), .B(G140), .Z(new_n438));
  XNOR2_X1  g252(.A(new_n437), .B(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n259), .B1(new_n256), .B2(new_n263), .ZN(new_n441));
  OAI211_X1 g255(.A(new_n194), .B(new_n441), .C1(new_n212), .C2(new_n218), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT10), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT64), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n444), .B1(new_n251), .B2(G146), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n251), .A2(G146), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n249), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(new_n263), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n443), .B1(new_n449), .B2(new_n259), .ZN(new_n450));
  AOI22_X1  g264(.A1(new_n442), .A2(new_n443), .B1(new_n236), .B2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT79), .ZN(new_n452));
  INV_X1    g266(.A(new_n244), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n254), .B1(new_n447), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n228), .A2(new_n454), .ZN(new_n455));
  NOR3_X1   g269(.A1(new_n224), .A2(new_n452), .A3(new_n455), .ZN(new_n456));
  AND2_X1   g270(.A1(new_n228), .A2(new_n454), .ZN(new_n457));
  AOI21_X1  g271(.A(KEYINPUT79), .B1(new_n232), .B2(new_n457), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n451), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  OAI21_X1  g273(.A(KEYINPUT11), .B1(new_n301), .B2(G137), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT11), .ZN(new_n461));
  INV_X1    g275(.A(G137), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n461), .A2(new_n462), .A3(G134), .ZN(new_n463));
  AND2_X1   g277(.A1(new_n460), .A2(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(KEYINPUT65), .B1(new_n462), .B2(G134), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT65), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n466), .A2(new_n301), .A3(G137), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  OAI21_X1  g282(.A(G131), .B1(new_n464), .B2(new_n468), .ZN(new_n469));
  AND2_X1   g283(.A1(new_n465), .A2(new_n467), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n460), .A2(new_n463), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n470), .A2(new_n393), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n459), .A2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n473), .ZN(new_n475));
  OAI211_X1 g289(.A(new_n451), .B(new_n475), .C1(new_n456), .C2(new_n458), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n440), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n475), .A2(KEYINPUT81), .ZN(new_n478));
  AND3_X1   g292(.A1(new_n280), .A2(new_n194), .A3(new_n441), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n449), .A2(new_n259), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n480), .B1(new_n280), .B2(new_n194), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n478), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(KEYINPUT12), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT12), .ZN(new_n484));
  OAI211_X1 g298(.A(new_n484), .B(new_n478), .C1(new_n479), .C2(new_n481), .ZN(new_n485));
  AND4_X1   g299(.A1(new_n476), .A2(new_n483), .A3(new_n485), .A4(new_n440), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n436), .B(new_n270), .C1(new_n477), .C2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(KEYINPUT82), .ZN(new_n488));
  INV_X1    g302(.A(new_n476), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n452), .B1(new_n224), .B2(new_n455), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n232), .A2(new_n457), .A3(KEYINPUT79), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n475), .B1(new_n492), .B2(new_n451), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n439), .B1(new_n489), .B2(new_n493), .ZN(new_n494));
  NAND4_X1  g308(.A1(new_n476), .A2(new_n483), .A3(new_n485), .A4(new_n440), .ZN(new_n495));
  AOI21_X1  g309(.A(G902), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT82), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n496), .A2(new_n497), .A3(new_n436), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n488), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n474), .A2(new_n476), .A3(new_n440), .ZN(new_n500));
  AND3_X1   g314(.A1(new_n476), .A2(new_n483), .A3(new_n485), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n500), .B1(new_n501), .B2(new_n440), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(new_n270), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(G469), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n435), .B1(new_n499), .B2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT70), .ZN(new_n506));
  NOR3_X1   g320(.A1(new_n464), .A2(G131), .A3(new_n468), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n393), .B1(new_n470), .B2(new_n471), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n454), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n301), .A2(G137), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n462), .A2(G134), .ZN(new_n511));
  OAI21_X1  g325(.A(G131), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n263), .B1(new_n249), .B2(new_n248), .ZN(new_n513));
  AND3_X1   g327(.A1(new_n258), .A2(new_n247), .A3(new_n252), .ZN(new_n514));
  OAI211_X1 g328(.A(new_n472), .B(new_n512), .C1(new_n513), .C2(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n509), .A2(new_n515), .A3(new_n234), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT66), .ZN(new_n518));
  OAI211_X1 g332(.A(new_n454), .B(new_n518), .C1(new_n507), .C2(new_n508), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n518), .B1(new_n473), .B2(new_n454), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n515), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT30), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n509), .A2(KEYINPUT30), .A3(new_n515), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(new_n225), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n517), .B1(new_n524), .B2(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n367), .A2(G210), .A3(new_n362), .ZN(new_n529));
  XNOR2_X1  g343(.A(new_n529), .B(KEYINPUT27), .ZN(new_n530));
  XNOR2_X1  g344(.A(KEYINPUT26), .B(G101), .ZN(new_n531));
  XNOR2_X1  g345(.A(new_n530), .B(new_n531), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n506), .B1(new_n528), .B2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT29), .ZN(new_n534));
  INV_X1    g348(.A(new_n531), .ZN(new_n535));
  XNOR2_X1  g349(.A(new_n530), .B(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n526), .B1(new_n522), .B2(new_n523), .ZN(new_n537));
  OAI211_X1 g351(.A(KEYINPUT70), .B(new_n536), .C1(new_n537), .C2(new_n517), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT28), .ZN(new_n539));
  AND3_X1   g353(.A1(new_n516), .A2(KEYINPUT69), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(KEYINPUT69), .B1(new_n516), .B2(new_n539), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n517), .B1(new_n522), .B2(new_n225), .ZN(new_n543));
  OAI211_X1 g357(.A(new_n542), .B(new_n532), .C1(new_n543), .C2(new_n539), .ZN(new_n544));
  NAND4_X1  g358(.A1(new_n533), .A2(new_n534), .A3(new_n538), .A4(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n234), .B1(new_n509), .B2(new_n515), .ZN(new_n546));
  OAI21_X1  g360(.A(KEYINPUT28), .B1(new_n517), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n542), .A2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n536), .A2(new_n534), .ZN(new_n550));
  AOI21_X1  g364(.A(G902), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n545), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(G472), .ZN(new_n553));
  NOR2_X1   g367(.A1(G472), .A2(G902), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n542), .B1(new_n543), .B2(new_n539), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n532), .A2(new_n516), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n537), .A2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT31), .ZN(new_n559));
  AOI22_X1  g373(.A1(new_n556), .A2(new_n536), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  OAI21_X1  g374(.A(KEYINPUT68), .B1(new_n537), .B2(new_n557), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT68), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n536), .A2(new_n517), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n509), .A2(KEYINPUT66), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(new_n519), .ZN(new_n565));
  AOI21_X1  g379(.A(KEYINPUT30), .B1(new_n565), .B2(new_n515), .ZN(new_n566));
  OAI211_X1 g380(.A(new_n562), .B(new_n563), .C1(new_n566), .C2(new_n526), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n561), .A2(KEYINPUT31), .A3(new_n567), .ZN(new_n568));
  AOI211_X1 g382(.A(KEYINPUT32), .B(new_n555), .C1(new_n560), .C2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT32), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n556), .A2(new_n536), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n558), .A2(new_n559), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n568), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n570), .B1(new_n573), .B2(new_n554), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n553), .B1(new_n569), .B2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(G119), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(G128), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n257), .A2(G119), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT71), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT24), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n582), .A2(G110), .ZN(new_n583));
  INV_X1    g397(.A(G110), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n584), .A2(KEYINPUT24), .ZN(new_n585));
  OAI21_X1  g399(.A(KEYINPUT72), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n577), .A2(new_n578), .A3(KEYINPUT71), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n584), .A2(KEYINPUT24), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n582), .A2(G110), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT72), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n581), .A2(new_n586), .A3(new_n587), .A4(new_n591), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n592), .B1(new_n402), .B2(new_n401), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT23), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n594), .B1(new_n576), .B2(G128), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n257), .A2(KEYINPUT23), .A3(G119), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n595), .A2(new_n596), .A3(new_n577), .ZN(new_n597));
  AND3_X1   g411(.A1(new_n597), .A2(KEYINPUT73), .A3(G110), .ZN(new_n598));
  AOI21_X1  g412(.A(KEYINPUT73), .B1(new_n597), .B2(G110), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n597), .A2(G110), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n581), .A2(new_n587), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n586), .A2(new_n591), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n601), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n388), .A2(new_n407), .ZN(new_n605));
  OAI22_X1  g419(.A1(new_n593), .A2(new_n600), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n367), .A2(G221), .A3(G234), .ZN(new_n607));
  XNOR2_X1  g421(.A(KEYINPUT22), .B(G137), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n607), .B(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n606), .A2(new_n610), .ZN(new_n611));
  OAI221_X1 g425(.A(new_n592), .B1(new_n401), .B2(new_n402), .C1(new_n598), .C2(new_n599), .ZN(new_n612));
  AOI22_X1  g426(.A1(new_n581), .A2(new_n587), .B1(new_n586), .B2(new_n591), .ZN(new_n613));
  OAI211_X1 g427(.A(new_n407), .B(new_n388), .C1(new_n613), .C2(new_n601), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n612), .A2(new_n614), .A3(new_n609), .ZN(new_n615));
  OAI21_X1  g429(.A(G217), .B1(new_n361), .B2(G902), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(new_n270), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n611), .A2(new_n615), .A3(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  OR2_X1    g434(.A1(new_n620), .A2(KEYINPUT75), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n611), .A2(new_n270), .A3(new_n615), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n616), .B1(new_n622), .B2(KEYINPUT25), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT25), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n611), .A2(new_n624), .A3(new_n615), .A4(new_n270), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n620), .A2(KEYINPUT75), .ZN(new_n627));
  AND3_X1   g441(.A1(new_n621), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n433), .A2(new_n505), .A3(new_n575), .A4(new_n628), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(G101), .ZN(G3));
  INV_X1    g444(.A(G472), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n631), .B1(new_n573), .B2(new_n270), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n555), .B1(new_n560), .B2(new_n568), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n505), .A2(new_n628), .A3(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  AND3_X1   g450(.A1(new_n292), .A2(new_n293), .A3(new_n287), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n287), .B1(new_n292), .B2(new_n293), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n187), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  OAI22_X1  g453(.A1(new_n428), .A2(new_n430), .B1(new_n417), .B2(new_n416), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT94), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n351), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n352), .A2(new_n642), .A3(KEYINPUT33), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT33), .ZN(new_n644));
  OAI211_X1 g458(.A(new_n340), .B(new_n351), .C1(new_n641), .C2(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n643), .A2(G478), .A3(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n353), .A2(new_n270), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n647), .B1(new_n357), .B2(new_n353), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n640), .A2(new_n646), .A3(new_n648), .ZN(new_n649));
  NOR3_X1   g463(.A1(new_n639), .A2(new_n649), .A3(new_n370), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n636), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(KEYINPUT95), .ZN(new_n652));
  XOR2_X1   g466(.A(KEYINPUT34), .B(G104), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G6));
  INV_X1    g468(.A(KEYINPUT96), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n655), .B1(new_n431), .B2(new_n358), .ZN(new_n656));
  INV_X1    g470(.A(new_n187), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n288), .B1(new_n269), .B2(new_n285), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n657), .B1(new_n658), .B2(new_n296), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n412), .B1(new_n423), .B2(new_n392), .ZN(new_n660));
  AND3_X1   g474(.A1(new_n380), .A2(new_n390), .A3(new_n391), .ZN(new_n661));
  AND3_X1   g475(.A1(new_n397), .A2(new_n403), .A3(new_n408), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n377), .A2(G131), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT17), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n375), .A2(new_n376), .A3(new_n393), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n663), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n661), .B1(new_n662), .B2(new_n666), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n660), .B1(new_n667), .B2(new_n412), .ZN(new_n668));
  OAI21_X1  g482(.A(KEYINPUT20), .B1(new_n668), .B2(new_n429), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n426), .A2(new_n418), .A3(new_n427), .ZN(new_n670));
  INV_X1    g484(.A(new_n415), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n666), .A2(new_n397), .A3(new_n403), .A4(new_n408), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n412), .B1(new_n672), .B2(new_n392), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n270), .B1(new_n671), .B2(new_n673), .ZN(new_n674));
  AOI22_X1  g488(.A1(new_n669), .A2(new_n670), .B1(G475), .B2(new_n674), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n354), .B1(new_n352), .B2(new_n270), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n355), .A2(new_n354), .ZN(new_n677));
  AOI211_X1 g491(.A(G902), .B(new_n677), .C1(new_n340), .C2(new_n351), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n675), .A2(KEYINPUT96), .A3(new_n679), .A4(new_n371), .ZN(new_n680));
  AND3_X1   g494(.A1(new_n656), .A2(new_n659), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n636), .A2(new_n681), .ZN(new_n682));
  XOR2_X1   g496(.A(KEYINPUT35), .B(G107), .Z(new_n683));
  XNOR2_X1  g497(.A(new_n682), .B(new_n683), .ZN(G9));
  INV_X1    g498(.A(KEYINPUT36), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n609), .A2(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n687), .A2(new_n612), .A3(new_n614), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n606), .A2(new_n686), .ZN(new_n689));
  AND3_X1   g503(.A1(new_n688), .A2(new_n689), .A3(new_n618), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n626), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(KEYINPUT97), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n690), .B1(new_n623), .B2(new_n625), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT97), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  AND2_X1   g510(.A1(new_n693), .A2(new_n696), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n433), .A2(new_n505), .A3(new_n634), .A4(new_n697), .ZN(new_n698));
  XOR2_X1   g512(.A(KEYINPUT37), .B(G110), .Z(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(KEYINPUT98), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n698), .B(new_n700), .ZN(G12));
  AND2_X1   g515(.A1(new_n697), .A2(new_n659), .ZN(new_n702));
  INV_X1    g516(.A(G900), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n364), .B1(new_n368), .B2(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n675), .A2(new_n679), .A3(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n505), .A2(new_n575), .A3(new_n702), .A4(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G128), .ZN(G30));
  XOR2_X1   g523(.A(new_n704), .B(KEYINPUT39), .Z(new_n710));
  NAND2_X1  g524(.A1(new_n505), .A2(new_n710), .ZN(new_n711));
  OR2_X1    g525(.A1(new_n711), .A2(KEYINPUT40), .ZN(new_n712));
  XNOR2_X1  g526(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n713));
  XOR2_X1   g527(.A(new_n297), .B(new_n713), .Z(new_n714));
  NAND4_X1  g528(.A1(new_n640), .A2(new_n679), .A3(new_n187), .A4(new_n694), .ZN(new_n715));
  XOR2_X1   g529(.A(new_n715), .B(KEYINPUT102), .Z(new_n716));
  AND2_X1   g530(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n711), .A2(KEYINPUT40), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n573), .A2(new_n554), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(KEYINPUT32), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n633), .A2(new_n570), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT101), .ZN(new_n723));
  AND2_X1   g537(.A1(new_n561), .A2(new_n567), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n536), .B1(new_n517), .B2(new_n546), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(KEYINPUT100), .ZN(new_n726));
  AOI21_X1  g540(.A(G902), .B1(new_n724), .B2(new_n726), .ZN(new_n727));
  OAI211_X1 g541(.A(new_n722), .B(new_n723), .C1(new_n631), .C2(new_n727), .ZN(new_n728));
  OAI22_X1  g542(.A1(new_n569), .A2(new_n574), .B1(new_n727), .B2(new_n631), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(KEYINPUT101), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n712), .A2(new_n717), .A3(new_n718), .A4(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G143), .ZN(G45));
  NAND4_X1  g547(.A1(new_n640), .A2(new_n646), .A3(new_n648), .A4(new_n705), .ZN(new_n734));
  INV_X1    g548(.A(new_n734), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n505), .A2(new_n575), .A3(new_n702), .A4(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G146), .ZN(G48));
  OAI21_X1  g551(.A(new_n434), .B1(new_n496), .B2(new_n436), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n738), .B1(new_n498), .B2(new_n488), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n575), .A2(new_n650), .A3(new_n628), .A4(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(KEYINPUT103), .ZN(new_n741));
  XOR2_X1   g555(.A(KEYINPUT41), .B(G113), .Z(new_n742));
  XNOR2_X1  g556(.A(new_n741), .B(new_n742), .ZN(G15));
  NAND4_X1  g557(.A1(new_n681), .A2(new_n575), .A3(new_n628), .A4(new_n739), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G116), .ZN(G18));
  INV_X1    g559(.A(new_n738), .ZN(new_n746));
  AND3_X1   g560(.A1(new_n499), .A2(new_n746), .A3(new_n659), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n693), .A2(new_n358), .A3(new_n696), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n748), .A2(new_n431), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n747), .A2(new_n575), .A3(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G119), .ZN(G21));
  AOI22_X1  g565(.A1(new_n536), .A2(new_n548), .B1(new_n558), .B2(new_n559), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n555), .B1(new_n752), .B2(new_n568), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n632), .A2(new_n753), .ZN(new_n754));
  AND3_X1   g568(.A1(new_n739), .A2(new_n754), .A3(new_n628), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT105), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT104), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n757), .B1(new_n675), .B2(new_n358), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n640), .A2(new_n679), .A3(KEYINPUT104), .ZN(new_n759));
  AND4_X1   g573(.A1(new_n756), .A2(new_n758), .A3(new_n659), .A4(new_n759), .ZN(new_n760));
  AOI21_X1  g574(.A(KEYINPUT104), .B1(new_n640), .B2(new_n679), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n761), .A2(new_n639), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n756), .B1(new_n762), .B2(new_n759), .ZN(new_n763));
  OAI211_X1 g577(.A(new_n755), .B(new_n371), .C1(new_n760), .C2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G122), .ZN(G24));
  NOR4_X1   g579(.A1(new_n632), .A2(new_n734), .A3(new_n753), .A4(new_n694), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n747), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G125), .ZN(G27));
  AND2_X1   g582(.A1(new_n296), .A2(new_n187), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n295), .A2(new_n434), .A3(new_n769), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n770), .B1(new_n499), .B2(new_n504), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n734), .A2(KEYINPUT42), .ZN(new_n772));
  AND4_X1   g586(.A1(new_n575), .A2(new_n771), .A3(new_n628), .A4(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT106), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n720), .A2(new_n774), .A3(new_n721), .ZN(new_n775));
  OAI21_X1  g589(.A(KEYINPUT106), .B1(new_n569), .B2(new_n574), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n775), .A2(new_n776), .A3(new_n553), .ZN(new_n777));
  AOI22_X1  g591(.A1(new_n488), .A2(new_n498), .B1(G469), .B2(new_n503), .ZN(new_n778));
  NOR3_X1   g592(.A1(new_n778), .A2(new_n734), .A3(new_n770), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n777), .A2(new_n628), .A3(new_n779), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n773), .B1(new_n780), .B2(KEYINPUT42), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G131), .ZN(G33));
  NAND4_X1  g596(.A1(new_n771), .A2(new_n575), .A3(new_n628), .A4(new_n707), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G134), .ZN(G36));
  NAND2_X1  g598(.A1(new_n295), .A2(new_n769), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n646), .A2(new_n648), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n786), .A2(new_n640), .ZN(new_n787));
  INV_X1    g601(.A(new_n787), .ZN(new_n788));
  OR2_X1    g602(.A1(new_n788), .A2(KEYINPUT43), .ZN(new_n789));
  INV_X1    g603(.A(new_n634), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n788), .A2(KEYINPUT43), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n789), .A2(new_n790), .A3(new_n692), .A4(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT44), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n785), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n794), .B1(new_n793), .B2(new_n792), .ZN(new_n795));
  INV_X1    g609(.A(new_n434), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT45), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n436), .B1(new_n502), .B2(new_n797), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n798), .B1(new_n797), .B2(new_n502), .ZN(new_n799));
  NAND2_X1  g613(.A1(G469), .A2(G902), .ZN(new_n800));
  AOI21_X1  g614(.A(KEYINPUT46), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n801), .B1(new_n498), .B2(new_n488), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n799), .A2(KEYINPUT46), .A3(new_n800), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n796), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(new_n710), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n795), .A2(new_n805), .ZN(new_n806));
  XOR2_X1   g620(.A(KEYINPUT107), .B(G137), .Z(new_n807));
  XNOR2_X1  g621(.A(new_n806), .B(new_n807), .ZN(G39));
  INV_X1    g622(.A(KEYINPUT47), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n809), .A2(KEYINPUT108), .ZN(new_n810));
  INV_X1    g624(.A(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n804), .A2(new_n811), .ZN(new_n812));
  NOR4_X1   g626(.A1(new_n575), .A2(new_n628), .A3(new_n734), .A4(new_n785), .ZN(new_n813));
  XNOR2_X1  g627(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n814));
  OAI211_X1 g628(.A(new_n812), .B(new_n813), .C1(new_n804), .C2(new_n814), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(G140), .ZN(G42));
  INV_X1    g630(.A(KEYINPUT110), .ZN(new_n817));
  AND4_X1   g631(.A1(new_n817), .A2(new_n626), .A3(new_n691), .A4(new_n705), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n817), .B1(new_n694), .B2(new_n705), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n434), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n820), .B1(new_n499), .B2(new_n504), .ZN(new_n821));
  OAI211_X1 g635(.A(new_n729), .B(new_n821), .C1(new_n763), .C2(new_n760), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n822), .A2(new_n708), .A3(new_n736), .A4(new_n767), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT52), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n697), .A2(new_n659), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n826), .B1(new_n722), .B2(new_n553), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n778), .A2(new_n435), .A3(new_n706), .ZN(new_n828));
  AOI22_X1  g642(.A1(new_n827), .A2(new_n828), .B1(new_n747), .B2(new_n766), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n829), .A2(KEYINPUT52), .A3(new_n736), .A4(new_n822), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n825), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n780), .A2(KEYINPUT42), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n675), .A2(new_n705), .ZN(new_n833));
  NOR3_X1   g647(.A1(new_n785), .A2(new_n748), .A3(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n505), .A2(new_n834), .A3(new_n575), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n766), .A2(new_n771), .ZN(new_n836));
  AND3_X1   g650(.A1(new_n783), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(new_n773), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n832), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n675), .A2(new_n679), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n649), .A2(new_n840), .ZN(new_n841));
  AND4_X1   g655(.A1(new_n187), .A2(new_n841), .A3(new_n297), .A4(new_n371), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n842), .A2(new_n628), .A3(new_n505), .A4(new_n634), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n843), .A2(new_n629), .A3(new_n698), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n763), .A2(new_n760), .ZN(new_n845));
  INV_X1    g659(.A(new_n628), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n632), .A2(new_n846), .A3(new_n753), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n847), .A2(new_n371), .A3(new_n739), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n744), .B1(new_n845), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n750), .A2(new_n740), .ZN(new_n850));
  NOR3_X1   g664(.A1(new_n844), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n831), .A2(new_n839), .A3(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT53), .ZN(new_n853));
  OAI21_X1  g667(.A(KEYINPUT111), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n825), .A2(new_n830), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n849), .A2(new_n850), .ZN(new_n856));
  AND3_X1   g670(.A1(new_n843), .A2(new_n629), .A3(new_n698), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n856), .A2(new_n781), .A3(new_n857), .A4(new_n837), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n853), .B1(new_n855), .B2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(new_n859), .ZN(new_n860));
  OR2_X1    g674(.A1(new_n854), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n854), .A2(new_n860), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n861), .A2(KEYINPUT54), .A3(new_n862), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n812), .B1(new_n804), .B2(new_n814), .ZN(new_n864));
  INV_X1    g678(.A(new_n496), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n865), .A2(G469), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n499), .A2(new_n435), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n864), .A2(new_n867), .ZN(new_n868));
  AND3_X1   g682(.A1(new_n789), .A2(new_n364), .A3(new_n791), .ZN(new_n869));
  INV_X1    g683(.A(new_n785), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n869), .A2(new_n847), .A3(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n868), .A2(new_n872), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n714), .A2(new_n187), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n874), .A2(new_n755), .A3(new_n869), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT50), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n875), .B(new_n876), .ZN(new_n877));
  AND3_X1   g691(.A1(new_n869), .A2(new_n739), .A3(new_n870), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n878), .A2(new_n692), .A3(new_n754), .ZN(new_n879));
  INV_X1    g693(.A(new_n731), .ZN(new_n880));
  AND4_X1   g694(.A1(new_n628), .A2(new_n739), .A3(new_n364), .A4(new_n870), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n880), .A2(new_n675), .A3(new_n786), .A4(new_n881), .ZN(new_n882));
  AND2_X1   g696(.A1(new_n879), .A2(new_n882), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n873), .A2(KEYINPUT51), .A3(new_n877), .A4(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT51), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n883), .A2(new_n877), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n871), .B1(new_n864), .B2(new_n867), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n885), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n869), .A2(new_n747), .A3(new_n847), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT115), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n889), .B(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n880), .A2(new_n881), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n892), .A2(new_n649), .ZN(new_n893));
  AND2_X1   g707(.A1(new_n777), .A2(new_n628), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n878), .A2(new_n894), .ZN(new_n895));
  OR2_X1    g709(.A1(new_n895), .A2(KEYINPUT48), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n895), .A2(KEYINPUT48), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n893), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  AND4_X1   g712(.A1(new_n884), .A2(new_n888), .A3(new_n891), .A4(new_n898), .ZN(new_n899));
  AND2_X1   g713(.A1(new_n750), .A2(new_n740), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n900), .A2(KEYINPUT112), .A3(new_n764), .A4(new_n744), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT112), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n902), .B1(new_n849), .B2(new_n850), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n844), .A2(new_n853), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n904), .A2(new_n839), .A3(new_n831), .A4(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n859), .A2(new_n906), .ZN(new_n907));
  OAI21_X1  g721(.A(KEYINPUT113), .B1(new_n907), .B2(KEYINPUT54), .ZN(new_n908));
  OR3_X1    g722(.A1(new_n907), .A2(KEYINPUT113), .A3(KEYINPUT54), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n863), .A2(new_n899), .A3(new_n908), .A4(new_n909), .ZN(new_n910));
  OAI21_X1  g724(.A(G953), .B1(new_n910), .B2(KEYINPUT114), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT114), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n360), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  NOR3_X1   g727(.A1(new_n846), .A2(new_n435), .A3(new_n657), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n914), .B(KEYINPUT109), .ZN(new_n915));
  NOR3_X1   g729(.A1(new_n915), .A2(new_n714), .A3(new_n788), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n499), .A2(new_n866), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n917), .B(KEYINPUT49), .Z(new_n918));
  NAND3_X1  g732(.A1(new_n916), .A2(new_n918), .A3(new_n880), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n911), .A2(new_n913), .A3(new_n919), .ZN(G75));
  NOR2_X1   g734(.A1(new_n367), .A2(G952), .ZN(new_n921));
  INV_X1    g735(.A(new_n921), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n270), .B1(new_n859), .B2(new_n906), .ZN(new_n923));
  AOI21_X1  g737(.A(KEYINPUT56), .B1(new_n923), .B2(G210), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n239), .A2(new_n243), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n925), .B(new_n268), .ZN(new_n926));
  XOR2_X1   g740(.A(KEYINPUT116), .B(KEYINPUT55), .Z(new_n927));
  XNOR2_X1  g741(.A(new_n926), .B(new_n927), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n922), .B1(new_n924), .B2(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n929), .B1(new_n924), .B2(new_n928), .ZN(G51));
  XNOR2_X1  g744(.A(new_n907), .B(KEYINPUT54), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n800), .B(KEYINPUT57), .Z(new_n932));
  AOI22_X1  g746(.A1(new_n931), .A2(new_n932), .B1(new_n494), .B2(new_n495), .ZN(new_n933));
  OR2_X1    g747(.A1(new_n933), .A2(KEYINPUT117), .ZN(new_n934));
  AOI211_X1 g748(.A(new_n270), .B(new_n799), .C1(new_n859), .C2(new_n906), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n935), .B1(new_n933), .B2(KEYINPUT117), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n921), .B1(new_n934), .B2(new_n936), .ZN(G54));
  AND3_X1   g751(.A1(new_n923), .A2(KEYINPUT58), .A3(G475), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n922), .B1(new_n938), .B2(new_n426), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n939), .B1(new_n426), .B2(new_n938), .ZN(G60));
  NAND2_X1  g754(.A1(new_n643), .A2(new_n645), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n863), .A2(new_n908), .A3(new_n909), .ZN(new_n942));
  XOR2_X1   g756(.A(new_n647), .B(KEYINPUT59), .Z(new_n943));
  AOI21_X1  g757(.A(new_n941), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  AND2_X1   g758(.A1(new_n941), .A2(new_n943), .ZN(new_n945));
  AOI211_X1 g759(.A(KEYINPUT118), .B(new_n921), .C1(new_n931), .C2(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT118), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n931), .A2(new_n945), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n947), .B1(new_n948), .B2(new_n922), .ZN(new_n949));
  NOR3_X1   g763(.A1(new_n944), .A2(new_n946), .A3(new_n949), .ZN(G63));
  NAND2_X1  g764(.A1(G217), .A2(G902), .ZN(new_n951));
  XOR2_X1   g765(.A(new_n951), .B(KEYINPUT120), .Z(new_n952));
  XOR2_X1   g766(.A(new_n952), .B(KEYINPUT60), .Z(new_n953));
  NAND2_X1  g767(.A1(new_n907), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n611), .A2(new_n615), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n955), .B(KEYINPUT121), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(new_n953), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n958), .B1(new_n859), .B2(new_n906), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n959), .A2(new_n688), .A3(new_n689), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n957), .A2(new_n960), .A3(KEYINPUT61), .A4(new_n922), .ZN(new_n961));
  XOR2_X1   g775(.A(KEYINPUT119), .B(KEYINPUT61), .Z(new_n962));
  AOI21_X1  g776(.A(KEYINPUT122), .B1(new_n957), .B2(new_n922), .ZN(new_n963));
  INV_X1    g777(.A(new_n956), .ZN(new_n964));
  OAI211_X1 g778(.A(KEYINPUT122), .B(new_n922), .C1(new_n959), .C2(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n965), .A2(new_n960), .ZN(new_n966));
  OAI211_X1 g780(.A(KEYINPUT123), .B(new_n962), .C1(new_n963), .C2(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n922), .B1(new_n959), .B2(new_n964), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT122), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n971), .A2(new_n960), .A3(new_n965), .ZN(new_n972));
  AOI21_X1  g786(.A(KEYINPUT123), .B1(new_n972), .B2(new_n962), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n961), .B1(new_n968), .B2(new_n973), .ZN(G66));
  OAI21_X1  g788(.A(G953), .B1(new_n369), .B2(new_n266), .ZN(new_n975));
  INV_X1    g789(.A(new_n367), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n975), .B1(new_n851), .B2(new_n976), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n925), .B1(G898), .B2(new_n367), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n977), .B(new_n978), .ZN(G69));
  NAND2_X1  g793(.A1(new_n524), .A2(new_n525), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n420), .A2(new_n421), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n980), .B(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(new_n982), .ZN(new_n983));
  AND2_X1   g797(.A1(new_n829), .A2(new_n736), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n732), .A2(new_n984), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n985), .B(KEYINPUT62), .ZN(new_n986));
  INV_X1    g800(.A(new_n815), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n575), .A2(new_n628), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n870), .A2(new_n841), .ZN(new_n989));
  NOR3_X1   g803(.A1(new_n711), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n990), .B(KEYINPUT124), .ZN(new_n991));
  NOR4_X1   g805(.A1(new_n986), .A2(new_n806), .A3(new_n987), .A4(new_n991), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n983), .B1(new_n992), .B2(new_n976), .ZN(new_n993));
  NAND4_X1  g807(.A1(new_n815), .A2(new_n781), .A3(new_n783), .A4(new_n984), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n894), .B1(new_n760), .B2(new_n763), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n805), .B1(new_n795), .B2(new_n995), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n367), .B1(new_n994), .B2(new_n996), .ZN(new_n997));
  NOR2_X1   g811(.A1(new_n367), .A2(G900), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n998), .B(KEYINPUT125), .ZN(new_n999));
  AND2_X1   g813(.A1(new_n997), .A2(new_n999), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n993), .B1(new_n983), .B2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n367), .B1(G227), .B2(G900), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n1002), .B1(new_n983), .B2(KEYINPUT126), .ZN(new_n1003));
  INV_X1    g817(.A(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g818(.A(new_n1001), .B(new_n1004), .ZN(G72));
  NAND2_X1  g819(.A1(G472), .A2(G902), .ZN(new_n1006));
  XNOR2_X1  g820(.A(new_n1006), .B(KEYINPUT63), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n861), .A2(new_n862), .ZN(new_n1008));
  AND2_X1   g822(.A1(new_n533), .A2(new_n538), .ZN(new_n1009));
  AOI211_X1 g823(.A(new_n1007), .B(new_n1008), .C1(new_n724), .C2(new_n1009), .ZN(new_n1010));
  INV_X1    g824(.A(new_n851), .ZN(new_n1011));
  NOR3_X1   g825(.A1(new_n994), .A2(new_n1011), .A3(new_n996), .ZN(new_n1012));
  XOR2_X1   g826(.A(new_n1007), .B(KEYINPUT127), .Z(new_n1013));
  OAI211_X1 g827(.A(new_n536), .B(new_n528), .C1(new_n1012), .C2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n1013), .B1(new_n992), .B2(new_n851), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n532), .B1(new_n537), .B2(new_n517), .ZN(new_n1016));
  OAI211_X1 g830(.A(new_n922), .B(new_n1014), .C1(new_n1015), .C2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g831(.A1(new_n1010), .A2(new_n1017), .ZN(G57));
endmodule


