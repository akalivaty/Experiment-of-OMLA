

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580;

  NOR2_X2 U320 ( .A1(n514), .A2(n469), .ZN(n470) );
  NOR2_X2 U321 ( .A1(n570), .A2(n451), .ZN(n452) );
  XNOR2_X2 U322 ( .A(n291), .B(n302), .ZN(n430) );
  BUF_X1 U323 ( .A(n561), .Z(n288) );
  NOR2_X1 U324 ( .A1(n402), .A2(n401), .ZN(n479) );
  XOR2_X1 U325 ( .A(n441), .B(n440), .Z(n574) );
  NOR2_X1 U326 ( .A1(n563), .A2(n467), .ZN(n468) );
  XNOR2_X1 U327 ( .A(n445), .B(n444), .ZN(n495) );
  XOR2_X1 U328 ( .A(n373), .B(n372), .Z(n512) );
  XNOR2_X1 U329 ( .A(KEYINPUT93), .B(n400), .ZN(n537) );
  XOR2_X1 U330 ( .A(G211GAT), .B(KEYINPUT21), .Z(n289) );
  XOR2_X1 U331 ( .A(n410), .B(n409), .Z(n290) );
  XOR2_X1 U332 ( .A(KEYINPUT70), .B(G1GAT), .Z(n291) );
  XOR2_X1 U333 ( .A(n365), .B(n431), .Z(n292) );
  XNOR2_X1 U334 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U335 ( .A(n437), .B(n436), .ZN(n438) );
  NAND2_X1 U336 ( .A1(n442), .A2(n549), .ZN(n443) );
  XOR2_X1 U337 ( .A(n530), .B(KEYINPUT36), .Z(n578) );
  XNOR2_X1 U338 ( .A(n443), .B(KEYINPUT37), .ZN(n510) );
  INV_X1 U339 ( .A(G190GAT), .ZN(n471) );
  INV_X1 U340 ( .A(G36GAT), .ZN(n446) );
  XNOR2_X1 U341 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U342 ( .A(n446), .B(KEYINPUT104), .ZN(n447) );
  XNOR2_X1 U343 ( .A(n474), .B(n473), .ZN(G1351GAT) );
  XNOR2_X1 U344 ( .A(n448), .B(n447), .ZN(G1329GAT) );
  XOR2_X1 U345 ( .A(KEYINPUT38), .B(KEYINPUT103), .Z(n445) );
  XOR2_X1 U346 ( .A(KEYINPUT66), .B(KEYINPUT67), .Z(n294) );
  XNOR2_X1 U347 ( .A(G113GAT), .B(G8GAT), .ZN(n293) );
  XNOR2_X1 U348 ( .A(n294), .B(n293), .ZN(n310) );
  XOR2_X1 U349 ( .A(G197GAT), .B(G141GAT), .Z(n296) );
  XNOR2_X1 U350 ( .A(G169GAT), .B(G36GAT), .ZN(n295) );
  XNOR2_X1 U351 ( .A(n296), .B(n295), .ZN(n298) );
  XOR2_X1 U352 ( .A(G29GAT), .B(G43GAT), .Z(n297) );
  XNOR2_X1 U353 ( .A(n298), .B(n297), .ZN(n306) );
  XNOR2_X1 U354 ( .A(KEYINPUT29), .B(KEYINPUT69), .ZN(n299) );
  XNOR2_X1 U355 ( .A(n299), .B(KEYINPUT68), .ZN(n300) );
  XOR2_X1 U356 ( .A(n300), .B(KEYINPUT30), .Z(n304) );
  XNOR2_X1 U357 ( .A(G50GAT), .B(KEYINPUT7), .ZN(n301) );
  XNOR2_X1 U358 ( .A(n301), .B(KEYINPUT8), .ZN(n409) );
  XNOR2_X1 U359 ( .A(G22GAT), .B(G15GAT), .ZN(n302) );
  XNOR2_X1 U360 ( .A(n409), .B(n430), .ZN(n303) );
  XNOR2_X1 U361 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U362 ( .A(n306), .B(n305), .ZN(n308) );
  NAND2_X1 U363 ( .A1(G229GAT), .A2(G233GAT), .ZN(n307) );
  XNOR2_X1 U364 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U365 ( .A(n310), .B(n309), .Z(n540) );
  XOR2_X1 U366 ( .A(KEYINPUT31), .B(KEYINPUT32), .Z(n312) );
  NAND2_X1 U367 ( .A1(G230GAT), .A2(G233GAT), .ZN(n311) );
  XNOR2_X1 U368 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U369 ( .A(n313), .B(KEYINPUT33), .Z(n318) );
  XOR2_X1 U370 ( .A(G78GAT), .B(KEYINPUT72), .Z(n315) );
  XNOR2_X1 U371 ( .A(G106GAT), .B(KEYINPUT71), .ZN(n314) );
  XNOR2_X1 U372 ( .A(n315), .B(n314), .ZN(n351) );
  XNOR2_X1 U373 ( .A(G204GAT), .B(G92GAT), .ZN(n316) );
  XOR2_X1 U374 ( .A(n316), .B(G64GAT), .Z(n373) );
  XOR2_X1 U375 ( .A(n351), .B(n373), .Z(n317) );
  XNOR2_X1 U376 ( .A(n318), .B(n317), .ZN(n322) );
  XOR2_X1 U377 ( .A(KEYINPUT13), .B(G85GAT), .Z(n320) );
  XNOR2_X1 U378 ( .A(G176GAT), .B(G120GAT), .ZN(n319) );
  XNOR2_X1 U379 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U380 ( .A(n322), .B(n321), .ZN(n324) );
  XOR2_X1 U381 ( .A(G99GAT), .B(G71GAT), .Z(n384) );
  XOR2_X1 U382 ( .A(G148GAT), .B(G57GAT), .Z(n328) );
  XOR2_X1 U383 ( .A(n384), .B(n328), .Z(n323) );
  XNOR2_X1 U384 ( .A(n324), .B(n323), .ZN(n570) );
  NOR2_X1 U385 ( .A1(n540), .A2(n570), .ZN(n480) );
  XOR2_X1 U386 ( .A(KEYINPUT90), .B(KEYINPUT92), .Z(n326) );
  XNOR2_X1 U387 ( .A(G134GAT), .B(KEYINPUT1), .ZN(n325) );
  XNOR2_X1 U388 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U389 ( .A(n327), .B(KEYINPUT4), .Z(n330) );
  XNOR2_X1 U390 ( .A(G1GAT), .B(n328), .ZN(n329) );
  XNOR2_X1 U391 ( .A(n330), .B(n329), .ZN(n336) );
  XOR2_X1 U392 ( .A(G29GAT), .B(G85GAT), .Z(n410) );
  XOR2_X1 U393 ( .A(G120GAT), .B(G127GAT), .Z(n332) );
  XNOR2_X1 U394 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n331) );
  XNOR2_X1 U395 ( .A(n332), .B(n331), .ZN(n381) );
  XOR2_X1 U396 ( .A(n410), .B(n381), .Z(n334) );
  NAND2_X1 U397 ( .A1(G225GAT), .A2(G233GAT), .ZN(n333) );
  XNOR2_X1 U398 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U399 ( .A(n336), .B(n335), .Z(n345) );
  XNOR2_X1 U400 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n337) );
  XNOR2_X1 U401 ( .A(n337), .B(KEYINPUT2), .ZN(n338) );
  XOR2_X1 U402 ( .A(n338), .B(KEYINPUT87), .Z(n340) );
  XNOR2_X1 U403 ( .A(G141GAT), .B(G162GAT), .ZN(n339) );
  XNOR2_X1 U404 ( .A(n340), .B(n339), .ZN(n356) );
  XOR2_X1 U405 ( .A(KEYINPUT89), .B(KEYINPUT5), .Z(n342) );
  XNOR2_X1 U406 ( .A(KEYINPUT91), .B(KEYINPUT6), .ZN(n341) );
  XNOR2_X1 U407 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U408 ( .A(n356), .B(n343), .ZN(n344) );
  XNOR2_X1 U409 ( .A(n345), .B(n344), .ZN(n400) );
  XOR2_X1 U410 ( .A(KEYINPUT86), .B(KEYINPUT24), .Z(n347) );
  XNOR2_X1 U411 ( .A(KEYINPUT23), .B(KEYINPUT22), .ZN(n346) );
  XNOR2_X1 U412 ( .A(n347), .B(n346), .ZN(n360) );
  XNOR2_X1 U413 ( .A(G197GAT), .B(G218GAT), .ZN(n348) );
  XNOR2_X1 U414 ( .A(n289), .B(n348), .ZN(n362) );
  XOR2_X1 U415 ( .A(KEYINPUT88), .B(n362), .Z(n350) );
  XNOR2_X1 U416 ( .A(G50GAT), .B(G148GAT), .ZN(n349) );
  XNOR2_X1 U417 ( .A(n350), .B(n349), .ZN(n355) );
  XOR2_X1 U418 ( .A(G204GAT), .B(n351), .Z(n353) );
  NAND2_X1 U419 ( .A1(G228GAT), .A2(G233GAT), .ZN(n352) );
  XNOR2_X1 U420 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U421 ( .A(n355), .B(n354), .Z(n358) );
  XNOR2_X1 U422 ( .A(G22GAT), .B(n356), .ZN(n357) );
  XNOR2_X1 U423 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U424 ( .A(n360), .B(n359), .Z(n467) );
  XOR2_X1 U425 ( .A(n467), .B(KEYINPUT28), .Z(n517) );
  INV_X1 U426 ( .A(n517), .ZN(n361) );
  NOR2_X1 U427 ( .A1(n537), .A2(n361), .ZN(n376) );
  XNOR2_X1 U428 ( .A(KEYINPUT94), .B(n362), .ZN(n364) );
  AND2_X1 U429 ( .A1(G226GAT), .A2(G233GAT), .ZN(n363) );
  XNOR2_X1 U430 ( .A(n364), .B(n363), .ZN(n365) );
  XOR2_X1 U431 ( .A(G8GAT), .B(KEYINPUT76), .Z(n431) );
  XOR2_X1 U432 ( .A(KEYINPUT82), .B(KEYINPUT17), .Z(n367) );
  XNOR2_X1 U433 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n366) );
  XNOR2_X1 U434 ( .A(n367), .B(n366), .ZN(n368) );
  XOR2_X1 U435 ( .A(n368), .B(G183GAT), .Z(n370) );
  XNOR2_X1 U436 ( .A(G169GAT), .B(G176GAT), .ZN(n369) );
  XNOR2_X1 U437 ( .A(n370), .B(n369), .ZN(n380) );
  XOR2_X1 U438 ( .A(G36GAT), .B(G190GAT), .Z(n412) );
  XNOR2_X1 U439 ( .A(n380), .B(n412), .ZN(n371) );
  XNOR2_X1 U440 ( .A(n292), .B(n371), .ZN(n372) );
  XNOR2_X1 U441 ( .A(n512), .B(KEYINPUT95), .ZN(n374) );
  XOR2_X1 U442 ( .A(KEYINPUT27), .B(n374), .Z(n396) );
  INV_X1 U443 ( .A(n396), .ZN(n375) );
  NAND2_X1 U444 ( .A1(n376), .A2(n375), .ZN(n521) );
  XNOR2_X1 U445 ( .A(n521), .B(KEYINPUT96), .ZN(n391) );
  XOR2_X1 U446 ( .A(KEYINPUT83), .B(KEYINPUT20), .Z(n378) );
  XNOR2_X1 U447 ( .A(G15GAT), .B(KEYINPUT84), .ZN(n377) );
  XNOR2_X1 U448 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U449 ( .A(n380), .B(n379), .ZN(n389) );
  XOR2_X1 U450 ( .A(G43GAT), .B(G134GAT), .Z(n413) );
  XOR2_X1 U451 ( .A(n381), .B(n413), .Z(n383) );
  NAND2_X1 U452 ( .A1(G227GAT), .A2(G233GAT), .ZN(n382) );
  XNOR2_X1 U453 ( .A(n383), .B(n382), .ZN(n385) );
  XOR2_X1 U454 ( .A(n385), .B(n384), .Z(n387) );
  XNOR2_X1 U455 ( .A(G190GAT), .B(KEYINPUT81), .ZN(n386) );
  XNOR2_X1 U456 ( .A(n387), .B(n386), .ZN(n388) );
  XOR2_X1 U457 ( .A(n389), .B(n388), .Z(n522) );
  XOR2_X1 U458 ( .A(n522), .B(KEYINPUT85), .Z(n390) );
  NOR2_X1 U459 ( .A1(n391), .A2(n390), .ZN(n402) );
  INV_X1 U460 ( .A(n522), .ZN(n514) );
  NOR2_X1 U461 ( .A1(n514), .A2(n512), .ZN(n392) );
  NOR2_X1 U462 ( .A1(n467), .A2(n392), .ZN(n393) );
  XOR2_X1 U463 ( .A(n393), .B(KEYINPUT98), .Z(n394) );
  XNOR2_X1 U464 ( .A(KEYINPUT25), .B(n394), .ZN(n398) );
  NAND2_X1 U465 ( .A1(n467), .A2(n514), .ZN(n395) );
  XNOR2_X1 U466 ( .A(n395), .B(KEYINPUT26), .ZN(n564) );
  NOR2_X1 U467 ( .A1(n564), .A2(n396), .ZN(n539) );
  XOR2_X1 U468 ( .A(n539), .B(KEYINPUT97), .Z(n397) );
  NOR2_X1 U469 ( .A1(n398), .A2(n397), .ZN(n399) );
  NOR2_X1 U470 ( .A1(n400), .A2(n399), .ZN(n401) );
  XOR2_X1 U471 ( .A(KEYINPUT9), .B(KEYINPUT75), .Z(n404) );
  XNOR2_X1 U472 ( .A(KEYINPUT10), .B(KEYINPUT11), .ZN(n403) );
  XNOR2_X1 U473 ( .A(n404), .B(n403), .ZN(n408) );
  XOR2_X1 U474 ( .A(G92GAT), .B(KEYINPUT74), .Z(n406) );
  XNOR2_X1 U475 ( .A(KEYINPUT73), .B(KEYINPUT65), .ZN(n405) );
  XNOR2_X1 U476 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U477 ( .A(n408), .B(n407), .ZN(n421) );
  NAND2_X1 U478 ( .A1(G232GAT), .A2(G233GAT), .ZN(n411) );
  XNOR2_X1 U479 ( .A(n290), .B(n411), .ZN(n417) );
  XOR2_X1 U480 ( .A(n412), .B(G218GAT), .Z(n415) );
  XNOR2_X1 U481 ( .A(n413), .B(G162GAT), .ZN(n414) );
  XOR2_X1 U482 ( .A(n415), .B(n414), .Z(n416) );
  XNOR2_X1 U483 ( .A(n417), .B(n416), .ZN(n419) );
  XNOR2_X1 U484 ( .A(G99GAT), .B(G106GAT), .ZN(n418) );
  XNOR2_X1 U485 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X2 U486 ( .A(n421), .B(n420), .Z(n530) );
  NOR2_X1 U487 ( .A1(n479), .A2(n578), .ZN(n442) );
  XOR2_X1 U488 ( .A(KEYINPUT78), .B(G64GAT), .Z(n423) );
  XNOR2_X1 U489 ( .A(KEYINPUT14), .B(KEYINPUT12), .ZN(n422) );
  XNOR2_X1 U490 ( .A(n423), .B(n422), .ZN(n441) );
  XOR2_X1 U491 ( .A(G211GAT), .B(G78GAT), .Z(n425) );
  XNOR2_X1 U492 ( .A(G183GAT), .B(G155GAT), .ZN(n424) );
  XNOR2_X1 U493 ( .A(n425), .B(n424), .ZN(n429) );
  XOR2_X1 U494 ( .A(KEYINPUT80), .B(G57GAT), .Z(n427) );
  XNOR2_X1 U495 ( .A(G71GAT), .B(G127GAT), .ZN(n426) );
  XNOR2_X1 U496 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U497 ( .A(n429), .B(n428), .Z(n439) );
  XOR2_X1 U498 ( .A(n431), .B(n430), .Z(n437) );
  XOR2_X1 U499 ( .A(KEYINPUT15), .B(KEYINPUT79), .Z(n433) );
  XNOR2_X1 U500 ( .A(KEYINPUT77), .B(KEYINPUT13), .ZN(n432) );
  XNOR2_X1 U501 ( .A(n433), .B(n432), .ZN(n435) );
  NAND2_X1 U502 ( .A1(G231GAT), .A2(G233GAT), .ZN(n434) );
  XNOR2_X1 U503 ( .A(n439), .B(n438), .ZN(n440) );
  INV_X1 U504 ( .A(n574), .ZN(n549) );
  NAND2_X1 U505 ( .A1(n480), .A2(n510), .ZN(n444) );
  NOR2_X1 U506 ( .A1(n495), .A2(n512), .ZN(n448) );
  INV_X1 U507 ( .A(KEYINPUT113), .ZN(n453) );
  NOR2_X1 U508 ( .A1(n549), .A2(n578), .ZN(n449) );
  XNOR2_X1 U509 ( .A(n449), .B(KEYINPUT45), .ZN(n450) );
  NAND2_X1 U510 ( .A1(n450), .A2(n540), .ZN(n451) );
  XNOR2_X1 U511 ( .A(n453), .B(n452), .ZN(n462) );
  XOR2_X1 U512 ( .A(KEYINPUT46), .B(KEYINPUT111), .Z(n456) );
  XNOR2_X1 U513 ( .A(KEYINPUT41), .B(KEYINPUT64), .ZN(n454) );
  XNOR2_X1 U514 ( .A(n570), .B(n454), .ZN(n543) );
  INV_X1 U515 ( .A(n543), .ZN(n557) );
  INV_X1 U516 ( .A(n540), .ZN(n565) );
  NAND2_X1 U517 ( .A1(n557), .A2(n565), .ZN(n455) );
  XNOR2_X1 U518 ( .A(n456), .B(n455), .ZN(n458) );
  NOR2_X1 U519 ( .A1(n530), .A2(n574), .ZN(n457) );
  NAND2_X1 U520 ( .A1(n458), .A2(n457), .ZN(n459) );
  XNOR2_X1 U521 ( .A(KEYINPUT112), .B(n459), .ZN(n460) );
  XNOR2_X1 U522 ( .A(KEYINPUT47), .B(n460), .ZN(n461) );
  NOR2_X1 U523 ( .A1(n462), .A2(n461), .ZN(n463) );
  XNOR2_X1 U524 ( .A(n463), .B(KEYINPUT48), .ZN(n536) );
  XOR2_X1 U525 ( .A(n512), .B(KEYINPUT121), .Z(n464) );
  NOR2_X1 U526 ( .A1(n536), .A2(n464), .ZN(n465) );
  XNOR2_X1 U527 ( .A(n465), .B(KEYINPUT54), .ZN(n466) );
  NAND2_X1 U528 ( .A1(n466), .A2(n537), .ZN(n563) );
  XNOR2_X1 U529 ( .A(n468), .B(KEYINPUT55), .ZN(n469) );
  XNOR2_X1 U530 ( .A(KEYINPUT122), .B(n470), .ZN(n561) );
  NAND2_X1 U531 ( .A1(n288), .A2(n530), .ZN(n474) );
  XOR2_X1 U532 ( .A(KEYINPUT58), .B(KEYINPUT124), .Z(n472) );
  XOR2_X1 U533 ( .A(KEYINPUT99), .B(KEYINPUT100), .Z(n476) );
  XNOR2_X1 U534 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n475) );
  XNOR2_X1 U535 ( .A(n476), .B(n475), .ZN(n482) );
  NOR2_X1 U536 ( .A1(n530), .A2(n549), .ZN(n477) );
  XOR2_X1 U537 ( .A(KEYINPUT16), .B(n477), .Z(n478) );
  NOR2_X1 U538 ( .A1(n479), .A2(n478), .ZN(n498) );
  NAND2_X1 U539 ( .A1(n480), .A2(n498), .ZN(n488) );
  NOR2_X1 U540 ( .A1(n537), .A2(n488), .ZN(n481) );
  XOR2_X1 U541 ( .A(n482), .B(n481), .Z(G1324GAT) );
  NOR2_X1 U542 ( .A1(n512), .A2(n488), .ZN(n483) );
  XOR2_X1 U543 ( .A(G8GAT), .B(n483), .Z(G1325GAT) );
  NOR2_X1 U544 ( .A1(n488), .A2(n514), .ZN(n487) );
  XOR2_X1 U545 ( .A(KEYINPUT101), .B(KEYINPUT35), .Z(n485) );
  XNOR2_X1 U546 ( .A(G15GAT), .B(KEYINPUT102), .ZN(n484) );
  XNOR2_X1 U547 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U548 ( .A(n487), .B(n486), .ZN(G1326GAT) );
  NOR2_X1 U549 ( .A1(n517), .A2(n488), .ZN(n489) );
  XOR2_X1 U550 ( .A(G22GAT), .B(n489), .Z(G1327GAT) );
  NOR2_X1 U551 ( .A1(n495), .A2(n537), .ZN(n491) );
  XNOR2_X1 U552 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n490) );
  XNOR2_X1 U553 ( .A(n491), .B(n490), .ZN(G1328GAT) );
  XNOR2_X1 U554 ( .A(KEYINPUT40), .B(KEYINPUT105), .ZN(n493) );
  NOR2_X1 U555 ( .A1(n514), .A2(n495), .ZN(n492) );
  XNOR2_X1 U556 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U557 ( .A(G43GAT), .B(n494), .ZN(G1330GAT) );
  NOR2_X1 U558 ( .A1(n517), .A2(n495), .ZN(n496) );
  XOR2_X1 U559 ( .A(G50GAT), .B(n496), .Z(G1331GAT) );
  NAND2_X1 U560 ( .A1(n557), .A2(n540), .ZN(n497) );
  XOR2_X1 U561 ( .A(KEYINPUT106), .B(n497), .Z(n509) );
  NAND2_X1 U562 ( .A1(n509), .A2(n498), .ZN(n499) );
  XOR2_X1 U563 ( .A(KEYINPUT107), .B(n499), .Z(n506) );
  NOR2_X1 U564 ( .A1(n537), .A2(n506), .ZN(n501) );
  XNOR2_X1 U565 ( .A(KEYINPUT108), .B(KEYINPUT42), .ZN(n500) );
  XNOR2_X1 U566 ( .A(n501), .B(n500), .ZN(n502) );
  XOR2_X1 U567 ( .A(G57GAT), .B(n502), .Z(G1332GAT) );
  NOR2_X1 U568 ( .A1(n512), .A2(n506), .ZN(n503) );
  XOR2_X1 U569 ( .A(G64GAT), .B(n503), .Z(G1333GAT) );
  NOR2_X1 U570 ( .A1(n514), .A2(n506), .ZN(n505) );
  XNOR2_X1 U571 ( .A(G71GAT), .B(KEYINPUT109), .ZN(n504) );
  XNOR2_X1 U572 ( .A(n505), .B(n504), .ZN(G1334GAT) );
  NOR2_X1 U573 ( .A1(n517), .A2(n506), .ZN(n508) );
  XNOR2_X1 U574 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n507) );
  XNOR2_X1 U575 ( .A(n508), .B(n507), .ZN(G1335GAT) );
  NAND2_X1 U576 ( .A1(n510), .A2(n509), .ZN(n516) );
  NOR2_X1 U577 ( .A1(n537), .A2(n516), .ZN(n511) );
  XOR2_X1 U578 ( .A(G85GAT), .B(n511), .Z(G1336GAT) );
  NOR2_X1 U579 ( .A1(n512), .A2(n516), .ZN(n513) );
  XOR2_X1 U580 ( .A(G92GAT), .B(n513), .Z(G1337GAT) );
  NOR2_X1 U581 ( .A1(n514), .A2(n516), .ZN(n515) );
  XOR2_X1 U582 ( .A(G99GAT), .B(n515), .Z(G1338GAT) );
  NOR2_X1 U583 ( .A1(n517), .A2(n516), .ZN(n519) );
  XNOR2_X1 U584 ( .A(KEYINPUT44), .B(KEYINPUT110), .ZN(n518) );
  XNOR2_X1 U585 ( .A(n519), .B(n518), .ZN(n520) );
  XOR2_X1 U586 ( .A(G106GAT), .B(n520), .Z(G1339GAT) );
  NOR2_X1 U587 ( .A1(n536), .A2(n521), .ZN(n523) );
  NAND2_X1 U588 ( .A1(n523), .A2(n522), .ZN(n531) );
  NOR2_X1 U589 ( .A1(n540), .A2(n531), .ZN(n524) );
  XOR2_X1 U590 ( .A(G113GAT), .B(n524), .Z(G1340GAT) );
  NOR2_X1 U591 ( .A1(n543), .A2(n531), .ZN(n526) );
  XNOR2_X1 U592 ( .A(KEYINPUT49), .B(KEYINPUT114), .ZN(n525) );
  XNOR2_X1 U593 ( .A(n526), .B(n525), .ZN(n527) );
  XNOR2_X1 U594 ( .A(G120GAT), .B(n527), .ZN(G1341GAT) );
  NOR2_X1 U595 ( .A1(n549), .A2(n531), .ZN(n528) );
  XOR2_X1 U596 ( .A(KEYINPUT50), .B(n528), .Z(n529) );
  XNOR2_X1 U597 ( .A(G127GAT), .B(n529), .ZN(G1342GAT) );
  INV_X1 U598 ( .A(n530), .ZN(n552) );
  NOR2_X1 U599 ( .A1(n531), .A2(n552), .ZN(n535) );
  XOR2_X1 U600 ( .A(KEYINPUT115), .B(KEYINPUT51), .Z(n533) );
  XNOR2_X1 U601 ( .A(G134GAT), .B(KEYINPUT116), .ZN(n532) );
  XNOR2_X1 U602 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U603 ( .A(n535), .B(n534), .ZN(G1343GAT) );
  NOR2_X1 U604 ( .A1(n537), .A2(n536), .ZN(n538) );
  NAND2_X1 U605 ( .A1(n539), .A2(n538), .ZN(n551) );
  NOR2_X1 U606 ( .A1(n540), .A2(n551), .ZN(n542) );
  XNOR2_X1 U607 ( .A(G141GAT), .B(KEYINPUT117), .ZN(n541) );
  XNOR2_X1 U608 ( .A(n542), .B(n541), .ZN(G1344GAT) );
  NOR2_X1 U609 ( .A1(n543), .A2(n551), .ZN(n548) );
  XOR2_X1 U610 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n545) );
  XNOR2_X1 U611 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n544) );
  XNOR2_X1 U612 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U613 ( .A(KEYINPUT53), .B(n546), .ZN(n547) );
  XNOR2_X1 U614 ( .A(n548), .B(n547), .ZN(G1345GAT) );
  NOR2_X1 U615 ( .A1(n549), .A2(n551), .ZN(n550) );
  XOR2_X1 U616 ( .A(G155GAT), .B(n550), .Z(G1346GAT) );
  NOR2_X1 U617 ( .A1(n552), .A2(n551), .ZN(n553) );
  XOR2_X1 U618 ( .A(KEYINPUT120), .B(n553), .Z(n554) );
  XNOR2_X1 U619 ( .A(G162GAT), .B(n554), .ZN(G1347GAT) );
  XOR2_X1 U620 ( .A(G169GAT), .B(KEYINPUT123), .Z(n556) );
  NAND2_X1 U621 ( .A1(n288), .A2(n565), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n556), .B(n555), .ZN(G1348GAT) );
  NAND2_X1 U623 ( .A1(n288), .A2(n557), .ZN(n559) );
  XOR2_X1 U624 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n558) );
  XNOR2_X1 U625 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U626 ( .A(G176GAT), .B(n560), .ZN(G1349GAT) );
  NAND2_X1 U627 ( .A1(n288), .A2(n574), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n562), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U629 ( .A(G197GAT), .B(KEYINPUT60), .Z(n567) );
  NOR2_X1 U630 ( .A1(n564), .A2(n563), .ZN(n576) );
  NAND2_X1 U631 ( .A1(n576), .A2(n565), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n567), .B(n566), .ZN(n569) );
  XOR2_X1 U633 ( .A(KEYINPUT125), .B(KEYINPUT59), .Z(n568) );
  XNOR2_X1 U634 ( .A(n569), .B(n568), .ZN(G1352GAT) );
  XOR2_X1 U635 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n572) );
  NAND2_X1 U636 ( .A1(n576), .A2(n570), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U638 ( .A(G204GAT), .B(n573), .ZN(G1353GAT) );
  NAND2_X1 U639 ( .A1(n576), .A2(n574), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n575), .B(G211GAT), .ZN(G1354GAT) );
  INV_X1 U641 ( .A(n576), .ZN(n577) );
  NOR2_X1 U642 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U643 ( .A(KEYINPUT62), .B(n579), .Z(n580) );
  XNOR2_X1 U644 ( .A(G218GAT), .B(n580), .ZN(G1355GAT) );
endmodule

