//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 0 0 1 0 0 0 0 1 1 1 0 1 0 1 0 0 1 1 0 0 0 0 0 0 0 0 0 1 0 1 1 0 0 0 1 0 0 1 0 1 0 0 1 0 0 0 1 1 1 1 1 0 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n756, new_n757,
    new_n758, new_n760, new_n761, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n791, new_n792, new_n793, new_n794, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n846, new_n847, new_n848,
    new_n850, new_n851, new_n852, new_n853, new_n855, new_n856, new_n857,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n917, new_n918, new_n919, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n942, new_n943, new_n944, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n982, new_n983, new_n984, new_n985, new_n987, new_n988,
    new_n989, new_n990, new_n991;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(G1gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(KEYINPUT16), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n205), .B1(G1gat), .B2(new_n202), .ZN(new_n206));
  INV_X1    g005(.A(G8gat), .ZN(new_n207));
  XNOR2_X1  g006(.A(new_n206), .B(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(G43gat), .B(G50gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT15), .ZN(new_n210));
  XNOR2_X1  g009(.A(new_n209), .B(new_n210), .ZN(new_n211));
  OAI21_X1  g010(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT89), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT14), .ZN(new_n215));
  INV_X1    g014(.A(G29gat), .ZN(new_n216));
  INV_X1    g015(.A(G36gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n215), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n218), .A2(KEYINPUT90), .ZN(new_n219));
  NOR3_X1   g018(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT90), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n214), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  XNOR2_X1  g022(.A(KEYINPUT88), .B(G29gat), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n224), .A2(new_n217), .ZN(new_n225));
  INV_X1    g024(.A(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n218), .A2(KEYINPUT90), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n220), .A2(new_n221), .ZN(new_n228));
  NAND4_X1  g027(.A1(new_n227), .A2(new_n228), .A3(new_n213), .A4(new_n212), .ZN(new_n229));
  NAND4_X1  g028(.A1(new_n211), .A2(new_n223), .A3(new_n226), .A4(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT17), .ZN(new_n231));
  AND2_X1   g030(.A1(new_n209), .A2(KEYINPUT15), .ZN(new_n232));
  OAI211_X1 g031(.A(new_n232), .B(new_n218), .C1(new_n225), .C2(new_n212), .ZN(new_n233));
  AND3_X1   g032(.A1(new_n230), .A2(new_n231), .A3(new_n233), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n231), .B1(new_n230), .B2(new_n233), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n208), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(new_n208), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n230), .A2(new_n233), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(G229gat), .A2(G233gat), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n236), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT18), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  XOR2_X1   g042(.A(new_n238), .B(new_n208), .Z(new_n244));
  XOR2_X1   g043(.A(new_n240), .B(KEYINPUT13), .Z(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n236), .A2(KEYINPUT18), .A3(new_n239), .A4(new_n240), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n243), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(G113gat), .B(G141gat), .ZN(new_n249));
  INV_X1    g048(.A(G197gat), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g050(.A(KEYINPUT11), .B(G169gat), .ZN(new_n252));
  XNOR2_X1  g051(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n253), .B(KEYINPUT12), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n248), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT91), .ZN(new_n257));
  NAND4_X1  g056(.A1(new_n243), .A2(new_n246), .A3(new_n254), .A4(new_n247), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n256), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n257), .B1(new_n256), .B2(new_n258), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(G15gat), .B(G43gat), .ZN(new_n264));
  INV_X1    g063(.A(G71gat), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n264), .B(new_n265), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n266), .B(G99gat), .ZN(new_n267));
  INV_X1    g066(.A(G227gat), .ZN(new_n268));
  INV_X1    g067(.A(G233gat), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  XOR2_X1   g070(.A(G127gat), .B(G134gat), .Z(new_n272));
  XNOR2_X1  g071(.A(new_n272), .B(KEYINPUT69), .ZN(new_n273));
  XNOR2_X1  g072(.A(G113gat), .B(G120gat), .ZN(new_n274));
  AND2_X1   g073(.A1(new_n274), .A2(KEYINPUT68), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT1), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n276), .B1(new_n274), .B2(KEYINPUT68), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n274), .A2(KEYINPUT1), .ZN(new_n279));
  XNOR2_X1  g078(.A(G127gat), .B(G134gat), .ZN(new_n280));
  OAI21_X1  g079(.A(KEYINPUT67), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT67), .ZN(new_n282));
  OAI211_X1 g081(.A(new_n272), .B(new_n282), .C1(KEYINPUT1), .C2(new_n274), .ZN(new_n283));
  AOI22_X1  g082(.A1(new_n273), .A2(new_n278), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(G190gat), .ZN(new_n285));
  AND2_X1   g084(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n286));
  NOR2_X1   g085(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n285), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(KEYINPUT28), .ZN(new_n289));
  XNOR2_X1  g088(.A(KEYINPUT27), .B(G183gat), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT28), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n290), .A2(new_n291), .A3(new_n285), .ZN(new_n292));
  INV_X1    g091(.A(G169gat), .ZN(new_n293));
  INV_X1    g092(.A(G176gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  AOI21_X1  g094(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n296));
  AOI22_X1  g095(.A1(new_n295), .A2(new_n296), .B1(G183gat), .B2(G190gat), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n293), .A2(new_n294), .A3(KEYINPUT26), .ZN(new_n298));
  NAND4_X1  g097(.A1(new_n289), .A2(new_n292), .A3(new_n297), .A4(new_n298), .ZN(new_n299));
  OR3_X1    g098(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n300));
  OAI21_X1  g099(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n301));
  AOI22_X1  g100(.A1(new_n300), .A2(new_n301), .B1(G169gat), .B2(G176gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(G183gat), .A2(G190gat), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT24), .ZN(new_n304));
  OAI21_X1  g103(.A(KEYINPUT64), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  AOI21_X1  g104(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(G183gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(new_n285), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT64), .ZN(new_n310));
  NAND4_X1  g109(.A1(new_n310), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n311));
  NAND4_X1  g110(.A1(new_n305), .A2(new_n307), .A3(new_n309), .A4(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT25), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n302), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n299), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n303), .A2(KEYINPUT65), .ZN(new_n317));
  AOI22_X1  g116(.A1(new_n317), .A2(KEYINPUT24), .B1(new_n306), .B2(KEYINPUT65), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n309), .A2(KEYINPUT66), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT66), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n320), .A2(new_n308), .A3(new_n285), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n318), .A2(new_n319), .A3(new_n321), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n313), .B1(new_n322), .B2(new_n302), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n284), .A2(new_n316), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n273), .A2(new_n278), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n281), .A2(new_n283), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(new_n301), .ZN(new_n329));
  NOR3_X1   g128(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n330));
  OAI22_X1  g129(.A1(new_n329), .A2(new_n330), .B1(new_n293), .B2(new_n294), .ZN(new_n331));
  AND2_X1   g130(.A1(new_n319), .A2(new_n321), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n331), .B1(new_n332), .B2(new_n318), .ZN(new_n333));
  OAI211_X1 g132(.A(new_n299), .B(new_n314), .C1(new_n333), .C2(new_n313), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n328), .A2(new_n334), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n271), .B1(new_n325), .B2(new_n335), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n267), .B1(new_n336), .B2(KEYINPUT33), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT32), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n325), .A2(new_n335), .A3(new_n271), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT34), .ZN(new_n343));
  OR2_X1    g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT70), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n342), .A2(new_n343), .ZN(new_n346));
  AND3_X1   g145(.A1(new_n344), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n337), .A2(new_n339), .ZN(new_n348));
  AND3_X1   g147(.A1(new_n341), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n347), .B1(new_n341), .B2(new_n348), .ZN(new_n350));
  OAI21_X1  g149(.A(KEYINPUT36), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND4_X1  g150(.A1(new_n341), .A2(new_n348), .A3(new_n346), .A4(new_n344), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n344), .A2(new_n346), .ZN(new_n353));
  INV_X1    g152(.A(new_n348), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n353), .B1(new_n354), .B2(new_n340), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n352), .A2(new_n355), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n351), .B1(KEYINPUT36), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(G226gat), .A2(G233gat), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT29), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n359), .B1(new_n334), .B2(new_n360), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n358), .B1(new_n316), .B2(new_n324), .ZN(new_n362));
  XNOR2_X1  g161(.A(G197gat), .B(G204gat), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT22), .ZN(new_n364));
  INV_X1    g163(.A(G211gat), .ZN(new_n365));
  INV_X1    g164(.A(G218gat), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n364), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n363), .A2(new_n367), .ZN(new_n368));
  XNOR2_X1  g167(.A(G211gat), .B(G218gat), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n369), .A2(new_n363), .A3(new_n367), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n373), .ZN(new_n374));
  NOR3_X1   g173(.A1(new_n361), .A2(new_n362), .A3(new_n374), .ZN(new_n375));
  XNOR2_X1  g174(.A(new_n373), .B(KEYINPUT71), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n360), .B1(new_n315), .B2(new_n323), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(new_n358), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n334), .A2(new_n359), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n376), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  XNOR2_X1  g179(.A(G8gat), .B(G36gat), .ZN(new_n381));
  XNOR2_X1  g180(.A(G64gat), .B(G92gat), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n381), .B(new_n382), .ZN(new_n383));
  OR3_X1    g182(.A1(new_n375), .A2(new_n380), .A3(new_n383), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n383), .B1(new_n375), .B2(new_n380), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n384), .A2(new_n385), .A3(KEYINPUT30), .ZN(new_n386));
  OR4_X1    g185(.A1(KEYINPUT30), .A2(new_n375), .A3(new_n380), .A4(new_n383), .ZN(new_n387));
  AND2_X1   g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  XNOR2_X1  g187(.A(G1gat), .B(G29gat), .ZN(new_n389));
  XNOR2_X1  g188(.A(new_n389), .B(KEYINPUT79), .ZN(new_n390));
  XNOR2_X1  g189(.A(KEYINPUT78), .B(KEYINPUT0), .ZN(new_n391));
  XNOR2_X1  g190(.A(new_n390), .B(new_n391), .ZN(new_n392));
  XNOR2_X1  g191(.A(G57gat), .B(G85gat), .ZN(new_n393));
  XOR2_X1   g192(.A(new_n392), .B(new_n393), .Z(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  AND2_X1   g194(.A1(KEYINPUT73), .A2(G148gat), .ZN(new_n396));
  NOR2_X1   g195(.A1(KEYINPUT73), .A2(G148gat), .ZN(new_n397));
  OAI21_X1  g196(.A(G141gat), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(G141gat), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(G148gat), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(G155gat), .A2(G162gat), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(KEYINPUT2), .ZN(new_n403));
  XNOR2_X1  g202(.A(G155gat), .B(G162gat), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(KEYINPUT74), .ZN(new_n405));
  OR2_X1    g204(.A1(G155gat), .A2(G162gat), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT74), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n406), .A2(new_n407), .A3(new_n402), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n401), .A2(new_n403), .A3(new_n405), .A4(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n403), .A2(KEYINPUT72), .ZN(new_n410));
  INV_X1    g209(.A(G148gat), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(G141gat), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n400), .A2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT72), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n402), .A2(new_n414), .A3(KEYINPUT2), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n410), .A2(new_n413), .A3(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n404), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  AND3_X1   g217(.A1(new_n409), .A2(KEYINPUT75), .A3(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(KEYINPUT75), .B1(new_n409), .B2(new_n418), .ZN(new_n420));
  OAI21_X1  g219(.A(KEYINPUT3), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  XOR2_X1   g220(.A(KEYINPUT76), .B(KEYINPUT3), .Z(new_n422));
  NAND3_X1  g221(.A1(new_n409), .A2(new_n422), .A3(new_n418), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n421), .A2(new_n423), .A3(new_n328), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(KEYINPUT77), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT77), .ZN(new_n426));
  NAND4_X1  g225(.A1(new_n421), .A2(new_n426), .A3(new_n423), .A4(new_n328), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(G225gat), .A2(G233gat), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n409), .A2(new_n418), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n284), .A2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT4), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n284), .A2(new_n431), .A3(KEYINPUT4), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  AND4_X1   g236(.A1(KEYINPUT5), .A2(new_n428), .A3(new_n429), .A4(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT5), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT75), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n430), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n409), .A2(KEYINPUT75), .A3(new_n418), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(new_n328), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(new_n432), .ZN(new_n445));
  INV_X1    g244(.A(new_n429), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n439), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n436), .B1(new_n425), .B2(new_n427), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n447), .B1(new_n448), .B2(new_n429), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n395), .B1(new_n438), .B2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT6), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n284), .B1(new_n443), .B2(KEYINPUT3), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n426), .B1(new_n452), .B2(new_n423), .ZN(new_n453));
  INV_X1    g252(.A(new_n427), .ZN(new_n454));
  OAI211_X1 g253(.A(new_n429), .B(new_n437), .C1(new_n453), .C2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n447), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND4_X1  g256(.A1(new_n428), .A2(KEYINPUT5), .A3(new_n429), .A4(new_n437), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n457), .A2(new_n394), .A3(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n450), .A2(new_n451), .A3(new_n459), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n457), .A2(KEYINPUT6), .A3(new_n394), .A4(new_n458), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n388), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  XOR2_X1   g261(.A(G78gat), .B(G106gat), .Z(new_n463));
  XNOR2_X1  g262(.A(new_n463), .B(KEYINPUT31), .ZN(new_n464));
  XNOR2_X1  g263(.A(KEYINPUT80), .B(G50gat), .ZN(new_n465));
  XOR2_X1   g264(.A(new_n464), .B(new_n465), .Z(new_n466));
  INV_X1    g265(.A(G22gat), .ZN(new_n467));
  NAND2_X1  g266(.A1(G228gat), .A2(G233gat), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT71), .ZN(new_n469));
  XNOR2_X1  g268(.A(new_n373), .B(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n423), .A2(new_n360), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n468), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n373), .A2(new_n360), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  OAI22_X1  g273(.A1(new_n474), .A2(KEYINPUT3), .B1(new_n419), .B2(new_n420), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n431), .B1(new_n473), .B2(new_n422), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n373), .B1(new_n423), .B2(new_n360), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n468), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n467), .B1(new_n476), .B2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n476), .A2(new_n479), .A3(new_n467), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n466), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(new_n466), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n485), .B1(new_n482), .B2(KEYINPUT81), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT81), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n476), .A2(new_n479), .A3(new_n487), .A4(new_n467), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n486), .A2(new_n481), .A3(new_n488), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n489), .A2(KEYINPUT82), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT82), .ZN(new_n491));
  INV_X1    g290(.A(new_n482), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n480), .B1(new_n492), .B2(new_n487), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n491), .B1(new_n493), .B2(new_n486), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n484), .B1(new_n490), .B2(new_n494), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n357), .B1(new_n462), .B2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT84), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n428), .A2(new_n437), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT39), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n429), .A2(KEYINPUT83), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n499), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n444), .A2(new_n429), .A3(new_n432), .ZN(new_n503));
  INV_X1    g302(.A(new_n501), .ZN(new_n504));
  OAI211_X1 g303(.A(KEYINPUT39), .B(new_n503), .C1(new_n448), .C2(new_n504), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n502), .A2(new_n505), .A3(new_n395), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT40), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n498), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n502), .A2(new_n505), .A3(KEYINPUT40), .A4(new_n395), .ZN(new_n510));
  AND2_X1   g309(.A1(new_n510), .A2(new_n388), .ZN(new_n511));
  AOI211_X1 g310(.A(new_n446), .B(new_n436), .C1(new_n425), .C2(new_n427), .ZN(new_n512));
  OAI211_X1 g311(.A(new_n458), .B(KEYINPUT85), .C1(new_n512), .C2(new_n447), .ZN(new_n513));
  INV_X1    g312(.A(new_n513), .ZN(new_n514));
  AOI21_X1  g313(.A(KEYINPUT85), .B1(new_n457), .B2(new_n458), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n394), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n506), .A2(new_n498), .A3(new_n507), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n509), .A2(new_n511), .A3(new_n516), .A4(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT38), .ZN(new_n519));
  NOR3_X1   g318(.A1(new_n375), .A2(new_n380), .A3(KEYINPUT37), .ZN(new_n520));
  OAI21_X1  g319(.A(KEYINPUT37), .B1(new_n375), .B2(new_n380), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(new_n383), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT87), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n520), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n521), .A2(KEYINPUT87), .A3(new_n383), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n519), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n520), .A2(KEYINPUT38), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n378), .A2(new_n376), .A3(new_n379), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT86), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n374), .B1(new_n361), .B2(new_n362), .ZN(new_n531));
  NAND4_X1  g330(.A1(new_n378), .A2(KEYINPUT86), .A3(new_n376), .A4(new_n379), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(KEYINPUT37), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n527), .A2(new_n383), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(new_n384), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n526), .A2(new_n536), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n459), .A2(new_n451), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT85), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n540), .B1(new_n438), .B2(new_n449), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n395), .B1(new_n541), .B2(new_n513), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n450), .A2(new_n451), .ZN(new_n543));
  OAI211_X1 g342(.A(new_n537), .B(new_n539), .C1(new_n542), .C2(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n518), .A2(new_n544), .A3(new_n495), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n497), .A2(new_n545), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n539), .B1(new_n542), .B2(new_n543), .ZN(new_n547));
  INV_X1    g346(.A(new_n388), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n489), .A2(KEYINPUT82), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n493), .A2(new_n491), .A3(new_n486), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n483), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n356), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n547), .A2(new_n548), .A3(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT35), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n349), .A2(new_n350), .ZN(new_n556));
  NOR3_X1   g355(.A1(new_n551), .A2(new_n556), .A3(new_n555), .ZN(new_n557));
  AOI22_X1  g356(.A1(new_n554), .A2(new_n555), .B1(new_n462), .B2(new_n557), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n263), .B1(new_n546), .B2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(G57gat), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n560), .A2(G64gat), .ZN(new_n561));
  XNOR2_X1  g360(.A(KEYINPUT92), .B(G57gat), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n561), .B1(new_n562), .B2(G64gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(G71gat), .A2(G78gat), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  NOR2_X1   g364(.A1(G71gat), .A2(G78gat), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n565), .B1(KEYINPUT9), .B2(new_n566), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n563), .A2(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(G57gat), .B(G64gat), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT9), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  OR2_X1    g370(.A1(new_n565), .A2(new_n566), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n568), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(KEYINPUT21), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(new_n208), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n576), .B(new_n308), .ZN(new_n577));
  NAND2_X1  g376(.A1(G231gat), .A2(G233gat), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n577), .B(new_n578), .ZN(new_n579));
  XOR2_X1   g378(.A(G127gat), .B(G155gat), .Z(new_n580));
  XNOR2_X1  g379(.A(new_n580), .B(KEYINPUT20), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  OR2_X1    g381(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n574), .A2(KEYINPUT21), .ZN(new_n584));
  XNOR2_X1  g383(.A(KEYINPUT93), .B(KEYINPUT19), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(G211gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n584), .B(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n579), .A2(new_n582), .ZN(new_n588));
  AND3_X1   g387(.A1(new_n583), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n587), .B1(new_n583), .B2(new_n588), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  AND2_X1   g390(.A1(G232gat), .A2(G233gat), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n592), .A2(KEYINPUT41), .ZN(new_n593));
  XNOR2_X1  g392(.A(G134gat), .B(G162gat), .ZN(new_n594));
  XOR2_X1   g393(.A(new_n593), .B(new_n594), .Z(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n238), .A2(KEYINPUT17), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n230), .A2(new_n231), .A3(new_n233), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(G85gat), .A2(G92gat), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n600), .A2(KEYINPUT7), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(KEYINPUT94), .ZN(new_n602));
  OAI21_X1  g401(.A(KEYINPUT95), .B1(new_n600), .B2(KEYINPUT7), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT95), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT7), .ZN(new_n605));
  NAND4_X1  g404(.A1(new_n604), .A2(new_n605), .A3(G85gat), .A4(G92gat), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT94), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n600), .A2(new_n607), .A3(KEYINPUT7), .ZN(new_n608));
  NAND4_X1  g407(.A1(new_n602), .A2(new_n603), .A3(new_n606), .A4(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(G99gat), .B(G106gat), .ZN(new_n610));
  NAND2_X1  g409(.A1(G99gat), .A2(G106gat), .ZN(new_n611));
  INV_X1    g410(.A(G85gat), .ZN(new_n612));
  INV_X1    g411(.A(G92gat), .ZN(new_n613));
  AOI22_X1  g412(.A1(KEYINPUT8), .A2(new_n611), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n609), .A2(new_n610), .A3(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n610), .B1(new_n609), .B2(new_n614), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  AOI22_X1  g418(.A1(new_n599), .A2(new_n619), .B1(KEYINPUT41), .B2(new_n592), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT96), .ZN(new_n621));
  XOR2_X1   g420(.A(G190gat), .B(G218gat), .Z(new_n622));
  NAND2_X1  g421(.A1(new_n238), .A2(new_n618), .ZN(new_n623));
  NAND4_X1  g422(.A1(new_n620), .A2(new_n621), .A3(new_n622), .A4(new_n623), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n619), .B1(new_n234), .B2(new_n235), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n592), .A2(KEYINPUT41), .ZN(new_n626));
  NAND4_X1  g425(.A1(new_n625), .A2(new_n622), .A3(new_n623), .A4(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n627), .A2(KEYINPUT96), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n624), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n625), .A2(new_n623), .A3(new_n626), .ZN(new_n630));
  INV_X1    g429(.A(new_n622), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT98), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n630), .A2(KEYINPUT98), .A3(new_n631), .ZN(new_n635));
  AND4_X1   g434(.A1(new_n596), .A2(new_n629), .A3(new_n634), .A4(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n629), .A2(KEYINPUT97), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT97), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n624), .A2(new_n638), .A3(new_n628), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n637), .A2(new_n639), .A3(new_n632), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n636), .B1(new_n595), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n591), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(G120gat), .B(G148gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(G176gat), .B(G204gat), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n643), .B(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(G230gat), .A2(G233gat), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n609), .A2(new_n614), .ZN(new_n648));
  INV_X1    g447(.A(new_n610), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  OR2_X1    g449(.A1(new_n610), .A2(KEYINPUT99), .ZN(new_n651));
  NAND4_X1  g450(.A1(new_n574), .A2(new_n650), .A3(new_n615), .A4(new_n651), .ZN(new_n652));
  OAI221_X1 g451(.A(new_n651), .B1(new_n571), .B2(new_n572), .C1(new_n563), .C2(new_n567), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n653), .B1(new_n616), .B2(new_n617), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT10), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n652), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n618), .A2(KEYINPUT10), .A3(new_n574), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n647), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n646), .B1(new_n652), .B2(new_n654), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n645), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n658), .A2(new_n659), .ZN(new_n661));
  INV_X1    g460(.A(new_n645), .ZN(new_n662));
  AOI21_X1  g461(.A(KEYINPUT100), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT100), .ZN(new_n664));
  NOR4_X1   g463(.A1(new_n658), .A2(new_n664), .A3(new_n659), .A4(new_n645), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n660), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT101), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  OAI211_X1 g467(.A(KEYINPUT101), .B(new_n660), .C1(new_n663), .C2(new_n665), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n642), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n559), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n460), .A2(new_n461), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(new_n203), .ZN(G1324gat));
  NOR2_X1   g474(.A1(new_n672), .A2(new_n548), .ZN(new_n676));
  NAND2_X1  g475(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n677));
  OR2_X1    g476(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n676), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT42), .ZN(new_n680));
  OR2_X1    g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n679), .A2(new_n680), .ZN(new_n682));
  OAI211_X1 g481(.A(new_n681), .B(new_n682), .C1(new_n207), .C2(new_n676), .ZN(G1325gat));
  INV_X1    g482(.A(G15gat), .ZN(new_n684));
  NOR3_X1   g483(.A1(new_n672), .A2(new_n684), .A3(new_n357), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n559), .A2(new_n671), .A3(new_n356), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n685), .B1(new_n684), .B2(new_n686), .ZN(G1326gat));
  NOR2_X1   g486(.A1(new_n672), .A2(new_n495), .ZN(new_n688));
  XOR2_X1   g487(.A(KEYINPUT43), .B(G22gat), .Z(new_n689));
  XNOR2_X1  g488(.A(new_n688), .B(new_n689), .ZN(G1327gat));
  INV_X1    g489(.A(new_n641), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n591), .A2(new_n670), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n559), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n224), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n693), .A2(new_n673), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g494(.A(KEYINPUT102), .B(KEYINPUT45), .ZN(new_n696));
  INV_X1    g495(.A(new_n696), .ZN(new_n697));
  OR2_X1    g496(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  AND3_X1   g497(.A1(new_n506), .A2(new_n498), .A3(new_n507), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n699), .A2(new_n508), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n510), .A2(new_n388), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n542), .A2(new_n701), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n551), .B1(new_n700), .B2(new_n702), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n496), .B1(new_n703), .B2(new_n544), .ZN(new_n704));
  AND2_X1   g503(.A1(new_n450), .A2(new_n451), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n538), .B1(new_n516), .B2(new_n705), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n495), .A2(new_n548), .A3(new_n356), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n555), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n557), .A2(new_n462), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n691), .B1(new_n704), .B2(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT44), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n546), .A2(new_n558), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n714), .A2(KEYINPUT44), .A3(new_n691), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n256), .A2(new_n258), .ZN(new_n716));
  NAND4_X1  g515(.A1(new_n713), .A2(new_n715), .A3(new_n716), .A4(new_n692), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n694), .B1(new_n717), .B2(new_n673), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n695), .A2(new_n697), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n698), .A2(new_n718), .A3(new_n719), .ZN(G1328gat));
  OAI21_X1  g519(.A(G36gat), .B1(new_n717), .B2(new_n548), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT46), .ZN(new_n722));
  NOR3_X1   g521(.A1(new_n693), .A2(G36gat), .A3(new_n548), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT103), .ZN(new_n724));
  AND3_X1   g523(.A1(new_n723), .A2(new_n724), .A3(new_n722), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n724), .B1(new_n723), .B2(new_n722), .ZN(new_n726));
  OAI221_X1 g525(.A(new_n721), .B1(new_n722), .B2(new_n723), .C1(new_n725), .C2(new_n726), .ZN(G1329gat));
  OAI21_X1  g526(.A(G43gat), .B1(new_n717), .B2(new_n357), .ZN(new_n728));
  OR2_X1    g527(.A1(new_n552), .A2(G43gat), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n728), .B1(new_n693), .B2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT47), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n730), .B(new_n731), .ZN(G1330gat));
  OAI21_X1  g531(.A(G50gat), .B1(new_n717), .B2(new_n495), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(KEYINPUT104), .ZN(new_n734));
  OR3_X1    g533(.A1(new_n693), .A2(G50gat), .A3(new_n495), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n734), .A2(new_n736), .A3(KEYINPUT48), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT48), .ZN(new_n738));
  OAI211_X1 g537(.A(new_n733), .B(new_n735), .C1(KEYINPUT104), .C2(new_n738), .ZN(new_n739));
  AND2_X1   g538(.A1(new_n737), .A2(new_n739), .ZN(G1331gat));
  AOI21_X1  g539(.A(new_n642), .B1(new_n546), .B2(new_n558), .ZN(new_n741));
  INV_X1    g540(.A(new_n670), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n742), .A2(new_n716), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n744), .A2(new_n673), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(new_n562), .ZN(G1332gat));
  INV_X1    g545(.A(new_n744), .ZN(new_n747));
  NAND2_X1  g546(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n747), .A2(new_n388), .A3(new_n748), .ZN(new_n749));
  OR2_X1    g548(.A1(new_n749), .A2(KEYINPUT105), .ZN(new_n750));
  NOR2_X1   g549(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n749), .A2(KEYINPUT105), .ZN(new_n752));
  AND3_X1   g551(.A1(new_n750), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n751), .B1(new_n750), .B2(new_n752), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n753), .A2(new_n754), .ZN(G1333gat));
  OAI21_X1  g554(.A(G71gat), .B1(new_n744), .B2(new_n357), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n356), .A2(new_n265), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n756), .B1(new_n744), .B2(new_n757), .ZN(new_n758));
  XOR2_X1   g557(.A(new_n758), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g558(.A1(new_n744), .A2(new_n495), .ZN(new_n760));
  XOR2_X1   g559(.A(KEYINPUT106), .B(G78gat), .Z(new_n761));
  XNOR2_X1  g560(.A(new_n760), .B(new_n761), .ZN(G1335gat));
  INV_X1    g561(.A(new_n591), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n713), .A2(new_n715), .A3(new_n763), .A4(new_n743), .ZN(new_n764));
  NOR3_X1   g563(.A1(new_n764), .A2(new_n612), .A3(new_n673), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n591), .A2(new_n716), .ZN(new_n766));
  OAI211_X1 g565(.A(new_n691), .B(new_n766), .C1(new_n704), .C2(new_n710), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT51), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n714), .A2(KEYINPUT51), .A3(new_n691), .A4(new_n766), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n771), .A2(new_n461), .A3(new_n460), .A4(new_n670), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n765), .B1(new_n612), .B2(new_n772), .ZN(G1336gat));
  NAND3_X1  g572(.A1(new_n769), .A2(KEYINPUT108), .A3(new_n770), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT108), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n767), .A2(new_n775), .A3(new_n768), .ZN(new_n776));
  NOR3_X1   g575(.A1(new_n742), .A2(G92gat), .A3(new_n548), .ZN(new_n777));
  XOR2_X1   g576(.A(new_n777), .B(KEYINPUT107), .Z(new_n778));
  NAND3_X1  g577(.A1(new_n774), .A2(new_n776), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(KEYINPUT109), .ZN(new_n780));
  OAI21_X1  g579(.A(G92gat), .B1(new_n764), .B2(new_n548), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT109), .ZN(new_n782));
  NAND4_X1  g581(.A1(new_n774), .A2(new_n782), .A3(new_n776), .A4(new_n778), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n780), .A2(new_n781), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(KEYINPUT52), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT52), .ZN(new_n786));
  AND3_X1   g585(.A1(new_n771), .A2(KEYINPUT110), .A3(new_n777), .ZN(new_n787));
  AOI21_X1  g586(.A(KEYINPUT110), .B1(new_n771), .B2(new_n777), .ZN(new_n788));
  OAI211_X1 g587(.A(new_n786), .B(new_n781), .C1(new_n787), .C2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n785), .A2(new_n789), .ZN(G1337gat));
  XNOR2_X1  g589(.A(KEYINPUT111), .B(G99gat), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n791), .B1(new_n764), .B2(new_n357), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n552), .A2(new_n791), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n771), .A2(new_n670), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n792), .A2(new_n794), .ZN(G1338gat));
  OAI21_X1  g594(.A(G106gat), .B1(new_n764), .B2(new_n495), .ZN(new_n796));
  NOR3_X1   g595(.A1(new_n742), .A2(new_n495), .A3(G106gat), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n774), .A2(new_n776), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(KEYINPUT53), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n771), .A2(new_n797), .ZN(new_n801));
  XNOR2_X1  g600(.A(KEYINPUT112), .B(KEYINPUT53), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n796), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n800), .A2(new_n803), .ZN(G1339gat));
  NOR3_X1   g603(.A1(new_n642), .A2(new_n670), .A3(new_n716), .ZN(new_n805));
  INV_X1    g604(.A(new_n805), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n244), .A2(new_n245), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n240), .B1(new_n236), .B2(new_n239), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n253), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n258), .A2(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(new_n658), .ZN(new_n812));
  INV_X1    g611(.A(new_n659), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n812), .A2(new_n813), .A3(new_n662), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(new_n664), .ZN(new_n815));
  INV_X1    g614(.A(new_n665), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT55), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT54), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n662), .B1(new_n658), .B2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n656), .A2(new_n647), .A3(new_n657), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(KEYINPUT54), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n823), .A2(new_n658), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n818), .B1(new_n821), .B2(new_n824), .ZN(new_n825));
  OAI211_X1 g624(.A(new_n820), .B(KEYINPUT55), .C1(new_n658), .C2(new_n823), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n817), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n691), .A2(new_n811), .A3(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(new_n829), .ZN(new_n830));
  AOI22_X1  g629(.A1(new_n670), .A2(new_n811), .B1(new_n828), .B2(new_n716), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n831), .A2(new_n691), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n763), .B1(new_n830), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n806), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n673), .A2(new_n388), .ZN(new_n835));
  AND2_X1   g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(new_n553), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT113), .ZN(new_n838));
  XNOR2_X1  g637(.A(new_n837), .B(new_n838), .ZN(new_n839));
  OAI21_X1  g638(.A(G113gat), .B1(new_n839), .B2(new_n263), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n551), .A2(new_n556), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n836), .A2(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(new_n716), .ZN(new_n843));
  OR3_X1    g642(.A1(new_n842), .A2(G113gat), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n840), .A2(new_n844), .ZN(G1340gat));
  OAI21_X1  g644(.A(G120gat), .B1(new_n839), .B2(new_n742), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n742), .A2(G120gat), .ZN(new_n847));
  XNOR2_X1  g646(.A(new_n847), .B(KEYINPUT114), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n846), .B1(new_n842), .B2(new_n848), .ZN(G1341gat));
  INV_X1    g648(.A(G127gat), .ZN(new_n850));
  NOR3_X1   g649(.A1(new_n839), .A2(new_n850), .A3(new_n763), .ZN(new_n851));
  INV_X1    g650(.A(new_n842), .ZN(new_n852));
  AOI21_X1  g651(.A(G127gat), .B1(new_n852), .B2(new_n591), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n851), .A2(new_n853), .ZN(G1342gat));
  NOR3_X1   g653(.A1(new_n842), .A2(G134gat), .A3(new_n641), .ZN(new_n855));
  XNOR2_X1  g654(.A(new_n855), .B(KEYINPUT56), .ZN(new_n856));
  OAI21_X1  g655(.A(G134gat), .B1(new_n839), .B2(new_n641), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(G1343gat));
  XOR2_X1   g657(.A(KEYINPUT115), .B(KEYINPUT55), .Z(new_n859));
  OAI21_X1  g658(.A(new_n859), .B1(new_n821), .B2(new_n824), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n817), .A2(new_n860), .A3(new_n826), .ZN(new_n861));
  NOR3_X1   g660(.A1(new_n260), .A2(new_n861), .A3(new_n261), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n810), .B1(new_n668), .B2(new_n669), .ZN(new_n863));
  NOR3_X1   g662(.A1(new_n862), .A2(new_n863), .A3(KEYINPUT116), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT116), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n670), .A2(new_n811), .ZN(new_n866));
  AND3_X1   g665(.A1(new_n817), .A2(new_n860), .A3(new_n826), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n716), .A2(KEYINPUT91), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n867), .A2(new_n868), .A3(new_n259), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n865), .B1(new_n866), .B2(new_n869), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n641), .B1(new_n864), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n591), .B1(new_n871), .B2(new_n829), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n551), .B1(new_n872), .B2(new_n805), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(KEYINPUT57), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n835), .A2(new_n357), .ZN(new_n875));
  INV_X1    g674(.A(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT57), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n834), .A2(new_n877), .A3(new_n551), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n874), .A2(new_n876), .A3(new_n878), .ZN(new_n879));
  OAI21_X1  g678(.A(G141gat), .B1(new_n879), .B2(new_n263), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT58), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n357), .A2(new_n551), .ZN(new_n882));
  OAI211_X1 g681(.A(new_n834), .B(new_n835), .C1(KEYINPUT117), .C2(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n883), .B1(KEYINPUT117), .B2(new_n882), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n884), .A2(new_n399), .A3(new_n262), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n880), .A2(new_n881), .A3(new_n885), .ZN(new_n886));
  OAI21_X1  g685(.A(G141gat), .B1(new_n879), .B2(new_n843), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n887), .A2(new_n885), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n886), .B1(new_n888), .B2(new_n881), .ZN(G1344gat));
  AOI21_X1  g688(.A(new_n877), .B1(new_n834), .B2(new_n551), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT119), .ZN(new_n891));
  OAI21_X1  g690(.A(KEYINPUT116), .B1(new_n862), .B2(new_n863), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n866), .A2(new_n869), .A3(new_n865), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n691), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  OAI21_X1  g693(.A(KEYINPUT118), .B1(new_n641), .B2(new_n827), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT118), .ZN(new_n896));
  AOI22_X1  g695(.A1(new_n629), .A2(KEYINPUT97), .B1(new_n631), .B2(new_n630), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n596), .B1(new_n897), .B2(new_n639), .ZN(new_n898));
  OAI211_X1 g697(.A(new_n828), .B(new_n896), .C1(new_n898), .C2(new_n636), .ZN(new_n899));
  AND3_X1   g698(.A1(new_n895), .A2(new_n899), .A3(new_n811), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n891), .B1(new_n894), .B2(new_n900), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n895), .A2(new_n899), .A3(new_n811), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n871), .A2(KEYINPUT119), .A3(new_n902), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n901), .A2(new_n903), .A3(new_n763), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n671), .A2(new_n263), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n495), .A2(KEYINPUT57), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n890), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n908), .A2(new_n670), .A3(new_n876), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n909), .A2(KEYINPUT59), .A3(G148gat), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n396), .A2(new_n397), .ZN(new_n911));
  INV_X1    g710(.A(new_n911), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n884), .A2(new_n912), .A3(new_n670), .ZN(new_n913));
  INV_X1    g712(.A(new_n879), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n912), .B1(new_n914), .B2(new_n670), .ZN(new_n915));
  OAI211_X1 g714(.A(new_n910), .B(new_n913), .C1(new_n915), .C2(KEYINPUT59), .ZN(G1345gat));
  AOI21_X1  g715(.A(G155gat), .B1(new_n884), .B2(new_n591), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n591), .A2(G155gat), .ZN(new_n918));
  XNOR2_X1  g717(.A(new_n918), .B(KEYINPUT120), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n917), .B1(new_n914), .B2(new_n919), .ZN(G1346gat));
  OAI21_X1  g719(.A(G162gat), .B1(new_n879), .B2(new_n641), .ZN(new_n921));
  INV_X1    g720(.A(G162gat), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n884), .A2(new_n922), .A3(new_n691), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT121), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n921), .A2(KEYINPUT121), .A3(new_n923), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(G1347gat));
  NAND2_X1  g727(.A1(new_n673), .A2(new_n388), .ZN(new_n929));
  INV_X1    g728(.A(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(new_n832), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n591), .B1(new_n931), .B2(new_n829), .ZN(new_n932));
  OAI211_X1 g731(.A(new_n553), .B(new_n930), .C1(new_n932), .C2(new_n805), .ZN(new_n933));
  OAI21_X1  g732(.A(G169gat), .B1(new_n933), .B2(new_n263), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n929), .B1(new_n806), .B2(new_n833), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(new_n841), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n716), .A2(new_n293), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n934), .B1(new_n936), .B2(new_n937), .ZN(G1348gat));
  NOR3_X1   g737(.A1(new_n933), .A2(new_n294), .A3(new_n742), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n935), .A2(new_n670), .A3(new_n841), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n939), .B1(new_n294), .B2(new_n940), .ZN(G1349gat));
  OAI21_X1  g740(.A(G183gat), .B1(new_n933), .B2(new_n763), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n591), .A2(new_n290), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n942), .B1(new_n936), .B2(new_n943), .ZN(new_n944));
  XNOR2_X1  g743(.A(new_n944), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g744(.A(G190gat), .B1(new_n933), .B2(new_n641), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT123), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  OAI211_X1 g747(.A(KEYINPUT123), .B(G190gat), .C1(new_n933), .C2(new_n641), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n948), .A2(KEYINPUT61), .A3(new_n949), .ZN(new_n950));
  NAND4_X1  g749(.A1(new_n935), .A2(new_n285), .A3(new_n691), .A4(new_n841), .ZN(new_n951));
  XNOR2_X1  g750(.A(new_n951), .B(KEYINPUT122), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT61), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n946), .A2(new_n947), .A3(new_n953), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n950), .A2(new_n952), .A3(new_n954), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT124), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND4_X1  g756(.A1(new_n950), .A2(new_n952), .A3(KEYINPUT124), .A4(new_n954), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(G1351gat));
  NAND2_X1  g758(.A1(new_n930), .A2(new_n357), .ZN(new_n960));
  INV_X1    g759(.A(new_n960), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n908), .A2(new_n262), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n962), .A2(KEYINPUT125), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT125), .ZN(new_n964));
  NAND4_X1  g763(.A1(new_n908), .A2(new_n964), .A3(new_n262), .A4(new_n961), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n963), .A2(G197gat), .A3(new_n965), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n935), .A2(new_n551), .A3(new_n357), .ZN(new_n967));
  INV_X1    g766(.A(new_n967), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n968), .A2(new_n250), .A3(new_n716), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n966), .A2(new_n969), .ZN(G1352gat));
  INV_X1    g769(.A(G204gat), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n968), .A2(new_n971), .A3(new_n670), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n972), .A2(KEYINPUT126), .A3(KEYINPUT62), .ZN(new_n973));
  NAND2_X1  g772(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n974));
  NOR3_X1   g773(.A1(new_n967), .A2(G204gat), .A3(new_n742), .ZN(new_n975));
  NOR2_X1   g774(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n974), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  INV_X1    g776(.A(new_n907), .ZN(new_n978));
  AOI21_X1  g777(.A(new_n978), .B1(new_n904), .B2(new_n905), .ZN(new_n979));
  NOR4_X1   g778(.A1(new_n979), .A2(new_n742), .A3(new_n890), .A4(new_n960), .ZN(new_n980));
  OAI211_X1 g779(.A(new_n973), .B(new_n977), .C1(new_n971), .C2(new_n980), .ZN(G1353gat));
  NAND3_X1  g780(.A1(new_n968), .A2(new_n365), .A3(new_n591), .ZN(new_n982));
  NAND3_X1  g781(.A1(new_n908), .A2(new_n591), .A3(new_n961), .ZN(new_n983));
  AND3_X1   g782(.A1(new_n983), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n984));
  AOI21_X1  g783(.A(KEYINPUT63), .B1(new_n983), .B2(G211gat), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n982), .B1(new_n984), .B2(new_n985), .ZN(G1354gat));
  NAND3_X1  g785(.A1(new_n968), .A2(new_n366), .A3(new_n691), .ZN(new_n987));
  INV_X1    g786(.A(KEYINPUT127), .ZN(new_n988));
  AOI21_X1  g787(.A(new_n988), .B1(new_n908), .B2(new_n961), .ZN(new_n989));
  NOR4_X1   g788(.A1(new_n979), .A2(KEYINPUT127), .A3(new_n890), .A4(new_n960), .ZN(new_n990));
  NOR3_X1   g789(.A1(new_n989), .A2(new_n990), .A3(new_n641), .ZN(new_n991));
  OAI21_X1  g790(.A(new_n987), .B1(new_n991), .B2(new_n366), .ZN(G1355gat));
endmodule


