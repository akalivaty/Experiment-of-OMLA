//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 1 0 1 0 0 0 0 1 0 0 1 0 0 0 1 0 0 0 1 1 0 1 0 1 0 0 1 1 0 1 0 1 1 1 0 1 1 0 0 1 1 0 0 1 0 0 0 1 1 1 0 1 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n765, new_n766, new_n767, new_n768, new_n770, new_n771,
    new_n772, new_n773, new_n775, new_n776, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n811, new_n812, new_n813, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n861, new_n862,
    new_n863, new_n865, new_n866, new_n867, new_n868, new_n870, new_n871,
    new_n872, new_n873, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n917, new_n918, new_n920, new_n921, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n932, new_n933, new_n934,
    new_n936, new_n937, new_n938, new_n939, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n962, new_n963;
  INV_X1    g000(.A(G50gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(G43gat), .ZN(new_n203));
  INV_X1    g002(.A(G43gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G50gat), .ZN(new_n205));
  AND3_X1   g004(.A1(new_n203), .A2(new_n205), .A3(KEYINPUT15), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT86), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n203), .A2(new_n205), .A3(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT15), .ZN(new_n209));
  OAI211_X1 g008(.A(new_n208), .B(new_n209), .C1(new_n207), .C2(new_n205), .ZN(new_n210));
  INV_X1    g009(.A(G29gat), .ZN(new_n211));
  AND2_X1   g010(.A1(new_n211), .A2(KEYINPUT14), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(G36gat), .ZN(new_n213));
  INV_X1    g012(.A(G36gat), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n214), .B1(new_n211), .B2(KEYINPUT14), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n213), .B1(new_n215), .B2(new_n212), .ZN(new_n216));
  AOI21_X1  g015(.A(new_n206), .B1(new_n210), .B2(new_n216), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n217), .B1(new_n206), .B2(new_n216), .ZN(new_n218));
  XNOR2_X1  g017(.A(G15gat), .B(G22gat), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT16), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n219), .B1(new_n220), .B2(G1gat), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n221), .B1(G1gat), .B2(new_n219), .ZN(new_n222));
  XNOR2_X1  g021(.A(new_n222), .B(G8gat), .ZN(new_n223));
  AND2_X1   g022(.A1(new_n218), .A2(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(new_n218), .B(KEYINPUT17), .ZN(new_n225));
  INV_X1    g024(.A(new_n223), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n224), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(G229gat), .A2(G233gat), .ZN(new_n228));
  AND2_X1   g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OR2_X1    g028(.A1(new_n229), .A2(KEYINPUT18), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(KEYINPUT18), .ZN(new_n231));
  XNOR2_X1  g030(.A(new_n218), .B(new_n223), .ZN(new_n232));
  XOR2_X1   g031(.A(new_n228), .B(KEYINPUT13), .Z(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n230), .A2(new_n231), .A3(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(G113gat), .B(G141gat), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n236), .B(G197gat), .ZN(new_n237));
  XOR2_X1   g036(.A(KEYINPUT11), .B(G169gat), .Z(new_n238));
  XNOR2_X1  g037(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g038(.A(new_n239), .B(KEYINPUT12), .Z(new_n240));
  NAND2_X1  g039(.A1(new_n235), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(new_n240), .ZN(new_n242));
  NAND4_X1  g041(.A1(new_n230), .A2(new_n242), .A3(new_n231), .A4(new_n234), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT73), .ZN(new_n246));
  XOR2_X1   g045(.A(G141gat), .B(G148gat), .Z(new_n247));
  INV_X1    g046(.A(G155gat), .ZN(new_n248));
  INV_X1    g047(.A(G162gat), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(G155gat), .A2(G162gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(KEYINPUT2), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n247), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  XNOR2_X1  g053(.A(G141gat), .B(G148gat), .ZN(new_n255));
  AND2_X1   g054(.A1(KEYINPUT72), .A2(KEYINPUT2), .ZN(new_n256));
  NOR2_X1   g055(.A1(KEYINPUT72), .A2(KEYINPUT2), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n255), .B1(new_n251), .B2(new_n258), .ZN(new_n259));
  AND2_X1   g058(.A1(G155gat), .A2(G162gat), .ZN(new_n260));
  NOR2_X1   g059(.A1(G155gat), .A2(G162gat), .ZN(new_n261));
  OAI21_X1  g060(.A(KEYINPUT71), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT71), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n250), .A2(new_n263), .A3(new_n251), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n254), .B1(new_n259), .B2(new_n265), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n246), .B1(new_n266), .B2(KEYINPUT3), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n266), .A2(new_n246), .A3(KEYINPUT3), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT3), .ZN(new_n270));
  OAI211_X1 g069(.A(new_n270), .B(new_n254), .C1(new_n259), .C2(new_n265), .ZN(new_n271));
  XNOR2_X1  g070(.A(G127gat), .B(G134gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(G113gat), .A2(G120gat), .ZN(new_n273));
  INV_X1    g072(.A(G113gat), .ZN(new_n274));
  INV_X1    g073(.A(G120gat), .ZN(new_n275));
  AOI21_X1  g074(.A(KEYINPUT1), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n272), .A2(new_n273), .A3(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(G127gat), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n278), .A2(G134gat), .ZN(new_n279));
  INV_X1    g078(.A(G134gat), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n280), .A2(G127gat), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT1), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n282), .B1(G113gat), .B2(G120gat), .ZN(new_n283));
  INV_X1    g082(.A(new_n273), .ZN(new_n284));
  OAI22_X1  g083(.A1(new_n279), .A2(new_n281), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n277), .A2(new_n285), .ZN(new_n286));
  AND2_X1   g085(.A1(new_n271), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n268), .A2(new_n269), .A3(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT4), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n289), .B1(new_n266), .B2(new_n286), .ZN(new_n290));
  OAI21_X1  g089(.A(KEYINPUT74), .B1(new_n266), .B2(new_n286), .ZN(new_n291));
  INV_X1    g090(.A(new_n286), .ZN(new_n292));
  NOR3_X1   g091(.A1(new_n260), .A2(new_n256), .A3(new_n257), .ZN(new_n293));
  OAI211_X1 g092(.A(new_n262), .B(new_n264), .C1(new_n293), .C2(new_n255), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT74), .ZN(new_n295));
  NAND4_X1  g094(.A1(new_n292), .A2(new_n294), .A3(new_n295), .A4(new_n254), .ZN(new_n296));
  AND2_X1   g095(.A1(new_n291), .A2(new_n296), .ZN(new_n297));
  OAI211_X1 g096(.A(new_n288), .B(new_n290), .C1(new_n297), .C2(new_n289), .ZN(new_n298));
  AND2_X1   g097(.A1(G225gat), .A2(G233gat), .ZN(new_n299));
  NOR3_X1   g098(.A1(new_n298), .A2(KEYINPUT5), .A3(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT76), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n266), .A2(new_n286), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n291), .A2(new_n296), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(new_n299), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(KEYINPUT5), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(KEYINPUT75), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT75), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n305), .A2(new_n308), .A3(KEYINPUT5), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n297), .A2(new_n289), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n266), .A2(new_n286), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n299), .B1(new_n312), .B2(KEYINPUT4), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n311), .A2(new_n288), .A3(new_n313), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n302), .B1(new_n310), .B2(new_n314), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n308), .B1(new_n305), .B2(KEYINPUT5), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT5), .ZN(new_n317));
  AOI211_X1 g116(.A(KEYINPUT75), .B(new_n317), .C1(new_n304), .C2(new_n299), .ZN(new_n318));
  OAI211_X1 g117(.A(new_n302), .B(new_n314), .C1(new_n316), .C2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n301), .B1(new_n315), .B2(new_n320), .ZN(new_n321));
  XOR2_X1   g120(.A(G1gat), .B(G29gat), .Z(new_n322));
  XNOR2_X1  g121(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n323));
  XNOR2_X1  g122(.A(new_n322), .B(new_n323), .ZN(new_n324));
  XNOR2_X1  g123(.A(G57gat), .B(G85gat), .ZN(new_n325));
  XNOR2_X1  g124(.A(new_n324), .B(new_n325), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n321), .A2(KEYINPUT6), .A3(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT6), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n314), .B1(new_n316), .B2(new_n318), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(KEYINPUT76), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n300), .B1(new_n330), .B2(new_n319), .ZN(new_n331));
  INV_X1    g130(.A(new_n326), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n328), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  AOI211_X1 g132(.A(new_n326), .B(new_n300), .C1(new_n330), .C2(new_n319), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n327), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT84), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n327), .A2(KEYINPUT84), .ZN(new_n338));
  AOI21_X1  g137(.A(KEYINPUT35), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT28), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT66), .ZN(new_n341));
  XNOR2_X1  g140(.A(KEYINPUT27), .B(G183gat), .ZN(new_n342));
  INV_X1    g141(.A(G190gat), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n341), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(G183gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(KEYINPUT27), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT27), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(G183gat), .ZN(new_n348));
  AND4_X1   g147(.A1(new_n341), .A2(new_n346), .A3(new_n348), .A4(new_n343), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n340), .B1(new_n344), .B2(new_n349), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n346), .A2(new_n348), .A3(new_n343), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(KEYINPUT66), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n342), .A2(new_n341), .A3(new_n343), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n352), .A2(new_n353), .A3(KEYINPUT28), .ZN(new_n354));
  INV_X1    g153(.A(G169gat), .ZN(new_n355));
  INV_X1    g154(.A(G176gat), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NOR2_X1   g156(.A1(G169gat), .A2(G176gat), .ZN(new_n358));
  NOR3_X1   g157(.A1(new_n357), .A2(KEYINPUT26), .A3(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(G183gat), .A2(G190gat), .ZN(new_n360));
  INV_X1    g159(.A(new_n358), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT26), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n360), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n359), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n350), .A2(new_n354), .A3(new_n364), .ZN(new_n365));
  XNOR2_X1  g164(.A(KEYINPUT64), .B(KEYINPUT23), .ZN(new_n366));
  OAI21_X1  g165(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(new_n360), .ZN(new_n368));
  NAND3_X1  g167(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n369));
  AOI22_X1  g168(.A1(new_n361), .A2(new_n366), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT65), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n357), .B1(KEYINPUT23), .B2(new_n358), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n370), .A2(new_n371), .A3(KEYINPUT25), .A4(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n368), .A2(new_n369), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT23), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(KEYINPUT64), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT64), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(KEYINPUT23), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n361), .A2(new_n377), .A3(new_n379), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n375), .A2(KEYINPUT65), .A3(new_n380), .ZN(new_n381));
  AOI22_X1  g180(.A1(KEYINPUT25), .A2(new_n381), .B1(new_n370), .B2(new_n372), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n365), .B1(new_n374), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(new_n286), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n381), .A2(KEYINPUT25), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n370), .A2(new_n372), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(new_n373), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n388), .A2(new_n292), .A3(new_n365), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n384), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n390), .A2(G227gat), .A3(G233gat), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT33), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  XOR2_X1   g192(.A(G15gat), .B(G43gat), .Z(new_n394));
  XNOR2_X1  g193(.A(G71gat), .B(G99gat), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n394), .B(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n393), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(G227gat), .A2(G233gat), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n384), .A2(new_n398), .A3(new_n389), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(KEYINPUT34), .ZN(new_n400));
  OR2_X1    g199(.A1(new_n399), .A2(KEYINPUT34), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n397), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  AND2_X1   g201(.A1(new_n391), .A2(KEYINPUT32), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n401), .A2(new_n400), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n404), .A2(new_n393), .A3(new_n396), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n402), .A2(new_n403), .A3(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n403), .B1(new_n402), .B2(new_n405), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  XNOR2_X1  g208(.A(KEYINPUT31), .B(G50gat), .ZN(new_n410));
  XOR2_X1   g209(.A(new_n410), .B(G106gat), .Z(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(G22gat), .ZN(new_n413));
  NAND2_X1  g212(.A1(G228gat), .A2(G233gat), .ZN(new_n414));
  AOI21_X1  g213(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n415));
  NOR2_X1   g214(.A1(G197gat), .A2(G204gat), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(G197gat), .A2(G204gat), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n415), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(G211gat), .ZN(new_n420));
  INV_X1    g219(.A(G218gat), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT79), .ZN(new_n423));
  NAND2_X1  g222(.A1(G211gat), .A2(G218gat), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n422), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(new_n424), .ZN(new_n426));
  NOR2_X1   g225(.A1(G211gat), .A2(G218gat), .ZN(new_n427));
  OAI21_X1  g226(.A(KEYINPUT79), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n419), .A2(new_n425), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n422), .A2(new_n424), .ZN(new_n430));
  AND2_X1   g229(.A1(G197gat), .A2(G204gat), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n431), .A2(new_n416), .ZN(new_n432));
  OAI211_X1 g231(.A(KEYINPUT79), .B(new_n430), .C1(new_n432), .C2(new_n415), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT29), .ZN(new_n434));
  AND3_X1   g233(.A1(new_n429), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n266), .B1(new_n435), .B2(KEYINPUT3), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n422), .A2(KEYINPUT67), .A3(new_n424), .ZN(new_n437));
  XNOR2_X1  g236(.A(new_n419), .B(new_n437), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n438), .B1(new_n271), .B2(new_n434), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT80), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n436), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  AOI211_X1 g240(.A(KEYINPUT80), .B(new_n438), .C1(new_n434), .C2(new_n271), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n414), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT81), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  OAI211_X1 g244(.A(KEYINPUT81), .B(new_n414), .C1(new_n441), .C2(new_n442), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n438), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n270), .B1(new_n448), .B2(KEYINPUT29), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n414), .B1(new_n449), .B2(new_n266), .ZN(new_n450));
  INV_X1    g249(.A(new_n271), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n448), .B1(new_n451), .B2(KEYINPUT29), .ZN(new_n452));
  AND2_X1   g251(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n413), .B1(new_n447), .B2(new_n454), .ZN(new_n455));
  AOI211_X1 g254(.A(G22gat), .B(new_n453), .C1(new_n445), .C2(new_n446), .ZN(new_n456));
  NOR3_X1   g255(.A1(new_n455), .A2(new_n456), .A3(G78gat), .ZN(new_n457));
  INV_X1    g256(.A(G78gat), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n452), .A2(KEYINPUT80), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n439), .A2(new_n440), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n459), .A2(new_n460), .A3(new_n436), .ZN(new_n461));
  AOI21_X1  g260(.A(KEYINPUT81), .B1(new_n461), .B2(new_n414), .ZN(new_n462));
  INV_X1    g261(.A(new_n446), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n454), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(G22gat), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n447), .A2(new_n413), .A3(new_n454), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n458), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n412), .B1(new_n457), .B2(new_n467), .ZN(new_n468));
  OAI21_X1  g267(.A(G78gat), .B1(new_n455), .B2(new_n456), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n465), .A2(new_n458), .A3(new_n466), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n469), .A2(new_n470), .A3(new_n411), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n409), .A2(new_n468), .A3(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT30), .ZN(new_n473));
  XOR2_X1   g272(.A(G8gat), .B(G36gat), .Z(new_n474));
  XNOR2_X1  g273(.A(G64gat), .B(G92gat), .ZN(new_n475));
  XNOR2_X1  g274(.A(new_n474), .B(new_n475), .ZN(new_n476));
  XOR2_X1   g275(.A(new_n476), .B(KEYINPUT70), .Z(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(G226gat), .ZN(new_n479));
  INV_X1    g278(.A(G233gat), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n481), .A2(KEYINPUT29), .ZN(new_n482));
  INV_X1    g281(.A(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT68), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n383), .A2(new_n484), .ZN(new_n485));
  OAI211_X1 g284(.A(KEYINPUT68), .B(new_n365), .C1(new_n374), .C2(new_n382), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n483), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n388), .A2(new_n481), .A3(new_n365), .ZN(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  OAI211_X1 g288(.A(KEYINPUT69), .B(new_n438), .C1(new_n487), .C2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n383), .A2(new_n482), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n485), .A2(new_n486), .ZN(new_n492));
  INV_X1    g291(.A(new_n481), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n448), .B(new_n491), .C1(new_n492), .C2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n490), .A2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(new_n486), .ZN(new_n496));
  AOI21_X1  g295(.A(KEYINPUT68), .B1(new_n388), .B2(new_n365), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n482), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(new_n488), .ZN(new_n499));
  AOI21_X1  g298(.A(KEYINPUT69), .B1(new_n499), .B2(new_n438), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n478), .B1(new_n495), .B2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT69), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n489), .B1(new_n492), .B2(new_n482), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n502), .B1(new_n503), .B2(new_n448), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n504), .A2(new_n476), .A3(new_n490), .A4(new_n494), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n473), .B1(new_n501), .B2(new_n505), .ZN(new_n506));
  AND2_X1   g305(.A1(new_n505), .A2(new_n473), .ZN(new_n507));
  OR2_X1    g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n472), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n339), .A2(new_n509), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n506), .A2(new_n507), .ZN(new_n511));
  AND3_X1   g310(.A1(new_n335), .A2(KEYINPUT78), .A3(new_n511), .ZN(new_n512));
  AOI21_X1  g311(.A(KEYINPUT78), .B1(new_n335), .B2(new_n511), .ZN(new_n513));
  NOR3_X1   g312(.A1(new_n512), .A2(new_n513), .A3(new_n472), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT35), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n510), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n495), .A2(new_n500), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT37), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n504), .A2(new_n490), .A3(new_n494), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n476), .B1(new_n520), .B2(KEYINPUT37), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n519), .B1(new_n521), .B2(KEYINPUT85), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT85), .ZN(new_n523));
  AOI211_X1 g322(.A(new_n523), .B(new_n476), .C1(new_n520), .C2(KEYINPUT37), .ZN(new_n524));
  OAI21_X1  g323(.A(KEYINPUT38), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n518), .B1(new_n499), .B2(new_n448), .ZN(new_n526));
  OAI211_X1 g325(.A(new_n438), .B(new_n491), .C1(new_n492), .C2(new_n493), .ZN(new_n527));
  AOI211_X1 g326(.A(KEYINPUT38), .B(new_n477), .C1(new_n526), .C2(new_n527), .ZN(new_n528));
  AOI22_X1  g327(.A1(new_n519), .A2(new_n528), .B1(new_n476), .B2(new_n517), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n337), .A2(new_n525), .A3(new_n338), .A4(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n468), .A2(new_n471), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT39), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n288), .A2(new_n290), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n297), .A2(new_n289), .ZN(new_n534));
  OAI211_X1 g333(.A(new_n532), .B(new_n299), .C1(new_n533), .C2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(new_n332), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT82), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n535), .A2(KEYINPUT82), .A3(new_n332), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n298), .A2(new_n299), .ZN(new_n540));
  OAI211_X1 g339(.A(new_n540), .B(KEYINPUT39), .C1(new_n299), .C2(new_n304), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n538), .A2(new_n539), .A3(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT40), .ZN(new_n543));
  AND3_X1   g342(.A1(new_n542), .A2(KEYINPUT83), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n543), .B1(new_n542), .B2(KEYINPUT83), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n331), .A2(new_n332), .ZN(new_n546));
  NOR3_X1   g345(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n531), .B1(new_n508), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n530), .A2(new_n548), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n531), .B1(new_n512), .B2(new_n513), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n409), .B(KEYINPUT36), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n245), .B1(new_n516), .B2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT97), .ZN(new_n554));
  NAND2_X1  g353(.A1(G230gat), .A2(G233gat), .ZN(new_n555));
  XOR2_X1   g354(.A(new_n555), .B(KEYINPUT96), .Z(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(G85gat), .A2(G92gat), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n558), .A2(KEYINPUT7), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(KEYINPUT91), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT92), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n561), .B1(new_n558), .B2(KEYINPUT7), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT7), .ZN(new_n563));
  NAND4_X1  g362(.A1(new_n563), .A2(KEYINPUT92), .A3(G85gat), .A4(G92gat), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT91), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n558), .A2(new_n565), .A3(KEYINPUT7), .ZN(new_n566));
  NAND4_X1  g365(.A1(new_n560), .A2(new_n562), .A3(new_n564), .A4(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(G99gat), .A2(G106gat), .ZN(new_n568));
  INV_X1    g367(.A(G85gat), .ZN(new_n569));
  INV_X1    g368(.A(G92gat), .ZN(new_n570));
  AOI22_X1  g369(.A1(KEYINPUT8), .A2(new_n568), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n567), .A2(new_n571), .ZN(new_n572));
  XOR2_X1   g371(.A(G99gat), .B(G106gat), .Z(new_n573));
  OR2_X1    g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT93), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n572), .A2(new_n573), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(G71gat), .B(G78gat), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n578), .A2(KEYINPUT87), .ZN(new_n579));
  AOI21_X1  g378(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n580));
  XNOR2_X1  g379(.A(G57gat), .B(G64gat), .ZN(new_n581));
  NOR3_X1   g380(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n578), .A2(KEYINPUT87), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  OAI211_X1 g383(.A(KEYINPUT87), .B(new_n578), .C1(new_n581), .C2(new_n580), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n572), .A2(KEYINPUT93), .A3(new_n573), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n577), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT10), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n586), .A2(new_n574), .A3(new_n576), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT94), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND4_X1  g393(.A1(new_n589), .A2(KEYINPUT94), .A3(new_n590), .A4(new_n591), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n577), .A2(new_n588), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n587), .A2(new_n590), .ZN(new_n597));
  AOI22_X1  g396(.A1(new_n594), .A2(new_n595), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n557), .B1(new_n598), .B2(KEYINPUT95), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n594), .A2(new_n595), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n597), .A2(new_n596), .ZN(new_n601));
  AND3_X1   g400(.A1(new_n600), .A2(KEYINPUT95), .A3(new_n601), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n554), .B1(new_n599), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n600), .A2(new_n601), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT95), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n598), .A2(KEYINPUT95), .ZN(new_n607));
  NAND4_X1  g406(.A1(new_n606), .A2(KEYINPUT97), .A3(new_n557), .A4(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n603), .A2(new_n608), .ZN(new_n609));
  XOR2_X1   g408(.A(G120gat), .B(G148gat), .Z(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(KEYINPUT98), .ZN(new_n611));
  XNOR2_X1  g410(.A(G176gat), .B(G204gat), .ZN(new_n612));
  XOR2_X1   g411(.A(new_n611), .B(new_n612), .Z(new_n613));
  NAND2_X1  g412(.A1(new_n589), .A2(new_n591), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n613), .B1(new_n614), .B2(new_n556), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n609), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT100), .ZN(new_n617));
  XOR2_X1   g416(.A(new_n556), .B(KEYINPUT99), .Z(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n604), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n614), .A2(new_n556), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n622), .A2(new_n613), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n616), .A2(new_n617), .A3(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n617), .B1(new_n616), .B2(new_n623), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n225), .A2(new_n588), .A3(new_n577), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n596), .A2(new_n218), .ZN(new_n630));
  NAND3_X1  g429(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n629), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(G190gat), .B(G218gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(G134gat), .B(G162gat), .ZN(new_n635));
  AOI21_X1  g434(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(new_n637));
  AND2_X1   g436(.A1(new_n634), .A2(new_n637), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n634), .A2(new_n637), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n223), .B1(KEYINPUT21), .B2(new_n586), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(KEYINPUT90), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n586), .A2(KEYINPUT21), .ZN(new_n643));
  XNOR2_X1  g442(.A(KEYINPUT89), .B(KEYINPUT19), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n642), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(G127gat), .B(G155gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(KEYINPUT20), .ZN(new_n648));
  NAND2_X1  g447(.A1(G231gat), .A2(G233gat), .ZN(new_n649));
  XOR2_X1   g448(.A(new_n649), .B(KEYINPUT88), .Z(new_n650));
  XNOR2_X1  g449(.A(new_n648), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(G183gat), .B(G211gat), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n651), .B(new_n652), .ZN(new_n653));
  OR2_X1    g452(.A1(new_n646), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n646), .A2(new_n653), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n640), .A2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n628), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n553), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  NOR3_X1   g460(.A1(new_n331), .A2(new_n328), .A3(new_n332), .ZN(new_n662));
  AOI21_X1  g461(.A(KEYINPUT6), .B1(new_n321), .B2(new_n326), .ZN(new_n663));
  INV_X1    g462(.A(new_n334), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n662), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n661), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(G1gat), .ZN(G1324gat));
  INV_X1    g466(.A(KEYINPUT42), .ZN(new_n668));
  XOR2_X1   g467(.A(KEYINPUT16), .B(G8gat), .Z(new_n669));
  NAND3_X1  g468(.A1(new_n661), .A2(new_n508), .A3(new_n669), .ZN(new_n670));
  OAI21_X1  g469(.A(G8gat), .B1(new_n660), .B2(new_n511), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n668), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n672), .B1(new_n668), .B2(new_n670), .ZN(new_n673));
  XOR2_X1   g472(.A(new_n673), .B(KEYINPUT101), .Z(G1325gat));
  OAI21_X1  g473(.A(G15gat), .B1(new_n660), .B2(new_n551), .ZN(new_n675));
  OR2_X1    g474(.A1(new_n407), .A2(new_n408), .ZN(new_n676));
  OR2_X1    g475(.A1(new_n676), .A2(G15gat), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n675), .B1(new_n660), .B2(new_n677), .ZN(G1326gat));
  NAND2_X1  g477(.A1(new_n661), .A2(new_n531), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(KEYINPUT102), .ZN(new_n680));
  XNOR2_X1  g479(.A(KEYINPUT43), .B(G22gat), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n680), .B(new_n681), .ZN(G1327gat));
  AND4_X1   g481(.A1(new_n553), .A2(new_n656), .A3(new_n640), .A4(new_n627), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n683), .A2(new_n211), .A3(new_n665), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(KEYINPUT45), .ZN(new_n685));
  AND3_X1   g484(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT78), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n687), .B1(new_n665), .B2(new_n508), .ZN(new_n688));
  INV_X1    g487(.A(new_n472), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n335), .A2(KEYINPUT78), .A3(new_n511), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n688), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  AOI22_X1  g490(.A1(new_n691), .A2(KEYINPUT35), .B1(new_n509), .B2(new_n339), .ZN(new_n692));
  OAI211_X1 g491(.A(KEYINPUT105), .B(new_n640), .C1(new_n686), .C2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT44), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(new_n640), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n696), .B1(new_n516), .B2(new_n552), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n697), .A2(KEYINPUT105), .A3(KEYINPUT44), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n244), .B(KEYINPUT103), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n656), .B(KEYINPUT104), .ZN(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  NOR3_X1   g500(.A1(new_n628), .A2(new_n699), .A3(new_n701), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n695), .A2(new_n698), .A3(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT106), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND4_X1  g504(.A1(new_n695), .A2(KEYINPUT106), .A3(new_n698), .A4(new_n702), .ZN(new_n706));
  AND3_X1   g505(.A1(new_n705), .A2(new_n665), .A3(new_n706), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n685), .B1(new_n707), .B2(new_n211), .ZN(G1328gat));
  INV_X1    g507(.A(KEYINPUT46), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n709), .A2(KEYINPUT108), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n683), .A2(new_n214), .A3(new_n508), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT107), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n710), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n713), .B1(new_n712), .B2(new_n711), .ZN(new_n714));
  AND2_X1   g513(.A1(new_n709), .A2(KEYINPUT108), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n714), .B(new_n715), .ZN(new_n716));
  AND3_X1   g515(.A1(new_n705), .A2(new_n508), .A3(new_n706), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n716), .B1(new_n214), .B2(new_n717), .ZN(G1329gat));
  NOR2_X1   g517(.A1(new_n676), .A2(G43gat), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n683), .A2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT47), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(new_n551), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n705), .A2(new_n723), .A3(new_n706), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n722), .B1(new_n724), .B2(G43gat), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT110), .ZN(new_n727));
  NAND4_X1  g526(.A1(new_n695), .A2(new_n723), .A3(new_n698), .A4(new_n702), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT109), .ZN(new_n729));
  OR2_X1    g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n204), .B1(new_n728), .B2(new_n729), .ZN(new_n731));
  AOI22_X1  g530(.A1(new_n730), .A2(new_n731), .B1(new_n683), .B2(new_n719), .ZN(new_n732));
  OAI211_X1 g531(.A(new_n726), .B(new_n727), .C1(new_n721), .C2(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n730), .A2(new_n731), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n721), .B1(new_n734), .B2(new_n720), .ZN(new_n735));
  OAI21_X1  g534(.A(KEYINPUT110), .B1(new_n735), .B2(new_n725), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n733), .A2(new_n736), .ZN(G1330gat));
  INV_X1    g536(.A(KEYINPUT112), .ZN(new_n738));
  NAND4_X1  g537(.A1(new_n695), .A2(new_n531), .A3(new_n698), .A4(new_n702), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n202), .B1(new_n739), .B2(KEYINPUT111), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n516), .A2(new_n552), .ZN(new_n741));
  AND4_X1   g540(.A1(KEYINPUT105), .A2(new_n741), .A3(KEYINPUT44), .A4(new_n640), .ZN(new_n742));
  AOI21_X1  g541(.A(KEYINPUT44), .B1(new_n697), .B2(KEYINPUT105), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT111), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n744), .A2(new_n745), .A3(new_n531), .A4(new_n702), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n740), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n683), .A2(new_n202), .A3(new_n531), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(KEYINPUT48), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT48), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n748), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n705), .A2(new_n531), .A3(new_n706), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n752), .B1(new_n753), .B2(G50gat), .ZN(new_n754));
  INV_X1    g553(.A(new_n754), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n738), .B1(new_n750), .B2(new_n755), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n751), .B1(new_n747), .B2(new_n748), .ZN(new_n757));
  NOR3_X1   g556(.A1(new_n757), .A2(new_n754), .A3(KEYINPUT112), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n756), .A2(new_n758), .ZN(G1331gat));
  NAND3_X1  g558(.A1(new_n628), .A2(new_n657), .A3(new_n699), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(KEYINPUT113), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(new_n741), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n762), .A2(new_n335), .ZN(new_n763));
  XOR2_X1   g562(.A(new_n763), .B(G57gat), .Z(G1332gat));
  NOR2_X1   g563(.A1(new_n762), .A2(new_n511), .ZN(new_n765));
  NOR2_X1   g564(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n766));
  AND2_X1   g565(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n765), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n768), .B1(new_n765), .B2(new_n766), .ZN(G1333gat));
  OAI21_X1  g568(.A(G71gat), .B1(new_n762), .B2(new_n551), .ZN(new_n770));
  OR2_X1    g569(.A1(new_n676), .A2(G71gat), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n770), .B1(new_n762), .B2(new_n771), .ZN(new_n772));
  XNOR2_X1  g571(.A(KEYINPUT114), .B(KEYINPUT50), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n772), .B(new_n773), .ZN(G1334gat));
  INV_X1    g573(.A(new_n531), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n762), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(new_n458), .ZN(G1335gat));
  INV_X1    g576(.A(KEYINPUT51), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT116), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n697), .A2(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT103), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n244), .B(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(new_n656), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  AND2_X1   g583(.A1(new_n780), .A2(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(new_n785), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n697), .A2(new_n779), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n778), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  OAI211_X1 g587(.A(new_n785), .B(KEYINPUT51), .C1(new_n779), .C2(new_n697), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(new_n628), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n665), .A2(new_n569), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n628), .A2(new_n784), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n793), .B(KEYINPUT115), .ZN(new_n794));
  AND2_X1   g593(.A1(new_n744), .A2(new_n794), .ZN(new_n795));
  AND2_X1   g594(.A1(new_n795), .A2(new_n665), .ZN(new_n796));
  OAI22_X1  g595(.A1(new_n791), .A2(new_n792), .B1(new_n569), .B2(new_n796), .ZN(G1336gat));
  INV_X1    g596(.A(KEYINPUT52), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n744), .A2(new_n508), .A3(new_n794), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT117), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(G92gat), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n799), .A2(new_n800), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n511), .A2(G92gat), .ZN(new_n804));
  INV_X1    g603(.A(new_n804), .ZN(new_n805));
  OAI221_X1 g604(.A(new_n798), .B1(new_n802), .B2(new_n803), .C1(new_n791), .C2(new_n805), .ZN(new_n806));
  AOI211_X1 g605(.A(new_n627), .B(new_n805), .C1(new_n788), .C2(new_n789), .ZN(new_n807));
  AND2_X1   g606(.A1(new_n799), .A2(G92gat), .ZN(new_n808));
  OAI21_X1  g607(.A(KEYINPUT52), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n806), .A2(new_n809), .ZN(G1337gat));
  NAND3_X1  g609(.A1(new_n790), .A2(new_n409), .A3(new_n628), .ZN(new_n811));
  INV_X1    g610(.A(G99gat), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n551), .A2(new_n812), .ZN(new_n813));
  AOI22_X1  g612(.A1(new_n811), .A2(new_n812), .B1(new_n795), .B2(new_n813), .ZN(G1338gat));
  NOR2_X1   g613(.A1(new_n775), .A2(G106gat), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n790), .A2(new_n628), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n795), .A2(new_n531), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(G106gat), .ZN(new_n818));
  XNOR2_X1  g617(.A(KEYINPUT118), .B(KEYINPUT53), .ZN(new_n819));
  AND3_X1   g618(.A1(new_n816), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n819), .B1(new_n816), .B2(new_n818), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n820), .A2(new_n821), .ZN(G1339gat));
  OAI21_X1  g621(.A(new_n613), .B1(new_n620), .B2(KEYINPUT54), .ZN(new_n823));
  AND3_X1   g622(.A1(new_n598), .A2(KEYINPUT120), .A3(new_n618), .ZN(new_n824));
  AOI21_X1  g623(.A(KEYINPUT120), .B1(new_n598), .B2(new_n618), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT54), .ZN(new_n826));
  NOR3_X1   g625(.A1(new_n824), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n823), .B1(new_n609), .B2(new_n827), .ZN(new_n828));
  AOI22_X1  g627(.A1(new_n828), .A2(KEYINPUT55), .B1(new_n609), .B2(new_n615), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n609), .A2(new_n827), .ZN(new_n830));
  INV_X1    g629(.A(new_n823), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT55), .ZN(new_n833));
  AOI21_X1  g632(.A(KEYINPUT121), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT121), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n828), .A2(new_n835), .A3(KEYINPUT55), .ZN(new_n836));
  OAI211_X1 g635(.A(new_n782), .B(new_n829), .C1(new_n834), .C2(new_n836), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n227), .A2(new_n228), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n232), .A2(new_n233), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n239), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  OAI211_X1 g639(.A(new_n243), .B(new_n840), .C1(new_n625), .C2(new_n626), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n640), .B1(new_n837), .B2(new_n841), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n832), .A2(KEYINPUT121), .A3(new_n833), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n835), .B1(new_n828), .B2(KEYINPUT55), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  AND3_X1   g644(.A1(new_n640), .A2(new_n243), .A3(new_n840), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n845), .A2(new_n829), .A3(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(new_n847), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n700), .B1(new_n842), .B2(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(new_n626), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n699), .A2(new_n850), .A3(new_n657), .A4(new_n624), .ZN(new_n851));
  XOR2_X1   g650(.A(new_n851), .B(KEYINPUT119), .Z(new_n852));
  AOI21_X1  g651(.A(new_n335), .B1(new_n849), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(new_n509), .ZN(new_n854));
  INV_X1    g653(.A(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n855), .A2(new_n274), .A3(new_n782), .ZN(new_n856));
  OAI21_X1  g655(.A(G113gat), .B1(new_n854), .B2(new_n245), .ZN(new_n857));
  AND2_X1   g656(.A1(new_n857), .A2(KEYINPUT122), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n857), .A2(KEYINPUT122), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n856), .B1(new_n858), .B2(new_n859), .ZN(G1340gat));
  OAI21_X1  g659(.A(G120gat), .B1(new_n854), .B2(new_n627), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n627), .A2(G120gat), .ZN(new_n862));
  XNOR2_X1  g661(.A(new_n862), .B(KEYINPUT123), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n861), .B1(new_n854), .B2(new_n863), .ZN(G1341gat));
  NOR3_X1   g663(.A1(new_n854), .A2(new_n278), .A3(new_n700), .ZN(new_n865));
  AND2_X1   g664(.A1(new_n865), .A2(KEYINPUT124), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n865), .A2(KEYINPUT124), .ZN(new_n867));
  AOI21_X1  g666(.A(G127gat), .B1(new_n855), .B2(new_n783), .ZN(new_n868));
  NOR3_X1   g667(.A1(new_n866), .A2(new_n867), .A3(new_n868), .ZN(G1342gat));
  NAND2_X1  g668(.A1(new_n855), .A2(new_n640), .ZN(new_n870));
  OR3_X1    g669(.A1(new_n870), .A2(KEYINPUT56), .A3(G134gat), .ZN(new_n871));
  OAI21_X1  g670(.A(KEYINPUT56), .B1(new_n870), .B2(G134gat), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n870), .A2(G134gat), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n871), .A2(new_n872), .A3(new_n873), .ZN(G1343gat));
  INV_X1    g673(.A(G141gat), .ZN(new_n875));
  NOR3_X1   g674(.A1(new_n723), .A2(new_n335), .A3(new_n508), .ZN(new_n876));
  INV_X1    g675(.A(new_n876), .ZN(new_n877));
  OAI211_X1 g676(.A(new_n829), .B(new_n244), .C1(KEYINPUT55), .C2(new_n828), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(new_n841), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(new_n696), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n783), .B1(new_n880), .B2(new_n847), .ZN(new_n881));
  XNOR2_X1  g680(.A(new_n851), .B(KEYINPUT119), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n531), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n877), .B1(new_n883), .B2(KEYINPUT57), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n775), .B1(new_n849), .B2(new_n852), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT57), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n875), .B1(new_n888), .B2(new_n782), .ZN(new_n889));
  NOR3_X1   g688(.A1(new_n723), .A2(new_n775), .A3(new_n508), .ZN(new_n890));
  AND2_X1   g689(.A1(new_n853), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n891), .A2(new_n875), .A3(new_n244), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT125), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  OAI21_X1  g693(.A(KEYINPUT58), .B1(new_n889), .B2(new_n894), .ZN(new_n895));
  AOI211_X1 g694(.A(KEYINPUT58), .B(new_n875), .C1(new_n888), .C2(new_n244), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT58), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n892), .B1(new_n893), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n895), .B1(new_n896), .B2(new_n898), .ZN(G1344gat));
  INV_X1    g698(.A(G148gat), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n891), .A2(new_n900), .A3(new_n628), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n775), .A2(KEYINPUT57), .ZN(new_n902));
  NOR3_X1   g701(.A1(new_n628), .A2(new_n244), .A3(new_n658), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n902), .B1(new_n881), .B2(new_n903), .ZN(new_n904));
  OAI211_X1 g703(.A(new_n904), .B(new_n628), .C1(new_n885), .C2(new_n886), .ZN(new_n905));
  OAI21_X1  g704(.A(G148gat), .B1(new_n905), .B2(new_n877), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n906), .A2(KEYINPUT59), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n884), .A2(new_n628), .A3(new_n887), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n900), .A2(KEYINPUT59), .ZN(new_n909));
  AND2_X1   g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  OAI211_X1 g709(.A(KEYINPUT126), .B(new_n901), .C1(new_n907), .C2(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT126), .ZN(new_n912));
  AOI22_X1  g711(.A1(new_n906), .A2(KEYINPUT59), .B1(new_n908), .B2(new_n909), .ZN(new_n913));
  INV_X1    g712(.A(new_n901), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n912), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n911), .A2(new_n915), .ZN(G1345gat));
  NAND3_X1  g715(.A1(new_n891), .A2(new_n248), .A3(new_n783), .ZN(new_n917));
  AND2_X1   g716(.A1(new_n888), .A2(new_n701), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n917), .B1(new_n918), .B2(new_n248), .ZN(G1346gat));
  AOI21_X1  g718(.A(G162gat), .B1(new_n891), .B2(new_n640), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n696), .A2(new_n249), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n920), .B1(new_n888), .B2(new_n921), .ZN(G1347gat));
  AOI21_X1  g721(.A(new_n665), .B1(new_n849), .B2(new_n852), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n472), .A2(new_n511), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NOR3_X1   g724(.A1(new_n925), .A2(new_n355), .A3(new_n245), .ZN(new_n926));
  INV_X1    g725(.A(new_n925), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(new_n782), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n926), .B1(new_n355), .B2(new_n928), .ZN(G1348gat));
  NOR2_X1   g728(.A1(new_n925), .A2(new_n627), .ZN(new_n930));
  XNOR2_X1  g729(.A(new_n930), .B(new_n356), .ZN(G1349gat));
  OAI21_X1  g730(.A(G183gat), .B1(new_n925), .B2(new_n700), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n783), .A2(new_n342), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n932), .B1(new_n925), .B2(new_n933), .ZN(new_n934));
  XNOR2_X1  g733(.A(new_n934), .B(KEYINPUT60), .ZN(G1350gat));
  NOR2_X1   g734(.A1(new_n925), .A2(new_n696), .ZN(new_n936));
  NAND2_X1  g735(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  XOR2_X1   g737(.A(KEYINPUT61), .B(G190gat), .Z(new_n939));
  OAI21_X1  g738(.A(new_n938), .B1(new_n936), .B2(new_n939), .ZN(G1351gat));
  AND4_X1   g739(.A1(new_n531), .A2(new_n923), .A3(new_n508), .A4(new_n551), .ZN(new_n941));
  AND2_X1   g740(.A1(new_n941), .A2(new_n782), .ZN(new_n942));
  NOR3_X1   g741(.A1(new_n723), .A2(new_n665), .A3(new_n511), .ZN(new_n943));
  OAI211_X1 g742(.A(new_n904), .B(new_n943), .C1(new_n885), .C2(new_n886), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n244), .A2(G197gat), .ZN(new_n945));
  OAI22_X1  g744(.A1(new_n942), .A2(G197gat), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  INV_X1    g745(.A(new_n946), .ZN(G1352gat));
  INV_X1    g746(.A(G204gat), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n941), .A2(new_n948), .A3(new_n628), .ZN(new_n949));
  OR2_X1    g748(.A1(new_n949), .A2(KEYINPUT62), .ZN(new_n950));
  INV_X1    g749(.A(new_n943), .ZN(new_n951));
  OAI21_X1  g750(.A(G204gat), .B1(new_n905), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n949), .A2(KEYINPUT62), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n950), .A2(new_n952), .A3(new_n953), .ZN(G1353gat));
  OAI221_X1 g753(.A(G211gat), .B1(KEYINPUT127), .B2(KEYINPUT63), .C1(new_n944), .C2(new_n656), .ZN(new_n955));
  NAND2_X1  g754(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n956));
  INV_X1    g755(.A(new_n956), .ZN(new_n957));
  OR2_X1    g756(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n955), .A2(new_n957), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n941), .A2(new_n420), .A3(new_n783), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n958), .A2(new_n959), .A3(new_n960), .ZN(G1354gat));
  NAND3_X1  g760(.A1(new_n941), .A2(new_n421), .A3(new_n640), .ZN(new_n962));
  OAI21_X1  g761(.A(G218gat), .B1(new_n944), .B2(new_n696), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n962), .A2(new_n963), .ZN(G1355gat));
endmodule


