//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 1 0 0 0 1 0 1 1 1 1 0 0 1 1 0 0 1 0 0 1 0 1 0 1 1 0 1 1 0 0 0 1 1 0 0 0 1 1 1 0 1 0 1 1 1 1 1 1 1 0 0 1 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:11 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n677, new_n678, new_n679, new_n680, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n734, new_n735, new_n736, new_n737, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n914, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978;
  INV_X1    g000(.A(G116), .ZN(new_n187));
  OAI21_X1  g001(.A(KEYINPUT70), .B1(new_n187), .B2(G119), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT70), .ZN(new_n189));
  INV_X1    g003(.A(G119), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n189), .A2(new_n190), .A3(G116), .ZN(new_n191));
  AND2_X1   g005(.A1(new_n188), .A2(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT71), .B(G116), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G119), .ZN(new_n194));
  XNOR2_X1  g008(.A(KEYINPUT2), .B(G113), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  AND3_X1   g010(.A1(new_n192), .A2(new_n194), .A3(new_n196), .ZN(new_n197));
  AOI21_X1  g011(.A(new_n196), .B1(new_n192), .B2(new_n194), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT11), .ZN(new_n201));
  INV_X1    g015(.A(G134), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n201), .B1(new_n202), .B2(G137), .ZN(new_n203));
  INV_X1    g017(.A(G137), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n204), .A2(KEYINPUT11), .A3(G134), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n202), .A2(G137), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n203), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(KEYINPUT68), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT68), .ZN(new_n209));
  NAND4_X1  g023(.A1(new_n203), .A2(new_n205), .A3(new_n209), .A4(new_n206), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n208), .A2(G131), .A3(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G131), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n203), .A2(new_n205), .A3(new_n212), .A4(new_n206), .ZN(new_n213));
  AND2_X1   g027(.A1(new_n213), .A2(KEYINPUT69), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n211), .A2(new_n214), .ZN(new_n215));
  AND2_X1   g029(.A1(KEYINPUT66), .A2(G143), .ZN(new_n216));
  NOR2_X1   g030(.A1(KEYINPUT66), .A2(G143), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  XNOR2_X1  g032(.A(KEYINPUT67), .B(G146), .ZN(new_n219));
  AOI22_X1  g033(.A1(new_n218), .A2(G146), .B1(new_n219), .B2(G143), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT0), .ZN(new_n221));
  INV_X1    g035(.A(G128), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G146), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n224), .B1(new_n216), .B2(new_n217), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n225), .B1(new_n219), .B2(G143), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT65), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n227), .B1(KEYINPUT0), .B2(G128), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n221), .A2(new_n222), .A3(KEYINPUT65), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n223), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  AOI22_X1  g044(.A1(new_n220), .A2(new_n223), .B1(new_n226), .B2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT69), .ZN(new_n232));
  NAND4_X1  g046(.A1(new_n208), .A2(new_n232), .A3(G131), .A4(new_n210), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n215), .A2(new_n231), .A3(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n224), .A2(KEYINPUT67), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT67), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G146), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n235), .A2(new_n237), .A3(G143), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n222), .A2(KEYINPUT1), .ZN(new_n239));
  XNOR2_X1  g053(.A(KEYINPUT66), .B(G143), .ZN(new_n240));
  OAI211_X1 g054(.A(new_n238), .B(new_n239), .C1(new_n224), .C2(new_n240), .ZN(new_n241));
  OR2_X1    g055(.A1(KEYINPUT66), .A2(G143), .ZN(new_n242));
  NAND2_X1  g056(.A1(KEYINPUT66), .A2(G143), .ZN(new_n243));
  AOI21_X1  g057(.A(G146), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(G143), .B1(new_n235), .B2(new_n237), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n222), .B1(new_n238), .B2(KEYINPUT1), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n241), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(new_n206), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n202), .A2(G137), .ZN(new_n250));
  OAI21_X1  g064(.A(G131), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n248), .A2(new_n213), .A3(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n234), .A2(new_n252), .ZN(new_n253));
  AOI21_X1  g067(.A(KEYINPUT30), .B1(new_n253), .B2(KEYINPUT64), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT64), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT30), .ZN(new_n256));
  AOI211_X1 g070(.A(new_n255), .B(new_n256), .C1(new_n234), .C2(new_n252), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n200), .B1(new_n254), .B2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(G237), .ZN(new_n259));
  INV_X1    g073(.A(G953), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n259), .A2(new_n260), .A3(G210), .ZN(new_n261));
  XOR2_X1   g075(.A(new_n261), .B(KEYINPUT27), .Z(new_n262));
  XNOR2_X1  g076(.A(KEYINPUT26), .B(G101), .ZN(new_n263));
  XOR2_X1   g077(.A(new_n262), .B(new_n263), .Z(new_n264));
  NAND3_X1  g078(.A1(new_n234), .A2(new_n199), .A3(new_n252), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n258), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(KEYINPUT31), .ZN(new_n267));
  INV_X1    g081(.A(new_n264), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT72), .ZN(new_n269));
  AND3_X1   g083(.A1(new_n234), .A2(new_n199), .A3(new_n252), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n199), .B1(new_n234), .B2(new_n252), .ZN(new_n271));
  OAI211_X1 g085(.A(new_n269), .B(KEYINPUT28), .C1(new_n270), .C2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT28), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n265), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n253), .A2(new_n200), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(new_n265), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n269), .B1(new_n277), .B2(KEYINPUT28), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n268), .B1(new_n275), .B2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT31), .ZN(new_n280));
  NAND4_X1  g094(.A1(new_n258), .A2(new_n280), .A3(new_n264), .A4(new_n265), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n267), .A2(new_n279), .A3(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT74), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT32), .ZN(new_n284));
  NOR3_X1   g098(.A1(new_n284), .A2(G472), .A3(G902), .ZN(new_n285));
  AND3_X1   g099(.A1(new_n282), .A2(new_n283), .A3(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n283), .B1(new_n282), .B2(new_n285), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NOR2_X1   g102(.A1(G472), .A2(G902), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n282), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(new_n284), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT73), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT29), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n277), .A2(KEYINPUT28), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(KEYINPUT72), .ZN(new_n295));
  INV_X1    g109(.A(new_n274), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n273), .B1(new_n276), .B2(new_n265), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n296), .B1(new_n297), .B2(new_n269), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n268), .B1(new_n295), .B2(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n258), .A2(new_n268), .A3(new_n265), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n293), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n297), .A2(new_n296), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n268), .A2(new_n293), .ZN(new_n304));
  AOI21_X1  g118(.A(G902), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n302), .A2(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n292), .B1(new_n306), .B2(G472), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n264), .B1(new_n275), .B2(new_n278), .ZN(new_n308));
  AOI21_X1  g122(.A(KEYINPUT29), .B1(new_n308), .B2(new_n300), .ZN(new_n309));
  INV_X1    g123(.A(new_n305), .ZN(new_n310));
  OAI211_X1 g124(.A(new_n292), .B(G472), .C1(new_n309), .C2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  OAI211_X1 g126(.A(new_n288), .B(new_n291), .C1(new_n307), .C2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(G140), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(G125), .ZN(new_n315));
  INV_X1    g129(.A(G125), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(G140), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT76), .ZN(new_n318));
  NAND4_X1  g132(.A1(new_n315), .A2(new_n317), .A3(new_n318), .A4(KEYINPUT16), .ZN(new_n319));
  AND3_X1   g133(.A1(new_n315), .A2(new_n317), .A3(KEYINPUT16), .ZN(new_n320));
  OAI21_X1  g134(.A(KEYINPUT76), .B1(new_n315), .B2(KEYINPUT16), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n319), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(G146), .ZN(new_n323));
  OAI211_X1 g137(.A(new_n224), .B(new_n319), .C1(new_n320), .C2(new_n321), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  OAI21_X1  g139(.A(KEYINPUT75), .B1(new_n190), .B2(G128), .ZN(new_n326));
  AOI22_X1  g140(.A1(new_n326), .A2(KEYINPUT23), .B1(new_n190), .B2(G128), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n327), .B1(KEYINPUT23), .B2(new_n326), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(G110), .ZN(new_n329));
  XOR2_X1   g143(.A(G119), .B(G128), .Z(new_n330));
  XNOR2_X1  g144(.A(KEYINPUT24), .B(G110), .ZN(new_n331));
  OAI211_X1 g145(.A(new_n325), .B(new_n329), .C1(new_n330), .C2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT77), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n323), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n322), .A2(KEYINPUT77), .A3(G146), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n316), .A2(G140), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n314), .A2(G125), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(new_n219), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n330), .A2(new_n331), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n340), .B1(new_n328), .B2(G110), .ZN(new_n341));
  NAND4_X1  g155(.A1(new_n334), .A2(new_n335), .A3(new_n339), .A4(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n332), .A2(new_n342), .ZN(new_n343));
  XNOR2_X1  g157(.A(KEYINPUT22), .B(G137), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n260), .A2(G221), .A3(G234), .ZN(new_n345));
  XNOR2_X1  g159(.A(new_n344), .B(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n343), .A2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(G902), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n332), .A2(new_n342), .A3(new_n346), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n348), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT78), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n352), .A2(KEYINPUT25), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(new_n353), .ZN(new_n355));
  NAND4_X1  g169(.A1(new_n348), .A2(new_n349), .A3(new_n350), .A4(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(G217), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n358), .B1(G234), .B2(new_n349), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  AND2_X1   g174(.A1(new_n348), .A2(new_n350), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n359), .A2(G902), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n360), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  OAI21_X1  g179(.A(G214), .B1(G237), .B2(G902), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT3), .ZN(new_n368));
  INV_X1    g182(.A(G104), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n368), .B1(new_n369), .B2(G107), .ZN(new_n370));
  INV_X1    g184(.A(G107), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n371), .A2(KEYINPUT3), .A3(G104), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n369), .A2(G107), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  XOR2_X1   g189(.A(KEYINPUT81), .B(KEYINPUT4), .Z(new_n376));
  NAND3_X1  g190(.A1(new_n375), .A2(G101), .A3(new_n376), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n377), .B1(new_n197), .B2(new_n198), .ZN(new_n378));
  INV_X1    g192(.A(G101), .ZN(new_n379));
  AND3_X1   g193(.A1(new_n371), .A2(KEYINPUT3), .A3(G104), .ZN(new_n380));
  AOI21_X1  g194(.A(KEYINPUT3), .B1(new_n371), .B2(G104), .ZN(new_n381));
  OAI211_X1 g195(.A(new_n379), .B(new_n374), .C1(new_n380), .C2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(KEYINPUT4), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n379), .B1(new_n373), .B2(new_n374), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n192), .A2(new_n194), .A3(KEYINPUT5), .ZN(new_n386));
  NOR3_X1   g200(.A1(new_n187), .A2(KEYINPUT5), .A3(G119), .ZN(new_n387));
  INV_X1    g201(.A(G113), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n188), .A2(new_n191), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n391), .B1(G119), .B2(new_n193), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(new_n196), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n390), .A2(new_n393), .ZN(new_n394));
  OAI21_X1  g208(.A(KEYINPUT83), .B1(new_n371), .B2(G104), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT83), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n396), .A2(new_n369), .A3(G107), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n371), .A2(G104), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n395), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(G101), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(new_n382), .ZN(new_n401));
  OAI22_X1  g215(.A1(new_n378), .A2(new_n385), .B1(new_n394), .B2(new_n401), .ZN(new_n402));
  XNOR2_X1  g216(.A(G110), .B(G122), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  AOI22_X1  g219(.A1(new_n386), .A2(new_n389), .B1(new_n392), .B2(new_n196), .ZN(new_n406));
  AND2_X1   g220(.A1(new_n400), .A2(new_n382), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  OAI211_X1 g222(.A(new_n408), .B(new_n403), .C1(new_n385), .C2(new_n378), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n405), .A2(KEYINPUT6), .A3(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT6), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n402), .A2(new_n411), .A3(new_n404), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT1), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n413), .B1(new_n219), .B2(G143), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n226), .B1(new_n414), .B2(new_n222), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n415), .A2(new_n316), .A3(new_n241), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n416), .B1(new_n231), .B2(new_n316), .ZN(new_n417));
  INV_X1    g231(.A(G224), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n418), .A2(G953), .ZN(new_n419));
  XNOR2_X1  g233(.A(new_n417), .B(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n410), .A2(new_n412), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n192), .A2(new_n194), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(new_n195), .ZN(new_n423));
  AOI22_X1  g237(.A1(new_n393), .A2(new_n423), .B1(new_n384), .B2(new_n376), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n375), .A2(G101), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n425), .A2(KEYINPUT4), .A3(new_n382), .ZN(new_n426));
  AOI22_X1  g240(.A1(new_n424), .A2(new_n426), .B1(new_n407), .B2(new_n406), .ZN(new_n427));
  OAI21_X1  g241(.A(KEYINPUT7), .B1(new_n418), .B2(G953), .ZN(new_n428));
  AOI22_X1  g242(.A1(new_n427), .A2(new_n403), .B1(new_n417), .B2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(new_n417), .ZN(new_n430));
  INV_X1    g244(.A(new_n428), .ZN(new_n431));
  XOR2_X1   g245(.A(new_n403), .B(KEYINPUT8), .Z(new_n432));
  INV_X1    g246(.A(KEYINPUT87), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n407), .A2(new_n433), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n432), .B1(new_n434), .B2(new_n406), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n394), .A2(new_n433), .A3(new_n407), .ZN(new_n436));
  AOI22_X1  g250(.A1(new_n430), .A2(new_n431), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  AOI21_X1  g251(.A(G902), .B1(new_n429), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n421), .A2(new_n438), .ZN(new_n439));
  OAI21_X1  g253(.A(G210), .B1(G237), .B2(G902), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n421), .A2(new_n438), .A3(new_n440), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n367), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(G234), .A2(G237), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n445), .A2(G952), .A3(new_n260), .ZN(new_n446));
  XOR2_X1   g260(.A(KEYINPUT21), .B(G898), .Z(new_n447));
  NAND3_X1  g261(.A1(new_n445), .A2(G902), .A3(G953), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n446), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n444), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n242), .A2(G128), .A3(new_n243), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n222), .A2(G143), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n451), .A2(KEYINPUT13), .A3(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT13), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n218), .A2(new_n454), .A3(G128), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n453), .A2(G134), .A3(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n451), .A2(new_n202), .A3(new_n452), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n187), .A2(KEYINPUT71), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT71), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(G116), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n458), .A2(new_n460), .A3(G122), .ZN(new_n461));
  OR2_X1    g275(.A1(new_n187), .A2(G122), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n461), .A2(new_n371), .A3(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n371), .B1(new_n461), .B2(new_n462), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n456), .B(new_n457), .C1(new_n464), .C2(new_n465), .ZN(new_n466));
  NOR3_X1   g280(.A1(new_n216), .A2(new_n217), .A3(new_n222), .ZN(new_n467));
  INV_X1    g281(.A(new_n452), .ZN(new_n468));
  OAI21_X1  g282(.A(G134), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(new_n457), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT14), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n461), .A2(new_n471), .A3(new_n462), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n193), .A2(KEYINPUT14), .A3(G122), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n472), .A2(G107), .A3(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n470), .A2(new_n463), .A3(new_n474), .ZN(new_n475));
  XNOR2_X1  g289(.A(KEYINPUT9), .B(G234), .ZN(new_n476));
  XNOR2_X1  g290(.A(new_n476), .B(KEYINPUT79), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n358), .A2(G953), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n466), .A2(new_n475), .A3(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT90), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n466), .A2(new_n475), .A3(new_n480), .A4(KEYINPUT90), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n466), .A2(new_n475), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(new_n479), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n483), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(new_n349), .ZN(new_n488));
  INV_X1    g302(.A(G478), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n489), .A2(KEYINPUT15), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  OAI211_X1 g305(.A(new_n487), .B(new_n349), .C1(KEYINPUT15), .C2(new_n489), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  NOR2_X1   g308(.A1(G475), .A2(G902), .ZN(new_n495));
  XNOR2_X1  g309(.A(G113), .B(G122), .ZN(new_n496));
  XNOR2_X1  g310(.A(new_n496), .B(new_n369), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n259), .A2(new_n260), .A3(G143), .A4(G214), .ZN(new_n498));
  INV_X1    g312(.A(G214), .ZN(new_n499));
  NOR3_X1   g313(.A1(new_n499), .A2(G237), .A3(G953), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n498), .B1(new_n240), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(G131), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n259), .A2(new_n260), .A3(G214), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n503), .A2(new_n242), .A3(new_n243), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n504), .A2(new_n212), .A3(new_n498), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT19), .ZN(new_n507));
  OAI21_X1  g321(.A(KEYINPUT89), .B1(new_n336), .B2(new_n337), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT89), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n315), .A2(new_n317), .A3(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n507), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n338), .A2(KEYINPUT19), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n219), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND4_X1  g327(.A1(new_n334), .A2(new_n335), .A3(new_n506), .A4(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n508), .A2(G146), .A3(new_n510), .ZN(new_n515));
  AND4_X1   g329(.A1(G143), .A2(new_n259), .A3(new_n260), .A4(G214), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n516), .B1(new_n218), .B2(new_n503), .ZN(new_n517));
  NAND2_X1  g331(.A1(KEYINPUT88), .A2(KEYINPUT18), .ZN(new_n518));
  AOI22_X1  g332(.A1(new_n339), .A2(new_n515), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n518), .ZN(new_n520));
  AND3_X1   g334(.A1(new_n504), .A2(new_n212), .A3(new_n498), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n212), .B1(new_n504), .B2(new_n498), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n519), .A2(new_n523), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n497), .B1(new_n514), .B2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT17), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n502), .A2(new_n526), .A3(new_n505), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n522), .A2(KEYINPUT17), .ZN(new_n528));
  NAND4_X1  g342(.A1(new_n527), .A2(new_n324), .A3(new_n323), .A4(new_n528), .ZN(new_n529));
  AND3_X1   g343(.A1(new_n529), .A2(new_n497), .A3(new_n524), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n495), .B1(new_n525), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(KEYINPUT20), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT20), .ZN(new_n533));
  OAI211_X1 g347(.A(new_n533), .B(new_n495), .C1(new_n525), .C2(new_n530), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n497), .B1(new_n529), .B2(new_n524), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n349), .B1(new_n530), .B2(new_n535), .ZN(new_n536));
  AOI22_X1  g350(.A1(new_n532), .A2(new_n534), .B1(new_n536), .B2(G475), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n494), .A2(new_n537), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n450), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n477), .A2(new_n349), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(G221), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n541), .B(KEYINPUT80), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT85), .ZN(new_n543));
  OAI21_X1  g357(.A(KEYINPUT84), .B1(new_n248), .B2(new_n407), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT84), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n415), .A2(new_n401), .A3(new_n545), .A4(new_n241), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n222), .B1(new_n225), .B2(KEYINPUT1), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n241), .B1(new_n220), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(new_n407), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n544), .A2(new_n546), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n215), .A2(new_n233), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  AND3_X1   g366(.A1(new_n550), .A2(new_n552), .A3(KEYINPUT12), .ZN(new_n553));
  AOI21_X1  g367(.A(KEYINPUT12), .B1(new_n550), .B2(new_n552), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n543), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n550), .A2(new_n552), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT12), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n550), .A2(new_n552), .A3(KEYINPUT12), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n558), .A2(KEYINPUT85), .A3(new_n559), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n230), .B1(new_n244), .B2(new_n245), .ZN(new_n561));
  OAI211_X1 g375(.A(new_n238), .B(new_n223), .C1(new_n224), .C2(new_n240), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n377), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  OAI21_X1  g377(.A(KEYINPUT82), .B1(new_n563), .B2(new_n385), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT82), .ZN(new_n565));
  NAND4_X1  g379(.A1(new_n231), .A2(new_n426), .A3(new_n565), .A4(new_n377), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT10), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n548), .A2(new_n568), .A3(new_n407), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n401), .B1(new_n415), .B2(new_n241), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n569), .B1(new_n570), .B2(new_n568), .ZN(new_n571));
  AND3_X1   g385(.A1(new_n567), .A2(new_n551), .A3(new_n571), .ZN(new_n572));
  XNOR2_X1  g386(.A(G110), .B(G140), .ZN(new_n573));
  AND2_X1   g387(.A1(new_n260), .A2(G227), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n573), .B(new_n574), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n555), .A2(new_n560), .A3(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n551), .B1(new_n567), .B2(new_n571), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n575), .B1(new_n572), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(KEYINPUT86), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT86), .ZN(new_n581));
  OAI211_X1 g395(.A(new_n581), .B(new_n575), .C1(new_n572), .C2(new_n578), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n577), .A2(new_n580), .A3(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(G469), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n583), .A2(new_n584), .A3(new_n349), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n584), .A2(new_n349), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n567), .A2(new_n551), .A3(new_n571), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n587), .B1(new_n553), .B2(new_n554), .ZN(new_n588));
  INV_X1    g402(.A(new_n578), .ZN(new_n589));
  AOI22_X1  g403(.A1(new_n588), .A2(new_n575), .B1(new_n576), .B2(new_n589), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n586), .B1(new_n590), .B2(G469), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n542), .B1(new_n585), .B2(new_n591), .ZN(new_n592));
  AND4_X1   g406(.A1(new_n313), .A2(new_n365), .A3(new_n539), .A4(new_n592), .ZN(new_n593));
  XNOR2_X1  g407(.A(KEYINPUT91), .B(G101), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n593), .B(new_n594), .ZN(G3));
  NAND2_X1  g409(.A1(new_n282), .A2(new_n349), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(G472), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT92), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n599), .B1(new_n282), .B2(new_n289), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n487), .A2(new_n489), .A3(new_n349), .ZN(new_n601));
  OR2_X1    g415(.A1(new_n487), .A2(KEYINPUT33), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT93), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n486), .B1(new_n603), .B2(new_n481), .ZN(new_n604));
  AND2_X1   g418(.A1(new_n481), .A2(new_n603), .ZN(new_n605));
  OAI21_X1  g419(.A(KEYINPUT33), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(G902), .B1(new_n602), .B2(new_n606), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n601), .B1(new_n607), .B2(new_n489), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(KEYINPUT94), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT94), .ZN(new_n610));
  OAI211_X1 g424(.A(new_n610), .B(new_n601), .C1(new_n607), .C2(new_n489), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n537), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n614), .A2(new_n450), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n597), .A2(new_n598), .ZN(new_n616));
  AND2_X1   g430(.A1(new_n592), .A2(new_n365), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n600), .A2(new_n615), .A3(new_n616), .A4(new_n617), .ZN(new_n618));
  XOR2_X1   g432(.A(KEYINPUT34), .B(G104), .Z(new_n619));
  XNOR2_X1  g433(.A(new_n618), .B(new_n619), .ZN(G6));
  NOR2_X1   g434(.A1(new_n613), .A2(new_n494), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n450), .A2(new_n622), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n600), .A2(new_n616), .A3(new_n617), .A4(new_n623), .ZN(new_n624));
  XOR2_X1   g438(.A(KEYINPUT35), .B(G107), .Z(new_n625));
  XNOR2_X1  g439(.A(new_n624), .B(new_n625), .ZN(G9));
  NOR2_X1   g440(.A1(new_n347), .A2(KEYINPUT36), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n343), .B(new_n627), .ZN(new_n628));
  AOI22_X1  g442(.A1(new_n357), .A2(new_n359), .B1(new_n362), .B2(new_n628), .ZN(new_n629));
  AOI211_X1 g443(.A(new_n542), .B(new_n629), .C1(new_n585), .C2(new_n591), .ZN(new_n630));
  NAND4_X1  g444(.A1(new_n600), .A2(new_n539), .A3(new_n616), .A4(new_n630), .ZN(new_n631));
  XOR2_X1   g445(.A(KEYINPUT37), .B(G110), .Z(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(G12));
  NAND2_X1  g447(.A1(new_n532), .A2(new_n534), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n536), .A2(G475), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n446), .B(KEYINPUT95), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n636), .B1(G900), .B2(new_n448), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n493), .A2(new_n634), .A3(new_n635), .A4(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(KEYINPUT96), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT96), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n537), .A2(new_n640), .A3(new_n493), .A4(new_n637), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n639), .A2(new_n444), .A3(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT97), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n639), .A2(new_n444), .A3(KEYINPUT97), .A4(new_n641), .ZN(new_n645));
  AND3_X1   g459(.A1(new_n630), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(new_n313), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(G128), .ZN(G30));
  INV_X1    g462(.A(new_n629), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n613), .A2(new_n493), .ZN(new_n650));
  NOR3_X1   g464(.A1(new_n649), .A2(new_n650), .A3(new_n367), .ZN(new_n651));
  XOR2_X1   g465(.A(new_n651), .B(KEYINPUT101), .Z(new_n652));
  XNOR2_X1  g466(.A(new_n637), .B(KEYINPUT39), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n592), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n654), .A2(KEYINPUT40), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n442), .A2(new_n443), .ZN(new_n656));
  XOR2_X1   g470(.A(KEYINPUT98), .B(KEYINPUT38), .Z(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(KEYINPUT99), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n656), .B(new_n658), .ZN(new_n659));
  NOR3_X1   g473(.A1(new_n652), .A2(new_n655), .A3(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n287), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n282), .A2(new_n283), .A3(new_n285), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n258), .A2(new_n265), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n264), .ZN(new_n664));
  OAI211_X1 g478(.A(new_n664), .B(new_n349), .C1(new_n264), .C2(new_n277), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(G472), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n661), .A2(new_n291), .A3(new_n662), .A4(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(KEYINPUT100), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT100), .ZN(new_n669));
  AOI22_X1  g483(.A1(new_n290), .A2(new_n284), .B1(G472), .B2(new_n665), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n288), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n654), .A2(KEYINPUT40), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n660), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  XOR2_X1   g488(.A(new_n674), .B(KEYINPUT102), .Z(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(new_n240), .ZN(G45));
  NAND3_X1  g490(.A1(new_n612), .A2(new_n613), .A3(new_n637), .ZN(new_n677));
  INV_X1    g491(.A(new_n444), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n313), .A2(new_n679), .A3(new_n630), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G146), .ZN(G48));
  INV_X1    g495(.A(new_n313), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n682), .A2(new_n364), .ZN(new_n683));
  INV_X1    g497(.A(new_n541), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n583), .A2(new_n349), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(G469), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT103), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n686), .A2(new_n687), .A3(new_n585), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n685), .A2(KEYINPUT103), .A3(G469), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n684), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n683), .A2(new_n615), .A3(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(KEYINPUT41), .B(G113), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(G15));
  NAND3_X1  g507(.A1(new_n683), .A2(new_n623), .A3(new_n690), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G116), .ZN(G18));
  INV_X1    g509(.A(new_n538), .ZN(new_n696));
  INV_X1    g510(.A(new_n450), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n690), .A2(new_n696), .A3(new_n697), .A4(new_n649), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n698), .A2(new_n682), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(KEYINPUT104), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G119), .ZN(G21));
  OAI211_X1 g515(.A(new_n267), .B(new_n281), .C1(new_n264), .C2(new_n303), .ZN(new_n702));
  AOI22_X1  g516(.A1(new_n596), .A2(G472), .B1(new_n289), .B2(new_n702), .ZN(new_n703));
  AND2_X1   g517(.A1(new_n703), .A2(new_n365), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT105), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n650), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n613), .A2(KEYINPUT105), .A3(new_n493), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n704), .A2(new_n690), .A3(new_n697), .A4(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G122), .ZN(G24));
  NAND2_X1  g524(.A1(new_n702), .A2(new_n289), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n597), .A2(new_n649), .A3(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT106), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n703), .A2(KEYINPUT106), .A3(new_n649), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(new_n677), .ZN(new_n717));
  AOI211_X1 g531(.A(new_n678), .B(new_n684), .C1(new_n688), .C2(new_n689), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n716), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G125), .ZN(G27));
  OAI21_X1  g534(.A(G472), .B1(new_n309), .B2(new_n310), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(KEYINPUT73), .ZN(new_n722));
  AOI22_X1  g536(.A1(new_n722), .A2(new_n311), .B1(new_n284), .B2(new_n290), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n282), .A2(new_n285), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n364), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n585), .A2(new_n591), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n656), .A2(new_n367), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n726), .A2(new_n541), .A3(new_n727), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n677), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n725), .A2(KEYINPUT42), .A3(new_n729), .ZN(new_n730));
  NOR4_X1   g544(.A1(new_n682), .A2(new_n364), .A3(new_n677), .A4(new_n728), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n730), .B1(new_n731), .B2(KEYINPUT42), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G131), .ZN(G33));
  INV_X1    g547(.A(new_n728), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n639), .A2(new_n641), .ZN(new_n735));
  XOR2_X1   g549(.A(new_n735), .B(KEYINPUT107), .Z(new_n736));
  NAND3_X1  g550(.A1(new_n683), .A2(new_n734), .A3(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G134), .ZN(G36));
  INV_X1    g552(.A(new_n727), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n600), .A2(new_n616), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n612), .A2(new_n537), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT43), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n741), .B1(KEYINPUT108), .B2(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(KEYINPUT108), .B(KEYINPUT43), .ZN(new_n744));
  OAI21_X1  g558(.A(new_n743), .B1(new_n741), .B2(new_n744), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n740), .A2(new_n649), .A3(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT44), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n739), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n748), .B1(new_n747), .B2(new_n746), .ZN(new_n749));
  OR2_X1    g563(.A1(new_n749), .A2(KEYINPUT109), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(KEYINPUT109), .ZN(new_n751));
  AND2_X1   g565(.A1(new_n590), .A2(KEYINPUT45), .ZN(new_n752));
  OAI21_X1  g566(.A(G469), .B1(new_n590), .B2(KEYINPUT45), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(new_n586), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n755), .A2(KEYINPUT46), .A3(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT46), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n758), .B1(new_n754), .B2(new_n586), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n757), .A2(new_n585), .A3(new_n759), .ZN(new_n760));
  AND3_X1   g574(.A1(new_n760), .A2(new_n541), .A3(new_n653), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n750), .A2(new_n751), .A3(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G137), .ZN(G39));
  NAND2_X1  g577(.A1(new_n760), .A2(new_n541), .ZN(new_n764));
  NAND2_X1  g578(.A1(KEYINPUT110), .A2(KEYINPUT47), .ZN(new_n765));
  NOR2_X1   g579(.A1(KEYINPUT110), .A2(KEYINPUT47), .ZN(new_n766));
  INV_X1    g580(.A(new_n766), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n764), .B1(new_n765), .B2(new_n767), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n768), .B1(new_n764), .B2(new_n767), .ZN(new_n769));
  NOR4_X1   g583(.A1(new_n313), .A2(new_n365), .A3(new_n677), .A4(new_n739), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G140), .ZN(G42));
  INV_X1    g586(.A(new_n542), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n659), .A2(new_n365), .A3(new_n366), .A4(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n688), .A2(new_n689), .ZN(new_n775));
  INV_X1    g589(.A(new_n775), .ZN(new_n776));
  AOI211_X1 g590(.A(new_n741), .B(new_n774), .C1(new_n776), .C2(KEYINPUT49), .ZN(new_n777));
  INV_X1    g591(.A(new_n672), .ZN(new_n778));
  OAI211_X1 g592(.A(new_n777), .B(new_n778), .C1(KEYINPUT49), .C2(new_n776), .ZN(new_n779));
  INV_X1    g593(.A(new_n636), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n745), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n781), .A2(new_n704), .ZN(new_n782));
  INV_X1    g596(.A(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n690), .A2(new_n367), .A3(new_n659), .ZN(new_n784));
  INV_X1    g598(.A(new_n784), .ZN(new_n785));
  OAI211_X1 g599(.A(new_n783), .B(new_n785), .C1(KEYINPUT119), .C2(KEYINPUT50), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT119), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT50), .ZN(new_n788));
  OAI211_X1 g602(.A(new_n787), .B(new_n788), .C1(new_n782), .C2(new_n784), .ZN(new_n789));
  OAI211_X1 g603(.A(new_n786), .B(new_n789), .C1(new_n787), .C2(new_n788), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n776), .A2(new_n773), .ZN(new_n791));
  OAI211_X1 g605(.A(new_n727), .B(new_n783), .C1(new_n769), .C2(new_n791), .ZN(new_n792));
  AND2_X1   g606(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  AND2_X1   g607(.A1(new_n690), .A2(new_n727), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n364), .A2(new_n446), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n778), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(KEYINPUT120), .ZN(new_n797));
  NOR3_X1   g611(.A1(new_n797), .A2(new_n613), .A3(new_n612), .ZN(new_n798));
  AND2_X1   g612(.A1(new_n781), .A2(new_n794), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n798), .B1(new_n716), .B2(new_n799), .ZN(new_n800));
  AOI21_X1  g614(.A(KEYINPUT51), .B1(new_n793), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n799), .A2(new_n725), .ZN(new_n802));
  XOR2_X1   g616(.A(new_n802), .B(KEYINPUT48), .Z(new_n803));
  NAND2_X1  g617(.A1(new_n260), .A2(G952), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n804), .B1(new_n783), .B2(new_n718), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n805), .B1(new_n797), .B2(new_n614), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n801), .A2(new_n803), .A3(new_n806), .ZN(new_n807));
  OR2_X1    g621(.A1(new_n800), .A2(KEYINPUT121), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n800), .A2(KEYINPUT121), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n808), .A2(KEYINPUT51), .A3(new_n809), .A4(new_n793), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n807), .A2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT54), .ZN(new_n812));
  INV_X1    g626(.A(new_n637), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n739), .A2(new_n538), .A3(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n313), .A2(new_n630), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n716), .A2(new_n729), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n732), .A2(new_n815), .A3(new_n737), .A4(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n618), .A2(new_n624), .A3(new_n631), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT111), .ZN(new_n820));
  OR3_X1    g634(.A1(new_n819), .A2(new_n820), .A3(new_n593), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n820), .B1(new_n819), .B2(new_n593), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n700), .A2(new_n694), .ZN(new_n824));
  AND2_X1   g638(.A1(new_n691), .A2(new_n709), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n818), .A2(new_n823), .A3(new_n824), .A4(new_n825), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n678), .B1(new_n706), .B2(new_n707), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n649), .A2(new_n684), .A3(new_n813), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n827), .A2(new_n726), .A3(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(new_n829), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n667), .A2(KEYINPUT100), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n669), .B1(new_n288), .B2(new_n670), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n830), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n833), .A2(KEYINPUT113), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT113), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n672), .A2(new_n835), .A3(new_n830), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  AND3_X1   g651(.A1(new_n719), .A2(new_n647), .A3(new_n680), .ZN(new_n838));
  AOI21_X1  g652(.A(KEYINPUT52), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n712), .A2(new_n713), .ZN(new_n840));
  AOI21_X1  g654(.A(KEYINPUT106), .B1(new_n703), .B2(new_n649), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n690), .A2(new_n717), .A3(new_n444), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n647), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n680), .A2(KEYINPUT52), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n846), .B1(new_n834), .B2(new_n836), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n839), .B1(new_n845), .B2(new_n847), .ZN(new_n848));
  XOR2_X1   g662(.A(KEYINPUT117), .B(KEYINPUT53), .Z(new_n849));
  NOR3_X1   g663(.A1(new_n826), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  AND2_X1   g664(.A1(new_n821), .A2(new_n822), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n825), .A2(new_n700), .A3(new_n694), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n851), .A2(new_n852), .A3(new_n817), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT115), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n844), .A2(KEYINPUT112), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT112), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n719), .A2(new_n856), .A3(new_n647), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  AND2_X1   g672(.A1(new_n680), .A2(KEYINPUT52), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n835), .B1(new_n672), .B2(new_n830), .ZN(new_n860));
  AOI211_X1 g674(.A(KEYINPUT113), .B(new_n829), .C1(new_n668), .C2(new_n671), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n859), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  OAI21_X1  g676(.A(KEYINPUT114), .B1(new_n858), .B2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT114), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n847), .A2(new_n864), .A3(new_n855), .A4(new_n857), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(new_n839), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n854), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  AOI211_X1 g682(.A(KEYINPUT115), .B(new_n839), .C1(new_n863), .C2(new_n865), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n853), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT53), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT116), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n850), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n870), .A2(KEYINPUT116), .A3(new_n871), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n812), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  OR2_X1    g690(.A1(new_n870), .A2(new_n871), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n849), .B1(new_n826), .B2(new_n848), .ZN(new_n878));
  AND3_X1   g692(.A1(new_n877), .A2(new_n878), .A3(new_n812), .ZN(new_n879));
  OAI21_X1  g693(.A(KEYINPUT118), .B1(new_n876), .B2(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT118), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n877), .A2(new_n878), .A3(new_n812), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n870), .A2(KEYINPUT116), .A3(new_n871), .ZN(new_n883));
  AOI21_X1  g697(.A(KEYINPUT116), .B1(new_n870), .B2(new_n871), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n883), .A2(new_n884), .A3(new_n850), .ZN(new_n885));
  OAI211_X1 g699(.A(new_n881), .B(new_n882), .C1(new_n885), .C2(new_n812), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n811), .B1(new_n880), .B2(new_n886), .ZN(new_n887));
  NOR2_X1   g701(.A1(G952), .A2(G953), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n779), .B1(new_n887), .B2(new_n888), .ZN(G75));
  AOI21_X1  g703(.A(new_n349), .B1(new_n877), .B2(new_n878), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n890), .A2(KEYINPUT122), .A3(G210), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT56), .ZN(new_n892));
  AND2_X1   g706(.A1(new_n410), .A2(new_n412), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n893), .B(new_n420), .ZN(new_n894));
  XOR2_X1   g708(.A(new_n894), .B(KEYINPUT55), .Z(new_n895));
  NAND3_X1  g709(.A1(new_n891), .A2(new_n892), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g710(.A(KEYINPUT122), .B1(new_n890), .B2(G210), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n260), .A2(G952), .ZN(new_n899));
  INV_X1    g713(.A(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(KEYINPUT56), .B1(new_n890), .B2(G210), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n900), .B1(new_n901), .B2(new_n895), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n898), .A2(new_n902), .ZN(G51));
  AOI21_X1  g717(.A(new_n812), .B1(new_n877), .B2(new_n878), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n879), .A2(new_n904), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n586), .B(KEYINPUT123), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(KEYINPUT57), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n583), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n890), .A2(new_n754), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n899), .B1(new_n908), .B2(new_n909), .ZN(G54));
  AND3_X1   g724(.A1(new_n890), .A2(KEYINPUT58), .A3(G475), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n525), .A2(new_n530), .ZN(new_n912));
  INV_X1    g726(.A(new_n912), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n900), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n914), .B1(new_n913), .B2(new_n911), .ZN(G60));
  NAND2_X1  g729(.A1(new_n602), .A2(new_n606), .ZN(new_n916));
  NAND2_X1  g730(.A1(G478), .A2(G902), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(KEYINPUT59), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n900), .B1(new_n905), .B2(new_n919), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n880), .A2(new_n886), .A3(new_n918), .ZN(new_n921));
  INV_X1    g735(.A(new_n916), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n920), .B1(new_n921), .B2(new_n922), .ZN(G63));
  NAND2_X1  g737(.A1(new_n877), .A2(new_n878), .ZN(new_n924));
  NAND2_X1  g738(.A1(G217), .A2(G902), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n925), .B(KEYINPUT60), .Z(new_n926));
  NAND2_X1  g740(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(new_n361), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n628), .B(KEYINPUT124), .Z(new_n930));
  NAND3_X1  g744(.A1(new_n924), .A2(new_n926), .A3(new_n930), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n929), .A2(new_n900), .A3(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT61), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n929), .A2(KEYINPUT61), .A3(new_n900), .A4(new_n931), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n934), .A2(new_n935), .ZN(G66));
  AOI21_X1  g750(.A(new_n260), .B1(new_n447), .B2(G224), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n823), .A2(new_n824), .A3(new_n825), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n937), .B1(new_n938), .B2(new_n260), .ZN(new_n939));
  INV_X1    g753(.A(G898), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n893), .B1(new_n940), .B2(G953), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n939), .B(new_n941), .ZN(G69));
  AOI21_X1  g756(.A(new_n260), .B1(G227), .B2(G900), .ZN(new_n943));
  INV_X1    g757(.A(new_n943), .ZN(new_n944));
  OR2_X1    g758(.A1(new_n944), .A2(KEYINPUT126), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n761), .A2(new_n725), .A3(new_n827), .ZN(new_n946));
  OR2_X1    g760(.A1(new_n946), .A2(KEYINPUT125), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n946), .A2(KEYINPUT125), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  AND3_X1   g763(.A1(new_n855), .A2(new_n680), .A3(new_n857), .ZN(new_n950));
  AND3_X1   g764(.A1(new_n949), .A2(new_n771), .A3(new_n950), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n762), .A2(new_n732), .A3(new_n737), .A4(new_n951), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n952), .A2(G953), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n254), .A2(new_n257), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n511), .A2(new_n512), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n954), .B(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(G900), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n956), .B1(new_n957), .B2(new_n260), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n675), .A2(new_n950), .ZN(new_n959));
  OR2_X1    g773(.A1(new_n959), .A2(KEYINPUT62), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n959), .A2(KEYINPUT62), .ZN(new_n961));
  AOI211_X1 g775(.A(new_n739), .B(new_n654), .C1(new_n614), .C2(new_n622), .ZN(new_n962));
  AOI22_X1  g776(.A1(new_n769), .A2(new_n770), .B1(new_n683), .B2(new_n962), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n960), .A2(new_n762), .A3(new_n961), .A4(new_n963), .ZN(new_n964));
  AND2_X1   g778(.A1(new_n964), .A2(new_n260), .ZN(new_n965));
  OAI221_X1 g779(.A(new_n945), .B1(new_n953), .B2(new_n958), .C1(new_n965), .C2(new_n956), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n944), .A2(KEYINPUT126), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n966), .B(new_n967), .ZN(G72));
  NAND2_X1  g782(.A1(G472), .A2(G902), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n969), .B(KEYINPUT63), .Z(new_n970));
  OAI21_X1  g784(.A(new_n970), .B1(new_n964), .B2(new_n938), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n971), .A2(new_n264), .A3(new_n663), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n970), .B1(new_n952), .B2(new_n938), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n300), .B(KEYINPUT127), .Z(new_n974));
  AOI21_X1  g788(.A(new_n899), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n972), .A2(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(new_n885), .ZN(new_n977));
  AND3_X1   g791(.A1(new_n664), .A2(new_n300), .A3(new_n970), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n976), .B1(new_n977), .B2(new_n978), .ZN(G57));
endmodule


