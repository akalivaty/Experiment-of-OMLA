//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 1 0 0 0 1 0 0 0 1 0 0 0 1 1 1 0 1 0 1 1 1 0 1 1 1 1 0 1 0 0 0 1 0 1 1 1 0 1 0 0 1 0 1 1 0 1 0 1 1 1 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:30 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n622,
    new_n623, new_n624, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n777, new_n778, new_n779, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n888, new_n889, new_n890, new_n891,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956;
  XOR2_X1   g000(.A(KEYINPUT9), .B(G234), .Z(new_n187));
  XNOR2_X1  g001(.A(new_n187), .B(KEYINPUT76), .ZN(new_n188));
  OAI21_X1  g002(.A(G221), .B1(new_n188), .B2(G902), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n189), .B(KEYINPUT77), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT78), .ZN(new_n191));
  INV_X1    g005(.A(G104), .ZN(new_n192));
  OAI21_X1  g006(.A(new_n191), .B1(new_n192), .B2(G107), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(G107), .ZN(new_n194));
  INV_X1    g008(.A(G107), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n195), .A2(KEYINPUT78), .A3(G104), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n193), .A2(new_n194), .A3(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G101), .ZN(new_n198));
  OAI21_X1  g012(.A(KEYINPUT3), .B1(new_n192), .B2(G107), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT3), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n200), .A2(new_n195), .A3(G104), .ZN(new_n201));
  INV_X1    g015(.A(G101), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n199), .A2(new_n201), .A3(new_n202), .A4(new_n194), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n198), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(KEYINPUT79), .ZN(new_n205));
  INV_X1    g019(.A(G143), .ZN(new_n206));
  OAI21_X1  g020(.A(KEYINPUT1), .B1(new_n206), .B2(G146), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G128), .ZN(new_n208));
  XNOR2_X1  g022(.A(G143), .B(G146), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n206), .A2(G146), .ZN(new_n211));
  INV_X1    g025(.A(G146), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n212), .A2(G143), .ZN(new_n213));
  OAI211_X1 g027(.A(G128), .B(new_n207), .C1(new_n211), .C2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n210), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT79), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n198), .A2(new_n216), .A3(new_n203), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n205), .A2(new_n215), .A3(new_n217), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n198), .A2(new_n210), .A3(new_n214), .A4(new_n203), .ZN(new_n219));
  AND2_X1   g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(G134), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G137), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n221), .A2(G137), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT11), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n224), .A2(KEYINPUT64), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n222), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G137), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(G134), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT64), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(KEYINPUT11), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n224), .A2(KEYINPUT64), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n228), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  NOR3_X1   g046(.A1(new_n226), .A2(new_n232), .A3(G131), .ZN(new_n233));
  INV_X1    g047(.A(G131), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n227), .A2(G134), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n235), .B1(new_n228), .B2(new_n230), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n229), .A2(KEYINPUT11), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n223), .B1(new_n225), .B2(new_n237), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n234), .B1(new_n236), .B2(new_n238), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n233), .A2(new_n239), .ZN(new_n240));
  OAI21_X1  g054(.A(KEYINPUT12), .B1(new_n220), .B2(new_n240), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n240), .B1(new_n218), .B2(new_n219), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT12), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n210), .A2(KEYINPUT10), .A3(new_n214), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n217), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n216), .B1(new_n198), .B2(new_n203), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n246), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT10), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n219), .A2(new_n250), .ZN(new_n251));
  AND2_X1   g065(.A1(KEYINPUT0), .A2(G128), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n209), .A2(new_n252), .ZN(new_n253));
  XNOR2_X1  g067(.A(KEYINPUT0), .B(G128), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n253), .B1(new_n209), .B2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n199), .A2(new_n201), .A3(new_n194), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G101), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n258), .A2(KEYINPUT4), .A3(new_n203), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n257), .A2(new_n260), .A3(G101), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n256), .A2(new_n259), .A3(new_n261), .ZN(new_n262));
  NAND4_X1  g076(.A1(new_n249), .A2(new_n240), .A3(new_n251), .A4(new_n262), .ZN(new_n263));
  XNOR2_X1  g077(.A(G110), .B(G140), .ZN(new_n264));
  INV_X1    g078(.A(G227), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n265), .A2(G953), .ZN(new_n266));
  XNOR2_X1  g080(.A(new_n264), .B(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  NAND4_X1  g082(.A1(new_n241), .A2(new_n244), .A3(new_n263), .A4(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(new_n240), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n262), .A2(new_n251), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n245), .B1(new_n205), .B2(new_n217), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n270), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT80), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n273), .A2(new_n263), .A3(new_n274), .ZN(new_n275));
  OAI211_X1 g089(.A(KEYINPUT80), .B(new_n270), .C1(new_n271), .C2(new_n272), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n275), .A2(new_n267), .A3(new_n276), .ZN(new_n277));
  AOI211_X1 g091(.A(G469), .B(G902), .C1(new_n269), .C2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(G469), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n275), .A2(new_n276), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(new_n268), .ZN(new_n281));
  INV_X1    g095(.A(new_n244), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n263), .B1(new_n242), .B2(new_n243), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n267), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n281), .A2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(G902), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n279), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT81), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n278), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(G902), .B1(new_n281), .B2(new_n284), .ZN(new_n290));
  OAI21_X1  g104(.A(KEYINPUT81), .B1(new_n290), .B2(new_n279), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n190), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT89), .ZN(new_n293));
  INV_X1    g107(.A(G237), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(KEYINPUT68), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT68), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(G237), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(G953), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n298), .A2(G214), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(new_n206), .ZN(new_n301));
  AOI21_X1  g115(.A(G953), .B1(new_n295), .B2(new_n297), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n302), .A2(G143), .A3(G214), .ZN(new_n303));
  NAND2_X1  g117(.A1(KEYINPUT18), .A2(G131), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n301), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT85), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND4_X1  g121(.A1(new_n301), .A2(KEYINPUT85), .A3(new_n303), .A4(new_n304), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n301), .A2(new_n303), .ZN(new_n310));
  INV_X1    g124(.A(new_n304), .ZN(new_n311));
  INV_X1    g125(.A(G140), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(G125), .ZN(new_n313));
  INV_X1    g127(.A(G125), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(G140), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n313), .A2(new_n315), .A3(new_n212), .ZN(new_n316));
  AND3_X1   g130(.A1(new_n314), .A2(KEYINPUT73), .A3(G140), .ZN(new_n317));
  AOI21_X1  g131(.A(KEYINPUT73), .B1(new_n314), .B2(G140), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n313), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G146), .ZN(new_n320));
  AOI22_X1  g134(.A1(new_n310), .A2(new_n311), .B1(new_n316), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n309), .A2(new_n321), .ZN(new_n322));
  AND4_X1   g136(.A1(G143), .A2(new_n298), .A3(G214), .A4(new_n299), .ZN(new_n323));
  AOI21_X1  g137(.A(G143), .B1(new_n302), .B2(G214), .ZN(new_n324));
  OAI21_X1  g138(.A(G131), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT17), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n301), .A2(new_n234), .A3(new_n303), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n325), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n319), .A2(KEYINPUT16), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT16), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n313), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n212), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n314), .A2(G140), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT73), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n334), .B1(new_n312), .B2(G125), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n314), .A2(KEYINPUT73), .A3(G140), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n333), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  OAI211_X1 g151(.A(new_n212), .B(new_n331), .C1(new_n337), .C2(new_n330), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n332), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n310), .A2(KEYINPUT17), .A3(G131), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n328), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n322), .A2(new_n342), .ZN(new_n343));
  XNOR2_X1  g157(.A(G113), .B(G122), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n344), .B(new_n192), .ZN(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n343), .A2(new_n346), .ZN(new_n347));
  AOI211_X1 g161(.A(new_n326), .B(new_n234), .C1(new_n301), .C2(new_n303), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n331), .B1(new_n337), .B2(new_n330), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(G146), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(new_n338), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n348), .A2(new_n351), .ZN(new_n352));
  AOI22_X1  g166(.A1(new_n352), .A2(new_n328), .B1(new_n309), .B2(new_n321), .ZN(new_n353));
  OAI21_X1  g167(.A(KEYINPUT88), .B1(new_n353), .B2(new_n345), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT88), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n343), .A2(new_n355), .A3(new_n346), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n347), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n293), .B1(new_n357), .B2(G902), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n353), .A2(new_n345), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n355), .B1(new_n343), .B2(new_n346), .ZN(new_n360));
  AOI211_X1 g174(.A(KEYINPUT88), .B(new_n345), .C1(new_n322), .C2(new_n342), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n359), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n362), .A2(KEYINPUT89), .A3(new_n286), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n358), .A2(new_n363), .A3(G475), .ZN(new_n364));
  NOR2_X1   g178(.A1(G475), .A2(G902), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n325), .A2(new_n327), .ZN(new_n366));
  XOR2_X1   g180(.A(KEYINPUT86), .B(KEYINPUT19), .Z(new_n367));
  NAND3_X1  g181(.A1(new_n367), .A2(new_n313), .A3(new_n315), .ZN(new_n368));
  OR2_X1    g182(.A1(new_n368), .A2(KEYINPUT87), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n319), .A2(KEYINPUT19), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n368), .A2(KEYINPUT87), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n369), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  OAI211_X1 g186(.A(new_n366), .B(new_n350), .C1(new_n372), .C2(G146), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n345), .B1(new_n322), .B2(new_n373), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n365), .B1(new_n347), .B2(new_n374), .ZN(new_n375));
  XNOR2_X1  g189(.A(new_n375), .B(KEYINPUT20), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n364), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(G128), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n378), .A2(G143), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n206), .A2(G128), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  XNOR2_X1  g195(.A(new_n381), .B(new_n221), .ZN(new_n382));
  INV_X1    g196(.A(G116), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n383), .A2(KEYINPUT14), .A3(G122), .ZN(new_n384));
  XNOR2_X1  g198(.A(G116), .B(G122), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  OAI211_X1 g200(.A(G107), .B(new_n384), .C1(new_n386), .C2(KEYINPUT14), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n385), .A2(new_n195), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n382), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT90), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n382), .A2(KEYINPUT90), .A3(new_n387), .A4(new_n388), .ZN(new_n392));
  XNOR2_X1  g206(.A(new_n385), .B(new_n195), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n381), .A2(new_n221), .ZN(new_n394));
  AND2_X1   g208(.A1(new_n379), .A2(KEYINPUT13), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n379), .A2(KEYINPUT13), .ZN(new_n396));
  NOR3_X1   g210(.A1(new_n395), .A2(new_n396), .A3(new_n380), .ZN(new_n397));
  OAI211_X1 g211(.A(new_n393), .B(new_n394), .C1(new_n397), .C2(new_n221), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n391), .A2(new_n392), .A3(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(G217), .ZN(new_n400));
  NOR3_X1   g214(.A1(new_n188), .A2(new_n400), .A3(G953), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n399), .A2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT91), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n391), .A2(new_n392), .A3(new_n398), .A4(new_n401), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n403), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n399), .A2(KEYINPUT91), .A3(new_n402), .ZN(new_n407));
  NAND4_X1  g221(.A1(new_n406), .A2(KEYINPUT92), .A3(new_n286), .A4(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(G478), .ZN(new_n409));
  OR2_X1    g223(.A1(new_n409), .A2(KEYINPUT15), .ZN(new_n410));
  XNOR2_X1  g224(.A(new_n408), .B(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n377), .A2(new_n412), .ZN(new_n413));
  AND2_X1   g227(.A1(new_n299), .A2(G952), .ZN(new_n414));
  NAND2_X1  g228(.A1(G234), .A2(G237), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n416), .B(KEYINPUT93), .ZN(new_n417));
  XNOR2_X1  g231(.A(KEYINPUT21), .B(G898), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n415), .A2(G902), .A3(G953), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n417), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  OAI21_X1  g235(.A(G214), .B1(G237), .B2(G902), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n383), .A2(G119), .ZN(new_n424));
  INV_X1    g238(.A(G119), .ZN(new_n425));
  OAI21_X1  g239(.A(KEYINPUT65), .B1(new_n425), .B2(G116), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT65), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n427), .A2(new_n383), .A3(G119), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n424), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  AND2_X1   g243(.A1(new_n429), .A2(KEYINPUT5), .ZN(new_n430));
  INV_X1    g244(.A(new_n424), .ZN(new_n431));
  OAI21_X1  g245(.A(G113), .B1(new_n431), .B2(KEYINPUT5), .ZN(new_n432));
  OR2_X1    g246(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  XNOR2_X1  g247(.A(KEYINPUT2), .B(G113), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n429), .A2(new_n435), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n433), .B(new_n436), .C1(new_n247), .C2(new_n248), .ZN(new_n437));
  XNOR2_X1  g251(.A(G110), .B(G122), .ZN(new_n438));
  AND2_X1   g252(.A1(new_n429), .A2(new_n435), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n429), .A2(new_n435), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT66), .ZN(new_n441));
  NOR3_X1   g255(.A1(new_n439), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n426), .A2(new_n428), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(new_n431), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(new_n434), .ZN(new_n445));
  AOI21_X1  g259(.A(KEYINPUT66), .B1(new_n445), .B2(new_n436), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n442), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n259), .A2(new_n261), .ZN(new_n448));
  OAI211_X1 g262(.A(new_n437), .B(new_n438), .C1(new_n447), .C2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(new_n438), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n436), .B1(new_n430), .B2(new_n432), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n451), .B1(new_n205), .B2(new_n217), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n441), .B1(new_n439), .B2(new_n440), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n445), .A2(KEYINPUT66), .A3(new_n436), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n448), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n450), .B1(new_n452), .B2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT82), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT6), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n449), .A2(new_n456), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n299), .A2(G224), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n461), .B(KEYINPUT84), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n462), .B(KEYINPUT83), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n210), .A2(new_n314), .A3(new_n214), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n464), .B1(new_n255), .B2(new_n314), .ZN(new_n465));
  XNOR2_X1  g279(.A(new_n463), .B(new_n465), .ZN(new_n466));
  OAI221_X1 g280(.A(new_n450), .B1(new_n457), .B2(new_n458), .C1(new_n452), .C2(new_n455), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n460), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  AND2_X1   g282(.A1(new_n462), .A2(KEYINPUT7), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n465), .B(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n451), .A2(new_n204), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n437), .A2(new_n471), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n438), .B(KEYINPUT8), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n470), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(G902), .B1(new_n474), .B2(new_n449), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n468), .A2(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(G210), .B1(G237), .B2(G902), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n468), .A2(new_n475), .A3(new_n477), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n423), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  AND4_X1   g295(.A1(new_n292), .A2(new_n413), .A3(new_n421), .A4(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT75), .ZN(new_n483));
  XNOR2_X1  g297(.A(KEYINPUT22), .B(G137), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n299), .A2(G221), .A3(G234), .ZN(new_n485));
  XNOR2_X1  g299(.A(new_n484), .B(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n378), .A2(G119), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n425), .A2(G128), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT71), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(KEYINPUT71), .B1(new_n425), .B2(G128), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n488), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  XNOR2_X1  g307(.A(KEYINPUT24), .B(G110), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(G110), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n425), .A2(G128), .ZN(new_n497));
  OAI21_X1  g311(.A(KEYINPUT23), .B1(new_n378), .B2(G119), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT72), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NOR3_X1   g314(.A1(new_n488), .A2(KEYINPUT72), .A3(KEYINPUT23), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n496), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n495), .A2(new_n502), .ZN(new_n503));
  AND3_X1   g317(.A1(new_n503), .A2(new_n350), .A3(new_n316), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT23), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n497), .A2(new_n499), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(KEYINPUT72), .B1(new_n489), .B2(KEYINPUT23), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n506), .B1(new_n507), .B2(new_n497), .ZN(new_n508));
  OAI22_X1  g322(.A1(new_n508), .A2(new_n496), .B1(new_n493), .B2(new_n494), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n509), .B1(new_n338), .B2(new_n350), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n487), .B1(new_n504), .B2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(new_n509), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n351), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n503), .A2(new_n350), .A3(new_n316), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n513), .A2(new_n514), .A3(new_n486), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n511), .A2(new_n286), .A3(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT74), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n517), .A2(KEYINPUT25), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n518), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n511), .A2(new_n286), .A3(new_n515), .A4(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n400), .B1(G234), .B2(new_n286), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n483), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(new_n523), .ZN(new_n525));
  AOI211_X1 g339(.A(KEYINPUT75), .B(new_n525), .C1(new_n519), .C2(new_n521), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  AND2_X1   g341(.A1(new_n511), .A2(new_n515), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n523), .A2(G902), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n527), .A2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(G472), .ZN(new_n532));
  INV_X1    g346(.A(new_n447), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n236), .A2(new_n238), .A3(new_n234), .ZN(new_n534));
  OAI21_X1  g348(.A(G131), .B1(new_n223), .B2(new_n235), .ZN(new_n535));
  AND4_X1   g349(.A1(new_n534), .A2(new_n210), .A3(new_n214), .A4(new_n535), .ZN(new_n536));
  OAI21_X1  g350(.A(G131), .B1(new_n226), .B2(new_n232), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n255), .B1(new_n537), .B2(new_n534), .ZN(new_n538));
  NOR3_X1   g352(.A1(new_n536), .A2(new_n538), .A3(KEYINPUT30), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT30), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n256), .B1(new_n233), .B2(new_n239), .ZN(new_n541));
  NAND4_X1  g355(.A1(new_n534), .A2(new_n210), .A3(new_n214), .A4(new_n535), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n533), .B1(new_n539), .B2(new_n543), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n536), .A2(new_n538), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT67), .ZN(new_n546));
  NOR3_X1   g360(.A1(new_n442), .A2(new_n446), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g361(.A(KEYINPUT67), .B1(new_n453), .B2(new_n454), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n545), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n302), .A2(G210), .ZN(new_n550));
  XNOR2_X1  g364(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n551));
  XNOR2_X1  g365(.A(new_n550), .B(new_n551), .ZN(new_n552));
  XNOR2_X1  g366(.A(KEYINPUT26), .B(G101), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n552), .B(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n544), .A2(new_n549), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(KEYINPUT31), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT31), .ZN(new_n557));
  NAND4_X1  g371(.A1(new_n544), .A2(new_n549), .A3(new_n557), .A4(new_n554), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n541), .A2(new_n542), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n546), .B1(new_n442), .B2(new_n446), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n453), .A2(KEYINPUT67), .A3(new_n454), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n560), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n545), .A2(new_n447), .ZN(new_n564));
  OAI21_X1  g378(.A(KEYINPUT28), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT28), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n547), .A2(new_n548), .ZN(new_n567));
  OAI21_X1  g381(.A(KEYINPUT70), .B1(new_n536), .B2(new_n538), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT70), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n541), .A2(new_n569), .A3(new_n542), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n566), .B1(new_n567), .B2(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n554), .B1(new_n565), .B2(new_n572), .ZN(new_n573));
  OAI211_X1 g387(.A(new_n532), .B(new_n286), .C1(new_n559), .C2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(KEYINPUT32), .ZN(new_n575));
  INV_X1    g389(.A(new_n554), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n533), .A2(new_n560), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n566), .B1(new_n549), .B2(new_n577), .ZN(new_n578));
  AND2_X1   g392(.A1(new_n568), .A2(new_n570), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n561), .A2(new_n562), .ZN(new_n580));
  AOI21_X1  g394(.A(KEYINPUT28), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n576), .B1(new_n578), .B2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n582), .A2(new_n556), .A3(new_n558), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT32), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n583), .A2(new_n584), .A3(new_n532), .A4(new_n286), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n575), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT29), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n576), .B1(new_n565), .B2(new_n572), .ZN(new_n588));
  INV_X1    g402(.A(new_n544), .ZN(new_n589));
  NOR3_X1   g403(.A1(new_n589), .A2(new_n563), .A3(new_n554), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n587), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n561), .A2(new_n560), .A3(new_n562), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n566), .B1(new_n549), .B2(new_n592), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n593), .A2(new_n581), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n576), .A2(new_n587), .ZN(new_n595));
  AOI21_X1  g409(.A(G902), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n591), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(G472), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n531), .B1(new_n586), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n482), .A2(new_n599), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n600), .B(G101), .ZN(G3));
  NAND2_X1  g415(.A1(new_n574), .A2(KEYINPUT94), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n286), .B1(new_n559), .B2(new_n573), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(G472), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n602), .B(new_n604), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n605), .A2(new_n531), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT33), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n406), .A2(new_n607), .A3(new_n407), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n403), .A2(KEYINPUT33), .A3(new_n405), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n409), .A2(G902), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n406), .A2(new_n286), .A3(new_n407), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(new_n409), .ZN(new_n613));
  AND2_X1   g427(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n614), .B1(new_n364), .B2(new_n376), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n481), .A2(new_n421), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n606), .A2(new_n292), .A3(new_n618), .ZN(new_n619));
  XOR2_X1   g433(.A(KEYINPUT34), .B(G104), .Z(new_n620));
  XNOR2_X1  g434(.A(new_n619), .B(new_n620), .ZN(G6));
  NOR3_X1   g435(.A1(new_n617), .A2(new_n377), .A3(new_n411), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n606), .A2(new_n292), .A3(new_n622), .ZN(new_n623));
  XOR2_X1   g437(.A(KEYINPUT35), .B(G107), .Z(new_n624));
  XNOR2_X1  g438(.A(new_n623), .B(new_n624), .ZN(G9));
  INV_X1    g439(.A(new_n605), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n513), .A2(new_n514), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n487), .A2(KEYINPUT36), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n627), .B(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(new_n529), .ZN(new_n630));
  AOI21_X1  g444(.A(KEYINPUT95), .B1(new_n527), .B2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT95), .ZN(new_n632));
  INV_X1    g446(.A(new_n630), .ZN(new_n633));
  NOR4_X1   g447(.A1(new_n524), .A2(new_n526), .A3(new_n632), .A4(new_n633), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n626), .A2(KEYINPUT96), .A3(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT96), .ZN(new_n637));
  INV_X1    g451(.A(new_n635), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n637), .B1(new_n638), .B2(new_n605), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n636), .A2(new_n639), .A3(new_n482), .ZN(new_n640));
  XOR2_X1   g454(.A(KEYINPUT37), .B(G110), .Z(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(G12));
  NAND2_X1  g456(.A1(new_n586), .A2(new_n598), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n635), .A2(new_n292), .A3(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n377), .ZN(new_n645));
  INV_X1    g459(.A(G900), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n415), .A2(new_n646), .A3(G902), .A4(G953), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(KEYINPUT97), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n417), .A2(new_n648), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n645), .A2(new_n412), .A3(new_n481), .A4(new_n649), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n644), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(new_n378), .ZN(G30));
  XOR2_X1   g466(.A(KEYINPUT99), .B(KEYINPUT39), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n649), .B(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n292), .A2(new_n654), .ZN(new_n655));
  OR2_X1    g469(.A1(new_n655), .A2(KEYINPUT40), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n589), .A2(new_n563), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n657), .A2(new_n576), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n576), .A2(new_n549), .A3(new_n592), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(new_n286), .ZN(new_n660));
  OAI21_X1  g474(.A(G472), .B1(new_n658), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n586), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n645), .A2(new_n411), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n479), .A2(new_n480), .ZN(new_n664));
  XNOR2_X1  g478(.A(KEYINPUT98), .B(KEYINPUT38), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n522), .A2(new_n523), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(KEYINPUT75), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n522), .A2(new_n483), .A3(new_n523), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n668), .A2(new_n669), .A3(new_n630), .ZN(new_n670));
  NOR3_X1   g484(.A1(new_n666), .A2(new_n423), .A3(new_n670), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n656), .A2(new_n662), .A3(new_n663), .A4(new_n671), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n672), .B1(KEYINPUT40), .B2(new_n655), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT100), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(new_n206), .ZN(G45));
  INV_X1    g490(.A(KEYINPUT102), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT101), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n615), .A2(new_n678), .A3(new_n481), .A4(new_n649), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n679), .A2(new_n643), .A3(new_n292), .A4(new_n635), .ZN(new_n680));
  INV_X1    g494(.A(new_n649), .ZN(new_n681));
  AOI211_X1 g495(.A(new_n681), .B(new_n614), .C1(new_n364), .C2(new_n376), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n678), .B1(new_n682), .B2(new_n481), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n677), .B1(new_n680), .B2(new_n683), .ZN(new_n684));
  AND3_X1   g498(.A1(new_n635), .A2(new_n292), .A3(new_n643), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n615), .A2(new_n481), .A3(new_n649), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(KEYINPUT101), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n685), .A2(KEYINPUT102), .A3(new_n687), .A4(new_n679), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n684), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(KEYINPUT103), .B(G146), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(G48));
  INV_X1    g505(.A(new_n531), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n643), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n269), .A2(new_n277), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n279), .B1(new_n694), .B2(new_n286), .ZN(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(new_n190), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n694), .A2(new_n279), .A3(new_n286), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n696), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n693), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(new_n618), .ZN(new_n701));
  XNOR2_X1  g515(.A(KEYINPUT41), .B(G113), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n701), .B(new_n702), .ZN(G15));
  NAND2_X1  g517(.A1(new_n700), .A2(new_n622), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G116), .ZN(G18));
  AND2_X1   g519(.A1(new_n413), .A2(new_n421), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT104), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n664), .A2(new_n422), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n707), .B1(new_n708), .B2(new_n699), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n695), .A2(new_n278), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n481), .A2(new_n710), .A3(KEYINPUT104), .A4(new_n697), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n706), .A2(new_n643), .A3(new_n712), .A4(new_n635), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G119), .ZN(G21));
  OAI211_X1 g528(.A(new_n556), .B(new_n558), .C1(new_n594), .C2(new_n554), .ZN(new_n715));
  NOR2_X1   g529(.A1(G472), .A2(G902), .ZN(new_n716));
  AOI22_X1  g530(.A1(new_n603), .A2(G472), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  AND3_X1   g531(.A1(new_n717), .A2(new_n527), .A3(new_n530), .ZN(new_n718));
  INV_X1    g532(.A(new_n699), .ZN(new_n719));
  AND3_X1   g533(.A1(new_n718), .A2(new_n421), .A3(new_n719), .ZN(new_n720));
  AND3_X1   g534(.A1(new_n377), .A2(new_n412), .A3(new_n481), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G122), .ZN(G24));
  INV_X1    g537(.A(KEYINPUT106), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n715), .A2(new_n716), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n670), .A2(new_n604), .A3(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT105), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  AOI21_X1  g542(.A(KEYINPUT105), .B1(new_n717), .B2(new_n670), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n682), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  AND2_X1   g544(.A1(new_n709), .A2(new_n711), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n724), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n726), .B(new_n727), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n733), .A2(KEYINPUT106), .A3(new_n682), .A4(new_n712), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G125), .ZN(G27));
  NAND2_X1  g550(.A1(new_n285), .A2(KEYINPUT107), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT107), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n281), .A2(new_n738), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n737), .A2(G469), .A3(new_n739), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n279), .A2(new_n286), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n278), .A2(new_n741), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n190), .B1(new_n740), .B2(new_n742), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n664), .A2(new_n423), .ZN(new_n744));
  AND2_X1   g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n745), .A2(new_n599), .A3(new_n682), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT108), .ZN(new_n747));
  AND3_X1   g561(.A1(new_n746), .A2(new_n747), .A3(KEYINPUT42), .ZN(new_n748));
  AOI21_X1  g562(.A(KEYINPUT42), .B1(new_n746), .B2(new_n747), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G131), .ZN(G33));
  NAND3_X1  g565(.A1(new_n645), .A2(new_n412), .A3(new_n649), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT109), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n645), .A2(KEYINPUT109), .A3(new_n412), .A4(new_n649), .ZN(new_n755));
  AND4_X1   g569(.A1(new_n599), .A2(new_n754), .A3(new_n745), .A4(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(new_n221), .ZN(G36));
  INV_X1    g571(.A(new_n744), .ZN(new_n758));
  INV_X1    g572(.A(new_n614), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n645), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(KEYINPUT43), .ZN(new_n761));
  AOI211_X1 g575(.A(new_n626), .B(new_n761), .C1(new_n527), .C2(new_n630), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n758), .B1(new_n762), .B2(KEYINPUT44), .ZN(new_n763));
  AND2_X1   g577(.A1(new_n281), .A2(new_n284), .ZN(new_n764));
  OAI21_X1  g578(.A(G469), .B1(new_n764), .B2(KEYINPUT45), .ZN(new_n765));
  AND2_X1   g579(.A1(new_n737), .A2(new_n739), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n765), .B1(new_n766), .B2(KEYINPUT45), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n767), .A2(new_n741), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n768), .A2(KEYINPUT46), .ZN(new_n769));
  OR2_X1    g583(.A1(new_n769), .A2(KEYINPUT110), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(KEYINPUT110), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n278), .B1(new_n768), .B2(KEYINPUT46), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n770), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  AND3_X1   g587(.A1(new_n773), .A2(new_n697), .A3(new_n654), .ZN(new_n774));
  OAI211_X1 g588(.A(new_n763), .B(new_n774), .C1(KEYINPUT44), .C2(new_n762), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G137), .ZN(G39));
  NAND2_X1  g590(.A1(new_n773), .A2(new_n697), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT47), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NOR3_X1   g593(.A1(new_n643), .A2(new_n758), .A3(new_n692), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n779), .A2(new_n682), .A3(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G140), .ZN(G42));
  INV_X1    g596(.A(KEYINPUT53), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n527), .A2(new_n630), .A3(new_n649), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n784), .B1(new_n586), .B2(new_n661), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n721), .A2(new_n785), .A3(new_n743), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(KEYINPUT112), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT112), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n721), .A2(new_n785), .A3(new_n788), .A4(new_n743), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n651), .B1(new_n787), .B2(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n689), .A2(new_n735), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(KEYINPUT52), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT52), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n689), .A2(new_n735), .A3(new_n790), .A4(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  NOR3_X1   g609(.A1(new_n756), .A2(new_n748), .A3(new_n749), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n640), .A2(new_n623), .A3(new_n713), .ZN(new_n797));
  INV_X1    g611(.A(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n701), .A2(new_n704), .A3(new_n722), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n600), .A2(new_n619), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n685), .A2(new_n413), .A3(new_n649), .A4(new_n744), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n733), .A2(new_n682), .A3(new_n745), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n796), .A2(new_n798), .A3(new_n801), .A4(new_n804), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n783), .B1(new_n795), .B2(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT113), .ZN(new_n807));
  AND3_X1   g621(.A1(new_n792), .A2(new_n807), .A3(new_n794), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n807), .B1(new_n792), .B2(new_n794), .ZN(new_n809));
  NOR3_X1   g623(.A1(new_n808), .A2(new_n809), .A3(new_n805), .ZN(new_n810));
  INV_X1    g624(.A(new_n810), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n806), .B1(new_n811), .B2(new_n783), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n812), .A2(KEYINPUT54), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n761), .A2(new_n417), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(new_n718), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n666), .A2(new_n719), .A3(new_n423), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(KEYINPUT50), .ZN(new_n818));
  INV_X1    g632(.A(new_n662), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n758), .A2(new_n699), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n531), .A2(new_n417), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n819), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n822), .A2(new_n377), .A3(new_n759), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n814), .A2(new_n820), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n823), .B1(new_n824), .B2(new_n733), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n818), .A2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT114), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n815), .A2(new_n758), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n695), .A2(new_n278), .A3(new_n697), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n829), .B1(new_n779), .B2(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n818), .A2(KEYINPUT114), .A3(new_n825), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n828), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT51), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT54), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n795), .A2(new_n805), .A3(new_n783), .ZN(new_n837));
  INV_X1    g651(.A(new_n837), .ZN(new_n838));
  OAI211_X1 g652(.A(new_n836), .B(new_n838), .C1(new_n810), .C2(KEYINPUT53), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n815), .A2(new_n731), .ZN(new_n840));
  XOR2_X1   g654(.A(new_n840), .B(KEYINPUT115), .Z(new_n841));
  NAND2_X1  g655(.A1(new_n824), .A2(new_n599), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n842), .B(KEYINPUT48), .ZN(new_n843));
  OR2_X1    g657(.A1(new_n822), .A2(new_n616), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n841), .A2(new_n843), .A3(new_n414), .A4(new_n844), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n826), .A2(new_n834), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n845), .B1(new_n846), .B2(new_n831), .ZN(new_n847));
  AND4_X1   g661(.A1(new_n813), .A2(new_n835), .A3(new_n839), .A4(new_n847), .ZN(new_n848));
  NOR2_X1   g662(.A1(G952), .A2(G953), .ZN(new_n849));
  NOR4_X1   g663(.A1(new_n760), .A2(new_n531), .A3(new_n190), .A4(new_n423), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n850), .A2(KEYINPUT111), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(KEYINPUT111), .ZN(new_n852));
  XNOR2_X1  g666(.A(new_n710), .B(KEYINPUT49), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n852), .A2(new_n819), .A3(new_n666), .A4(new_n853), .ZN(new_n854));
  OAI22_X1  g668(.A1(new_n848), .A2(new_n849), .B1(new_n851), .B2(new_n854), .ZN(G75));
  NOR2_X1   g669(.A1(new_n299), .A2(G952), .ZN(new_n856));
  INV_X1    g670(.A(new_n856), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n805), .B1(new_n795), .B2(KEYINPUT113), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n792), .A2(new_n807), .A3(new_n794), .ZN(new_n859));
  AOI21_X1  g673(.A(KEYINPUT53), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n860), .A2(new_n837), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n861), .A2(new_n286), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n862), .A2(G210), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT56), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n460), .A2(new_n467), .ZN(new_n866));
  XNOR2_X1  g680(.A(new_n866), .B(new_n466), .ZN(new_n867));
  XOR2_X1   g681(.A(new_n867), .B(KEYINPUT55), .Z(new_n868));
  OAI21_X1  g682(.A(new_n857), .B1(new_n865), .B2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT116), .ZN(new_n870));
  AOI21_X1  g684(.A(KEYINPUT56), .B1(new_n862), .B2(G210), .ZN(new_n871));
  INV_X1    g685(.A(new_n868), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n870), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n865), .A2(KEYINPUT116), .A3(new_n868), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n869), .B1(new_n873), .B2(new_n874), .ZN(G51));
  OAI21_X1  g689(.A(KEYINPUT54), .B1(new_n860), .B2(new_n837), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n876), .A2(new_n839), .A3(KEYINPUT117), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT117), .ZN(new_n878));
  OAI211_X1 g692(.A(new_n878), .B(KEYINPUT54), .C1(new_n860), .C2(new_n837), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n741), .B(KEYINPUT57), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n877), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT118), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n877), .A2(KEYINPUT118), .A3(new_n879), .A4(new_n880), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n883), .A2(new_n694), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n862), .A2(new_n767), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n856), .B1(new_n885), .B2(new_n886), .ZN(G54));
  NAND3_X1  g701(.A1(new_n862), .A2(KEYINPUT58), .A3(G475), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n347), .A2(new_n374), .ZN(new_n889));
  AND2_X1   g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n888), .A2(new_n889), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n890), .A2(new_n891), .A3(new_n856), .ZN(G60));
  NAND2_X1  g706(.A1(G478), .A2(G902), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n893), .B(KEYINPUT59), .Z(new_n894));
  AOI21_X1  g708(.A(new_n894), .B1(new_n813), .B2(new_n839), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n608), .A2(new_n609), .ZN(new_n896));
  INV_X1    g710(.A(new_n896), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n857), .B1(new_n895), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n877), .A2(new_n879), .ZN(new_n899));
  NOR3_X1   g713(.A1(new_n899), .A2(new_n896), .A3(new_n894), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n898), .A2(new_n900), .ZN(G63));
  NAND2_X1  g715(.A1(G217), .A2(G902), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(KEYINPUT60), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n861), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(new_n629), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n528), .B(KEYINPUT119), .Z(new_n906));
  INV_X1    g720(.A(new_n906), .ZN(new_n907));
  OAI211_X1 g721(.A(new_n905), .B(new_n857), .C1(new_n904), .C2(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT61), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n908), .B(new_n909), .ZN(G66));
  INV_X1    g724(.A(G224), .ZN(new_n911));
  OAI21_X1  g725(.A(G953), .B1(new_n418), .B2(new_n911), .ZN(new_n912));
  AOI22_X1  g726(.A1(new_n700), .A2(new_n618), .B1(new_n720), .B2(new_n721), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n913), .A2(new_n600), .A3(new_n619), .A4(new_n704), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n914), .A2(new_n797), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n912), .B1(new_n915), .B2(G953), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n866), .B1(G898), .B2(new_n299), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n916), .B(new_n917), .ZN(G69));
  AOI21_X1  g732(.A(new_n615), .B1(new_n645), .B2(new_n412), .ZN(new_n919));
  NOR4_X1   g733(.A1(new_n693), .A2(new_n655), .A3(new_n919), .A4(new_n758), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n920), .B(KEYINPUT123), .Z(new_n921));
  OAI211_X1 g735(.A(new_n689), .B(new_n735), .C1(new_n644), .C2(new_n650), .ZN(new_n922));
  OR2_X1    g736(.A1(new_n675), .A2(new_n922), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n921), .B1(new_n923), .B2(KEYINPUT62), .ZN(new_n924));
  AND2_X1   g738(.A1(new_n781), .A2(new_n775), .ZN(new_n925));
  OAI211_X1 g739(.A(new_n924), .B(new_n925), .C1(KEYINPUT62), .C2(new_n923), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n539), .A2(new_n543), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n372), .B(KEYINPUT122), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n927), .B(new_n928), .ZN(new_n929));
  XNOR2_X1  g743(.A(KEYINPUT120), .B(KEYINPUT121), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n929), .B(new_n930), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n931), .A2(G953), .ZN(new_n932));
  OAI21_X1  g746(.A(G953), .B1(new_n265), .B2(new_n646), .ZN(new_n933));
  AOI22_X1  g747(.A1(new_n926), .A2(new_n932), .B1(KEYINPUT124), .B2(new_n933), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n774), .A2(new_n599), .A3(new_n721), .ZN(new_n935));
  INV_X1    g749(.A(new_n796), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n936), .A2(new_n922), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n925), .A2(new_n935), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(new_n299), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n646), .A2(G953), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n939), .A2(new_n940), .A3(new_n931), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n934), .A2(new_n941), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n933), .A2(KEYINPUT124), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(KEYINPUT125), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n942), .B(new_n944), .ZN(G72));
  NAND2_X1  g759(.A1(G472), .A2(G902), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n946), .B(KEYINPUT63), .Z(new_n947));
  INV_X1    g761(.A(new_n915), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n947), .B1(new_n926), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(new_n658), .ZN(new_n950));
  INV_X1    g764(.A(new_n590), .ZN(new_n951));
  INV_X1    g765(.A(new_n658), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n812), .A2(new_n951), .A3(new_n952), .A4(new_n947), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n947), .B1(new_n938), .B2(new_n948), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n590), .B(KEYINPUT126), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n856), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  AND3_X1   g770(.A1(new_n950), .A2(new_n953), .A3(new_n956), .ZN(G57));
endmodule


