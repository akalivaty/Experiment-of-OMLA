

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X1 U555 ( .A1(n938), .A2(n634), .ZN(n633) );
  OR2_X1 U556 ( .A1(n705), .A2(n704), .ZN(n522) );
  INV_X1 U557 ( .A(KEYINPUT27), .ZN(n638) );
  XNOR2_X1 U558 ( .A(n639), .B(n638), .ZN(n640) );
  NOR2_X1 U559 ( .A1(n939), .A2(n645), .ZN(n646) );
  XNOR2_X1 U560 ( .A(KEYINPUT102), .B(n682), .ZN(n701) );
  AND2_X1 U561 ( .A1(n706), .A2(n522), .ZN(n707) );
  NOR2_X1 U562 ( .A1(G2104), .A2(G2105), .ZN(n523) );
  NOR2_X1 U563 ( .A1(G651), .A2(n595), .ZN(n798) );
  XOR2_X2 U564 ( .A(KEYINPUT17), .B(n523), .Z(n892) );
  NAND2_X1 U565 ( .A1(G137), .A2(n892), .ZN(n524) );
  XNOR2_X1 U566 ( .A(n524), .B(KEYINPUT64), .ZN(n533) );
  INV_X1 U567 ( .A(G2105), .ZN(n525) );
  NOR2_X1 U568 ( .A1(G2104), .A2(n525), .ZN(n888) );
  NAND2_X1 U569 ( .A1(G125), .A2(n888), .ZN(n527) );
  INV_X1 U570 ( .A(G2104), .ZN(n528) );
  NOR2_X1 U571 ( .A1(n528), .A2(n525), .ZN(n889) );
  NAND2_X1 U572 ( .A1(G113), .A2(n889), .ZN(n526) );
  AND2_X1 U573 ( .A1(n527), .A2(n526), .ZN(n531) );
  NOR2_X2 U574 ( .A1(G2105), .A2(n528), .ZN(n893) );
  NAND2_X1 U575 ( .A1(G101), .A2(n893), .ZN(n529) );
  XOR2_X1 U576 ( .A(KEYINPUT23), .B(n529), .Z(n530) );
  AND2_X1 U577 ( .A1(n531), .A2(n530), .ZN(n532) );
  AND2_X1 U578 ( .A1(n533), .A2(n532), .ZN(G160) );
  NOR2_X1 U579 ( .A1(G543), .A2(G651), .ZN(n793) );
  NAND2_X1 U580 ( .A1(n793), .A2(G86), .ZN(n534) );
  XNOR2_X1 U581 ( .A(n534), .B(KEYINPUT78), .ZN(n537) );
  INV_X1 U582 ( .A(G651), .ZN(n538) );
  NOR2_X1 U583 ( .A1(G543), .A2(n538), .ZN(n535) );
  XOR2_X1 U584 ( .A(KEYINPUT1), .B(n535), .Z(n794) );
  NAND2_X1 U585 ( .A1(G61), .A2(n794), .ZN(n536) );
  NAND2_X1 U586 ( .A1(n537), .A2(n536), .ZN(n542) );
  XOR2_X1 U587 ( .A(G543), .B(KEYINPUT0), .Z(n595) );
  NOR2_X1 U588 ( .A1(n595), .A2(n538), .ZN(n797) );
  NAND2_X1 U589 ( .A1(G73), .A2(n797), .ZN(n539) );
  XNOR2_X1 U590 ( .A(n539), .B(KEYINPUT79), .ZN(n540) );
  XNOR2_X1 U591 ( .A(n540), .B(KEYINPUT2), .ZN(n541) );
  NOR2_X1 U592 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U593 ( .A(n543), .B(KEYINPUT80), .ZN(n545) );
  NAND2_X1 U594 ( .A1(G48), .A2(n798), .ZN(n544) );
  NAND2_X1 U595 ( .A1(n545), .A2(n544), .ZN(G305) );
  NAND2_X1 U596 ( .A1(G138), .A2(n892), .ZN(n547) );
  NAND2_X1 U597 ( .A1(G102), .A2(n893), .ZN(n546) );
  NAND2_X1 U598 ( .A1(n547), .A2(n546), .ZN(n551) );
  NAND2_X1 U599 ( .A1(G126), .A2(n888), .ZN(n549) );
  NAND2_X1 U600 ( .A1(G114), .A2(n889), .ZN(n548) );
  NAND2_X1 U601 ( .A1(n549), .A2(n548), .ZN(n550) );
  NOR2_X1 U602 ( .A1(n551), .A2(n550), .ZN(G164) );
  NAND2_X1 U603 ( .A1(G53), .A2(n798), .ZN(n553) );
  NAND2_X1 U604 ( .A1(G65), .A2(n794), .ZN(n552) );
  NAND2_X1 U605 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U606 ( .A(KEYINPUT68), .B(n554), .ZN(n557) );
  NAND2_X1 U607 ( .A1(G91), .A2(n793), .ZN(n555) );
  XNOR2_X1 U608 ( .A(KEYINPUT67), .B(n555), .ZN(n556) );
  NOR2_X1 U609 ( .A1(n557), .A2(n556), .ZN(n559) );
  NAND2_X1 U610 ( .A1(n797), .A2(G78), .ZN(n558) );
  NAND2_X1 U611 ( .A1(n559), .A2(n558), .ZN(G299) );
  NAND2_X1 U612 ( .A1(G52), .A2(n798), .ZN(n561) );
  NAND2_X1 U613 ( .A1(G64), .A2(n794), .ZN(n560) );
  NAND2_X1 U614 ( .A1(n561), .A2(n560), .ZN(n567) );
  NAND2_X1 U615 ( .A1(G77), .A2(n797), .ZN(n563) );
  NAND2_X1 U616 ( .A1(G90), .A2(n793), .ZN(n562) );
  NAND2_X1 U617 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U618 ( .A(KEYINPUT66), .B(n564), .Z(n565) );
  XNOR2_X1 U619 ( .A(KEYINPUT9), .B(n565), .ZN(n566) );
  NOR2_X1 U620 ( .A1(n567), .A2(n566), .ZN(G171) );
  NAND2_X1 U621 ( .A1(n798), .A2(G51), .ZN(n568) );
  XOR2_X1 U622 ( .A(KEYINPUT73), .B(n568), .Z(n570) );
  NAND2_X1 U623 ( .A1(n794), .A2(G63), .ZN(n569) );
  NAND2_X1 U624 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U625 ( .A(KEYINPUT6), .B(n571), .ZN(n579) );
  NAND2_X1 U626 ( .A1(n797), .A2(G76), .ZN(n572) );
  XNOR2_X1 U627 ( .A(KEYINPUT72), .B(n572), .ZN(n576) );
  XOR2_X1 U628 ( .A(KEYINPUT4), .B(KEYINPUT71), .Z(n574) );
  NAND2_X1 U629 ( .A1(G89), .A2(n793), .ZN(n573) );
  XNOR2_X1 U630 ( .A(n574), .B(n573), .ZN(n575) );
  NAND2_X1 U631 ( .A1(n576), .A2(n575), .ZN(n577) );
  XOR2_X1 U632 ( .A(n577), .B(KEYINPUT5), .Z(n578) );
  NOR2_X1 U633 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U634 ( .A(KEYINPUT7), .B(n580), .Z(n582) );
  XOR2_X1 U635 ( .A(KEYINPUT74), .B(KEYINPUT75), .Z(n581) );
  XNOR2_X1 U636 ( .A(n582), .B(n581), .ZN(G168) );
  XOR2_X1 U637 ( .A(KEYINPUT76), .B(KEYINPUT8), .Z(n583) );
  XNOR2_X1 U638 ( .A(G168), .B(n583), .ZN(G286) );
  NAND2_X1 U639 ( .A1(n794), .A2(G62), .ZN(n584) );
  XOR2_X1 U640 ( .A(KEYINPUT81), .B(n584), .Z(n586) );
  NAND2_X1 U641 ( .A1(n798), .A2(G50), .ZN(n585) );
  NAND2_X1 U642 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U643 ( .A(KEYINPUT82), .B(n587), .ZN(n591) );
  NAND2_X1 U644 ( .A1(G75), .A2(n797), .ZN(n589) );
  NAND2_X1 U645 ( .A1(G88), .A2(n793), .ZN(n588) );
  NAND2_X1 U646 ( .A1(n589), .A2(n588), .ZN(n590) );
  NOR2_X1 U647 ( .A1(n591), .A2(n590), .ZN(G166) );
  XOR2_X1 U648 ( .A(KEYINPUT90), .B(G166), .Z(G303) );
  NAND2_X1 U649 ( .A1(G49), .A2(n798), .ZN(n593) );
  NAND2_X1 U650 ( .A1(G74), .A2(G651), .ZN(n592) );
  NAND2_X1 U651 ( .A1(n593), .A2(n592), .ZN(n594) );
  NOR2_X1 U652 ( .A1(n794), .A2(n594), .ZN(n597) );
  NAND2_X1 U653 ( .A1(n595), .A2(G87), .ZN(n596) );
  NAND2_X1 U654 ( .A1(n597), .A2(n596), .ZN(G288) );
  NAND2_X1 U655 ( .A1(G72), .A2(n797), .ZN(n599) );
  NAND2_X1 U656 ( .A1(G85), .A2(n793), .ZN(n598) );
  NAND2_X1 U657 ( .A1(n599), .A2(n598), .ZN(n602) );
  NAND2_X1 U658 ( .A1(G60), .A2(n794), .ZN(n600) );
  XNOR2_X1 U659 ( .A(KEYINPUT65), .B(n600), .ZN(n601) );
  NOR2_X1 U660 ( .A1(n602), .A2(n601), .ZN(n604) );
  NAND2_X1 U661 ( .A1(n798), .A2(G47), .ZN(n603) );
  NAND2_X1 U662 ( .A1(n604), .A2(n603), .ZN(G290) );
  XNOR2_X1 U663 ( .A(G1981), .B(G305), .ZN(n953) );
  NAND2_X1 U664 ( .A1(G66), .A2(n794), .ZN(n611) );
  NAND2_X1 U665 ( .A1(G79), .A2(n797), .ZN(n606) );
  NAND2_X1 U666 ( .A1(G54), .A2(n798), .ZN(n605) );
  NAND2_X1 U667 ( .A1(n606), .A2(n605), .ZN(n609) );
  NAND2_X1 U668 ( .A1(n793), .A2(G92), .ZN(n607) );
  XOR2_X1 U669 ( .A(KEYINPUT70), .B(n607), .Z(n608) );
  NOR2_X1 U670 ( .A1(n609), .A2(n608), .ZN(n610) );
  NAND2_X1 U671 ( .A1(n611), .A2(n610), .ZN(n612) );
  XNOR2_X1 U672 ( .A(n612), .B(KEYINPUT15), .ZN(n938) );
  INV_X1 U673 ( .A(G1348), .ZN(n614) );
  NAND2_X1 U674 ( .A1(G160), .A2(G40), .ZN(n710) );
  NOR2_X1 U675 ( .A1(G164), .A2(G1384), .ZN(n711) );
  INV_X1 U676 ( .A(n711), .ZN(n613) );
  NOR2_X4 U677 ( .A1(n710), .A2(n613), .ZN(n650) );
  OR2_X1 U678 ( .A1(n614), .A2(n650), .ZN(n616) );
  NAND2_X1 U679 ( .A1(G2067), .A2(n650), .ZN(n615) );
  NAND2_X1 U680 ( .A1(n616), .A2(n615), .ZN(n617) );
  XNOR2_X1 U681 ( .A(KEYINPUT99), .B(n617), .ZN(n634) );
  NAND2_X1 U682 ( .A1(G56), .A2(n794), .ZN(n618) );
  XOR2_X1 U683 ( .A(KEYINPUT14), .B(n618), .Z(n624) );
  NAND2_X1 U684 ( .A1(n793), .A2(G81), .ZN(n619) );
  XNOR2_X1 U685 ( .A(n619), .B(KEYINPUT12), .ZN(n621) );
  NAND2_X1 U686 ( .A1(G68), .A2(n797), .ZN(n620) );
  NAND2_X1 U687 ( .A1(n621), .A2(n620), .ZN(n622) );
  XOR2_X1 U688 ( .A(KEYINPUT13), .B(n622), .Z(n623) );
  NOR2_X1 U689 ( .A1(n624), .A2(n623), .ZN(n626) );
  NAND2_X1 U690 ( .A1(n798), .A2(G43), .ZN(n625) );
  NAND2_X1 U691 ( .A1(n626), .A2(n625), .ZN(n943) );
  NAND2_X1 U692 ( .A1(n650), .A2(G1996), .ZN(n628) );
  INV_X1 U693 ( .A(KEYINPUT26), .ZN(n627) );
  XOR2_X1 U694 ( .A(n628), .B(n627), .Z(n630) );
  INV_X1 U695 ( .A(n650), .ZN(n665) );
  NAND2_X1 U696 ( .A1(n665), .A2(G1341), .ZN(n629) );
  NAND2_X1 U697 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U698 ( .A1(n943), .A2(n631), .ZN(n632) );
  NAND2_X1 U699 ( .A1(n633), .A2(n632), .ZN(n636) );
  NAND2_X1 U700 ( .A1(n634), .A2(n938), .ZN(n635) );
  NAND2_X1 U701 ( .A1(n636), .A2(n635), .ZN(n637) );
  XOR2_X1 U702 ( .A(n637), .B(KEYINPUT100), .Z(n644) );
  INV_X1 U703 ( .A(G299), .ZN(n939) );
  NAND2_X1 U704 ( .A1(G1956), .A2(n665), .ZN(n641) );
  NAND2_X1 U705 ( .A1(n650), .A2(G2072), .ZN(n639) );
  NAND2_X1 U706 ( .A1(n641), .A2(n640), .ZN(n642) );
  XOR2_X1 U707 ( .A(KEYINPUT98), .B(n642), .Z(n645) );
  NAND2_X1 U708 ( .A1(n939), .A2(n645), .ZN(n643) );
  NAND2_X1 U709 ( .A1(n644), .A2(n643), .ZN(n648) );
  XOR2_X1 U710 ( .A(n646), .B(KEYINPUT28), .Z(n647) );
  NAND2_X1 U711 ( .A1(n648), .A2(n647), .ZN(n649) );
  XNOR2_X1 U712 ( .A(n649), .B(KEYINPUT29), .ZN(n654) );
  XNOR2_X1 U713 ( .A(G2078), .B(KEYINPUT25), .ZN(n915) );
  NOR2_X1 U714 ( .A1(n665), .A2(n915), .ZN(n652) );
  INV_X1 U715 ( .A(G1961), .ZN(n935) );
  NOR2_X1 U716 ( .A1(n650), .A2(n935), .ZN(n651) );
  NOR2_X1 U717 ( .A1(n652), .A2(n651), .ZN(n659) );
  AND2_X1 U718 ( .A1(G171), .A2(n659), .ZN(n653) );
  NOR2_X2 U719 ( .A1(n654), .A2(n653), .ZN(n655) );
  XNOR2_X1 U720 ( .A(n655), .B(KEYINPUT101), .ZN(n664) );
  NAND2_X1 U721 ( .A1(G8), .A2(n665), .ZN(n705) );
  NOR2_X1 U722 ( .A1(G1966), .A2(n705), .ZN(n677) );
  NOR2_X1 U723 ( .A1(G2084), .A2(n665), .ZN(n673) );
  NOR2_X1 U724 ( .A1(n677), .A2(n673), .ZN(n656) );
  NAND2_X1 U725 ( .A1(G8), .A2(n656), .ZN(n657) );
  XNOR2_X1 U726 ( .A(KEYINPUT30), .B(n657), .ZN(n658) );
  NOR2_X1 U727 ( .A1(G168), .A2(n658), .ZN(n661) );
  NOR2_X1 U728 ( .A1(G171), .A2(n659), .ZN(n660) );
  NOR2_X1 U729 ( .A1(n661), .A2(n660), .ZN(n662) );
  XOR2_X1 U730 ( .A(KEYINPUT31), .B(n662), .Z(n663) );
  NAND2_X1 U731 ( .A1(n664), .A2(n663), .ZN(n675) );
  NAND2_X1 U732 ( .A1(n675), .A2(G286), .ZN(n670) );
  NOR2_X1 U733 ( .A1(G1971), .A2(n705), .ZN(n667) );
  NOR2_X1 U734 ( .A1(G2090), .A2(n665), .ZN(n666) );
  NOR2_X1 U735 ( .A1(n667), .A2(n666), .ZN(n668) );
  NAND2_X1 U736 ( .A1(G303), .A2(n668), .ZN(n669) );
  NAND2_X1 U737 ( .A1(n670), .A2(n669), .ZN(n671) );
  NAND2_X1 U738 ( .A1(n671), .A2(G8), .ZN(n672) );
  XNOR2_X1 U739 ( .A(n672), .B(KEYINPUT32), .ZN(n681) );
  NAND2_X1 U740 ( .A1(G8), .A2(n673), .ZN(n674) );
  XOR2_X1 U741 ( .A(KEYINPUT97), .B(n674), .Z(n679) );
  INV_X1 U742 ( .A(n675), .ZN(n676) );
  NOR2_X1 U743 ( .A1(n677), .A2(n676), .ZN(n678) );
  NAND2_X1 U744 ( .A1(n679), .A2(n678), .ZN(n680) );
  NAND2_X1 U745 ( .A1(n681), .A2(n680), .ZN(n682) );
  NOR2_X1 U746 ( .A1(G1976), .A2(G288), .ZN(n685) );
  NOR2_X1 U747 ( .A1(G303), .A2(G1971), .ZN(n683) );
  NOR2_X1 U748 ( .A1(n685), .A2(n683), .ZN(n959) );
  NAND2_X1 U749 ( .A1(n701), .A2(n959), .ZN(n691) );
  NAND2_X1 U750 ( .A1(G288), .A2(G1976), .ZN(n684) );
  XNOR2_X1 U751 ( .A(n684), .B(KEYINPUT103), .ZN(n937) );
  NOR2_X1 U752 ( .A1(n937), .A2(n705), .ZN(n689) );
  INV_X1 U753 ( .A(KEYINPUT33), .ZN(n693) );
  INV_X1 U754 ( .A(n705), .ZN(n686) );
  NAND2_X1 U755 ( .A1(n686), .A2(n685), .ZN(n687) );
  NOR2_X1 U756 ( .A1(n693), .A2(n687), .ZN(n688) );
  XOR2_X1 U757 ( .A(n688), .B(KEYINPUT104), .Z(n692) );
  AND2_X1 U758 ( .A1(n689), .A2(n692), .ZN(n690) );
  NAND2_X1 U759 ( .A1(n691), .A2(n690), .ZN(n696) );
  INV_X1 U760 ( .A(n692), .ZN(n694) );
  OR2_X1 U761 ( .A1(n694), .A2(n693), .ZN(n695) );
  AND2_X1 U762 ( .A1(n696), .A2(n695), .ZN(n697) );
  NOR2_X1 U763 ( .A1(n953), .A2(n697), .ZN(n698) );
  INV_X1 U764 ( .A(n698), .ZN(n708) );
  NOR2_X1 U765 ( .A1(G303), .A2(G2090), .ZN(n699) );
  NAND2_X1 U766 ( .A1(G8), .A2(n699), .ZN(n700) );
  NAND2_X1 U767 ( .A1(n701), .A2(n700), .ZN(n702) );
  NAND2_X1 U768 ( .A1(n702), .A2(n705), .ZN(n706) );
  NOR2_X1 U769 ( .A1(G1981), .A2(G305), .ZN(n703) );
  XOR2_X1 U770 ( .A(n703), .B(KEYINPUT24), .Z(n704) );
  NAND2_X1 U771 ( .A1(n708), .A2(n707), .ZN(n743) );
  XOR2_X1 U772 ( .A(G1986), .B(KEYINPUT91), .Z(n709) );
  XNOR2_X1 U773 ( .A(G290), .B(n709), .ZN(n949) );
  NOR2_X1 U774 ( .A1(n711), .A2(n710), .ZN(n755) );
  NAND2_X1 U775 ( .A1(n949), .A2(n755), .ZN(n741) );
  XOR2_X1 U776 ( .A(G2067), .B(KEYINPUT37), .Z(n712) );
  XNOR2_X1 U777 ( .A(KEYINPUT92), .B(n712), .ZN(n752) );
  NAND2_X1 U778 ( .A1(n889), .A2(G116), .ZN(n713) );
  XNOR2_X1 U779 ( .A(KEYINPUT94), .B(n713), .ZN(n716) );
  NAND2_X1 U780 ( .A1(n888), .A2(G128), .ZN(n714) );
  XOR2_X1 U781 ( .A(KEYINPUT93), .B(n714), .Z(n715) );
  NAND2_X1 U782 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U783 ( .A(n717), .B(KEYINPUT35), .ZN(n722) );
  NAND2_X1 U784 ( .A1(G140), .A2(n892), .ZN(n719) );
  NAND2_X1 U785 ( .A1(G104), .A2(n893), .ZN(n718) );
  NAND2_X1 U786 ( .A1(n719), .A2(n718), .ZN(n720) );
  XOR2_X1 U787 ( .A(KEYINPUT34), .B(n720), .Z(n721) );
  NAND2_X1 U788 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U789 ( .A(n723), .B(KEYINPUT36), .ZN(n885) );
  NAND2_X1 U790 ( .A1(n752), .A2(n885), .ZN(n724) );
  XNOR2_X1 U791 ( .A(n724), .B(KEYINPUT95), .ZN(n1019) );
  NAND2_X1 U792 ( .A1(n1019), .A2(n755), .ZN(n725) );
  XNOR2_X1 U793 ( .A(n725), .B(KEYINPUT96), .ZN(n750) );
  NAND2_X1 U794 ( .A1(G131), .A2(n892), .ZN(n727) );
  NAND2_X1 U795 ( .A1(G119), .A2(n888), .ZN(n726) );
  NAND2_X1 U796 ( .A1(n727), .A2(n726), .ZN(n731) );
  NAND2_X1 U797 ( .A1(G95), .A2(n893), .ZN(n729) );
  NAND2_X1 U798 ( .A1(G107), .A2(n889), .ZN(n728) );
  NAND2_X1 U799 ( .A1(n729), .A2(n728), .ZN(n730) );
  OR2_X1 U800 ( .A1(n731), .A2(n730), .ZN(n873) );
  AND2_X1 U801 ( .A1(n873), .A2(G1991), .ZN(n994) );
  NAND2_X1 U802 ( .A1(G141), .A2(n892), .ZN(n733) );
  NAND2_X1 U803 ( .A1(G129), .A2(n888), .ZN(n732) );
  NAND2_X1 U804 ( .A1(n733), .A2(n732), .ZN(n736) );
  NAND2_X1 U805 ( .A1(n893), .A2(G105), .ZN(n734) );
  XOR2_X1 U806 ( .A(KEYINPUT38), .B(n734), .Z(n735) );
  NOR2_X1 U807 ( .A1(n736), .A2(n735), .ZN(n738) );
  NAND2_X1 U808 ( .A1(n889), .A2(G117), .ZN(n737) );
  NAND2_X1 U809 ( .A1(n738), .A2(n737), .ZN(n874) );
  AND2_X1 U810 ( .A1(n874), .A2(G1996), .ZN(n996) );
  OR2_X1 U811 ( .A1(n994), .A2(n996), .ZN(n739) );
  NAND2_X1 U812 ( .A1(n755), .A2(n739), .ZN(n744) );
  AND2_X1 U813 ( .A1(n750), .A2(n744), .ZN(n740) );
  AND2_X1 U814 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U815 ( .A1(n743), .A2(n742), .ZN(n758) );
  NOR2_X1 U816 ( .A1(G1996), .A2(n874), .ZN(n1000) );
  INV_X1 U817 ( .A(n744), .ZN(n747) );
  NOR2_X1 U818 ( .A1(G1986), .A2(G290), .ZN(n745) );
  NOR2_X1 U819 ( .A1(G1991), .A2(n873), .ZN(n995) );
  NOR2_X1 U820 ( .A1(n745), .A2(n995), .ZN(n746) );
  NOR2_X1 U821 ( .A1(n747), .A2(n746), .ZN(n748) );
  NOR2_X1 U822 ( .A1(n1000), .A2(n748), .ZN(n749) );
  XNOR2_X1 U823 ( .A(n749), .B(KEYINPUT39), .ZN(n751) );
  NAND2_X1 U824 ( .A1(n751), .A2(n750), .ZN(n754) );
  NOR2_X1 U825 ( .A1(n752), .A2(n885), .ZN(n753) );
  XNOR2_X1 U826 ( .A(n753), .B(KEYINPUT105), .ZN(n1016) );
  NAND2_X1 U827 ( .A1(n754), .A2(n1016), .ZN(n756) );
  NAND2_X1 U828 ( .A1(n756), .A2(n755), .ZN(n757) );
  NAND2_X1 U829 ( .A1(n758), .A2(n757), .ZN(n759) );
  XNOR2_X1 U830 ( .A(n759), .B(KEYINPUT40), .ZN(G329) );
  INV_X1 U831 ( .A(G171), .ZN(G301) );
  XOR2_X1 U832 ( .A(G2438), .B(G2454), .Z(n761) );
  XNOR2_X1 U833 ( .A(G2435), .B(G2430), .ZN(n760) );
  XNOR2_X1 U834 ( .A(n761), .B(n760), .ZN(n762) );
  XOR2_X1 U835 ( .A(n762), .B(G2427), .Z(n764) );
  XNOR2_X1 U836 ( .A(G1341), .B(G1348), .ZN(n763) );
  XNOR2_X1 U837 ( .A(n764), .B(n763), .ZN(n768) );
  XOR2_X1 U838 ( .A(G2443), .B(G2446), .Z(n766) );
  XNOR2_X1 U839 ( .A(KEYINPUT106), .B(G2451), .ZN(n765) );
  XNOR2_X1 U840 ( .A(n766), .B(n765), .ZN(n767) );
  XOR2_X1 U841 ( .A(n768), .B(n767), .Z(n769) );
  AND2_X1 U842 ( .A1(G14), .A2(n769), .ZN(G401) );
  AND2_X1 U843 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U844 ( .A(G57), .ZN(G237) );
  INV_X1 U845 ( .A(G132), .ZN(G219) );
  INV_X1 U846 ( .A(G82), .ZN(G220) );
  NAND2_X1 U847 ( .A1(G7), .A2(G661), .ZN(n770) );
  XOR2_X1 U848 ( .A(n770), .B(KEYINPUT10), .Z(n914) );
  NAND2_X1 U849 ( .A1(n914), .A2(G567), .ZN(n771) );
  XNOR2_X1 U850 ( .A(n771), .B(KEYINPUT11), .ZN(n772) );
  XNOR2_X1 U851 ( .A(KEYINPUT69), .B(n772), .ZN(G234) );
  INV_X1 U852 ( .A(G860), .ZN(n778) );
  OR2_X1 U853 ( .A1(n943), .A2(n778), .ZN(G153) );
  NAND2_X1 U854 ( .A1(G868), .A2(G301), .ZN(n774) );
  OR2_X1 U855 ( .A1(n938), .A2(G868), .ZN(n773) );
  NAND2_X1 U856 ( .A1(n774), .A2(n773), .ZN(G284) );
  INV_X1 U857 ( .A(G868), .ZN(n819) );
  NOR2_X1 U858 ( .A1(G286), .A2(n819), .ZN(n775) );
  XOR2_X1 U859 ( .A(KEYINPUT77), .B(n775), .Z(n777) );
  NOR2_X1 U860 ( .A1(G868), .A2(G299), .ZN(n776) );
  NOR2_X1 U861 ( .A1(n777), .A2(n776), .ZN(G297) );
  NAND2_X1 U862 ( .A1(n778), .A2(G559), .ZN(n779) );
  NAND2_X1 U863 ( .A1(n779), .A2(n938), .ZN(n780) );
  XNOR2_X1 U864 ( .A(n780), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U865 ( .A1(G868), .A2(n943), .ZN(n783) );
  NAND2_X1 U866 ( .A1(G868), .A2(n938), .ZN(n781) );
  NOR2_X1 U867 ( .A1(G559), .A2(n781), .ZN(n782) );
  NOR2_X1 U868 ( .A1(n783), .A2(n782), .ZN(G282) );
  NAND2_X1 U869 ( .A1(G123), .A2(n888), .ZN(n784) );
  XNOR2_X1 U870 ( .A(n784), .B(KEYINPUT18), .ZN(n786) );
  NAND2_X1 U871 ( .A1(n893), .A2(G99), .ZN(n785) );
  NAND2_X1 U872 ( .A1(n786), .A2(n785), .ZN(n790) );
  NAND2_X1 U873 ( .A1(G135), .A2(n892), .ZN(n788) );
  NAND2_X1 U874 ( .A1(G111), .A2(n889), .ZN(n787) );
  NAND2_X1 U875 ( .A1(n788), .A2(n787), .ZN(n789) );
  NOR2_X1 U876 ( .A1(n790), .A2(n789), .ZN(n993) );
  XNOR2_X1 U877 ( .A(G2096), .B(n993), .ZN(n791) );
  INV_X1 U878 ( .A(G2100), .ZN(n849) );
  NAND2_X1 U879 ( .A1(n791), .A2(n849), .ZN(G156) );
  NAND2_X1 U880 ( .A1(n938), .A2(G559), .ZN(n814) );
  XNOR2_X1 U881 ( .A(n943), .B(n814), .ZN(n792) );
  NOR2_X1 U882 ( .A1(n792), .A2(G860), .ZN(n803) );
  NAND2_X1 U883 ( .A1(G93), .A2(n793), .ZN(n796) );
  NAND2_X1 U884 ( .A1(G67), .A2(n794), .ZN(n795) );
  NAND2_X1 U885 ( .A1(n796), .A2(n795), .ZN(n802) );
  NAND2_X1 U886 ( .A1(G80), .A2(n797), .ZN(n800) );
  NAND2_X1 U887 ( .A1(G55), .A2(n798), .ZN(n799) );
  NAND2_X1 U888 ( .A1(n800), .A2(n799), .ZN(n801) );
  OR2_X1 U889 ( .A1(n802), .A2(n801), .ZN(n818) );
  XOR2_X1 U890 ( .A(n803), .B(n818), .Z(G145) );
  XNOR2_X1 U891 ( .A(KEYINPUT84), .B(KEYINPUT83), .ZN(n805) );
  XNOR2_X1 U892 ( .A(G288), .B(KEYINPUT19), .ZN(n804) );
  XNOR2_X1 U893 ( .A(n805), .B(n804), .ZN(n806) );
  XOR2_X1 U894 ( .A(n806), .B(KEYINPUT86), .Z(n808) );
  XOR2_X1 U895 ( .A(G299), .B(KEYINPUT85), .Z(n807) );
  XNOR2_X1 U896 ( .A(n808), .B(n807), .ZN(n811) );
  XOR2_X1 U897 ( .A(n818), .B(G290), .Z(n809) );
  XNOR2_X1 U898 ( .A(n809), .B(n943), .ZN(n810) );
  XNOR2_X1 U899 ( .A(n811), .B(n810), .ZN(n812) );
  XNOR2_X1 U900 ( .A(n812), .B(G305), .ZN(n813) );
  XNOR2_X1 U901 ( .A(G166), .B(n813), .ZN(n840) );
  XNOR2_X1 U902 ( .A(KEYINPUT87), .B(n840), .ZN(n815) );
  XNOR2_X1 U903 ( .A(n815), .B(n814), .ZN(n816) );
  NAND2_X1 U904 ( .A1(n816), .A2(G868), .ZN(n817) );
  XNOR2_X1 U905 ( .A(n817), .B(KEYINPUT88), .ZN(n821) );
  NAND2_X1 U906 ( .A1(n819), .A2(n818), .ZN(n820) );
  NAND2_X1 U907 ( .A1(n821), .A2(n820), .ZN(G295) );
  NAND2_X1 U908 ( .A1(G2084), .A2(G2078), .ZN(n822) );
  XNOR2_X1 U909 ( .A(n822), .B(KEYINPUT20), .ZN(n823) );
  XNOR2_X1 U910 ( .A(KEYINPUT89), .B(n823), .ZN(n824) );
  NAND2_X1 U911 ( .A1(n824), .A2(G2090), .ZN(n825) );
  XNOR2_X1 U912 ( .A(KEYINPUT21), .B(n825), .ZN(n826) );
  NAND2_X1 U913 ( .A1(n826), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U914 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U915 ( .A1(G220), .A2(G219), .ZN(n827) );
  XOR2_X1 U916 ( .A(KEYINPUT22), .B(n827), .Z(n828) );
  NOR2_X1 U917 ( .A1(G218), .A2(n828), .ZN(n829) );
  NAND2_X1 U918 ( .A1(G96), .A2(n829), .ZN(n838) );
  NAND2_X1 U919 ( .A1(n838), .A2(G2106), .ZN(n833) );
  NAND2_X1 U920 ( .A1(G69), .A2(G120), .ZN(n830) );
  NOR2_X1 U921 ( .A1(G237), .A2(n830), .ZN(n831) );
  NAND2_X1 U922 ( .A1(G108), .A2(n831), .ZN(n839) );
  NAND2_X1 U923 ( .A1(n839), .A2(G567), .ZN(n832) );
  NAND2_X1 U924 ( .A1(n833), .A2(n832), .ZN(n913) );
  NAND2_X1 U925 ( .A1(G661), .A2(G483), .ZN(n834) );
  NOR2_X1 U926 ( .A1(n913), .A2(n834), .ZN(n837) );
  NAND2_X1 U927 ( .A1(n837), .A2(G36), .ZN(G176) );
  NAND2_X1 U928 ( .A1(G2106), .A2(n914), .ZN(G217) );
  AND2_X1 U929 ( .A1(G15), .A2(G2), .ZN(n835) );
  NAND2_X1 U930 ( .A1(G661), .A2(n835), .ZN(G259) );
  NAND2_X1 U931 ( .A1(G3), .A2(G1), .ZN(n836) );
  NAND2_X1 U932 ( .A1(n837), .A2(n836), .ZN(G188) );
  INV_X1 U934 ( .A(G120), .ZN(G236) );
  INV_X1 U935 ( .A(G96), .ZN(G221) );
  INV_X1 U936 ( .A(G69), .ZN(G235) );
  NOR2_X1 U937 ( .A1(n839), .A2(n838), .ZN(G325) );
  INV_X1 U938 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U939 ( .A(n938), .B(G286), .ZN(n841) );
  XNOR2_X1 U940 ( .A(n841), .B(n840), .ZN(n842) );
  XOR2_X1 U941 ( .A(n842), .B(G301), .Z(n843) );
  NOR2_X1 U942 ( .A1(G37), .A2(n843), .ZN(G397) );
  XOR2_X1 U943 ( .A(KEYINPUT42), .B(G2084), .Z(n845) );
  XNOR2_X1 U944 ( .A(G2067), .B(G2078), .ZN(n844) );
  XNOR2_X1 U945 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U946 ( .A(n846), .B(G2096), .Z(n848) );
  XNOR2_X1 U947 ( .A(G2090), .B(G2072), .ZN(n847) );
  XNOR2_X1 U948 ( .A(n848), .B(n847), .ZN(n853) );
  XOR2_X1 U949 ( .A(KEYINPUT43), .B(G2678), .Z(n851) );
  XOR2_X1 U950 ( .A(KEYINPUT107), .B(n849), .Z(n850) );
  XNOR2_X1 U951 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U952 ( .A(n853), .B(n852), .Z(G227) );
  XOR2_X1 U953 ( .A(KEYINPUT108), .B(G1956), .Z(n855) );
  XNOR2_X1 U954 ( .A(G1996), .B(G1991), .ZN(n854) );
  XNOR2_X1 U955 ( .A(n855), .B(n854), .ZN(n856) );
  XOR2_X1 U956 ( .A(n856), .B(KEYINPUT41), .Z(n858) );
  XNOR2_X1 U957 ( .A(G1971), .B(G1976), .ZN(n857) );
  XNOR2_X1 U958 ( .A(n858), .B(n857), .ZN(n862) );
  XNOR2_X1 U959 ( .A(G1981), .B(n935), .ZN(n860) );
  XNOR2_X1 U960 ( .A(G1986), .B(G1966), .ZN(n859) );
  XNOR2_X1 U961 ( .A(n860), .B(n859), .ZN(n861) );
  XOR2_X1 U962 ( .A(n862), .B(n861), .Z(n864) );
  XNOR2_X1 U963 ( .A(G2474), .B(KEYINPUT109), .ZN(n863) );
  XNOR2_X1 U964 ( .A(n864), .B(n863), .ZN(G229) );
  NAND2_X1 U965 ( .A1(G124), .A2(n888), .ZN(n865) );
  XNOR2_X1 U966 ( .A(n865), .B(KEYINPUT44), .ZN(n866) );
  XNOR2_X1 U967 ( .A(n866), .B(KEYINPUT110), .ZN(n868) );
  NAND2_X1 U968 ( .A1(G100), .A2(n893), .ZN(n867) );
  NAND2_X1 U969 ( .A1(n868), .A2(n867), .ZN(n872) );
  NAND2_X1 U970 ( .A1(G136), .A2(n892), .ZN(n870) );
  NAND2_X1 U971 ( .A1(G112), .A2(n889), .ZN(n869) );
  NAND2_X1 U972 ( .A1(n870), .A2(n869), .ZN(n871) );
  NOR2_X1 U973 ( .A1(n872), .A2(n871), .ZN(G162) );
  XOR2_X1 U974 ( .A(n993), .B(G162), .Z(n876) );
  XNOR2_X1 U975 ( .A(n874), .B(n873), .ZN(n875) );
  XNOR2_X1 U976 ( .A(n876), .B(n875), .ZN(n884) );
  NAND2_X1 U977 ( .A1(G139), .A2(n892), .ZN(n878) );
  NAND2_X1 U978 ( .A1(G103), .A2(n893), .ZN(n877) );
  NAND2_X1 U979 ( .A1(n878), .A2(n877), .ZN(n883) );
  NAND2_X1 U980 ( .A1(G127), .A2(n888), .ZN(n880) );
  NAND2_X1 U981 ( .A1(G115), .A2(n889), .ZN(n879) );
  NAND2_X1 U982 ( .A1(n880), .A2(n879), .ZN(n881) );
  XOR2_X1 U983 ( .A(KEYINPUT47), .B(n881), .Z(n882) );
  NOR2_X1 U984 ( .A1(n883), .A2(n882), .ZN(n1007) );
  XOR2_X1 U985 ( .A(n884), .B(n1007), .Z(n887) );
  XNOR2_X1 U986 ( .A(G160), .B(n885), .ZN(n886) );
  XNOR2_X1 U987 ( .A(n887), .B(n886), .ZN(n905) );
  XOR2_X1 U988 ( .A(KEYINPUT112), .B(KEYINPUT46), .Z(n902) );
  NAND2_X1 U989 ( .A1(G130), .A2(n888), .ZN(n891) );
  NAND2_X1 U990 ( .A1(G118), .A2(n889), .ZN(n890) );
  NAND2_X1 U991 ( .A1(n891), .A2(n890), .ZN(n899) );
  NAND2_X1 U992 ( .A1(G142), .A2(n892), .ZN(n895) );
  NAND2_X1 U993 ( .A1(G106), .A2(n893), .ZN(n894) );
  NAND2_X1 U994 ( .A1(n895), .A2(n894), .ZN(n896) );
  XNOR2_X1 U995 ( .A(KEYINPUT45), .B(n896), .ZN(n897) );
  XNOR2_X1 U996 ( .A(KEYINPUT111), .B(n897), .ZN(n898) );
  NOR2_X1 U997 ( .A1(n899), .A2(n898), .ZN(n900) );
  XNOR2_X1 U998 ( .A(KEYINPUT48), .B(n900), .ZN(n901) );
  XNOR2_X1 U999 ( .A(n902), .B(n901), .ZN(n903) );
  XNOR2_X1 U1000 ( .A(G164), .B(n903), .ZN(n904) );
  XNOR2_X1 U1001 ( .A(n905), .B(n904), .ZN(n906) );
  NOR2_X1 U1002 ( .A1(G37), .A2(n906), .ZN(G395) );
  NOR2_X1 U1003 ( .A1(G401), .A2(n913), .ZN(n910) );
  NOR2_X1 U1004 ( .A1(G227), .A2(G229), .ZN(n907) );
  XNOR2_X1 U1005 ( .A(KEYINPUT49), .B(n907), .ZN(n908) );
  NOR2_X1 U1006 ( .A1(G397), .A2(n908), .ZN(n909) );
  NAND2_X1 U1007 ( .A1(n910), .A2(n909), .ZN(n911) );
  NOR2_X1 U1008 ( .A1(n911), .A2(G395), .ZN(n912) );
  XNOR2_X1 U1009 ( .A(n912), .B(KEYINPUT113), .ZN(G225) );
  XOR2_X1 U1010 ( .A(KEYINPUT114), .B(G225), .Z(G308) );
  INV_X1 U1011 ( .A(n913), .ZN(G319) );
  INV_X1 U1012 ( .A(G108), .ZN(G238) );
  INV_X1 U1013 ( .A(n914), .ZN(G223) );
  INV_X1 U1014 ( .A(KEYINPUT55), .ZN(n1021) );
  XNOR2_X1 U1015 ( .A(G27), .B(n915), .ZN(n926) );
  XNOR2_X1 U1016 ( .A(G32), .B(G1996), .ZN(n916) );
  XNOR2_X1 U1017 ( .A(n916), .B(KEYINPUT121), .ZN(n921) );
  XOR2_X1 U1018 ( .A(G25), .B(G1991), .Z(n917) );
  NAND2_X1 U1019 ( .A1(n917), .A2(G28), .ZN(n919) );
  XNOR2_X1 U1020 ( .A(G33), .B(G2072), .ZN(n918) );
  NOR2_X1 U1021 ( .A1(n919), .A2(n918), .ZN(n920) );
  NAND2_X1 U1022 ( .A1(n921), .A2(n920), .ZN(n924) );
  XNOR2_X1 U1023 ( .A(KEYINPUT120), .B(G2067), .ZN(n922) );
  XNOR2_X1 U1024 ( .A(G26), .B(n922), .ZN(n923) );
  NOR2_X1 U1025 ( .A1(n924), .A2(n923), .ZN(n925) );
  NAND2_X1 U1026 ( .A1(n926), .A2(n925), .ZN(n927) );
  XNOR2_X1 U1027 ( .A(n927), .B(KEYINPUT53), .ZN(n930) );
  XOR2_X1 U1028 ( .A(G2084), .B(G34), .Z(n928) );
  XNOR2_X1 U1029 ( .A(KEYINPUT54), .B(n928), .ZN(n929) );
  NAND2_X1 U1030 ( .A1(n930), .A2(n929), .ZN(n932) );
  XNOR2_X1 U1031 ( .A(G35), .B(G2090), .ZN(n931) );
  NOR2_X1 U1032 ( .A1(n932), .A2(n931), .ZN(n933) );
  XNOR2_X1 U1033 ( .A(n1021), .B(n933), .ZN(n934) );
  NOR2_X1 U1034 ( .A1(G29), .A2(n934), .ZN(n991) );
  INV_X1 U1035 ( .A(G16), .ZN(n986) );
  XOR2_X1 U1036 ( .A(n986), .B(KEYINPUT56), .Z(n961) );
  XOR2_X1 U1037 ( .A(G301), .B(n935), .Z(n936) );
  NOR2_X1 U1038 ( .A1(n937), .A2(n936), .ZN(n947) );
  XNOR2_X1 U1039 ( .A(n938), .B(G1348), .ZN(n942) );
  XNOR2_X1 U1040 ( .A(G1956), .B(KEYINPUT123), .ZN(n940) );
  XOR2_X1 U1041 ( .A(n940), .B(n939), .Z(n941) );
  NAND2_X1 U1042 ( .A1(n942), .A2(n941), .ZN(n945) );
  XNOR2_X1 U1043 ( .A(G1341), .B(n943), .ZN(n944) );
  NOR2_X1 U1044 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1045 ( .A1(n947), .A2(n946), .ZN(n948) );
  NOR2_X1 U1046 ( .A1(n949), .A2(n948), .ZN(n951) );
  NAND2_X1 U1047 ( .A1(G303), .A2(G1971), .ZN(n950) );
  NAND2_X1 U1048 ( .A1(n951), .A2(n950), .ZN(n957) );
  XOR2_X1 U1049 ( .A(G1966), .B(KEYINPUT122), .Z(n952) );
  XNOR2_X1 U1050 ( .A(G168), .B(n952), .ZN(n954) );
  NOR2_X1 U1051 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1052 ( .A(KEYINPUT57), .B(n955), .ZN(n956) );
  NOR2_X1 U1053 ( .A1(n957), .A2(n956), .ZN(n958) );
  NAND2_X1 U1054 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1055 ( .A1(n961), .A2(n960), .ZN(n988) );
  XNOR2_X1 U1056 ( .A(G1986), .B(KEYINPUT126), .ZN(n962) );
  XNOR2_X1 U1057 ( .A(n962), .B(G24), .ZN(n967) );
  XNOR2_X1 U1058 ( .A(G1971), .B(G22), .ZN(n964) );
  XNOR2_X1 U1059 ( .A(G23), .B(G1976), .ZN(n963) );
  NOR2_X1 U1060 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1061 ( .A(n965), .B(KEYINPUT125), .ZN(n966) );
  NOR2_X1 U1062 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1063 ( .A(KEYINPUT58), .B(n968), .ZN(n981) );
  XOR2_X1 U1064 ( .A(G1348), .B(KEYINPUT59), .Z(n969) );
  XNOR2_X1 U1065 ( .A(G4), .B(n969), .ZN(n971) );
  XNOR2_X1 U1066 ( .A(G20), .B(G1956), .ZN(n970) );
  NOR2_X1 U1067 ( .A1(n971), .A2(n970), .ZN(n975) );
  XNOR2_X1 U1068 ( .A(G1341), .B(G19), .ZN(n973) );
  XNOR2_X1 U1069 ( .A(G6), .B(G1981), .ZN(n972) );
  NOR2_X1 U1070 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1071 ( .A1(n975), .A2(n974), .ZN(n976) );
  XNOR2_X1 U1072 ( .A(n976), .B(KEYINPUT60), .ZN(n979) );
  XNOR2_X1 U1073 ( .A(G1961), .B(G5), .ZN(n977) );
  XNOR2_X1 U1074 ( .A(KEYINPUT124), .B(n977), .ZN(n978) );
  NOR2_X1 U1075 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1076 ( .A1(n981), .A2(n980), .ZN(n983) );
  XNOR2_X1 U1077 ( .A(G21), .B(G1966), .ZN(n982) );
  NOR2_X1 U1078 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1079 ( .A(KEYINPUT61), .B(n984), .ZN(n985) );
  NAND2_X1 U1080 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1081 ( .A1(n988), .A2(n987), .ZN(n989) );
  XOR2_X1 U1082 ( .A(n989), .B(KEYINPUT127), .Z(n990) );
  NOR2_X1 U1083 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1084 ( .A1(G11), .A2(n992), .ZN(n1026) );
  NOR2_X1 U1085 ( .A1(n994), .A2(n993), .ZN(n1006) );
  XNOR2_X1 U1086 ( .A(G160), .B(G2084), .ZN(n998) );
  NOR2_X1 U1087 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1088 ( .A1(n998), .A2(n997), .ZN(n1004) );
  XOR2_X1 U1089 ( .A(G2090), .B(G162), .Z(n999) );
  NOR2_X1 U1090 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XOR2_X1 U1091 ( .A(KEYINPUT51), .B(n1001), .Z(n1002) );
  XNOR2_X1 U1092 ( .A(n1002), .B(KEYINPUT115), .ZN(n1003) );
  NOR2_X1 U1093 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1094 ( .A1(n1006), .A2(n1005), .ZN(n1015) );
  XNOR2_X1 U1095 ( .A(G2072), .B(n1007), .ZN(n1010) );
  XNOR2_X1 U1096 ( .A(G164), .B(G2078), .ZN(n1008) );
  XNOR2_X1 U1097 ( .A(n1008), .B(KEYINPUT116), .ZN(n1009) );
  NAND2_X1 U1098 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1099 ( .A(n1011), .B(KEYINPUT50), .ZN(n1013) );
  XOR2_X1 U1100 ( .A(KEYINPUT117), .B(KEYINPUT118), .Z(n1012) );
  XNOR2_X1 U1101 ( .A(n1013), .B(n1012), .ZN(n1014) );
  NOR2_X1 U1102 ( .A1(n1015), .A2(n1014), .ZN(n1017) );
  NAND2_X1 U1103 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NOR2_X1 U1104 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1105 ( .A(n1020), .B(KEYINPUT52), .ZN(n1022) );
  NAND2_X1 U1106 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1107 ( .A1(G29), .A2(n1023), .ZN(n1024) );
  XNOR2_X1 U1108 ( .A(KEYINPUT119), .B(n1024), .ZN(n1025) );
  NOR2_X1 U1109 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XOR2_X1 U1110 ( .A(KEYINPUT62), .B(n1027), .Z(G150) );
  INV_X1 U1111 ( .A(G150), .ZN(G311) );
endmodule

