

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U561 ( .A(n918), .ZN(n697) );
  XNOR2_X1 U562 ( .A(n540), .B(KEYINPUT87), .ZN(n544) );
  AND2_X1 U563 ( .A1(n543), .A2(n542), .ZN(n526) );
  XNOR2_X1 U564 ( .A(n618), .B(KEYINPUT94), .ZN(n630) );
  OR2_X1 U565 ( .A1(n795), .A2(n643), .ZN(n644) );
  INV_X1 U566 ( .A(KEYINPUT29), .ZN(n656) );
  XNOR2_X1 U567 ( .A(n657), .B(n656), .ZN(n661) );
  NAND2_X1 U568 ( .A1(n698), .A2(n697), .ZN(n699) );
  NOR2_X2 U569 ( .A1(G2104), .A2(n541), .ZN(n884) );
  AND2_X2 U570 ( .A1(n541), .A2(G2104), .ZN(n890) );
  NOR2_X1 U571 ( .A1(G651), .A2(n587), .ZN(n803) );
  AND2_X1 U572 ( .A1(n544), .A2(n526), .ZN(G164) );
  XOR2_X1 U573 ( .A(G543), .B(KEYINPUT0), .Z(n587) );
  INV_X1 U574 ( .A(G651), .ZN(n529) );
  NOR2_X1 U575 ( .A1(n587), .A2(n529), .ZN(n799) );
  NAND2_X1 U576 ( .A1(G72), .A2(n799), .ZN(n528) );
  NOR2_X1 U577 ( .A1(G651), .A2(G543), .ZN(n797) );
  NAND2_X1 U578 ( .A1(G85), .A2(n797), .ZN(n527) );
  NAND2_X1 U579 ( .A1(n528), .A2(n527), .ZN(n533) );
  NOR2_X1 U580 ( .A1(G543), .A2(n529), .ZN(n530) );
  XOR2_X1 U581 ( .A(KEYINPUT1), .B(n530), .Z(n804) );
  NAND2_X1 U582 ( .A1(G60), .A2(n804), .ZN(n531) );
  XOR2_X1 U583 ( .A(KEYINPUT66), .B(n531), .Z(n532) );
  NOR2_X1 U584 ( .A1(n533), .A2(n532), .ZN(n535) );
  NAND2_X1 U585 ( .A1(n803), .A2(G47), .ZN(n534) );
  NAND2_X1 U586 ( .A1(n535), .A2(n534), .ZN(G290) );
  INV_X1 U587 ( .A(G2105), .ZN(n541) );
  NAND2_X1 U588 ( .A1(G102), .A2(n890), .ZN(n539) );
  XNOR2_X1 U589 ( .A(KEYINPUT65), .B(KEYINPUT17), .ZN(n537) );
  NOR2_X1 U590 ( .A1(G2105), .A2(G2104), .ZN(n536) );
  XNOR2_X2 U591 ( .A(n537), .B(n536), .ZN(n888) );
  NAND2_X1 U592 ( .A1(G138), .A2(n888), .ZN(n538) );
  NAND2_X1 U593 ( .A1(n539), .A2(n538), .ZN(n540) );
  NAND2_X1 U594 ( .A1(G126), .A2(n884), .ZN(n543) );
  AND2_X1 U595 ( .A1(G2105), .A2(G2104), .ZN(n885) );
  NAND2_X1 U596 ( .A1(G114), .A2(n885), .ZN(n542) );
  NAND2_X1 U597 ( .A1(G125), .A2(n884), .ZN(n545) );
  XNOR2_X1 U598 ( .A(n545), .B(KEYINPUT64), .ZN(n548) );
  NAND2_X1 U599 ( .A1(G101), .A2(n890), .ZN(n546) );
  XOR2_X1 U600 ( .A(KEYINPUT23), .B(n546), .Z(n547) );
  NAND2_X1 U601 ( .A1(n548), .A2(n547), .ZN(n552) );
  NAND2_X1 U602 ( .A1(G137), .A2(n888), .ZN(n550) );
  NAND2_X1 U603 ( .A1(G113), .A2(n885), .ZN(n549) );
  NAND2_X1 U604 ( .A1(n550), .A2(n549), .ZN(n551) );
  NOR2_X2 U605 ( .A1(n552), .A2(n551), .ZN(G160) );
  NAND2_X1 U606 ( .A1(G91), .A2(n797), .ZN(n554) );
  NAND2_X1 U607 ( .A1(G65), .A2(n804), .ZN(n553) );
  NAND2_X1 U608 ( .A1(n554), .A2(n553), .ZN(n558) );
  NAND2_X1 U609 ( .A1(G78), .A2(n799), .ZN(n556) );
  NAND2_X1 U610 ( .A1(G53), .A2(n803), .ZN(n555) );
  NAND2_X1 U611 ( .A1(n556), .A2(n555), .ZN(n557) );
  NOR2_X1 U612 ( .A1(n558), .A2(n557), .ZN(n559) );
  XOR2_X1 U613 ( .A(KEYINPUT68), .B(n559), .Z(G299) );
  NAND2_X1 U614 ( .A1(G64), .A2(n804), .ZN(n560) );
  XNOR2_X1 U615 ( .A(n560), .B(KEYINPUT67), .ZN(n567) );
  NAND2_X1 U616 ( .A1(G77), .A2(n799), .ZN(n562) );
  NAND2_X1 U617 ( .A1(G90), .A2(n797), .ZN(n561) );
  NAND2_X1 U618 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U619 ( .A(n563), .B(KEYINPUT9), .ZN(n565) );
  NAND2_X1 U620 ( .A1(G52), .A2(n803), .ZN(n564) );
  NAND2_X1 U621 ( .A1(n565), .A2(n564), .ZN(n566) );
  NOR2_X1 U622 ( .A1(n567), .A2(n566), .ZN(G171) );
  NAND2_X1 U623 ( .A1(G89), .A2(n797), .ZN(n568) );
  XNOR2_X1 U624 ( .A(n568), .B(KEYINPUT4), .ZN(n569) );
  XNOR2_X1 U625 ( .A(KEYINPUT72), .B(n569), .ZN(n572) );
  NAND2_X1 U626 ( .A1(n799), .A2(G76), .ZN(n570) );
  XOR2_X1 U627 ( .A(KEYINPUT73), .B(n570), .Z(n571) );
  NAND2_X1 U628 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U629 ( .A(n573), .B(KEYINPUT5), .ZN(n578) );
  NAND2_X1 U630 ( .A1(G51), .A2(n803), .ZN(n575) );
  NAND2_X1 U631 ( .A1(G63), .A2(n804), .ZN(n574) );
  NAND2_X1 U632 ( .A1(n575), .A2(n574), .ZN(n576) );
  XOR2_X1 U633 ( .A(KEYINPUT6), .B(n576), .Z(n577) );
  NAND2_X1 U634 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U635 ( .A(n579), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U636 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U637 ( .A1(G75), .A2(n799), .ZN(n581) );
  NAND2_X1 U638 ( .A1(G88), .A2(n797), .ZN(n580) );
  NAND2_X1 U639 ( .A1(n581), .A2(n580), .ZN(n586) );
  NAND2_X1 U640 ( .A1(G50), .A2(n803), .ZN(n583) );
  NAND2_X1 U641 ( .A1(G62), .A2(n804), .ZN(n582) );
  NAND2_X1 U642 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U643 ( .A(KEYINPUT79), .B(n584), .Z(n585) );
  NOR2_X1 U644 ( .A1(n586), .A2(n585), .ZN(G166) );
  INV_X1 U645 ( .A(G166), .ZN(G303) );
  NAND2_X1 U646 ( .A1(G87), .A2(n587), .ZN(n589) );
  NAND2_X1 U647 ( .A1(G74), .A2(G651), .ZN(n588) );
  NAND2_X1 U648 ( .A1(n589), .A2(n588), .ZN(n590) );
  NOR2_X1 U649 ( .A1(n804), .A2(n590), .ZN(n593) );
  NAND2_X1 U650 ( .A1(G49), .A2(n803), .ZN(n591) );
  XOR2_X1 U651 ( .A(KEYINPUT77), .B(n591), .Z(n592) );
  NAND2_X1 U652 ( .A1(n593), .A2(n592), .ZN(G288) );
  XOR2_X1 U653 ( .A(KEYINPUT2), .B(KEYINPUT78), .Z(n595) );
  NAND2_X1 U654 ( .A1(G73), .A2(n799), .ZN(n594) );
  XNOR2_X1 U655 ( .A(n595), .B(n594), .ZN(n599) );
  NAND2_X1 U656 ( .A1(G86), .A2(n797), .ZN(n597) );
  NAND2_X1 U657 ( .A1(G61), .A2(n804), .ZN(n596) );
  NAND2_X1 U658 ( .A1(n597), .A2(n596), .ZN(n598) );
  NOR2_X1 U659 ( .A1(n599), .A2(n598), .ZN(n601) );
  NAND2_X1 U660 ( .A1(n803), .A2(G48), .ZN(n600) );
  NAND2_X1 U661 ( .A1(n601), .A2(n600), .ZN(G305) );
  XNOR2_X1 U662 ( .A(G1986), .B(KEYINPUT88), .ZN(n602) );
  XNOR2_X1 U663 ( .A(n602), .B(G290), .ZN(n941) );
  NOR2_X1 U664 ( .A1(G164), .A2(G1384), .ZN(n606) );
  NAND2_X1 U665 ( .A1(G40), .A2(G160), .ZN(n603) );
  XOR2_X1 U666 ( .A(KEYINPUT89), .B(n603), .Z(n604) );
  NOR2_X1 U667 ( .A1(n606), .A2(n604), .ZN(n755) );
  NAND2_X1 U668 ( .A1(n941), .A2(n755), .ZN(n743) );
  INV_X1 U669 ( .A(n604), .ZN(n605) );
  NAND2_X2 U670 ( .A1(n606), .A2(n605), .ZN(n673) );
  INV_X1 U671 ( .A(n673), .ZN(n646) );
  INV_X1 U672 ( .A(KEYINPUT26), .ZN(n614) );
  NOR2_X1 U673 ( .A1(n646), .A2(n614), .ZN(n608) );
  XNOR2_X1 U674 ( .A(KEYINPUT93), .B(G1341), .ZN(n607) );
  NAND2_X1 U675 ( .A1(n608), .A2(n607), .ZN(n613) );
  INV_X1 U676 ( .A(G1996), .ZN(n615) );
  NOR2_X1 U677 ( .A1(n615), .A2(n614), .ZN(n609) );
  NOR2_X1 U678 ( .A1(n673), .A2(n609), .ZN(n611) );
  INV_X1 U679 ( .A(KEYINPUT93), .ZN(n610) );
  NAND2_X1 U680 ( .A1(n611), .A2(n610), .ZN(n612) );
  NAND2_X1 U681 ( .A1(n613), .A2(n612), .ZN(n617) );
  NAND2_X1 U682 ( .A1(n615), .A2(n614), .ZN(n616) );
  NAND2_X1 U683 ( .A1(n617), .A2(n616), .ZN(n618) );
  NAND2_X1 U684 ( .A1(n803), .A2(G43), .ZN(n619) );
  XNOR2_X1 U685 ( .A(KEYINPUT70), .B(n619), .ZN(n629) );
  XNOR2_X1 U686 ( .A(KEYINPUT13), .B(KEYINPUT69), .ZN(n624) );
  NAND2_X1 U687 ( .A1(n797), .A2(G81), .ZN(n620) );
  XNOR2_X1 U688 ( .A(n620), .B(KEYINPUT12), .ZN(n622) );
  NAND2_X1 U689 ( .A1(G68), .A2(n799), .ZN(n621) );
  NAND2_X1 U690 ( .A1(n622), .A2(n621), .ZN(n623) );
  XNOR2_X1 U691 ( .A(n624), .B(n623), .ZN(n627) );
  NAND2_X1 U692 ( .A1(n804), .A2(G56), .ZN(n625) );
  XOR2_X1 U693 ( .A(KEYINPUT14), .B(n625), .Z(n626) );
  NOR2_X1 U694 ( .A1(n627), .A2(n626), .ZN(n628) );
  NAND2_X1 U695 ( .A1(n629), .A2(n628), .ZN(n916) );
  NOR2_X1 U696 ( .A1(n630), .A2(n916), .ZN(n643) );
  NAND2_X1 U697 ( .A1(G92), .A2(n797), .ZN(n632) );
  NAND2_X1 U698 ( .A1(G66), .A2(n804), .ZN(n631) );
  NAND2_X1 U699 ( .A1(n632), .A2(n631), .ZN(n636) );
  NAND2_X1 U700 ( .A1(G79), .A2(n799), .ZN(n634) );
  NAND2_X1 U701 ( .A1(G54), .A2(n803), .ZN(n633) );
  NAND2_X1 U702 ( .A1(n634), .A2(n633), .ZN(n635) );
  NOR2_X1 U703 ( .A1(n636), .A2(n635), .ZN(n637) );
  XOR2_X1 U704 ( .A(KEYINPUT15), .B(n637), .Z(n795) );
  NAND2_X1 U705 ( .A1(n643), .A2(n795), .ZN(n642) );
  AND2_X1 U706 ( .A1(n673), .A2(G1348), .ZN(n638) );
  XNOR2_X1 U707 ( .A(n638), .B(KEYINPUT95), .ZN(n640) );
  NAND2_X1 U708 ( .A1(n646), .A2(G2067), .ZN(n639) );
  NAND2_X1 U709 ( .A1(n640), .A2(n639), .ZN(n641) );
  NAND2_X1 U710 ( .A1(n642), .A2(n641), .ZN(n645) );
  NAND2_X1 U711 ( .A1(n645), .A2(n644), .ZN(n651) );
  NAND2_X1 U712 ( .A1(n646), .A2(G2072), .ZN(n647) );
  XNOR2_X1 U713 ( .A(n647), .B(KEYINPUT27), .ZN(n649) );
  AND2_X1 U714 ( .A1(G1956), .A2(n673), .ZN(n648) );
  NOR2_X1 U715 ( .A1(n649), .A2(n648), .ZN(n652) );
  INV_X1 U716 ( .A(G299), .ZN(n937) );
  NAND2_X1 U717 ( .A1(n652), .A2(n937), .ZN(n650) );
  NAND2_X1 U718 ( .A1(n651), .A2(n650), .ZN(n655) );
  NOR2_X1 U719 ( .A1(n652), .A2(n937), .ZN(n653) );
  XOR2_X1 U720 ( .A(n653), .B(KEYINPUT28), .Z(n654) );
  NAND2_X1 U721 ( .A1(n655), .A2(n654), .ZN(n657) );
  XNOR2_X1 U722 ( .A(G2078), .B(KEYINPUT25), .ZN(n955) );
  NOR2_X1 U723 ( .A1(n673), .A2(n955), .ZN(n659) );
  AND2_X1 U724 ( .A1(n673), .A2(G1961), .ZN(n658) );
  NOR2_X1 U725 ( .A1(n659), .A2(n658), .ZN(n666) );
  NAND2_X1 U726 ( .A1(G171), .A2(n666), .ZN(n660) );
  NAND2_X1 U727 ( .A1(n661), .A2(n660), .ZN(n671) );
  NAND2_X1 U728 ( .A1(G8), .A2(n673), .ZN(n710) );
  NOR2_X1 U729 ( .A1(G1966), .A2(n710), .ZN(n684) );
  NOR2_X1 U730 ( .A1(G2084), .A2(n673), .ZN(n681) );
  NOR2_X1 U731 ( .A1(n684), .A2(n681), .ZN(n662) );
  NAND2_X1 U732 ( .A1(G8), .A2(n662), .ZN(n663) );
  XNOR2_X1 U733 ( .A(KEYINPUT30), .B(n663), .ZN(n664) );
  XNOR2_X1 U734 ( .A(KEYINPUT96), .B(n664), .ZN(n665) );
  NOR2_X1 U735 ( .A1(G168), .A2(n665), .ZN(n668) );
  NOR2_X1 U736 ( .A1(G171), .A2(n666), .ZN(n667) );
  NOR2_X1 U737 ( .A1(n668), .A2(n667), .ZN(n669) );
  XOR2_X1 U738 ( .A(KEYINPUT31), .B(n669), .Z(n670) );
  NAND2_X1 U739 ( .A1(n671), .A2(n670), .ZN(n682) );
  NAND2_X1 U740 ( .A1(n682), .A2(G286), .ZN(n678) );
  NOR2_X1 U741 ( .A1(G1971), .A2(n710), .ZN(n672) );
  XNOR2_X1 U742 ( .A(KEYINPUT97), .B(n672), .ZN(n676) );
  NOR2_X1 U743 ( .A1(G2090), .A2(n673), .ZN(n674) );
  NOR2_X1 U744 ( .A1(G166), .A2(n674), .ZN(n675) );
  NAND2_X1 U745 ( .A1(n676), .A2(n675), .ZN(n677) );
  NAND2_X1 U746 ( .A1(n678), .A2(n677), .ZN(n679) );
  NAND2_X1 U747 ( .A1(n679), .A2(G8), .ZN(n680) );
  XNOR2_X1 U748 ( .A(n680), .B(KEYINPUT32), .ZN(n688) );
  NAND2_X1 U749 ( .A1(G8), .A2(n681), .ZN(n686) );
  INV_X1 U750 ( .A(n682), .ZN(n683) );
  NOR2_X1 U751 ( .A1(n684), .A2(n683), .ZN(n685) );
  NAND2_X1 U752 ( .A1(n686), .A2(n685), .ZN(n687) );
  NAND2_X1 U753 ( .A1(n688), .A2(n687), .ZN(n703) );
  NOR2_X1 U754 ( .A1(G1971), .A2(G303), .ZN(n690) );
  NOR2_X1 U755 ( .A1(G1976), .A2(G288), .ZN(n689) );
  XOR2_X1 U756 ( .A(KEYINPUT98), .B(n689), .Z(n695) );
  INV_X1 U757 ( .A(n695), .ZN(n935) );
  NOR2_X1 U758 ( .A1(n690), .A2(n935), .ZN(n691) );
  NAND2_X1 U759 ( .A1(n703), .A2(n691), .ZN(n692) );
  NAND2_X1 U760 ( .A1(G1976), .A2(G288), .ZN(n932) );
  NAND2_X1 U761 ( .A1(n692), .A2(n932), .ZN(n693) );
  NOR2_X1 U762 ( .A1(n693), .A2(n710), .ZN(n694) );
  NOR2_X1 U763 ( .A1(KEYINPUT33), .A2(n694), .ZN(n700) );
  NOR2_X1 U764 ( .A1(n695), .A2(n710), .ZN(n696) );
  NAND2_X1 U765 ( .A1(KEYINPUT33), .A2(n696), .ZN(n698) );
  XNOR2_X1 U766 ( .A(G1981), .B(G305), .ZN(n918) );
  OR2_X1 U767 ( .A1(n700), .A2(n699), .ZN(n706) );
  NOR2_X1 U768 ( .A1(G2090), .A2(G303), .ZN(n701) );
  NAND2_X1 U769 ( .A1(G8), .A2(n701), .ZN(n702) );
  NAND2_X1 U770 ( .A1(n703), .A2(n702), .ZN(n704) );
  NAND2_X1 U771 ( .A1(n704), .A2(n710), .ZN(n705) );
  NAND2_X1 U772 ( .A1(n706), .A2(n705), .ZN(n713) );
  NOR2_X1 U773 ( .A1(G1981), .A2(G305), .ZN(n707) );
  XNOR2_X1 U774 ( .A(KEYINPUT24), .B(n707), .ZN(n708) );
  XNOR2_X1 U775 ( .A(KEYINPUT91), .B(n708), .ZN(n709) );
  NOR2_X1 U776 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U777 ( .A(n711), .B(KEYINPUT92), .ZN(n712) );
  NOR2_X1 U778 ( .A1(n713), .A2(n712), .ZN(n741) );
  XNOR2_X1 U779 ( .A(G2067), .B(KEYINPUT37), .ZN(n753) );
  NAND2_X1 U780 ( .A1(G104), .A2(n890), .ZN(n715) );
  NAND2_X1 U781 ( .A1(G140), .A2(n888), .ZN(n714) );
  NAND2_X1 U782 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U783 ( .A(KEYINPUT34), .B(n716), .ZN(n721) );
  NAND2_X1 U784 ( .A1(G128), .A2(n884), .ZN(n718) );
  NAND2_X1 U785 ( .A1(G116), .A2(n885), .ZN(n717) );
  NAND2_X1 U786 ( .A1(n718), .A2(n717), .ZN(n719) );
  XOR2_X1 U787 ( .A(KEYINPUT35), .B(n719), .Z(n720) );
  NOR2_X1 U788 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U789 ( .A(KEYINPUT36), .B(n722), .ZN(n898) );
  NOR2_X1 U790 ( .A1(n753), .A2(n898), .ZN(n1002) );
  NAND2_X1 U791 ( .A1(n755), .A2(n1002), .ZN(n751) );
  NAND2_X1 U792 ( .A1(G95), .A2(n890), .ZN(n724) );
  NAND2_X1 U793 ( .A1(G131), .A2(n888), .ZN(n723) );
  NAND2_X1 U794 ( .A1(n724), .A2(n723), .ZN(n728) );
  NAND2_X1 U795 ( .A1(G119), .A2(n884), .ZN(n726) );
  NAND2_X1 U796 ( .A1(G107), .A2(n885), .ZN(n725) );
  NAND2_X1 U797 ( .A1(n726), .A2(n725), .ZN(n727) );
  OR2_X1 U798 ( .A1(n728), .A2(n727), .ZN(n881) );
  AND2_X1 U799 ( .A1(n881), .A2(G1991), .ZN(n738) );
  XOR2_X1 U800 ( .A(KEYINPUT38), .B(KEYINPUT90), .Z(n730) );
  NAND2_X1 U801 ( .A1(G105), .A2(n890), .ZN(n729) );
  XNOR2_X1 U802 ( .A(n730), .B(n729), .ZN(n734) );
  NAND2_X1 U803 ( .A1(G141), .A2(n888), .ZN(n732) );
  NAND2_X1 U804 ( .A1(G129), .A2(n884), .ZN(n731) );
  NAND2_X1 U805 ( .A1(n732), .A2(n731), .ZN(n733) );
  NOR2_X1 U806 ( .A1(n734), .A2(n733), .ZN(n736) );
  NAND2_X1 U807 ( .A1(n885), .A2(G117), .ZN(n735) );
  NAND2_X1 U808 ( .A1(n736), .A2(n735), .ZN(n876) );
  AND2_X1 U809 ( .A1(n876), .A2(G1996), .ZN(n737) );
  NOR2_X1 U810 ( .A1(n738), .A2(n737), .ZN(n1000) );
  INV_X1 U811 ( .A(n1000), .ZN(n739) );
  NAND2_X1 U812 ( .A1(n739), .A2(n755), .ZN(n744) );
  NAND2_X1 U813 ( .A1(n751), .A2(n744), .ZN(n740) );
  NOR2_X1 U814 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U815 ( .A1(n743), .A2(n742), .ZN(n758) );
  NOR2_X1 U816 ( .A1(G1996), .A2(n876), .ZN(n997) );
  INV_X1 U817 ( .A(n744), .ZN(n748) );
  NOR2_X1 U818 ( .A1(G1991), .A2(n881), .ZN(n1001) );
  NOR2_X1 U819 ( .A1(G1986), .A2(G290), .ZN(n745) );
  NOR2_X1 U820 ( .A1(n1001), .A2(n745), .ZN(n746) );
  XOR2_X1 U821 ( .A(KEYINPUT99), .B(n746), .Z(n747) );
  NOR2_X1 U822 ( .A1(n748), .A2(n747), .ZN(n749) );
  NOR2_X1 U823 ( .A1(n997), .A2(n749), .ZN(n750) );
  XNOR2_X1 U824 ( .A(n750), .B(KEYINPUT39), .ZN(n752) );
  NAND2_X1 U825 ( .A1(n752), .A2(n751), .ZN(n754) );
  NAND2_X1 U826 ( .A1(n753), .A2(n898), .ZN(n1011) );
  NAND2_X1 U827 ( .A1(n754), .A2(n1011), .ZN(n756) );
  NAND2_X1 U828 ( .A1(n756), .A2(n755), .ZN(n757) );
  NAND2_X1 U829 ( .A1(n758), .A2(n757), .ZN(n760) );
  XNOR2_X1 U830 ( .A(KEYINPUT40), .B(KEYINPUT100), .ZN(n759) );
  XNOR2_X1 U831 ( .A(n760), .B(n759), .ZN(G329) );
  XOR2_X1 U832 ( .A(G2435), .B(G2454), .Z(n762) );
  XNOR2_X1 U833 ( .A(KEYINPUT101), .B(G2438), .ZN(n761) );
  XNOR2_X1 U834 ( .A(n762), .B(n761), .ZN(n769) );
  XOR2_X1 U835 ( .A(G2446), .B(G2430), .Z(n764) );
  XNOR2_X1 U836 ( .A(G2451), .B(G2443), .ZN(n763) );
  XNOR2_X1 U837 ( .A(n764), .B(n763), .ZN(n765) );
  XOR2_X1 U838 ( .A(n765), .B(G2427), .Z(n767) );
  XNOR2_X1 U839 ( .A(G1348), .B(G1341), .ZN(n766) );
  XNOR2_X1 U840 ( .A(n767), .B(n766), .ZN(n768) );
  XNOR2_X1 U841 ( .A(n769), .B(n768), .ZN(n770) );
  AND2_X1 U842 ( .A1(n770), .A2(G14), .ZN(G401) );
  AND2_X1 U843 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U844 ( .A(G57), .ZN(G237) );
  INV_X1 U845 ( .A(G132), .ZN(G219) );
  INV_X1 U846 ( .A(G82), .ZN(G220) );
  NAND2_X1 U847 ( .A1(G7), .A2(G661), .ZN(n771) );
  XNOR2_X1 U848 ( .A(n771), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U849 ( .A(G223), .ZN(n836) );
  NAND2_X1 U850 ( .A1(n836), .A2(G567), .ZN(n772) );
  XOR2_X1 U851 ( .A(KEYINPUT11), .B(n772), .Z(G234) );
  INV_X1 U852 ( .A(G860), .ZN(n779) );
  OR2_X1 U853 ( .A1(n916), .A2(n779), .ZN(n773) );
  XOR2_X1 U854 ( .A(KEYINPUT71), .B(n773), .Z(G153) );
  INV_X1 U855 ( .A(G171), .ZN(G301) );
  NAND2_X1 U856 ( .A1(G868), .A2(G301), .ZN(n775) );
  INV_X1 U857 ( .A(n795), .ZN(n924) );
  INV_X1 U858 ( .A(G868), .ZN(n776) );
  NAND2_X1 U859 ( .A1(n924), .A2(n776), .ZN(n774) );
  NAND2_X1 U860 ( .A1(n775), .A2(n774), .ZN(G284) );
  NOR2_X1 U861 ( .A1(G286), .A2(n776), .ZN(n778) );
  NOR2_X1 U862 ( .A1(G299), .A2(G868), .ZN(n777) );
  NOR2_X1 U863 ( .A1(n778), .A2(n777), .ZN(G297) );
  NAND2_X1 U864 ( .A1(n779), .A2(G559), .ZN(n780) );
  NAND2_X1 U865 ( .A1(n780), .A2(n795), .ZN(n781) );
  XNOR2_X1 U866 ( .A(n781), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U867 ( .A1(G868), .A2(n916), .ZN(n784) );
  NAND2_X1 U868 ( .A1(G868), .A2(n795), .ZN(n782) );
  NOR2_X1 U869 ( .A1(G559), .A2(n782), .ZN(n783) );
  NOR2_X1 U870 ( .A1(n784), .A2(n783), .ZN(G282) );
  NAND2_X1 U871 ( .A1(G123), .A2(n884), .ZN(n785) );
  XNOR2_X1 U872 ( .A(n785), .B(KEYINPUT18), .ZN(n788) );
  NAND2_X1 U873 ( .A1(G99), .A2(n890), .ZN(n786) );
  XNOR2_X1 U874 ( .A(n786), .B(KEYINPUT74), .ZN(n787) );
  NAND2_X1 U875 ( .A1(n788), .A2(n787), .ZN(n792) );
  NAND2_X1 U876 ( .A1(G135), .A2(n888), .ZN(n790) );
  NAND2_X1 U877 ( .A1(G111), .A2(n885), .ZN(n789) );
  NAND2_X1 U878 ( .A1(n790), .A2(n789), .ZN(n791) );
  NOR2_X1 U879 ( .A1(n792), .A2(n791), .ZN(n1005) );
  XNOR2_X1 U880 ( .A(n1005), .B(G2096), .ZN(n794) );
  INV_X1 U881 ( .A(G2100), .ZN(n793) );
  NAND2_X1 U882 ( .A1(n794), .A2(n793), .ZN(G156) );
  NAND2_X1 U883 ( .A1(G559), .A2(n795), .ZN(n796) );
  XNOR2_X1 U884 ( .A(n916), .B(n796), .ZN(n817) );
  NOR2_X1 U885 ( .A1(n817), .A2(G860), .ZN(n809) );
  NAND2_X1 U886 ( .A1(n797), .A2(G93), .ZN(n798) );
  XOR2_X1 U887 ( .A(KEYINPUT75), .B(n798), .Z(n801) );
  NAND2_X1 U888 ( .A1(n799), .A2(G80), .ZN(n800) );
  NAND2_X1 U889 ( .A1(n801), .A2(n800), .ZN(n802) );
  XNOR2_X1 U890 ( .A(KEYINPUT76), .B(n802), .ZN(n808) );
  NAND2_X1 U891 ( .A1(G55), .A2(n803), .ZN(n806) );
  NAND2_X1 U892 ( .A1(G67), .A2(n804), .ZN(n805) );
  NAND2_X1 U893 ( .A1(n806), .A2(n805), .ZN(n807) );
  NOR2_X1 U894 ( .A1(n808), .A2(n807), .ZN(n901) );
  XNOR2_X1 U895 ( .A(n809), .B(n901), .ZN(G145) );
  XOR2_X1 U896 ( .A(KEYINPUT80), .B(KEYINPUT82), .Z(n811) );
  XNOR2_X1 U897 ( .A(KEYINPUT19), .B(KEYINPUT81), .ZN(n810) );
  XNOR2_X1 U898 ( .A(n811), .B(n810), .ZN(n814) );
  XNOR2_X1 U899 ( .A(G299), .B(G290), .ZN(n812) );
  XNOR2_X1 U900 ( .A(n812), .B(G305), .ZN(n813) );
  XNOR2_X1 U901 ( .A(n814), .B(n813), .ZN(n816) );
  XNOR2_X1 U902 ( .A(G288), .B(G166), .ZN(n815) );
  XNOR2_X1 U903 ( .A(n816), .B(n815), .ZN(n902) );
  XOR2_X1 U904 ( .A(n902), .B(n817), .Z(n818) );
  NAND2_X1 U905 ( .A1(n818), .A2(G868), .ZN(n819) );
  XNOR2_X1 U906 ( .A(n819), .B(KEYINPUT83), .ZN(n820) );
  XNOR2_X1 U907 ( .A(n901), .B(n820), .ZN(G295) );
  NAND2_X1 U908 ( .A1(G2078), .A2(G2084), .ZN(n821) );
  XOR2_X1 U909 ( .A(KEYINPUT20), .B(n821), .Z(n822) );
  NAND2_X1 U910 ( .A1(G2090), .A2(n822), .ZN(n824) );
  XNOR2_X1 U911 ( .A(KEYINPUT21), .B(KEYINPUT84), .ZN(n823) );
  XNOR2_X1 U912 ( .A(n824), .B(n823), .ZN(n825) );
  NAND2_X1 U913 ( .A1(n825), .A2(G2072), .ZN(n826) );
  XOR2_X1 U914 ( .A(KEYINPUT85), .B(n826), .Z(G158) );
  XNOR2_X1 U915 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U916 ( .A1(G220), .A2(G219), .ZN(n827) );
  XOR2_X1 U917 ( .A(KEYINPUT22), .B(n827), .Z(n828) );
  NOR2_X1 U918 ( .A1(G218), .A2(n828), .ZN(n829) );
  NAND2_X1 U919 ( .A1(G96), .A2(n829), .ZN(n841) );
  NAND2_X1 U920 ( .A1(n841), .A2(G2106), .ZN(n834) );
  NAND2_X1 U921 ( .A1(G120), .A2(G69), .ZN(n830) );
  NOR2_X1 U922 ( .A1(G237), .A2(n830), .ZN(n831) );
  NAND2_X1 U923 ( .A1(n831), .A2(G108), .ZN(n832) );
  XNOR2_X1 U924 ( .A(n832), .B(KEYINPUT86), .ZN(n842) );
  NAND2_X1 U925 ( .A1(n842), .A2(G567), .ZN(n833) );
  NAND2_X1 U926 ( .A1(n834), .A2(n833), .ZN(n915) );
  NAND2_X1 U927 ( .A1(G661), .A2(G483), .ZN(n835) );
  NOR2_X1 U928 ( .A1(n915), .A2(n835), .ZN(n839) );
  NAND2_X1 U929 ( .A1(n839), .A2(G36), .ZN(G176) );
  NAND2_X1 U930 ( .A1(G2106), .A2(n836), .ZN(G217) );
  AND2_X1 U931 ( .A1(G15), .A2(G2), .ZN(n837) );
  NAND2_X1 U932 ( .A1(G661), .A2(n837), .ZN(G259) );
  NAND2_X1 U933 ( .A1(G3), .A2(G1), .ZN(n838) );
  XNOR2_X1 U934 ( .A(KEYINPUT102), .B(n838), .ZN(n840) );
  NAND2_X1 U935 ( .A1(n840), .A2(n839), .ZN(G188) );
  XNOR2_X1 U936 ( .A(G69), .B(KEYINPUT103), .ZN(G235) );
  INV_X1 U938 ( .A(G120), .ZN(G236) );
  INV_X1 U939 ( .A(G96), .ZN(G221) );
  NOR2_X1 U940 ( .A1(n842), .A2(n841), .ZN(G325) );
  INV_X1 U941 ( .A(G325), .ZN(G261) );
  XOR2_X1 U942 ( .A(G1956), .B(G1961), .Z(n844) );
  XNOR2_X1 U943 ( .A(G1986), .B(G1971), .ZN(n843) );
  XNOR2_X1 U944 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U945 ( .A(n845), .B(G2474), .Z(n847) );
  XNOR2_X1 U946 ( .A(G1981), .B(G1966), .ZN(n846) );
  XNOR2_X1 U947 ( .A(n847), .B(n846), .ZN(n851) );
  XOR2_X1 U948 ( .A(KEYINPUT41), .B(G1976), .Z(n849) );
  XNOR2_X1 U949 ( .A(G1996), .B(G1991), .ZN(n848) );
  XNOR2_X1 U950 ( .A(n849), .B(n848), .ZN(n850) );
  XNOR2_X1 U951 ( .A(n851), .B(n850), .ZN(G229) );
  XOR2_X1 U952 ( .A(G2100), .B(G2096), .Z(n853) );
  XNOR2_X1 U953 ( .A(KEYINPUT42), .B(G2678), .ZN(n852) );
  XNOR2_X1 U954 ( .A(n853), .B(n852), .ZN(n857) );
  XOR2_X1 U955 ( .A(KEYINPUT43), .B(G2090), .Z(n855) );
  XNOR2_X1 U956 ( .A(G2067), .B(G2072), .ZN(n854) );
  XNOR2_X1 U957 ( .A(n855), .B(n854), .ZN(n856) );
  XOR2_X1 U958 ( .A(n857), .B(n856), .Z(n859) );
  XNOR2_X1 U959 ( .A(G2078), .B(G2084), .ZN(n858) );
  XNOR2_X1 U960 ( .A(n859), .B(n858), .ZN(G227) );
  NAND2_X1 U961 ( .A1(G124), .A2(n884), .ZN(n860) );
  XNOR2_X1 U962 ( .A(n860), .B(KEYINPUT44), .ZN(n862) );
  NAND2_X1 U963 ( .A1(n890), .A2(G100), .ZN(n861) );
  NAND2_X1 U964 ( .A1(n862), .A2(n861), .ZN(n866) );
  NAND2_X1 U965 ( .A1(G136), .A2(n888), .ZN(n864) );
  NAND2_X1 U966 ( .A1(G112), .A2(n885), .ZN(n863) );
  NAND2_X1 U967 ( .A1(n864), .A2(n863), .ZN(n865) );
  NOR2_X1 U968 ( .A1(n866), .A2(n865), .ZN(G162) );
  XOR2_X1 U969 ( .A(KEYINPUT48), .B(KEYINPUT105), .Z(n875) );
  NAND2_X1 U970 ( .A1(G103), .A2(n890), .ZN(n868) );
  NAND2_X1 U971 ( .A1(G139), .A2(n888), .ZN(n867) );
  NAND2_X1 U972 ( .A1(n868), .A2(n867), .ZN(n873) );
  NAND2_X1 U973 ( .A1(G127), .A2(n884), .ZN(n870) );
  NAND2_X1 U974 ( .A1(G115), .A2(n885), .ZN(n869) );
  NAND2_X1 U975 ( .A1(n870), .A2(n869), .ZN(n871) );
  XOR2_X1 U976 ( .A(KEYINPUT47), .B(n871), .Z(n872) );
  NOR2_X1 U977 ( .A1(n873), .A2(n872), .ZN(n1013) );
  XNOR2_X1 U978 ( .A(n1013), .B(KEYINPUT46), .ZN(n874) );
  XNOR2_X1 U979 ( .A(n875), .B(n874), .ZN(n880) );
  XOR2_X1 U980 ( .A(G162), .B(n1005), .Z(n878) );
  XOR2_X1 U981 ( .A(G160), .B(n876), .Z(n877) );
  XNOR2_X1 U982 ( .A(n878), .B(n877), .ZN(n879) );
  XOR2_X1 U983 ( .A(n880), .B(n879), .Z(n883) );
  XOR2_X1 U984 ( .A(G164), .B(n881), .Z(n882) );
  XNOR2_X1 U985 ( .A(n883), .B(n882), .ZN(n897) );
  NAND2_X1 U986 ( .A1(G130), .A2(n884), .ZN(n887) );
  NAND2_X1 U987 ( .A1(G118), .A2(n885), .ZN(n886) );
  NAND2_X1 U988 ( .A1(n887), .A2(n886), .ZN(n895) );
  NAND2_X1 U989 ( .A1(n888), .A2(G142), .ZN(n889) );
  XNOR2_X1 U990 ( .A(n889), .B(KEYINPUT104), .ZN(n892) );
  NAND2_X1 U991 ( .A1(G106), .A2(n890), .ZN(n891) );
  NAND2_X1 U992 ( .A1(n892), .A2(n891), .ZN(n893) );
  XOR2_X1 U993 ( .A(n893), .B(KEYINPUT45), .Z(n894) );
  NOR2_X1 U994 ( .A1(n895), .A2(n894), .ZN(n896) );
  XOR2_X1 U995 ( .A(n897), .B(n896), .Z(n899) );
  XOR2_X1 U996 ( .A(n899), .B(n898), .Z(n900) );
  NOR2_X1 U997 ( .A1(G37), .A2(n900), .ZN(G395) );
  XNOR2_X1 U998 ( .A(n902), .B(n901), .ZN(n904) );
  XNOR2_X1 U999 ( .A(n916), .B(G286), .ZN(n903) );
  XNOR2_X1 U1000 ( .A(n904), .B(n903), .ZN(n906) );
  XOR2_X1 U1001 ( .A(n924), .B(G171), .Z(n905) );
  XNOR2_X1 U1002 ( .A(n906), .B(n905), .ZN(n907) );
  NOR2_X1 U1003 ( .A1(G37), .A2(n907), .ZN(G397) );
  NOR2_X1 U1004 ( .A1(G229), .A2(G227), .ZN(n908) );
  XNOR2_X1 U1005 ( .A(n908), .B(KEYINPUT49), .ZN(n911) );
  NOR2_X1 U1006 ( .A1(G395), .A2(G397), .ZN(n909) );
  XNOR2_X1 U1007 ( .A(n909), .B(KEYINPUT107), .ZN(n910) );
  NOR2_X1 U1008 ( .A1(n911), .A2(n910), .ZN(n914) );
  NOR2_X1 U1009 ( .A1(G401), .A2(n915), .ZN(n912) );
  XNOR2_X1 U1010 ( .A(n912), .B(KEYINPUT106), .ZN(n913) );
  NAND2_X1 U1011 ( .A1(n914), .A2(n913), .ZN(G225) );
  INV_X1 U1012 ( .A(G225), .ZN(G308) );
  INV_X1 U1013 ( .A(n915), .ZN(G319) );
  INV_X1 U1014 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1015 ( .A(n916), .B(G1341), .ZN(n922) );
  XOR2_X1 U1016 ( .A(G1966), .B(G168), .Z(n917) );
  NOR2_X1 U1017 ( .A1(n918), .A2(n917), .ZN(n919) );
  XOR2_X1 U1018 ( .A(KEYINPUT115), .B(n919), .Z(n920) );
  XNOR2_X1 U1019 ( .A(KEYINPUT57), .B(n920), .ZN(n921) );
  NOR2_X1 U1020 ( .A1(n922), .A2(n921), .ZN(n930) );
  XNOR2_X1 U1021 ( .A(G171), .B(G1961), .ZN(n923) );
  XNOR2_X1 U1022 ( .A(n923), .B(KEYINPUT117), .ZN(n927) );
  XNOR2_X1 U1023 ( .A(G1348), .B(KEYINPUT116), .ZN(n925) );
  XNOR2_X1 U1024 ( .A(n925), .B(n924), .ZN(n926) );
  NOR2_X1 U1025 ( .A1(n927), .A2(n926), .ZN(n928) );
  XNOR2_X1 U1026 ( .A(n928), .B(KEYINPUT118), .ZN(n929) );
  NAND2_X1 U1027 ( .A1(n930), .A2(n929), .ZN(n944) );
  XNOR2_X1 U1028 ( .A(G1971), .B(G303), .ZN(n931) );
  XNOR2_X1 U1029 ( .A(n931), .B(KEYINPUT119), .ZN(n933) );
  NAND2_X1 U1030 ( .A1(n933), .A2(n932), .ZN(n934) );
  NOR2_X1 U1031 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1032 ( .A(KEYINPUT120), .B(n936), .ZN(n939) );
  XNOR2_X1 U1033 ( .A(n937), .B(G1956), .ZN(n938) );
  NAND2_X1 U1034 ( .A1(n939), .A2(n938), .ZN(n940) );
  NOR2_X1 U1035 ( .A1(n941), .A2(n940), .ZN(n942) );
  XNOR2_X1 U1036 ( .A(KEYINPUT121), .B(n942), .ZN(n943) );
  NOR2_X1 U1037 ( .A1(n944), .A2(n943), .ZN(n945) );
  XOR2_X1 U1038 ( .A(KEYINPUT122), .B(n945), .Z(n947) );
  XNOR2_X1 U1039 ( .A(G16), .B(KEYINPUT56), .ZN(n946) );
  NAND2_X1 U1040 ( .A1(n947), .A2(n946), .ZN(n1030) );
  XNOR2_X1 U1041 ( .A(G1996), .B(G32), .ZN(n949) );
  XNOR2_X1 U1042 ( .A(G33), .B(G2072), .ZN(n948) );
  NOR2_X1 U1043 ( .A1(n949), .A2(n948), .ZN(n954) );
  XOR2_X1 U1044 ( .A(G25), .B(G1991), .Z(n950) );
  NAND2_X1 U1045 ( .A1(n950), .A2(G28), .ZN(n952) );
  XNOR2_X1 U1046 ( .A(G26), .B(G2067), .ZN(n951) );
  NOR2_X1 U1047 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1048 ( .A1(n954), .A2(n953), .ZN(n957) );
  XOR2_X1 U1049 ( .A(G27), .B(n955), .Z(n956) );
  NOR2_X1 U1050 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1051 ( .A(KEYINPUT113), .B(n958), .ZN(n959) );
  XNOR2_X1 U1052 ( .A(n959), .B(KEYINPUT53), .ZN(n963) );
  XOR2_X1 U1053 ( .A(KEYINPUT114), .B(G34), .Z(n961) );
  XNOR2_X1 U1054 ( .A(G2084), .B(KEYINPUT54), .ZN(n960) );
  XNOR2_X1 U1055 ( .A(n961), .B(n960), .ZN(n962) );
  NAND2_X1 U1056 ( .A1(n963), .A2(n962), .ZN(n965) );
  XNOR2_X1 U1057 ( .A(G35), .B(G2090), .ZN(n964) );
  NOR2_X1 U1058 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1059 ( .A(KEYINPUT55), .B(n966), .ZN(n968) );
  INV_X1 U1060 ( .A(G29), .ZN(n967) );
  NAND2_X1 U1061 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1062 ( .A1(n969), .A2(G11), .ZN(n1028) );
  XOR2_X1 U1063 ( .A(G5), .B(G1961), .Z(n990) );
  XOR2_X1 U1064 ( .A(G1986), .B(KEYINPUT126), .Z(n970) );
  XNOR2_X1 U1065 ( .A(G24), .B(n970), .ZN(n974) );
  XNOR2_X1 U1066 ( .A(G1976), .B(G23), .ZN(n972) );
  XNOR2_X1 U1067 ( .A(G1971), .B(G22), .ZN(n971) );
  NOR2_X1 U1068 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1069 ( .A1(n974), .A2(n973), .ZN(n975) );
  XNOR2_X1 U1070 ( .A(n975), .B(KEYINPUT58), .ZN(n988) );
  XNOR2_X1 U1071 ( .A(G1956), .B(G20), .ZN(n982) );
  XNOR2_X1 U1072 ( .A(G1981), .B(G6), .ZN(n976) );
  XNOR2_X1 U1073 ( .A(n976), .B(KEYINPUT124), .ZN(n979) );
  XOR2_X1 U1074 ( .A(G1341), .B(KEYINPUT123), .Z(n977) );
  XNOR2_X1 U1075 ( .A(G19), .B(n977), .ZN(n978) );
  NOR2_X1 U1076 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1077 ( .A(KEYINPUT125), .B(n980), .ZN(n981) );
  NOR2_X1 U1078 ( .A1(n982), .A2(n981), .ZN(n985) );
  XNOR2_X1 U1079 ( .A(G1348), .B(KEYINPUT59), .ZN(n983) );
  XNOR2_X1 U1080 ( .A(n983), .B(G4), .ZN(n984) );
  NAND2_X1 U1081 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1082 ( .A(KEYINPUT60), .B(n986), .ZN(n987) );
  NOR2_X1 U1083 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1084 ( .A1(n990), .A2(n989), .ZN(n992) );
  XNOR2_X1 U1085 ( .A(G21), .B(G1966), .ZN(n991) );
  NOR2_X1 U1086 ( .A1(n992), .A2(n991), .ZN(n993) );
  XOR2_X1 U1087 ( .A(KEYINPUT61), .B(n993), .Z(n994) );
  NOR2_X1 U1088 ( .A1(G16), .A2(n994), .ZN(n995) );
  XNOR2_X1 U1089 ( .A(KEYINPUT127), .B(n995), .ZN(n1026) );
  XOR2_X1 U1090 ( .A(G2090), .B(G162), .Z(n996) );
  NOR2_X1 U1091 ( .A1(n997), .A2(n996), .ZN(n998) );
  XOR2_X1 U1092 ( .A(KEYINPUT51), .B(n998), .Z(n999) );
  NAND2_X1 U1093 ( .A1(n1000), .A2(n999), .ZN(n1010) );
  NOR2_X1 U1094 ( .A1(n1002), .A2(n1001), .ZN(n1007) );
  XOR2_X1 U1095 ( .A(G2084), .B(G160), .Z(n1003) );
  XNOR2_X1 U1096 ( .A(KEYINPUT108), .B(n1003), .ZN(n1004) );
  NOR2_X1 U1097 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1098 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XOR2_X1 U1099 ( .A(KEYINPUT109), .B(n1008), .Z(n1009) );
  NOR2_X1 U1100 ( .A1(n1010), .A2(n1009), .ZN(n1012) );
  NAND2_X1 U1101 ( .A1(n1012), .A2(n1011), .ZN(n1020) );
  XNOR2_X1 U1102 ( .A(G164), .B(G2078), .ZN(n1016) );
  XNOR2_X1 U1103 ( .A(G2072), .B(n1013), .ZN(n1014) );
  XNOR2_X1 U1104 ( .A(n1014), .B(KEYINPUT110), .ZN(n1015) );
  NAND2_X1 U1105 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1106 ( .A(n1017), .B(KEYINPUT111), .ZN(n1018) );
  XOR2_X1 U1107 ( .A(KEYINPUT50), .B(n1018), .Z(n1019) );
  NOR2_X1 U1108 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XOR2_X1 U1109 ( .A(KEYINPUT52), .B(n1021), .Z(n1022) );
  NOR2_X1 U1110 ( .A1(KEYINPUT55), .A2(n1022), .ZN(n1023) );
  XOR2_X1 U1111 ( .A(KEYINPUT112), .B(n1023), .Z(n1024) );
  NAND2_X1 U1112 ( .A1(n1024), .A2(G29), .ZN(n1025) );
  NAND2_X1 U1113 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NOR2_X1 U1114 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NAND2_X1 U1115 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XOR2_X1 U1116 ( .A(KEYINPUT62), .B(n1031), .Z(G311) );
  INV_X1 U1117 ( .A(G311), .ZN(G150) );
endmodule

