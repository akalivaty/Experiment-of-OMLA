//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 0 0 1 0 1 1 0 0 0 1 0 1 0 1 1 0 1 0 0 0 0 1 1 1 0 1 1 0 1 1 0 1 0 0 1 0 0 1 1 1 1 0 0 0 1 0 0 1 0 1 0 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n778, new_n779, new_n780, new_n781, new_n783, new_n784, new_n785,
    new_n787, new_n788, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n815, new_n816, new_n817,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n869,
    new_n870, new_n871, new_n872, new_n874, new_n875, new_n876, new_n877,
    new_n879, new_n880, new_n881, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n922, new_n923,
    new_n925, new_n926, new_n927, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n940, new_n941,
    new_n942, new_n943, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n983, new_n984;
  INV_X1    g000(.A(KEYINPUT36), .ZN(new_n202));
  INV_X1    g001(.A(G127gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n203), .A2(G134gat), .ZN(new_n204));
  INV_X1    g003(.A(G134gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n205), .A2(G127gat), .ZN(new_n206));
  OAI21_X1  g005(.A(KEYINPUT70), .B1(new_n204), .B2(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n205), .A2(G127gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n203), .A2(G134gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT70), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n208), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT1), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n212), .B1(G113gat), .B2(G120gat), .ZN(new_n213));
  AND2_X1   g012(.A1(G113gat), .A2(G120gat), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n207), .A2(new_n211), .A3(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(G127gat), .B(G134gat), .ZN(new_n217));
  OAI211_X1 g016(.A(new_n217), .B(new_n210), .C1(new_n214), .C2(new_n213), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT25), .ZN(new_n220));
  INV_X1    g019(.A(G169gat), .ZN(new_n221));
  INV_X1    g020(.A(G176gat), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n221), .A2(new_n222), .A3(KEYINPUT23), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT65), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NOR2_X1   g024(.A1(G169gat), .A2(G176gat), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n226), .A2(KEYINPUT65), .A3(KEYINPUT23), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g027(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(G183gat), .A2(G190gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT64), .ZN(new_n232));
  NAND4_X1  g031(.A1(new_n232), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n233));
  NAND3_X1  g032(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(KEYINPUT64), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n231), .A2(new_n233), .A3(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT23), .ZN(new_n237));
  OAI211_X1 g036(.A(new_n237), .B(KEYINPUT66), .C1(G169gat), .C2(G176gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(G169gat), .A2(G176gat), .ZN(new_n239));
  AND2_X1   g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT66), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n241), .B1(new_n226), .B2(KEYINPUT23), .ZN(new_n242));
  NAND4_X1  g041(.A1(new_n228), .A2(new_n236), .A3(new_n240), .A4(new_n242), .ZN(new_n243));
  AND2_X1   g042(.A1(new_n240), .A2(new_n242), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n223), .A2(KEYINPUT25), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n245), .B1(new_n234), .B2(new_n231), .ZN(new_n246));
  AOI22_X1  g045(.A1(new_n220), .A2(new_n243), .B1(new_n244), .B2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(G183gat), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(KEYINPUT27), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT27), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(G183gat), .ZN(new_n251));
  INV_X1    g050(.A(G190gat), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n249), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n253), .A2(KEYINPUT67), .A3(KEYINPUT28), .ZN(new_n254));
  OAI21_X1  g053(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT68), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n255), .B(new_n256), .ZN(new_n257));
  OR2_X1    g056(.A1(KEYINPUT69), .A2(KEYINPUT26), .ZN(new_n258));
  NAND2_X1  g057(.A1(KEYINPUT69), .A2(KEYINPUT26), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n258), .A2(new_n226), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(new_n239), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n254), .B1(new_n257), .B2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT67), .ZN(new_n263));
  XNOR2_X1  g062(.A(KEYINPUT27), .B(G183gat), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n263), .B1(new_n264), .B2(new_n252), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n230), .B1(new_n265), .B2(KEYINPUT28), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n262), .A2(new_n266), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n219), .B1(new_n247), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n243), .A2(new_n220), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n244), .A2(new_n246), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  OR2_X1    g070(.A1(new_n265), .A2(KEYINPUT28), .ZN(new_n272));
  XNOR2_X1  g071(.A(new_n255), .B(KEYINPUT68), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n273), .A2(new_n239), .A3(new_n260), .ZN(new_n274));
  NAND4_X1  g073(.A1(new_n272), .A2(new_n274), .A3(new_n230), .A4(new_n254), .ZN(new_n275));
  INV_X1    g074(.A(new_n219), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n271), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(G227gat), .ZN(new_n278));
  INV_X1    g077(.A(G233gat), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n268), .A2(new_n277), .A3(new_n280), .ZN(new_n281));
  XOR2_X1   g080(.A(G71gat), .B(G99gat), .Z(new_n282));
  XNOR2_X1  g081(.A(G15gat), .B(G43gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n282), .B(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(KEYINPUT33), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n281), .A2(KEYINPUT32), .A3(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT71), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND4_X1  g087(.A1(new_n281), .A2(KEYINPUT71), .A3(KEYINPUT32), .A4(new_n285), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT34), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n268), .A2(new_n277), .ZN(new_n292));
  INV_X1    g091(.A(new_n280), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n291), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  AOI211_X1 g093(.A(KEYINPUT34), .B(new_n280), .C1(new_n268), .C2(new_n277), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n281), .A2(KEYINPUT32), .ZN(new_n297));
  INV_X1    g096(.A(new_n281), .ZN(new_n298));
  OAI211_X1 g097(.A(new_n297), .B(new_n284), .C1(new_n298), .C2(KEYINPUT33), .ZN(new_n299));
  AND3_X1   g098(.A1(new_n290), .A2(new_n296), .A3(new_n299), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n296), .B1(new_n290), .B2(new_n299), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n202), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n290), .A2(new_n299), .ZN(new_n303));
  INV_X1    g102(.A(new_n296), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n290), .A2(new_n296), .A3(new_n299), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n305), .A2(KEYINPUT36), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n302), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT81), .ZN(new_n309));
  XNOR2_X1  g108(.A(KEYINPUT78), .B(KEYINPUT31), .ZN(new_n310));
  INV_X1    g109(.A(G228gat), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n311), .A2(new_n279), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  AND2_X1   g112(.A1(G211gat), .A2(G218gat), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n314), .A2(KEYINPUT22), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(G197gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(KEYINPUT72), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT72), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(G197gat), .ZN(new_n320));
  AND3_X1   g119(.A1(new_n318), .A2(new_n320), .A3(G204gat), .ZN(new_n321));
  AOI21_X1  g120(.A(G204gat), .B1(new_n318), .B2(new_n320), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n316), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NOR2_X1   g122(.A1(G211gat), .A2(G218gat), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n314), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(G204gat), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n319), .A2(G197gat), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n317), .A2(KEYINPUT72), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n327), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n318), .A2(new_n320), .A3(G204gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(new_n325), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n332), .A2(new_n333), .A3(new_n316), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n326), .A2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT29), .ZN(new_n336));
  AND2_X1   g135(.A1(G155gat), .A2(G162gat), .ZN(new_n337));
  NOR2_X1   g136(.A1(G155gat), .A2(G162gat), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  XNOR2_X1  g138(.A(G141gat), .B(G148gat), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT2), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n341), .B1(G155gat), .B2(G162gat), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n339), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(G141gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(G148gat), .ZN(new_n345));
  INV_X1    g144(.A(G148gat), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(G141gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  XNOR2_X1  g147(.A(G155gat), .B(G162gat), .ZN(new_n349));
  INV_X1    g148(.A(G155gat), .ZN(new_n350));
  INV_X1    g149(.A(G162gat), .ZN(new_n351));
  OAI21_X1  g150(.A(KEYINPUT2), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n348), .A2(new_n349), .A3(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT3), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n343), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n335), .B1(new_n336), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n343), .A2(new_n353), .ZN(new_n357));
  AOI21_X1  g156(.A(KEYINPUT29), .B1(new_n326), .B2(new_n334), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n357), .B1(new_n358), .B2(KEYINPUT3), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n356), .B1(new_n359), .B2(KEYINPUT80), .ZN(new_n360));
  AND2_X1   g159(.A1(new_n343), .A2(new_n353), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n333), .B1(new_n332), .B2(new_n316), .ZN(new_n362));
  AOI211_X1 g161(.A(new_n325), .B(new_n315), .C1(new_n330), .C2(new_n331), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n336), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n361), .B1(new_n364), .B2(new_n354), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT80), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n313), .B1(new_n360), .B2(new_n367), .ZN(new_n368));
  AND3_X1   g167(.A1(new_n326), .A2(KEYINPUT79), .A3(new_n334), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n336), .B1(new_n326), .B2(KEYINPUT79), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n354), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  AOI211_X1 g170(.A(new_n312), .B(new_n356), .C1(new_n371), .C2(new_n357), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n310), .B1(new_n368), .B2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n335), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n355), .A2(new_n336), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n376), .B1(new_n365), .B2(new_n366), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n359), .A2(KEYINPUT80), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n312), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n371), .A2(new_n357), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n380), .A2(new_n313), .A3(new_n376), .ZN(new_n381));
  INV_X1    g180(.A(new_n310), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n379), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  XNOR2_X1  g182(.A(G78gat), .B(G106gat), .ZN(new_n384));
  INV_X1    g183(.A(G50gat), .ZN(new_n385));
  XNOR2_X1  g184(.A(new_n384), .B(new_n385), .ZN(new_n386));
  XNOR2_X1  g185(.A(new_n386), .B(G22gat), .ZN(new_n387));
  AND3_X1   g186(.A1(new_n373), .A2(new_n383), .A3(new_n387), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n387), .B1(new_n373), .B2(new_n383), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n309), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(new_n387), .ZN(new_n391));
  NOR3_X1   g190(.A1(new_n368), .A2(new_n372), .A3(new_n310), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n382), .B1(new_n379), .B2(new_n381), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n391), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n373), .A2(new_n383), .A3(new_n387), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n394), .A2(KEYINPUT81), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n390), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(G226gat), .A2(G233gat), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  NOR3_X1   g198(.A1(new_n247), .A2(new_n267), .A3(new_n399), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n399), .A2(KEYINPUT29), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n401), .B1(new_n271), .B2(new_n275), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n374), .B1(new_n400), .B2(new_n402), .ZN(new_n403));
  OAI22_X1  g202(.A1(new_n247), .A2(new_n267), .B1(KEYINPUT29), .B2(new_n399), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n271), .A2(new_n275), .A3(new_n398), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n404), .A2(new_n405), .A3(new_n335), .ZN(new_n406));
  XNOR2_X1  g205(.A(G8gat), .B(G36gat), .ZN(new_n407));
  XNOR2_X1  g206(.A(G64gat), .B(G92gat), .ZN(new_n408));
  XOR2_X1   g207(.A(new_n407), .B(new_n408), .Z(new_n409));
  NAND3_X1  g208(.A1(new_n403), .A2(new_n406), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(KEYINPUT73), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT30), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT73), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n403), .A2(new_n406), .A3(new_n413), .A4(new_n409), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n411), .A2(new_n412), .A3(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(new_n409), .ZN(new_n416));
  AND3_X1   g215(.A1(new_n404), .A2(new_n405), .A3(new_n335), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n335), .B1(new_n404), .B2(new_n405), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n416), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND4_X1  g218(.A1(new_n403), .A2(new_n406), .A3(KEYINPUT30), .A4(new_n409), .ZN(new_n420));
  AND2_X1   g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n415), .A2(new_n421), .ZN(new_n422));
  XOR2_X1   g221(.A(KEYINPUT76), .B(KEYINPUT6), .Z(new_n423));
  INV_X1    g222(.A(KEYINPUT4), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n219), .A2(new_n361), .A3(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT75), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n219), .A2(new_n361), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(KEYINPUT4), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n219), .A2(new_n361), .A3(KEYINPUT75), .A4(new_n424), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n427), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n355), .A2(new_n218), .A3(new_n216), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n354), .B1(new_n343), .B2(new_n353), .ZN(new_n433));
  OAI21_X1  g232(.A(KEYINPUT74), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n357), .A2(KEYINPUT3), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT74), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n276), .A2(new_n435), .A3(new_n436), .A4(new_n355), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n434), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(G225gat), .A2(G233gat), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n431), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n439), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n357), .A2(new_n218), .A3(new_n216), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n357), .B1(new_n218), .B2(new_n216), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n441), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(KEYINPUT5), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n440), .A2(new_n447), .ZN(new_n448));
  XNOR2_X1  g247(.A(G1gat), .B(G29gat), .ZN(new_n449));
  XNOR2_X1  g248(.A(new_n449), .B(KEYINPUT0), .ZN(new_n450));
  XNOR2_X1  g249(.A(G57gat), .B(G85gat), .ZN(new_n451));
  XNOR2_X1  g250(.A(new_n450), .B(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n441), .B1(new_n434), .B2(new_n437), .ZN(new_n453));
  AOI21_X1  g252(.A(KEYINPUT5), .B1(new_n429), .B2(new_n425), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n452), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n423), .B1(new_n448), .B2(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n446), .B1(new_n453), .B2(new_n431), .ZN(new_n457));
  AND2_X1   g256(.A1(new_n453), .A2(new_n454), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n452), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n456), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT77), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n456), .A2(new_n459), .A3(KEYINPUT77), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  OAI211_X1 g263(.A(new_n452), .B(new_n423), .C1(new_n457), .C2(new_n458), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n422), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n308), .B1(new_n397), .B2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT82), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NOR3_X1   g268(.A1(new_n417), .A2(new_n418), .A3(KEYINPUT85), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT85), .ZN(new_n471));
  OAI21_X1  g270(.A(KEYINPUT37), .B1(new_n406), .B2(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n409), .B1(new_n403), .B2(new_n406), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT37), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n409), .A2(new_n474), .ZN(new_n475));
  OAI22_X1  g274(.A1(new_n470), .A2(new_n472), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT38), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n419), .B1(new_n474), .B2(new_n409), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n403), .A2(new_n406), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n477), .B1(new_n479), .B2(KEYINPUT37), .ZN(new_n480));
  AOI22_X1  g279(.A1(new_n476), .A2(new_n477), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n460), .A2(new_n411), .A3(new_n414), .A4(new_n465), .ZN(new_n482));
  OAI211_X1 g281(.A(new_n395), .B(new_n394), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n428), .A2(new_n439), .A3(new_n442), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(KEYINPUT39), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(KEYINPUT83), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT83), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n484), .A2(new_n487), .A3(KEYINPUT39), .ZN(new_n488));
  AOI22_X1  g287(.A1(new_n434), .A2(new_n437), .B1(new_n429), .B2(new_n425), .ZN(new_n489));
  OAI211_X1 g288(.A(new_n486), .B(new_n488), .C1(new_n489), .C2(new_n439), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n429), .A2(new_n425), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n438), .A2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT39), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n492), .A2(new_n493), .A3(new_n441), .ZN(new_n494));
  INV_X1    g293(.A(new_n452), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n490), .A2(new_n494), .A3(KEYINPUT40), .A4(new_n495), .ZN(new_n496));
  AND2_X1   g295(.A1(new_n496), .A2(new_n459), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n439), .B1(new_n438), .B2(new_n491), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n452), .B1(new_n498), .B2(new_n493), .ZN(new_n499));
  AOI211_X1 g298(.A(KEYINPUT84), .B(KEYINPUT40), .C1(new_n499), .C2(new_n490), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT84), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n490), .A2(new_n495), .A3(new_n494), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT40), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n497), .B1(new_n500), .B2(new_n504), .ZN(new_n505));
  AND2_X1   g304(.A1(new_n415), .A2(new_n421), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  OAI21_X1  g306(.A(KEYINPUT86), .B1(new_n483), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n460), .A2(new_n465), .ZN(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  AND2_X1   g309(.A1(new_n411), .A2(new_n414), .ZN(new_n511));
  AND2_X1   g310(.A1(new_n476), .A2(new_n477), .ZN(new_n512));
  AND2_X1   g311(.A1(new_n478), .A2(new_n480), .ZN(new_n513));
  OAI211_X1 g312(.A(new_n510), .B(new_n511), .C1(new_n512), .C2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n394), .A2(new_n395), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  OAI211_X1 g315(.A(new_n422), .B(new_n497), .C1(new_n504), .C2(new_n500), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT86), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n514), .A2(new_n516), .A3(new_n517), .A4(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n508), .A2(new_n519), .ZN(new_n520));
  OAI211_X1 g319(.A(new_n308), .B(KEYINPUT82), .C1(new_n397), .C2(new_n466), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n469), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT87), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n305), .A2(new_n306), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n524), .A2(new_n515), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(new_n466), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(KEYINPUT35), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n506), .A2(new_n305), .A3(new_n306), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n528), .A2(new_n515), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT35), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n529), .A2(new_n530), .A3(new_n509), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n527), .A2(new_n531), .ZN(new_n532));
  AND3_X1   g331(.A1(new_n522), .A2(new_n523), .A3(new_n532), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n523), .B1(new_n522), .B2(new_n532), .ZN(new_n534));
  XNOR2_X1  g333(.A(G15gat), .B(G22gat), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT16), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n535), .B1(new_n536), .B2(G1gat), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n537), .B1(G1gat), .B2(new_n535), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n538), .B(G8gat), .ZN(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(G29gat), .A2(G36gat), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n541), .B(KEYINPUT89), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n542), .B(KEYINPUT90), .ZN(new_n543));
  XNOR2_X1  g342(.A(G43gat), .B(G50gat), .ZN(new_n544));
  AND2_X1   g343(.A1(new_n544), .A2(KEYINPUT15), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n544), .A2(KEYINPUT15), .ZN(new_n546));
  NOR2_X1   g345(.A1(G29gat), .A2(G36gat), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n547), .B(KEYINPUT14), .ZN(new_n548));
  NOR3_X1   g347(.A1(new_n545), .A2(new_n546), .A3(new_n548), .ZN(new_n549));
  OR2_X1    g348(.A1(new_n548), .A2(new_n542), .ZN(new_n550));
  AOI22_X1  g349(.A1(new_n543), .A2(new_n549), .B1(new_n550), .B2(new_n545), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(KEYINPUT17), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT91), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n543), .A2(new_n549), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n550), .A2(new_n545), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT17), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n553), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NOR3_X1   g357(.A1(new_n551), .A2(KEYINPUT91), .A3(KEYINPUT17), .ZN(new_n559));
  OAI211_X1 g358(.A(new_n540), .B(new_n552), .C1(new_n558), .C2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n556), .A2(new_n539), .ZN(new_n561));
  NAND2_X1  g360(.A1(G229gat), .A2(G233gat), .ZN(new_n562));
  NAND4_X1  g361(.A1(new_n560), .A2(KEYINPUT18), .A3(new_n561), .A4(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n551), .B(new_n539), .ZN(new_n564));
  XOR2_X1   g363(.A(new_n562), .B(KEYINPUT13), .Z(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  OR2_X1    g365(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(G113gat), .B(G141gat), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n568), .B(G197gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(KEYINPUT11), .B(G169gat), .ZN(new_n570));
  XOR2_X1   g369(.A(new_n569), .B(new_n570), .Z(new_n571));
  XNOR2_X1  g370(.A(new_n571), .B(KEYINPUT12), .ZN(new_n572));
  AND3_X1   g371(.A1(new_n563), .A2(new_n567), .A3(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n560), .A2(new_n561), .A3(new_n562), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT18), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT92), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n574), .A2(KEYINPUT92), .A3(new_n575), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n573), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n580), .A2(KEYINPUT93), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT93), .ZN(new_n582));
  NAND4_X1  g381(.A1(new_n573), .A2(new_n578), .A3(new_n582), .A4(new_n579), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n576), .A2(new_n567), .A3(new_n563), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n572), .B(KEYINPUT88), .ZN(new_n585));
  AOI22_X1  g384(.A1(new_n581), .A2(new_n583), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NOR3_X1   g385(.A1(new_n533), .A2(new_n534), .A3(new_n586), .ZN(new_n587));
  XOR2_X1   g386(.A(G57gat), .B(G64gat), .Z(new_n588));
  INV_X1    g387(.A(KEYINPUT9), .ZN(new_n589));
  INV_X1    g388(.A(G71gat), .ZN(new_n590));
  INV_X1    g389(.A(G78gat), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n589), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n588), .A2(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(G71gat), .B(G78gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n593), .B(new_n594), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n595), .A2(KEYINPUT21), .ZN(new_n596));
  NAND2_X1  g395(.A1(G231gat), .A2(G233gat), .ZN(new_n597));
  XOR2_X1   g396(.A(new_n596), .B(new_n597), .Z(new_n598));
  XOR2_X1   g397(.A(G127gat), .B(G155gat), .Z(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(KEYINPUT20), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n598), .B(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(G183gat), .B(G211gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n595), .B(KEYINPUT95), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n539), .B1(new_n604), .B2(KEYINPUT21), .ZN(new_n605));
  XOR2_X1   g404(.A(KEYINPUT94), .B(KEYINPUT19), .Z(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  OR2_X1    g406(.A1(new_n603), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n603), .A2(new_n607), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(G85gat), .A2(G92gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n611), .B(KEYINPUT7), .ZN(new_n612));
  INV_X1    g411(.A(G99gat), .ZN(new_n613));
  INV_X1    g412(.A(G106gat), .ZN(new_n614));
  OAI21_X1  g413(.A(KEYINPUT8), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(KEYINPUT96), .B(G85gat), .ZN(new_n616));
  OAI211_X1 g415(.A(new_n612), .B(new_n615), .C1(G92gat), .C2(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(G99gat), .B(G106gat), .ZN(new_n618));
  XOR2_X1   g417(.A(new_n617), .B(new_n618), .Z(new_n619));
  OAI211_X1 g418(.A(new_n552), .B(new_n619), .C1(new_n558), .C2(new_n559), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n617), .B(new_n618), .ZN(new_n621));
  AND2_X1   g420(.A1(G232gat), .A2(G233gat), .ZN(new_n622));
  AOI22_X1  g421(.A1(new_n556), .A2(new_n621), .B1(KEYINPUT41), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n620), .A2(new_n623), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n622), .A2(KEYINPUT41), .ZN(new_n625));
  XNOR2_X1  g424(.A(G134gat), .B(G162gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n624), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(G190gat), .B(G218gat), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n620), .A2(new_n623), .A3(new_n627), .ZN(new_n632));
  AND3_X1   g431(.A1(new_n629), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n631), .B1(new_n629), .B2(new_n632), .ZN(new_n634));
  XNOR2_X1  g433(.A(KEYINPUT97), .B(KEYINPUT98), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  OR3_X1    g435(.A1(new_n633), .A2(new_n634), .A3(new_n636), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n636), .B1(new_n633), .B2(new_n634), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n610), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n595), .A2(KEYINPUT99), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT99), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n595), .B(new_n643), .ZN(new_n644));
  MUX2_X1   g443(.A(new_n642), .B(new_n644), .S(new_n621), .Z(new_n645));
  NAND2_X1  g444(.A1(G230gat), .A2(G233gat), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n619), .A2(new_n641), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT10), .ZN(new_n650));
  OAI211_X1 g449(.A(new_n649), .B(new_n650), .C1(new_n644), .C2(new_n619), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n604), .A2(KEYINPUT10), .A3(new_n621), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n653), .A2(new_n646), .ZN(new_n654));
  XNOR2_X1  g453(.A(G120gat), .B(G148gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(G176gat), .B(G204gat), .ZN(new_n656));
  XOR2_X1   g455(.A(new_n655), .B(new_n656), .Z(new_n657));
  AND3_X1   g456(.A1(new_n648), .A2(new_n654), .A3(new_n657), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n657), .B1(new_n648), .B2(new_n654), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n640), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n464), .A2(new_n465), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  AND2_X1   g463(.A1(new_n664), .A2(KEYINPUT100), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n664), .A2(KEYINPUT100), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n587), .A2(new_n662), .A3(new_n667), .ZN(new_n668));
  XNOR2_X1  g467(.A(KEYINPUT101), .B(G1gat), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n668), .B(new_n669), .ZN(G1324gat));
  NAND3_X1  g469(.A1(new_n587), .A2(new_n422), .A3(new_n662), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT42), .ZN(new_n672));
  XNOR2_X1  g471(.A(KEYINPUT16), .B(G8gat), .ZN(new_n673));
  NOR3_X1   g472(.A1(new_n671), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(KEYINPUT103), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n672), .B1(new_n671), .B2(new_n673), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT102), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n676), .B(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n671), .A2(G8gat), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n675), .A2(new_n678), .A3(new_n679), .ZN(G1325gat));
  NAND2_X1  g479(.A1(new_n587), .A2(new_n662), .ZN(new_n681));
  OAI21_X1  g480(.A(G15gat), .B1(new_n681), .B2(new_n308), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n522), .A2(new_n532), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(KEYINPUT87), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n522), .A2(new_n523), .A3(new_n532), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n581), .A2(new_n583), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n584), .A2(new_n585), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n684), .A2(new_n685), .A3(new_n688), .ZN(new_n689));
  OR3_X1    g488(.A1(new_n661), .A2(G15gat), .A3(new_n524), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n682), .B1(new_n689), .B2(new_n690), .ZN(G1326gat));
  NOR2_X1   g490(.A1(new_n681), .A2(new_n397), .ZN(new_n692));
  XOR2_X1   g491(.A(KEYINPUT43), .B(G22gat), .Z(new_n693));
  XNOR2_X1  g492(.A(new_n692), .B(new_n693), .ZN(G1327gat));
  NAND2_X1  g493(.A1(new_n610), .A2(new_n660), .ZN(new_n695));
  INV_X1    g494(.A(new_n639), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND4_X1  g496(.A1(new_n684), .A2(new_n685), .A3(new_n688), .A4(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n667), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n699), .A2(G29gat), .ZN(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(KEYINPUT45), .ZN(new_n703));
  INV_X1    g502(.A(G29gat), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT44), .ZN(new_n705));
  INV_X1    g504(.A(new_n532), .ZN(new_n706));
  AND2_X1   g505(.A1(new_n390), .A2(new_n396), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n663), .A2(new_n506), .ZN(new_n708));
  AOI22_X1  g507(.A1(new_n707), .A2(new_n708), .B1(new_n307), .B2(new_n302), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n520), .A2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT105), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n520), .A2(new_n709), .A3(KEYINPUT105), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n706), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n705), .B1(new_n714), .B2(new_n696), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n639), .A2(KEYINPUT44), .ZN(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n684), .A2(new_n685), .A3(new_n717), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n695), .A2(new_n586), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(KEYINPUT104), .ZN(new_n720));
  AND3_X1   g519(.A1(new_n715), .A2(new_n718), .A3(new_n720), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n704), .B1(new_n721), .B2(new_n667), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT106), .ZN(new_n723));
  OR3_X1    g522(.A1(new_n703), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n723), .B1(new_n703), .B2(new_n722), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(G1328gat));
  INV_X1    g525(.A(G36gat), .ZN(new_n727));
  NAND4_X1  g526(.A1(new_n715), .A2(new_n422), .A3(new_n718), .A4(new_n720), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT108), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n727), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NOR3_X1   g529(.A1(new_n533), .A2(new_n534), .A3(new_n716), .ZN(new_n731));
  AND3_X1   g530(.A1(new_n520), .A2(new_n709), .A3(KEYINPUT105), .ZN(new_n732));
  AOI21_X1  g531(.A(KEYINPUT105), .B1(new_n520), .B2(new_n709), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n532), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  AOI21_X1  g533(.A(KEYINPUT44), .B1(new_n734), .B2(new_n639), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n731), .A2(new_n735), .ZN(new_n736));
  NAND4_X1  g535(.A1(new_n736), .A2(KEYINPUT108), .A3(new_n422), .A4(new_n720), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n730), .A2(new_n737), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n506), .A2(G36gat), .ZN(new_n739));
  INV_X1    g538(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n698), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g540(.A(KEYINPUT107), .B(KEYINPUT46), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n741), .B(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n738), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(KEYINPUT109), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT109), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n738), .A2(new_n746), .A3(new_n743), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n745), .A2(new_n747), .ZN(G1329gat));
  NOR2_X1   g547(.A1(new_n524), .A2(G43gat), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n587), .A2(KEYINPUT110), .A3(new_n697), .A4(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT110), .ZN(new_n751));
  INV_X1    g550(.A(new_n749), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n751), .B1(new_n698), .B2(new_n752), .ZN(new_n753));
  AND2_X1   g552(.A1(new_n750), .A2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(new_n308), .ZN(new_n755));
  NAND4_X1  g554(.A1(new_n715), .A2(new_n755), .A3(new_n718), .A4(new_n720), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(G43gat), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n754), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(KEYINPUT111), .A2(KEYINPUT47), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT111), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT47), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n758), .A2(new_n759), .A3(new_n762), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n754), .A2(new_n760), .A3(new_n761), .A4(new_n757), .ZN(new_n764));
  AND2_X1   g563(.A1(new_n763), .A2(new_n764), .ZN(G1330gat));
  AOI21_X1  g564(.A(new_n385), .B1(new_n721), .B2(new_n707), .ZN(new_n766));
  INV_X1    g565(.A(new_n698), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n397), .A2(G50gat), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n766), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n385), .B1(new_n721), .B2(new_n515), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n767), .A2(new_n768), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(KEYINPUT48), .ZN(new_n772));
  OAI22_X1  g571(.A1(new_n769), .A2(KEYINPUT48), .B1(new_n770), .B2(new_n772), .ZN(G1331gat));
  INV_X1    g572(.A(new_n660), .ZN(new_n774));
  AND4_X1   g573(.A1(new_n586), .A2(new_n734), .A3(new_n640), .A4(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(new_n667), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g576(.A(new_n506), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n775), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n779), .B(KEYINPUT112), .ZN(new_n780));
  NOR2_X1   g579(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n780), .B(new_n781), .ZN(G1333gat));
  AOI21_X1  g581(.A(new_n590), .B1(new_n775), .B2(new_n755), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n524), .A2(G71gat), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n783), .B1(new_n775), .B2(new_n784), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n785), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g585(.A1(new_n775), .A2(new_n707), .ZN(new_n787));
  XOR2_X1   g586(.A(KEYINPUT113), .B(G78gat), .Z(new_n788));
  XNOR2_X1  g587(.A(new_n787), .B(new_n788), .ZN(G1335gat));
  INV_X1    g588(.A(new_n736), .ZN(new_n790));
  INV_X1    g589(.A(new_n610), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n791), .A2(new_n688), .ZN(new_n792));
  INV_X1    g591(.A(new_n792), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n793), .A2(new_n660), .ZN(new_n794));
  INV_X1    g593(.A(new_n794), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n790), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(new_n667), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(new_n616), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n734), .A2(new_n639), .A3(new_n792), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n799), .A2(KEYINPUT114), .A3(KEYINPUT51), .ZN(new_n800));
  XOR2_X1   g599(.A(KEYINPUT114), .B(KEYINPUT51), .Z(new_n801));
  NAND4_X1  g600(.A1(new_n734), .A2(new_n639), .A3(new_n792), .A4(new_n801), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n699), .A2(new_n616), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n800), .A2(new_n774), .A3(new_n802), .A4(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n798), .A2(new_n804), .ZN(G1336gat));
  INV_X1    g604(.A(KEYINPUT52), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n715), .A2(new_n422), .A3(new_n718), .A4(new_n794), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(G92gat), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n806), .B1(new_n808), .B2(KEYINPUT116), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n660), .A2(G92gat), .A3(new_n506), .ZN(new_n810));
  XOR2_X1   g609(.A(new_n810), .B(KEYINPUT115), .Z(new_n811));
  NAND3_X1  g610(.A1(new_n800), .A2(new_n802), .A3(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n808), .A2(new_n812), .ZN(new_n813));
  XNOR2_X1  g612(.A(new_n809), .B(new_n813), .ZN(G1337gat));
  NOR2_X1   g613(.A1(new_n524), .A2(G99gat), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n800), .A2(new_n774), .A3(new_n802), .A4(new_n815), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n790), .A2(new_n308), .A3(new_n795), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n816), .B1(new_n817), .B2(new_n613), .ZN(G1338gat));
  NAND4_X1  g617(.A1(new_n715), .A2(new_n707), .A3(new_n718), .A4(new_n794), .ZN(new_n819));
  AND3_X1   g618(.A1(new_n819), .A2(KEYINPUT117), .A3(G106gat), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n516), .A2(G106gat), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n800), .A2(new_n774), .A3(new_n802), .A4(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(new_n822), .ZN(new_n823));
  AOI21_X1  g622(.A(KEYINPUT117), .B1(new_n819), .B2(G106gat), .ZN(new_n824));
  NOR3_X1   g623(.A1(new_n820), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT53), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n614), .B1(new_n796), .B2(new_n515), .ZN(new_n827));
  XNOR2_X1  g626(.A(KEYINPUT118), .B(KEYINPUT53), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n822), .A2(new_n828), .ZN(new_n829));
  OAI22_X1  g628(.A1(new_n825), .A2(new_n826), .B1(new_n827), .B2(new_n829), .ZN(G1339gat));
  AND2_X1   g629(.A1(new_n653), .A2(new_n646), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT54), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n657), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  OR2_X1    g632(.A1(new_n653), .A2(new_n646), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n834), .A2(KEYINPUT54), .A3(new_n654), .ZN(new_n835));
  AOI21_X1  g634(.A(KEYINPUT55), .B1(new_n833), .B2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(new_n836), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n833), .A2(new_n835), .A3(KEYINPUT55), .ZN(new_n838));
  INV_X1    g637(.A(new_n658), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(new_n840), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n688), .A2(new_n837), .A3(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(new_n571), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n564), .A2(new_n566), .ZN(new_n844));
  XNOR2_X1  g643(.A(new_n844), .B(KEYINPUT119), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n560), .A2(new_n561), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n846), .A2(G229gat), .A3(G233gat), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n843), .B1(new_n845), .B2(new_n847), .ZN(new_n848));
  AOI211_X1 g647(.A(new_n848), .B(new_n660), .C1(new_n581), .C2(new_n583), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n639), .B1(new_n842), .B2(new_n850), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n840), .A2(new_n836), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n848), .B1(new_n581), .B2(new_n583), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n852), .A2(new_n853), .A3(new_n639), .ZN(new_n854));
  INV_X1    g653(.A(new_n854), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n610), .B1(new_n851), .B2(new_n855), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n661), .A2(new_n688), .ZN(new_n857));
  INV_X1    g656(.A(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n707), .B1(new_n856), .B2(new_n858), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n699), .A2(new_n528), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(G113gat), .B1(new_n861), .B2(new_n586), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n856), .A2(new_n858), .ZN(new_n863));
  AND2_X1   g662(.A1(new_n667), .A2(new_n529), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n586), .A2(G113gat), .ZN(new_n866));
  XNOR2_X1  g665(.A(new_n866), .B(KEYINPUT120), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n862), .B1(new_n865), .B2(new_n867), .ZN(G1340gat));
  INV_X1    g667(.A(new_n865), .ZN(new_n869));
  AOI21_X1  g668(.A(G120gat), .B1(new_n869), .B2(new_n774), .ZN(new_n870));
  INV_X1    g669(.A(G120gat), .ZN(new_n871));
  NOR3_X1   g670(.A1(new_n861), .A2(new_n871), .A3(new_n660), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n870), .A2(new_n872), .ZN(G1341gat));
  NAND4_X1  g672(.A1(new_n859), .A2(G127gat), .A3(new_n791), .A4(new_n860), .ZN(new_n874));
  AND2_X1   g673(.A1(new_n874), .A2(KEYINPUT121), .ZN(new_n875));
  AOI21_X1  g674(.A(G127gat), .B1(new_n869), .B2(new_n791), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n874), .A2(KEYINPUT121), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(G1342gat));
  NOR3_X1   g677(.A1(new_n865), .A2(G134gat), .A3(new_n696), .ZN(new_n879));
  XNOR2_X1  g678(.A(new_n879), .B(KEYINPUT56), .ZN(new_n880));
  OAI21_X1  g679(.A(G134gat), .B1(new_n861), .B2(new_n696), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n881), .ZN(G1343gat));
  NOR3_X1   g681(.A1(new_n699), .A2(new_n422), .A3(new_n755), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n586), .A2(new_n344), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n707), .A2(KEYINPUT57), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n836), .A2(KEYINPUT123), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT123), .ZN(new_n887));
  AOI211_X1 g686(.A(new_n887), .B(KEYINPUT55), .C1(new_n833), .C2(new_n835), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n889), .A2(new_n688), .A3(new_n841), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n639), .B1(new_n890), .B2(new_n850), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n610), .B1(new_n891), .B2(new_n855), .ZN(new_n892));
  OR2_X1    g691(.A1(new_n892), .A2(KEYINPUT124), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n857), .B1(new_n892), .B2(KEYINPUT124), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n885), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n516), .B1(new_n856), .B2(new_n858), .ZN(new_n896));
  XNOR2_X1  g695(.A(KEYINPUT122), .B(KEYINPUT57), .ZN(new_n897));
  INV_X1    g696(.A(new_n897), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  OAI211_X1 g698(.A(new_n883), .B(new_n884), .C1(new_n895), .C2(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n896), .A2(new_n883), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n344), .B1(new_n901), .B2(new_n586), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT58), .ZN(new_n904));
  XNOR2_X1  g703(.A(new_n903), .B(new_n904), .ZN(G1344gat));
  OR2_X1    g704(.A1(new_n895), .A2(new_n899), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT59), .ZN(new_n907));
  NAND4_X1  g706(.A1(new_n906), .A2(new_n907), .A3(new_n774), .A4(new_n883), .ZN(new_n908));
  AND3_X1   g707(.A1(new_n896), .A2(new_n774), .A3(new_n883), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n346), .B1(new_n909), .B2(new_n907), .ZN(new_n910));
  NOR3_X1   g709(.A1(new_n586), .A2(new_n836), .A3(new_n840), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n696), .B1(new_n911), .B2(new_n849), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n791), .B1(new_n912), .B2(new_n854), .ZN(new_n913));
  OAI211_X1 g712(.A(new_n515), .B(new_n898), .C1(new_n913), .C2(new_n857), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n397), .B1(new_n892), .B2(new_n858), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n914), .B1(new_n915), .B2(KEYINPUT57), .ZN(new_n916));
  AND3_X1   g715(.A1(new_n916), .A2(new_n774), .A3(new_n883), .ZN(new_n917));
  NAND2_X1  g716(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n918));
  OAI211_X1 g717(.A(new_n908), .B(new_n910), .C1(new_n917), .C2(new_n918), .ZN(G1345gat));
  INV_X1    g718(.A(new_n901), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n920), .A2(new_n350), .A3(new_n791), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n906), .A2(new_n791), .A3(new_n883), .ZN(new_n922));
  INV_X1    g721(.A(new_n922), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n921), .B1(new_n923), .B2(new_n350), .ZN(G1346gat));
  NAND3_X1  g723(.A1(new_n920), .A2(new_n351), .A3(new_n639), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n906), .A2(new_n639), .A3(new_n883), .ZN(new_n926));
  INV_X1    g725(.A(new_n926), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n925), .B1(new_n927), .B2(new_n351), .ZN(G1347gat));
  NAND2_X1  g727(.A1(new_n699), .A2(new_n422), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n929), .B1(new_n856), .B2(new_n858), .ZN(new_n930));
  AND2_X1   g729(.A1(new_n930), .A2(new_n525), .ZN(new_n931));
  AOI21_X1  g730(.A(G169gat), .B1(new_n931), .B2(new_n688), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n929), .A2(new_n524), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n859), .A2(new_n933), .ZN(new_n934));
  NOR3_X1   g733(.A1(new_n934), .A2(new_n221), .A3(new_n586), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n932), .A2(new_n935), .ZN(G1348gat));
  NAND3_X1  g735(.A1(new_n931), .A2(new_n222), .A3(new_n774), .ZN(new_n937));
  OAI21_X1  g736(.A(G176gat), .B1(new_n934), .B2(new_n660), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(G1349gat));
  NAND3_X1  g738(.A1(new_n931), .A2(new_n264), .A3(new_n791), .ZN(new_n940));
  OAI21_X1  g739(.A(G183gat), .B1(new_n934), .B2(new_n610), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  XNOR2_X1  g741(.A(KEYINPUT125), .B(KEYINPUT60), .ZN(new_n943));
  XNOR2_X1  g742(.A(new_n942), .B(new_n943), .ZN(G1350gat));
  NAND3_X1  g743(.A1(new_n931), .A2(new_n252), .A3(new_n639), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n859), .A2(new_n639), .A3(new_n933), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT61), .ZN(new_n947));
  AND3_X1   g746(.A1(new_n946), .A2(new_n947), .A3(G190gat), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n947), .B1(new_n946), .B2(G190gat), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n945), .B1(new_n948), .B2(new_n949), .ZN(G1351gat));
  NOR2_X1   g749(.A1(new_n755), .A2(new_n516), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n930), .A2(new_n951), .ZN(new_n952));
  INV_X1    g751(.A(new_n952), .ZN(new_n953));
  AOI21_X1  g752(.A(G197gat), .B1(new_n953), .B2(new_n688), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n699), .A2(new_n422), .A3(new_n308), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT57), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n586), .A2(new_n840), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n849), .B1(new_n957), .B2(new_n889), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n854), .B1(new_n958), .B2(new_n639), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n857), .B1(new_n959), .B2(new_n610), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n956), .B1(new_n960), .B2(new_n397), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n955), .B1(new_n961), .B2(new_n914), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n586), .A2(new_n317), .ZN(new_n963));
  AOI21_X1  g762(.A(new_n954), .B1(new_n962), .B2(new_n963), .ZN(G1352gat));
  NOR3_X1   g763(.A1(new_n952), .A2(G204gat), .A3(new_n660), .ZN(new_n965));
  XNOR2_X1  g764(.A(new_n965), .B(KEYINPUT62), .ZN(new_n966));
  INV_X1    g765(.A(new_n955), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n916), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g767(.A(G204gat), .B1(new_n968), .B2(new_n660), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n966), .A2(new_n969), .ZN(G1353gat));
  NAND4_X1  g769(.A1(new_n916), .A2(KEYINPUT127), .A3(new_n791), .A4(new_n967), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n971), .A2(G211gat), .ZN(new_n972));
  AOI21_X1  g771(.A(KEYINPUT127), .B1(new_n962), .B2(new_n791), .ZN(new_n973));
  OAI21_X1  g772(.A(KEYINPUT63), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  INV_X1    g773(.A(KEYINPUT127), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n975), .B1(new_n968), .B2(new_n610), .ZN(new_n976));
  INV_X1    g775(.A(KEYINPUT63), .ZN(new_n977));
  NAND4_X1  g776(.A1(new_n976), .A2(new_n977), .A3(G211gat), .A4(new_n971), .ZN(new_n978));
  OR2_X1    g777(.A1(new_n610), .A2(G211gat), .ZN(new_n979));
  NOR2_X1   g778(.A1(new_n952), .A2(new_n979), .ZN(new_n980));
  XOR2_X1   g779(.A(new_n980), .B(KEYINPUT126), .Z(new_n981));
  NAND3_X1  g780(.A1(new_n974), .A2(new_n978), .A3(new_n981), .ZN(G1354gat));
  OAI21_X1  g781(.A(G218gat), .B1(new_n968), .B2(new_n696), .ZN(new_n983));
  OR2_X1    g782(.A1(new_n696), .A2(G218gat), .ZN(new_n984));
  OAI21_X1  g783(.A(new_n983), .B1(new_n952), .B2(new_n984), .ZN(G1355gat));
endmodule


