//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 1 1 1 1 0 1 0 0 1 0 1 1 0 1 1 1 1 0 0 1 1 1 0 1 1 1 1 1 1 0 0 0 0 0 1 0 1 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n741, new_n742, new_n743,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n775, new_n776, new_n777, new_n778, new_n779, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n819,
    new_n820, new_n821, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n864, new_n865, new_n866,
    new_n867, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n980, new_n981, new_n983, new_n984, new_n985, new_n986, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n999, new_n1000, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1036, new_n1037;
  INV_X1    g000(.A(KEYINPUT90), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT32), .ZN(new_n203));
  AND2_X1   g002(.A1(G183gat), .A2(G190gat), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT24), .ZN(new_n205));
  AOI22_X1  g004(.A1(new_n204), .A2(new_n205), .B1(G169gat), .B2(G176gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT23), .ZN(new_n207));
  INV_X1    g006(.A(G169gat), .ZN(new_n208));
  INV_X1    g007(.A(G176gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n207), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  OAI21_X1  g009(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G183gat), .ZN(new_n213));
  INV_X1    g012(.A(G190gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(G183gat), .A2(G190gat), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n215), .A2(KEYINPUT24), .A3(new_n216), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n206), .A2(new_n212), .A3(new_n217), .ZN(new_n218));
  XOR2_X1   g017(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(KEYINPUT65), .ZN(new_n221));
  NAND4_X1  g020(.A1(new_n206), .A2(new_n212), .A3(new_n217), .A4(KEYINPUT25), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT65), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n218), .A2(new_n223), .A3(new_n219), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n221), .A2(new_n222), .A3(new_n224), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n208), .A2(new_n209), .A3(KEYINPUT67), .ZN(new_n226));
  AOI22_X1  g025(.A1(new_n226), .A2(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT26), .ZN(new_n228));
  NAND4_X1  g027(.A1(new_n228), .A2(new_n208), .A3(new_n209), .A4(KEYINPUT67), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n204), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT66), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n213), .A2(KEYINPUT27), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT27), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n233), .A2(G183gat), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n231), .B1(new_n232), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n233), .A2(G183gat), .ZN(new_n236));
  AOI21_X1  g035(.A(G190gat), .B1(new_n236), .B2(KEYINPUT66), .ZN(new_n237));
  AOI21_X1  g036(.A(KEYINPUT28), .B1(new_n235), .B2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n214), .A2(KEYINPUT28), .ZN(new_n239));
  NOR3_X1   g038(.A1(new_n232), .A2(new_n234), .A3(new_n239), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n230), .B1(new_n238), .B2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(KEYINPUT68), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT68), .ZN(new_n243));
  OAI211_X1 g042(.A(new_n230), .B(new_n243), .C1(new_n238), .C2(new_n240), .ZN(new_n244));
  AND3_X1   g043(.A1(new_n225), .A2(new_n242), .A3(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(G127gat), .B(G134gat), .ZN(new_n246));
  XOR2_X1   g045(.A(G113gat), .B(G120gat), .Z(new_n247));
  INV_X1    g046(.A(KEYINPUT1), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n246), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n246), .A2(new_n248), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(G120gat), .ZN(new_n252));
  OAI21_X1  g051(.A(KEYINPUT70), .B1(new_n252), .B2(G113gat), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT70), .ZN(new_n254));
  INV_X1    g053(.A(G113gat), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n254), .A2(new_n255), .A3(G120gat), .ZN(new_n256));
  AND2_X1   g055(.A1(new_n253), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT69), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n258), .B1(new_n255), .B2(G120gat), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n252), .A2(KEYINPUT69), .A3(G113gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NOR3_X1   g060(.A1(new_n257), .A2(KEYINPUT71), .A3(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT71), .ZN(new_n263));
  AND2_X1   g062(.A1(new_n259), .A2(new_n260), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n253), .A2(new_n256), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n263), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n251), .B1(new_n262), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(KEYINPUT72), .ZN(new_n268));
  OAI21_X1  g067(.A(KEYINPUT71), .B1(new_n257), .B2(new_n261), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n264), .A2(new_n263), .A3(new_n265), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT72), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n271), .A2(new_n272), .A3(new_n251), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n249), .B1(new_n268), .B2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT73), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n245), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n249), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n272), .B1(new_n271), .B2(new_n251), .ZN(new_n278));
  AOI211_X1 g077(.A(KEYINPUT72), .B(new_n250), .C1(new_n269), .C2(new_n270), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n277), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n225), .A2(new_n242), .A3(new_n244), .ZN(new_n281));
  OAI21_X1  g080(.A(KEYINPUT73), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n280), .A2(new_n281), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n276), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(G227gat), .A2(G233gat), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n203), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  AOI21_X1  g086(.A(KEYINPUT33), .B1(new_n284), .B2(new_n286), .ZN(new_n288));
  XNOR2_X1  g087(.A(G15gat), .B(G43gat), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n289), .B(KEYINPUT74), .ZN(new_n290));
  XNOR2_X1  g089(.A(G71gat), .B(G99gat), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n290), .B(new_n291), .ZN(new_n292));
  NOR3_X1   g091(.A1(new_n287), .A2(new_n288), .A3(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n292), .ZN(new_n294));
  OR2_X1    g093(.A1(new_n294), .A2(KEYINPUT75), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(KEYINPUT75), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n295), .A2(KEYINPUT33), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n287), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  NAND4_X1  g098(.A1(new_n276), .A2(new_n282), .A3(new_n285), .A4(new_n283), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n300), .B(KEYINPUT34), .ZN(new_n301));
  NOR3_X1   g100(.A1(new_n293), .A2(new_n299), .A3(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT34), .ZN(new_n303));
  XNOR2_X1  g102(.A(new_n300), .B(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(new_n287), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n284), .A2(new_n286), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT33), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n305), .A2(new_n308), .A3(new_n294), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n304), .B1(new_n309), .B2(new_n298), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n202), .B1(new_n302), .B2(new_n310), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n301), .B1(new_n293), .B2(new_n299), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n309), .A2(new_n304), .A3(new_n298), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n312), .A2(KEYINPUT90), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n311), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(G226gat), .A2(G233gat), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n245), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n224), .A2(new_n222), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n223), .B1(new_n218), .B2(new_n219), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n241), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(KEYINPUT78), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n317), .A2(KEYINPUT29), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT78), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n225), .A2(new_n324), .A3(new_n241), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n322), .A2(new_n323), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n318), .A2(new_n326), .ZN(new_n327));
  XNOR2_X1  g126(.A(G197gat), .B(G204gat), .ZN(new_n328));
  INV_X1    g127(.A(G211gat), .ZN(new_n329));
  INV_X1    g128(.A(G218gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(KEYINPUT76), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT76), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(G218gat), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n329), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n328), .B1(new_n334), .B2(KEYINPUT22), .ZN(new_n335));
  XOR2_X1   g134(.A(G211gat), .B(G218gat), .Z(new_n336));
  NAND3_X1  g135(.A1(new_n335), .A2(KEYINPUT77), .A3(new_n336), .ZN(new_n337));
  XNOR2_X1  g136(.A(G211gat), .B(G218gat), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT77), .ZN(new_n339));
  OAI221_X1 g138(.A(new_n328), .B1(new_n338), .B2(new_n339), .C1(new_n334), .C2(KEYINPUT22), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n337), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n327), .A2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n341), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n281), .A2(new_n323), .ZN(new_n344));
  AND2_X1   g143(.A1(new_n322), .A2(new_n325), .ZN(new_n345));
  OAI211_X1 g144(.A(new_n343), .B(new_n344), .C1(new_n345), .C2(new_n316), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n342), .A2(new_n346), .A3(KEYINPUT79), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n316), .B1(new_n322), .B2(new_n325), .ZN(new_n348));
  AND2_X1   g147(.A1(new_n281), .A2(new_n323), .ZN(new_n349));
  NOR3_X1   g148(.A1(new_n348), .A2(new_n349), .A3(new_n341), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT79), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n347), .A2(new_n352), .ZN(new_n353));
  XNOR2_X1  g152(.A(G8gat), .B(G36gat), .ZN(new_n354));
  XNOR2_X1  g153(.A(G64gat), .B(G92gat), .ZN(new_n355));
  XOR2_X1   g154(.A(new_n354), .B(new_n355), .Z(new_n356));
  NAND2_X1  g155(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT30), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n356), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n347), .A2(new_n352), .A3(new_n360), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n343), .B1(new_n318), .B2(new_n326), .ZN(new_n362));
  NOR3_X1   g161(.A1(new_n350), .A2(new_n362), .A3(new_n351), .ZN(new_n363));
  NOR4_X1   g162(.A1(new_n348), .A2(new_n349), .A3(KEYINPUT79), .A4(new_n341), .ZN(new_n364));
  OAI211_X1 g163(.A(KEYINPUT30), .B(new_n356), .C1(new_n363), .C2(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n359), .A2(new_n361), .A3(new_n365), .ZN(new_n366));
  AND2_X1   g165(.A1(G155gat), .A2(G162gat), .ZN(new_n367));
  NOR2_X1   g166(.A1(G155gat), .A2(G162gat), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  XNOR2_X1  g168(.A(G141gat), .B(G148gat), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT2), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n371), .B1(G155gat), .B2(G162gat), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n369), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(G141gat), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(G148gat), .ZN(new_n375));
  INV_X1    g174(.A(G148gat), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(G141gat), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  XNOR2_X1  g177(.A(G155gat), .B(G162gat), .ZN(new_n379));
  INV_X1    g178(.A(G155gat), .ZN(new_n380));
  INV_X1    g179(.A(G162gat), .ZN(new_n381));
  OAI21_X1  g180(.A(KEYINPUT2), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n378), .A2(new_n379), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n373), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  OAI211_X1 g184(.A(new_n385), .B(new_n277), .C1(new_n278), .C2(new_n279), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT4), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n268), .A2(new_n273), .ZN(new_n389));
  NAND4_X1  g188(.A1(new_n389), .A2(KEYINPUT4), .A3(new_n385), .A4(new_n277), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT3), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n373), .A2(new_n383), .A3(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT81), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND4_X1  g193(.A1(new_n373), .A2(new_n383), .A3(KEYINPUT81), .A4(new_n391), .ZN(new_n395));
  AOI22_X1  g194(.A1(new_n394), .A2(new_n395), .B1(KEYINPUT3), .B2(new_n384), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n280), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(G225gat), .A2(G233gat), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n388), .A2(new_n390), .A3(new_n397), .A4(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n280), .A2(new_n384), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n398), .B1(new_n400), .B2(new_n386), .ZN(new_n401));
  XOR2_X1   g200(.A(KEYINPUT82), .B(KEYINPUT5), .Z(new_n402));
  OAI21_X1  g201(.A(new_n399), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  XNOR2_X1  g202(.A(G1gat), .B(G29gat), .ZN(new_n404));
  XNOR2_X1  g203(.A(new_n404), .B(KEYINPUT0), .ZN(new_n405));
  XNOR2_X1  g204(.A(G57gat), .B(G85gat), .ZN(new_n406));
  XOR2_X1   g205(.A(new_n405), .B(new_n406), .Z(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  AOI22_X1  g207(.A1(new_n386), .A2(new_n387), .B1(new_n280), .B2(new_n396), .ZN(new_n409));
  INV_X1    g208(.A(new_n402), .ZN(new_n410));
  NAND4_X1  g209(.A1(new_n409), .A2(new_n398), .A3(new_n390), .A4(new_n410), .ZN(new_n411));
  XNOR2_X1  g210(.A(KEYINPUT83), .B(KEYINPUT6), .ZN(new_n412));
  NAND4_X1  g211(.A1(new_n403), .A2(new_n408), .A3(new_n411), .A4(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n403), .A2(new_n408), .A3(new_n411), .ZN(new_n415));
  INV_X1    g214(.A(new_n412), .ZN(new_n416));
  AND2_X1   g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n408), .B1(new_n403), .B2(new_n411), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n414), .B1(new_n417), .B2(new_n419), .ZN(new_n420));
  OAI21_X1  g219(.A(KEYINPUT89), .B1(new_n366), .B2(new_n420), .ZN(new_n421));
  XOR2_X1   g220(.A(G78gat), .B(G106gat), .Z(new_n422));
  XNOR2_X1  g221(.A(new_n422), .B(KEYINPUT84), .ZN(new_n423));
  XNOR2_X1  g222(.A(KEYINPUT31), .B(G50gat), .ZN(new_n424));
  XOR2_X1   g223(.A(new_n423), .B(new_n424), .Z(new_n425));
  INV_X1    g224(.A(KEYINPUT29), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n341), .A2(new_n426), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n385), .B1(new_n427), .B2(new_n391), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n394), .A2(new_n395), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n341), .B1(new_n429), .B2(new_n426), .ZN(new_n430));
  NAND2_X1  g229(.A1(G228gat), .A2(G233gat), .ZN(new_n431));
  OR3_X1    g230(.A1(new_n428), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  AOI21_X1  g231(.A(KEYINPUT29), .B1(new_n394), .B2(new_n395), .ZN(new_n433));
  AOI21_X1  g232(.A(KEYINPUT29), .B1(new_n335), .B2(new_n338), .ZN(new_n434));
  OAI211_X1 g233(.A(new_n336), .B(new_n328), .C1(new_n334), .C2(KEYINPUT22), .ZN(new_n435));
  AOI21_X1  g234(.A(KEYINPUT3), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  OAI22_X1  g235(.A1(new_n433), .A2(new_n341), .B1(new_n436), .B2(new_n385), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT85), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n437), .A2(new_n438), .A3(new_n431), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n438), .B1(new_n437), .B2(new_n431), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n432), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(G22gat), .ZN(new_n443));
  NOR3_X1   g242(.A1(new_n428), .A2(new_n430), .A3(new_n431), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n434), .A2(new_n435), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n385), .B1(new_n445), .B2(new_n391), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n431), .B1(new_n430), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(KEYINPUT85), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n444), .B1(new_n448), .B2(new_n439), .ZN(new_n449));
  INV_X1    g248(.A(G22gat), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n425), .B1(new_n443), .B2(new_n451), .ZN(new_n452));
  OAI21_X1  g251(.A(KEYINPUT86), .B1(new_n449), .B2(new_n450), .ZN(new_n453));
  INV_X1    g252(.A(new_n425), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n454), .B1(new_n449), .B2(new_n450), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT86), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n442), .A2(new_n456), .A3(G22gat), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n453), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT87), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n453), .A2(new_n455), .A3(new_n457), .A4(KEYINPUT87), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n452), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n462), .A2(KEYINPUT35), .ZN(new_n463));
  AND3_X1   g262(.A1(new_n315), .A2(new_n421), .A3(new_n463), .ZN(new_n464));
  OR3_X1    g263(.A1(new_n366), .A2(KEYINPUT89), .A3(new_n420), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n460), .A2(new_n461), .ZN(new_n466));
  INV_X1    g265(.A(new_n452), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n302), .A2(new_n310), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n468), .A2(KEYINPUT91), .A3(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT91), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n312), .A2(new_n313), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n471), .B1(new_n462), .B2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT80), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n365), .A2(new_n474), .A3(new_n361), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n415), .A2(new_n416), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n413), .B1(new_n476), .B2(new_n418), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n475), .A2(new_n477), .A3(new_n359), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n474), .B1(new_n365), .B2(new_n361), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n470), .A2(new_n473), .A3(new_n480), .ZN(new_n481));
  AOI22_X1  g280(.A1(new_n464), .A2(new_n465), .B1(new_n481), .B2(KEYINPUT35), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n388), .A2(new_n390), .A3(new_n397), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT39), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n483), .A2(new_n484), .A3(G225gat), .A4(G233gat), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n398), .B1(new_n409), .B2(new_n390), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n400), .A2(new_n398), .A3(new_n386), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(KEYINPUT39), .ZN(new_n488));
  OAI211_X1 g287(.A(new_n485), .B(new_n407), .C1(new_n486), .C2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT40), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n408), .B1(new_n486), .B2(new_n484), .ZN(new_n492));
  OAI211_X1 g291(.A(new_n492), .B(KEYINPUT40), .C1(new_n486), .C2(new_n488), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n491), .A2(new_n493), .A3(new_n415), .ZN(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n366), .A2(new_n495), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n348), .A2(new_n349), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n351), .B1(new_n497), .B2(new_n343), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n364), .B1(new_n498), .B2(new_n342), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n360), .B1(new_n499), .B2(KEYINPUT37), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT37), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n353), .A2(new_n501), .ZN(new_n502));
  OAI21_X1  g301(.A(KEYINPUT38), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n503), .A2(new_n420), .A3(new_n357), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n501), .B1(new_n497), .B2(new_n341), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n327), .A2(new_n343), .ZN(new_n506));
  AOI21_X1  g305(.A(KEYINPUT38), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  OAI211_X1 g306(.A(new_n360), .B(new_n507), .C1(new_n499), .C2(KEYINPUT37), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT88), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n360), .A2(KEYINPUT37), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n361), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n512), .A2(KEYINPUT88), .A3(new_n507), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n496), .B1(new_n504), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(new_n468), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n480), .A2(new_n462), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n312), .A2(KEYINPUT36), .A3(new_n313), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT36), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n519), .B1(new_n302), .B2(new_n310), .ZN(new_n520));
  AOI22_X1  g319(.A1(new_n516), .A2(new_n517), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n482), .A2(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(G113gat), .B(G141gat), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n523), .B(G197gat), .ZN(new_n524));
  XOR2_X1   g323(.A(KEYINPUT11), .B(G169gat), .Z(new_n525));
  XNOR2_X1  g324(.A(new_n524), .B(new_n525), .ZN(new_n526));
  XNOR2_X1  g325(.A(KEYINPUT92), .B(KEYINPUT12), .ZN(new_n527));
  XOR2_X1   g326(.A(new_n526), .B(new_n527), .Z(new_n528));
  INV_X1    g327(.A(KEYINPUT94), .ZN(new_n529));
  NAND2_X1  g328(.A1(G43gat), .A2(G50gat), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  NOR2_X1   g330(.A1(G43gat), .A2(G50gat), .ZN(new_n532));
  OAI21_X1  g331(.A(KEYINPUT15), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(G43gat), .ZN(new_n534));
  INV_X1    g333(.A(G50gat), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT15), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n536), .A2(new_n537), .A3(new_n530), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT14), .ZN(new_n539));
  INV_X1    g338(.A(G29gat), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n542));
  AOI21_X1  g341(.A(G36gat), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(G36gat), .ZN(new_n544));
  NOR3_X1   g343(.A1(new_n539), .A2(new_n544), .A3(G29gat), .ZN(new_n545));
  OAI211_X1 g344(.A(new_n533), .B(new_n538), .C1(new_n543), .C2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT93), .ZN(new_n547));
  INV_X1    g346(.A(new_n545), .ZN(new_n548));
  INV_X1    g347(.A(new_n542), .ZN(new_n549));
  NOR2_X1   g348(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n544), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  OAI22_X1  g351(.A1(new_n546), .A2(new_n547), .B1(new_n552), .B2(new_n533), .ZN(new_n553));
  AND2_X1   g352(.A1(new_n533), .A2(new_n538), .ZN(new_n554));
  AOI21_X1  g353(.A(KEYINPUT93), .B1(new_n554), .B2(new_n552), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n529), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n554), .A2(new_n552), .A3(KEYINPUT93), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n546), .A2(new_n547), .ZN(new_n558));
  OR3_X1    g357(.A1(new_n533), .A2(new_n543), .A3(new_n545), .ZN(new_n559));
  NAND4_X1  g358(.A1(new_n557), .A2(new_n558), .A3(KEYINPUT94), .A4(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n556), .A2(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(G15gat), .B(G22gat), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT16), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n562), .B1(new_n563), .B2(G1gat), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n564), .B1(G1gat), .B2(new_n562), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(G8gat), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n561), .A2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT96), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n561), .A2(new_n567), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n561), .A2(KEYINPUT96), .A3(new_n567), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n570), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(G229gat), .A2(G233gat), .ZN(new_n575));
  XOR2_X1   g374(.A(new_n575), .B(KEYINPUT13), .Z(new_n576));
  NAND2_X1  g375(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  NAND4_X1  g376(.A1(new_n557), .A2(new_n558), .A3(KEYINPUT17), .A4(new_n559), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n567), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT17), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n556), .A2(new_n580), .A3(new_n560), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(KEYINPUT95), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT95), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n556), .A2(new_n583), .A3(new_n580), .A4(new_n560), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n579), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n575), .ZN(new_n586));
  NOR3_X1   g385(.A1(new_n585), .A2(new_n586), .A3(new_n571), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n577), .B1(new_n587), .B2(KEYINPUT18), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT18), .ZN(new_n589));
  NOR4_X1   g388(.A1(new_n585), .A2(new_n589), .A3(new_n586), .A4(new_n571), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n528), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n582), .A2(new_n584), .ZN(new_n592));
  INV_X1    g391(.A(new_n579), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n594), .A2(new_n575), .A3(new_n572), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n595), .A2(new_n589), .ZN(new_n596));
  INV_X1    g395(.A(new_n528), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n571), .B1(new_n592), .B2(new_n593), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n598), .A2(KEYINPUT18), .A3(new_n575), .ZN(new_n599));
  NAND4_X1  g398(.A1(new_n596), .A2(new_n597), .A3(new_n599), .A4(new_n577), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n591), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n522), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n603), .A2(new_n420), .ZN(new_n604));
  AND2_X1   g403(.A1(G232gat), .A2(G233gat), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n605), .A2(KEYINPUT41), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(KEYINPUT100), .ZN(new_n607));
  XNOR2_X1  g406(.A(G134gat), .B(G162gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  XOR2_X1   g409(.A(G190gat), .B(G218gat), .Z(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(G85gat), .A2(G92gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(KEYINPUT7), .ZN(new_n614));
  NAND2_X1  g413(.A1(G99gat), .A2(G106gat), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n615), .A2(KEYINPUT8), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT101), .ZN(new_n617));
  OR2_X1    g416(.A1(G85gat), .A2(G92gat), .ZN(new_n618));
  AND3_X1   g417(.A1(new_n616), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n617), .B1(new_n616), .B2(new_n618), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n614), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NOR2_X1   g420(.A1(G99gat), .A2(G106gat), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n623), .A2(KEYINPUT102), .A3(new_n615), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT102), .ZN(new_n625));
  INV_X1    g424(.A(new_n615), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n625), .B1(new_n626), .B2(new_n622), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n621), .A2(new_n629), .ZN(new_n630));
  OAI211_X1 g429(.A(new_n628), .B(new_n614), .C1(new_n619), .C2(new_n620), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n630), .A2(KEYINPUT103), .A3(new_n631), .ZN(new_n632));
  OR2_X1    g431(.A1(new_n619), .A2(new_n620), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT103), .ZN(new_n634));
  NAND4_X1  g433(.A1(new_n633), .A2(new_n634), .A3(new_n628), .A4(new_n614), .ZN(new_n635));
  AND2_X1   g434(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n636), .A2(new_n578), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n592), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n605), .A2(KEYINPUT41), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n640), .B1(new_n636), .B2(new_n561), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n612), .B1(new_n639), .B2(new_n642), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n637), .B1(new_n582), .B2(new_n584), .ZN(new_n644));
  NOR3_X1   g443(.A1(new_n644), .A2(new_n641), .A3(new_n611), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n610), .B1(new_n643), .B2(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n639), .A2(new_n612), .A3(new_n642), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n611), .B1(new_n644), .B2(new_n641), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n647), .A2(new_n609), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  XOR2_X1   g450(.A(G57gat), .B(G64gat), .Z(new_n652));
  NAND2_X1  g451(.A1(G71gat), .A2(G78gat), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT9), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g454(.A1(G71gat), .A2(G78gat), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  AND2_X1   g456(.A1(new_n657), .A2(new_n653), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT97), .ZN(new_n659));
  OAI211_X1 g458(.A(new_n652), .B(new_n655), .C1(new_n658), .C2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n652), .A2(new_n655), .ZN(new_n661));
  AOI22_X1  g460(.A1(new_n653), .A2(new_n657), .B1(new_n655), .B2(new_n659), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n664), .A2(KEYINPUT21), .ZN(new_n665));
  XOR2_X1   g464(.A(G127gat), .B(G155gat), .Z(new_n666));
  XNOR2_X1  g465(.A(new_n665), .B(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT99), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n664), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n660), .A2(new_n663), .A3(KEYINPUT99), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n566), .B1(new_n671), .B2(KEYINPUT21), .ZN(new_n672));
  XOR2_X1   g471(.A(new_n667), .B(new_n672), .Z(new_n673));
  NAND2_X1  g472(.A1(G231gat), .A2(G233gat), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(KEYINPUT98), .ZN(new_n675));
  XOR2_X1   g474(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n676));
  XNOR2_X1  g475(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g476(.A(G183gat), .B(G211gat), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n673), .B(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n664), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n632), .A2(new_n682), .A3(new_n635), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n664), .A2(new_n630), .A3(new_n631), .ZN(new_n684));
  XNOR2_X1  g483(.A(KEYINPUT104), .B(KEYINPUT10), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n683), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n632), .A2(new_n635), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n687), .A2(new_n671), .A3(KEYINPUT10), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(G230gat), .A2(G233gat), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g490(.A(G120gat), .B(G148gat), .ZN(new_n692));
  XNOR2_X1  g491(.A(G176gat), .B(G204gat), .ZN(new_n693));
  XOR2_X1   g492(.A(new_n692), .B(new_n693), .Z(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n683), .A2(new_n684), .ZN(new_n696));
  INV_X1    g495(.A(new_n690), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n695), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n691), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  XOR2_X1   g499(.A(new_n690), .B(KEYINPUT105), .Z(new_n701));
  INV_X1    g500(.A(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n689), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n696), .A2(new_n697), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n700), .B1(new_n705), .B2(new_n695), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n651), .A2(new_n681), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(KEYINPUT106), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n650), .A2(new_n680), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT106), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n709), .A2(new_n710), .A3(new_n706), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n708), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n604), .A2(new_n712), .ZN(new_n713));
  XOR2_X1   g512(.A(new_n713), .B(G1gat), .Z(G1324gat));
  NAND2_X1  g513(.A1(new_n603), .A2(new_n366), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n715), .A2(new_n712), .ZN(new_n716));
  XNOR2_X1  g515(.A(KEYINPUT16), .B(G8gat), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT107), .ZN(new_n718));
  AOI21_X1  g517(.A(KEYINPUT42), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n719), .B1(new_n718), .B2(new_n717), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n716), .A2(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT42), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n721), .B1(new_n722), .B2(G8gat), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n717), .A2(new_n722), .ZN(new_n724));
  AOI21_X1  g523(.A(KEYINPUT108), .B1(new_n716), .B2(new_n724), .ZN(new_n725));
  AND3_X1   g524(.A1(new_n716), .A2(KEYINPUT108), .A3(new_n724), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n723), .B1(new_n725), .B2(new_n726), .ZN(G1325gat));
  INV_X1    g526(.A(new_n603), .ZN(new_n728));
  INV_X1    g527(.A(new_n315), .ZN(new_n729));
  OR4_X1    g528(.A1(G15gat), .A2(new_n728), .A3(new_n712), .A4(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(G15gat), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT109), .ZN(new_n732));
  AND3_X1   g531(.A1(new_n312), .A2(KEYINPUT36), .A3(new_n313), .ZN(new_n733));
  AOI21_X1  g532(.A(KEYINPUT36), .B1(new_n312), .B2(new_n313), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n732), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n520), .A2(KEYINPUT109), .A3(new_n518), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(new_n737), .ZN(new_n738));
  NOR3_X1   g537(.A1(new_n728), .A2(new_n712), .A3(new_n738), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n730), .B1(new_n731), .B2(new_n739), .ZN(G1326gat));
  OAI211_X1 g539(.A(new_n462), .B(new_n601), .C1(new_n482), .C2(new_n521), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n741), .A2(new_n712), .ZN(new_n742));
  XOR2_X1   g541(.A(KEYINPUT43), .B(G22gat), .Z(new_n743));
  XNOR2_X1  g542(.A(new_n742), .B(new_n743), .ZN(G1327gat));
  INV_X1    g543(.A(KEYINPUT45), .ZN(new_n745));
  INV_X1    g544(.A(new_n706), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n681), .A2(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n748), .A2(new_n651), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(new_n540), .ZN(new_n750));
  OR3_X1    g549(.A1(new_n604), .A2(new_n745), .A3(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT44), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n651), .A2(new_n752), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n753), .B1(new_n482), .B2(new_n521), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n748), .A2(new_n602), .ZN(new_n755));
  AND2_X1   g554(.A1(new_n365), .A2(new_n361), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n494), .B1(new_n756), .B2(new_n359), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT38), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n499), .A2(KEYINPUT37), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n758), .B1(new_n512), .B2(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(new_n357), .ZN(new_n761));
  NOR3_X1   g560(.A1(new_n760), .A2(new_n477), .A3(new_n761), .ZN(new_n762));
  AND2_X1   g561(.A1(new_n510), .A2(new_n513), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n757), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n517), .B1(new_n764), .B2(new_n462), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(new_n738), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n481), .A2(KEYINPUT35), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n465), .A2(new_n315), .A3(new_n421), .A4(new_n463), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n651), .B1(new_n766), .B2(new_n769), .ZN(new_n770));
  OAI211_X1 g569(.A(new_n754), .B(new_n755), .C1(new_n770), .C2(KEYINPUT44), .ZN(new_n771));
  OAI21_X1  g570(.A(G29gat), .B1(new_n771), .B2(new_n477), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n745), .B1(new_n604), .B2(new_n750), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n751), .A2(new_n772), .A3(new_n773), .ZN(G1328gat));
  NAND2_X1  g573(.A1(new_n749), .A2(new_n544), .ZN(new_n775));
  OR3_X1    g574(.A1(new_n715), .A2(KEYINPUT46), .A3(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(new_n366), .ZN(new_n777));
  OAI21_X1  g576(.A(G36gat), .B1(new_n771), .B2(new_n777), .ZN(new_n778));
  OAI21_X1  g577(.A(KEYINPUT46), .B1(new_n715), .B2(new_n775), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n776), .A2(new_n778), .A3(new_n779), .ZN(G1329gat));
  OAI21_X1  g579(.A(G43gat), .B1(new_n771), .B2(new_n738), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n749), .A2(new_n534), .ZN(new_n782));
  NOR4_X1   g581(.A1(new_n522), .A2(new_n729), .A3(new_n602), .A4(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n781), .A2(new_n784), .ZN(new_n785));
  AOI21_X1  g584(.A(KEYINPUT47), .B1(new_n785), .B2(KEYINPUT110), .ZN(new_n786));
  AOI22_X1  g585(.A1(new_n765), .A2(new_n738), .B1(new_n767), .B2(new_n768), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n752), .B1(new_n787), .B2(new_n651), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n788), .A2(new_n737), .A3(new_n754), .A4(new_n755), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n783), .B1(new_n789), .B2(G43gat), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT110), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT47), .ZN(new_n792));
  NOR3_X1   g591(.A1(new_n790), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n786), .A2(new_n793), .ZN(G1330gat));
  NAND2_X1  g593(.A1(new_n749), .A2(new_n535), .ZN(new_n795));
  OAI21_X1  g594(.A(KEYINPUT111), .B1(new_n741), .B2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT48), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(KEYINPUT112), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT112), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n796), .A2(new_n800), .A3(new_n797), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n741), .A2(new_n795), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n788), .A2(new_n462), .A3(new_n754), .A4(new_n755), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n803), .B1(new_n804), .B2(G50gat), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n802), .A2(new_n805), .ZN(new_n806));
  AND2_X1   g605(.A1(new_n804), .A2(G50gat), .ZN(new_n807));
  OAI211_X1 g606(.A(new_n799), .B(new_n801), .C1(new_n807), .C2(new_n803), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n806), .A2(new_n808), .ZN(G1331gat));
  NAND3_X1  g608(.A1(new_n602), .A2(new_n709), .A3(new_n746), .ZN(new_n810));
  OAI21_X1  g609(.A(KEYINPUT113), .B1(new_n787), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n766), .A2(new_n769), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT113), .ZN(new_n813));
  INV_X1    g612(.A(new_n810), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n812), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n811), .A2(new_n815), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n816), .A2(new_n477), .ZN(new_n817));
  XOR2_X1   g616(.A(new_n817), .B(G57gat), .Z(G1332gat));
  NAND3_X1  g617(.A1(new_n811), .A2(new_n815), .A3(new_n366), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n819), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n820));
  XOR2_X1   g619(.A(KEYINPUT49), .B(G64gat), .Z(new_n821));
  OAI21_X1  g620(.A(new_n820), .B1(new_n819), .B2(new_n821), .ZN(G1333gat));
  OAI21_X1  g621(.A(G71gat), .B1(new_n816), .B2(new_n738), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n729), .A2(G71gat), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n811), .A2(new_n815), .A3(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT50), .ZN(new_n827));
  XNOR2_X1  g626(.A(new_n826), .B(new_n827), .ZN(G1334gat));
  OAI21_X1  g627(.A(KEYINPUT115), .B1(new_n816), .B2(new_n468), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT115), .ZN(new_n830));
  NAND4_X1  g629(.A1(new_n811), .A2(new_n815), .A3(new_n830), .A4(new_n462), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  XNOR2_X1  g631(.A(KEYINPUT114), .B(G78gat), .ZN(new_n833));
  XNOR2_X1  g632(.A(new_n832), .B(new_n833), .ZN(G1335gat));
  NOR3_X1   g633(.A1(new_n601), .A2(new_n681), .A3(new_n706), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n788), .A2(new_n754), .A3(new_n835), .ZN(new_n836));
  OAI21_X1  g635(.A(G85gat), .B1(new_n836), .B2(new_n477), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n601), .A2(new_n681), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n737), .B1(new_n516), .B2(new_n517), .ZN(new_n839));
  OAI211_X1 g638(.A(new_n650), .B(new_n838), .C1(new_n482), .C2(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT51), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT116), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n812), .A2(KEYINPUT51), .A3(new_n650), .A4(new_n838), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n842), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n840), .A2(KEYINPUT116), .A3(new_n841), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  OR3_X1    g646(.A1(new_n477), .A2(G85gat), .A3(new_n706), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n837), .B1(new_n847), .B2(new_n848), .ZN(G1336gat));
  NOR3_X1   g648(.A1(new_n777), .A2(G92gat), .A3(new_n706), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n845), .A2(new_n846), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(KEYINPUT117), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT117), .ZN(new_n853));
  NAND4_X1  g652(.A1(new_n845), .A2(new_n846), .A3(new_n853), .A4(new_n850), .ZN(new_n854));
  XNOR2_X1  g653(.A(KEYINPUT118), .B(KEYINPUT52), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n788), .A2(new_n366), .A3(new_n754), .A4(new_n835), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n855), .B1(new_n856), .B2(G92gat), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n852), .A2(new_n854), .A3(new_n857), .ZN(new_n858));
  AND2_X1   g657(.A1(new_n856), .A2(G92gat), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n842), .A2(new_n844), .ZN(new_n860));
  AND2_X1   g659(.A1(new_n860), .A2(new_n850), .ZN(new_n861));
  OAI21_X1  g660(.A(KEYINPUT52), .B1(new_n859), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n858), .A2(new_n862), .ZN(G1337gat));
  OAI21_X1  g662(.A(G99gat), .B1(new_n836), .B2(new_n738), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n729), .A2(new_n706), .ZN(new_n865));
  INV_X1    g664(.A(new_n865), .ZN(new_n866));
  OR2_X1    g665(.A1(new_n866), .A2(G99gat), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n864), .B1(new_n847), .B2(new_n867), .ZN(G1338gat));
  NAND4_X1  g667(.A1(new_n788), .A2(new_n462), .A3(new_n754), .A4(new_n835), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(G106gat), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT53), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NOR3_X1   g671(.A1(new_n468), .A2(G106gat), .A3(new_n706), .ZN(new_n873));
  AND3_X1   g672(.A1(new_n845), .A2(new_n846), .A3(new_n873), .ZN(new_n874));
  AOI22_X1  g673(.A1(G106gat), .A2(new_n869), .B1(new_n860), .B2(new_n873), .ZN(new_n875));
  OAI22_X1  g674(.A1(new_n872), .A2(new_n874), .B1(new_n875), .B2(new_n871), .ZN(G1339gat));
  NOR2_X1   g675(.A1(new_n707), .A2(new_n601), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT120), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n695), .B1(new_n703), .B2(KEYINPUT54), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n686), .A2(new_n701), .A3(new_n688), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n691), .A2(KEYINPUT54), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(KEYINPUT119), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT54), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n883), .B1(new_n689), .B2(new_n690), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT119), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n884), .A2(new_n885), .A3(new_n880), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n879), .B1(new_n882), .B2(new_n886), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n878), .B1(new_n887), .B2(KEYINPUT55), .ZN(new_n888));
  INV_X1    g687(.A(new_n879), .ZN(new_n889));
  AND3_X1   g688(.A1(new_n884), .A2(new_n885), .A3(new_n880), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n885), .B1(new_n884), .B2(new_n880), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n889), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT55), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n892), .A2(KEYINPUT120), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n888), .A2(new_n894), .ZN(new_n895));
  OAI22_X1  g694(.A1(new_n598), .A2(new_n575), .B1(new_n574), .B2(new_n576), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(new_n526), .ZN(new_n897));
  AND3_X1   g696(.A1(new_n650), .A2(new_n600), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n700), .B1(new_n887), .B2(KEYINPUT55), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n895), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n895), .A2(new_n601), .A3(new_n899), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n600), .A2(new_n897), .A3(new_n746), .ZN(new_n902));
  AND2_X1   g701(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n900), .B1(new_n903), .B2(new_n650), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n877), .B1(new_n904), .B2(new_n680), .ZN(new_n905));
  INV_X1    g704(.A(new_n905), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n366), .A2(new_n477), .ZN(new_n907));
  NAND4_X1  g706(.A1(new_n906), .A2(new_n468), .A3(new_n315), .A4(new_n907), .ZN(new_n908));
  NOR3_X1   g707(.A1(new_n908), .A2(new_n255), .A3(new_n602), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n905), .A2(new_n477), .ZN(new_n910));
  AND2_X1   g709(.A1(new_n470), .A2(new_n473), .ZN(new_n911));
  AND2_X1   g710(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  AND2_X1   g711(.A1(new_n912), .A2(new_n777), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(new_n601), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n909), .B1(new_n914), .B2(new_n255), .ZN(G1340gat));
  NOR3_X1   g714(.A1(new_n908), .A2(new_n252), .A3(new_n706), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n913), .A2(new_n746), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n916), .B1(new_n917), .B2(new_n252), .ZN(G1341gat));
  INV_X1    g717(.A(G127gat), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n913), .A2(new_n919), .A3(new_n681), .ZN(new_n920));
  OAI21_X1  g719(.A(G127gat), .B1(new_n908), .B2(new_n680), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(G1342gat));
  NAND2_X1  g721(.A1(new_n777), .A2(new_n650), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n923), .A2(G134gat), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n912), .A2(new_n924), .ZN(new_n925));
  OR2_X1    g724(.A1(new_n925), .A2(KEYINPUT56), .ZN(new_n926));
  OAI21_X1  g725(.A(G134gat), .B1(new_n908), .B2(new_n651), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n925), .A2(KEYINPUT56), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n926), .A2(new_n927), .A3(new_n928), .ZN(G1343gat));
  NAND2_X1  g728(.A1(new_n738), .A2(new_n907), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT57), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n931), .B1(new_n905), .B2(new_n468), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n468), .A2(new_n931), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n892), .A2(new_n893), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n601), .A2(new_n899), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(new_n902), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n936), .A2(new_n651), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n681), .B1(new_n937), .B2(new_n900), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n933), .B1(new_n938), .B2(new_n877), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n930), .B1(new_n932), .B2(new_n939), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n374), .B1(new_n940), .B2(new_n601), .ZN(new_n941));
  INV_X1    g740(.A(new_n941), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n737), .A2(new_n468), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n602), .A2(G141gat), .ZN(new_n944));
  NAND4_X1  g743(.A1(new_n910), .A2(new_n777), .A3(new_n943), .A4(new_n944), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT121), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n947), .A2(KEYINPUT58), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n942), .A2(new_n945), .A3(new_n948), .ZN(new_n949));
  INV_X1    g748(.A(new_n945), .ZN(new_n950));
  OAI211_X1 g749(.A(KEYINPUT58), .B(new_n947), .C1(new_n941), .C2(new_n950), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n949), .A2(new_n951), .ZN(G1344gat));
  NOR2_X1   g751(.A1(new_n930), .A2(new_n706), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n937), .A2(KEYINPUT123), .A3(new_n900), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT123), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n650), .B1(new_n935), .B2(new_n902), .ZN(new_n956));
  AND3_X1   g755(.A1(new_n895), .A2(new_n898), .A3(new_n899), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n955), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n954), .A2(new_n958), .A3(new_n680), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n708), .A2(new_n711), .A3(new_n602), .ZN(new_n960));
  XNOR2_X1  g759(.A(new_n960), .B(KEYINPUT122), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  AOI21_X1  g761(.A(KEYINPUT57), .B1(new_n962), .B2(new_n462), .ZN(new_n963));
  INV_X1    g762(.A(new_n933), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n905), .A2(new_n964), .ZN(new_n965));
  OAI211_X1 g764(.A(KEYINPUT124), .B(new_n953), .C1(new_n963), .C2(new_n965), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n966), .A2(G148gat), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n468), .B1(new_n959), .B2(new_n961), .ZN(new_n968));
  OAI22_X1  g767(.A1(new_n968), .A2(KEYINPUT57), .B1(new_n905), .B2(new_n964), .ZN(new_n969));
  AOI21_X1  g768(.A(KEYINPUT124), .B1(new_n969), .B2(new_n953), .ZN(new_n970));
  OAI21_X1  g769(.A(KEYINPUT59), .B1(new_n967), .B2(new_n970), .ZN(new_n971));
  NOR2_X1   g770(.A1(new_n376), .A2(KEYINPUT59), .ZN(new_n972));
  INV_X1    g771(.A(new_n940), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n972), .B1(new_n973), .B2(new_n706), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n971), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n910), .A2(new_n943), .ZN(new_n976));
  NOR2_X1   g775(.A1(new_n976), .A2(new_n366), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n977), .A2(new_n376), .A3(new_n746), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n975), .A2(new_n978), .ZN(G1345gat));
  OAI21_X1  g778(.A(G155gat), .B1(new_n973), .B2(new_n680), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n977), .A2(new_n380), .A3(new_n681), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n980), .A2(new_n981), .ZN(G1346gat));
  AOI21_X1  g781(.A(new_n381), .B1(new_n940), .B2(new_n650), .ZN(new_n983));
  NOR3_X1   g782(.A1(new_n976), .A2(G162gat), .A3(new_n923), .ZN(new_n984));
  OR3_X1    g783(.A1(new_n983), .A2(KEYINPUT125), .A3(new_n984), .ZN(new_n985));
  OAI21_X1  g784(.A(KEYINPUT125), .B1(new_n983), .B2(new_n984), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n985), .A2(new_n986), .ZN(G1347gat));
  NOR3_X1   g786(.A1(new_n905), .A2(new_n420), .A3(new_n777), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n988), .A2(new_n911), .ZN(new_n989));
  INV_X1    g788(.A(new_n989), .ZN(new_n990));
  NAND3_X1  g789(.A1(new_n990), .A2(new_n208), .A3(new_n601), .ZN(new_n991));
  INV_X1    g790(.A(KEYINPUT126), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n315), .A2(new_n468), .ZN(new_n993));
  NOR4_X1   g792(.A1(new_n905), .A2(new_n420), .A3(new_n777), .A4(new_n993), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n994), .A2(new_n601), .ZN(new_n995));
  AOI21_X1  g794(.A(new_n992), .B1(new_n995), .B2(G169gat), .ZN(new_n996));
  AOI211_X1 g795(.A(KEYINPUT126), .B(new_n208), .C1(new_n994), .C2(new_n601), .ZN(new_n997));
  OAI21_X1  g796(.A(new_n991), .B1(new_n996), .B2(new_n997), .ZN(G1348gat));
  AOI21_X1  g797(.A(G176gat), .B1(new_n990), .B2(new_n746), .ZN(new_n999));
  NOR3_X1   g798(.A1(new_n866), .A2(new_n209), .A3(new_n462), .ZN(new_n1000));
  AOI21_X1  g799(.A(new_n999), .B1(new_n988), .B2(new_n1000), .ZN(G1349gat));
  OR3_X1    g800(.A1(new_n680), .A2(new_n232), .A3(new_n234), .ZN(new_n1002));
  NOR2_X1   g801(.A1(new_n989), .A2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g802(.A(new_n213), .B1(new_n994), .B2(new_n681), .ZN(new_n1004));
  NOR2_X1   g803(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g804(.A(KEYINPUT60), .ZN(new_n1006));
  XNOR2_X1  g805(.A(new_n1005), .B(new_n1006), .ZN(G1350gat));
  NAND3_X1  g806(.A1(new_n990), .A2(new_n214), .A3(new_n650), .ZN(new_n1008));
  INV_X1    g807(.A(KEYINPUT61), .ZN(new_n1009));
  NAND2_X1  g808(.A1(new_n994), .A2(new_n650), .ZN(new_n1010));
  AOI21_X1  g809(.A(new_n1009), .B1(new_n1010), .B2(G190gat), .ZN(new_n1011));
  AOI211_X1 g810(.A(KEYINPUT61), .B(new_n214), .C1(new_n994), .C2(new_n650), .ZN(new_n1012));
  OAI21_X1  g811(.A(new_n1008), .B1(new_n1011), .B2(new_n1012), .ZN(G1351gat));
  NOR3_X1   g812(.A1(new_n737), .A2(new_n420), .A3(new_n777), .ZN(new_n1014));
  INV_X1    g813(.A(new_n1014), .ZN(new_n1015));
  NOR3_X1   g814(.A1(new_n905), .A2(new_n1015), .A3(new_n468), .ZN(new_n1016));
  AOI21_X1  g815(.A(G197gat), .B1(new_n1016), .B2(new_n601), .ZN(new_n1017));
  AND2_X1   g816(.A1(new_n969), .A2(new_n1014), .ZN(new_n1018));
  AND2_X1   g817(.A1(new_n601), .A2(G197gat), .ZN(new_n1019));
  AOI21_X1  g818(.A(new_n1017), .B1(new_n1018), .B2(new_n1019), .ZN(G1352gat));
  NAND2_X1  g819(.A1(new_n1018), .A2(new_n746), .ZN(new_n1021));
  NAND2_X1  g820(.A1(new_n1021), .A2(G204gat), .ZN(new_n1022));
  INV_X1    g821(.A(KEYINPUT127), .ZN(new_n1023));
  NOR2_X1   g822(.A1(new_n706), .A2(G204gat), .ZN(new_n1024));
  AND3_X1   g823(.A1(new_n1016), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  AOI21_X1  g824(.A(new_n1023), .B1(new_n1016), .B2(new_n1024), .ZN(new_n1026));
  INV_X1    g825(.A(KEYINPUT62), .ZN(new_n1027));
  OR3_X1    g826(.A1(new_n1025), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  OAI21_X1  g827(.A(new_n1027), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1029));
  NAND3_X1  g828(.A1(new_n1022), .A2(new_n1028), .A3(new_n1029), .ZN(G1353gat));
  NAND3_X1  g829(.A1(new_n1016), .A2(new_n329), .A3(new_n681), .ZN(new_n1031));
  NAND3_X1  g830(.A1(new_n969), .A2(new_n681), .A3(new_n1014), .ZN(new_n1032));
  AND3_X1   g831(.A1(new_n1032), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1033));
  AOI21_X1  g832(.A(KEYINPUT63), .B1(new_n1032), .B2(G211gat), .ZN(new_n1034));
  OAI21_X1  g833(.A(new_n1031), .B1(new_n1033), .B2(new_n1034), .ZN(G1354gat));
  AOI21_X1  g834(.A(G218gat), .B1(new_n1016), .B2(new_n650), .ZN(new_n1036));
  AOI21_X1  g835(.A(new_n651), .B1(new_n331), .B2(new_n333), .ZN(new_n1037));
  AOI21_X1  g836(.A(new_n1036), .B1(new_n1018), .B2(new_n1037), .ZN(G1355gat));
endmodule


