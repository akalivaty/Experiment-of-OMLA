//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 0 1 1 0 1 0 0 0 1 1 1 1 1 1 0 1 0 0 1 1 1 1 1 0 0 0 0 1 1 0 1 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 0 0 0 1 0 1 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n755, new_n756, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n784, new_n785, new_n786, new_n787,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n815, new_n816, new_n817, new_n818, new_n820, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n901, new_n902, new_n903, new_n905,
    new_n906, new_n907, new_n908, new_n910, new_n911, new_n912, new_n913,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n967, new_n968, new_n969, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n982,
    new_n983, new_n985, new_n986, new_n987, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1021, new_n1022, new_n1023, new_n1024, new_n1026,
    new_n1027, new_n1028;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(G1gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(KEYINPUT16), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G8gat), .ZN(new_n206));
  OAI211_X1 g005(.A(new_n205), .B(new_n206), .C1(G1gat), .C2(new_n202), .ZN(new_n207));
  INV_X1    g006(.A(G15gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(G22gat), .ZN(new_n209));
  INV_X1    g008(.A(G22gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(G15gat), .ZN(new_n211));
  AND3_X1   g010(.A1(new_n204), .A2(new_n209), .A3(new_n211), .ZN(new_n212));
  AOI21_X1  g011(.A(G1gat), .B1(new_n209), .B2(new_n211), .ZN(new_n213));
  OAI21_X1  g012(.A(G8gat), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n207), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(G43gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(G50gat), .ZN(new_n217));
  INV_X1    g016(.A(G50gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(G43gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n217), .A2(new_n219), .A3(KEYINPUT15), .ZN(new_n220));
  AND2_X1   g019(.A1(G29gat), .A2(G36gat), .ZN(new_n221));
  NOR2_X1   g020(.A1(G29gat), .A2(G36gat), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n221), .B1(KEYINPUT14), .B2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT14), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n224), .B1(G29gat), .B2(G36gat), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n220), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(new_n220), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n222), .A2(KEYINPUT14), .ZN(new_n228));
  NAND2_X1  g027(.A1(G29gat), .A2(G36gat), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n228), .A2(new_n225), .A3(new_n229), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n227), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT84), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n232), .B1(new_n216), .B2(G50gat), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n218), .A2(KEYINPUT84), .A3(G43gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n233), .A2(new_n217), .A3(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT15), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n226), .B1(new_n231), .B2(new_n237), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n215), .B1(new_n238), .B2(KEYINPUT17), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT85), .ZN(new_n240));
  AND3_X1   g039(.A1(new_n228), .A2(new_n225), .A3(new_n229), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n237), .A2(new_n220), .A3(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n227), .A2(new_n230), .ZN(new_n243));
  AOI211_X1 g042(.A(new_n240), .B(KEYINPUT17), .C1(new_n242), .C2(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(KEYINPUT84), .B1(new_n218), .B2(G43gat), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n218), .A2(G43gat), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  AOI21_X1  g046(.A(KEYINPUT15), .B1(new_n247), .B2(new_n234), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n223), .A2(new_n220), .A3(new_n225), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n243), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT17), .ZN(new_n251));
  AOI21_X1  g050(.A(KEYINPUT85), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n239), .B1(new_n244), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(KEYINPUT86), .ZN(new_n254));
  NAND2_X1  g053(.A1(G229gat), .A2(G233gat), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n250), .A2(new_n215), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT86), .ZN(new_n257));
  OAI211_X1 g056(.A(new_n257), .B(new_n239), .C1(new_n244), .C2(new_n252), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n254), .A2(new_n255), .A3(new_n256), .A4(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT18), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  AND2_X1   g060(.A1(new_n258), .A2(new_n256), .ZN(new_n262));
  NAND4_X1  g061(.A1(new_n262), .A2(KEYINPUT18), .A3(new_n255), .A4(new_n254), .ZN(new_n263));
  OAI21_X1  g062(.A(KEYINPUT87), .B1(new_n250), .B2(new_n215), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n264), .B(new_n256), .ZN(new_n265));
  XOR2_X1   g064(.A(new_n255), .B(KEYINPUT13), .Z(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n261), .A2(new_n263), .A3(new_n267), .ZN(new_n268));
  XNOR2_X1  g067(.A(G113gat), .B(G141gat), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n269), .B(G197gat), .ZN(new_n270));
  XOR2_X1   g069(.A(KEYINPUT11), .B(G169gat), .Z(new_n271));
  XNOR2_X1  g070(.A(new_n270), .B(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(new_n272), .B(KEYINPUT12), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n268), .A2(new_n274), .ZN(new_n275));
  NAND4_X1  g074(.A1(new_n261), .A2(new_n263), .A3(new_n273), .A4(new_n267), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n275), .A2(KEYINPUT88), .A3(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT88), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n268), .A2(new_n278), .A3(new_n274), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(G190gat), .B(G218gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n282), .B(KEYINPUT96), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT97), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  OAI211_X1 g084(.A(KEYINPUT17), .B(new_n243), .C1(new_n248), .C2(new_n249), .ZN(new_n286));
  NOR2_X1   g085(.A1(KEYINPUT7), .A2(G85gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(KEYINPUT7), .A2(G85gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(G92gat), .ZN(new_n289));
  INV_X1    g088(.A(G92gat), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n290), .A2(KEYINPUT7), .A3(G85gat), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n287), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  XOR2_X1   g091(.A(G99gat), .B(G106gat), .Z(new_n293));
  NAND2_X1  g092(.A1(G99gat), .A2(G106gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(KEYINPUT94), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT94), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n296), .A2(G99gat), .A3(G106gat), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n295), .A2(new_n297), .A3(KEYINPUT8), .ZN(new_n298));
  AND3_X1   g097(.A1(new_n292), .A2(new_n293), .A3(new_n298), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n293), .B1(new_n292), .B2(new_n298), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  AND2_X1   g100(.A1(new_n286), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT95), .ZN(new_n303));
  OAI211_X1 g102(.A(new_n302), .B(new_n303), .C1(new_n244), .C2(new_n252), .ZN(new_n304));
  AND2_X1   g103(.A1(G232gat), .A2(G233gat), .ZN(new_n305));
  AND2_X1   g104(.A1(new_n305), .A2(KEYINPUT41), .ZN(new_n306));
  AND2_X1   g105(.A1(new_n283), .A2(new_n284), .ZN(new_n307));
  INV_X1    g106(.A(new_n301), .ZN(new_n308));
  AOI211_X1 g107(.A(new_n306), .B(new_n307), .C1(new_n308), .C2(new_n250), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n304), .A2(new_n309), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n240), .B1(new_n238), .B2(KEYINPUT17), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n250), .A2(KEYINPUT85), .A3(new_n251), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n303), .B1(new_n313), .B2(new_n302), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n285), .B1(new_n310), .B2(new_n314), .ZN(new_n315));
  XOR2_X1   g114(.A(G134gat), .B(G162gat), .Z(new_n316));
  NOR2_X1   g115(.A1(new_n305), .A2(KEYINPUT41), .ZN(new_n317));
  XNOR2_X1  g116(.A(new_n316), .B(new_n317), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n318), .A2(KEYINPUT98), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n302), .B1(new_n244), .B2(new_n252), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(KEYINPUT95), .ZN(new_n321));
  INV_X1    g120(.A(new_n285), .ZN(new_n322));
  NAND4_X1  g121(.A1(new_n321), .A2(new_n322), .A3(new_n304), .A4(new_n309), .ZN(new_n323));
  AND3_X1   g122(.A1(new_n315), .A2(new_n319), .A3(new_n323), .ZN(new_n324));
  XNOR2_X1  g123(.A(new_n318), .B(KEYINPUT98), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n325), .B1(new_n315), .B2(new_n323), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(G71gat), .A2(G78gat), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT9), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n328), .A2(KEYINPUT90), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(G57gat), .A2(G64gat), .ZN(new_n331));
  NOR2_X1   g130(.A1(G57gat), .A2(G64gat), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  AND3_X1   g132(.A1(new_n330), .A2(new_n331), .A3(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT91), .ZN(new_n335));
  XNOR2_X1  g134(.A(G71gat), .B(G78gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n328), .A2(new_n329), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT90), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND4_X1  g138(.A1(new_n334), .A2(new_n335), .A3(new_n336), .A4(new_n339), .ZN(new_n340));
  AND2_X1   g139(.A1(G57gat), .A2(G64gat), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n341), .A2(new_n332), .ZN(new_n342));
  NAND4_X1  g141(.A1(new_n339), .A2(new_n342), .A3(new_n336), .A4(new_n330), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(KEYINPUT91), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n340), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n334), .A2(new_n339), .ZN(new_n346));
  OR3_X1    g145(.A1(KEYINPUT89), .A2(G71gat), .A3(G78gat), .ZN(new_n347));
  OAI21_X1  g146(.A(KEYINPUT89), .B1(G71gat), .B2(G78gat), .ZN(new_n348));
  AOI22_X1  g147(.A1(new_n347), .A2(new_n348), .B1(G71gat), .B2(G78gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n346), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n345), .A2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT21), .ZN(new_n352));
  OAI211_X1 g151(.A(new_n214), .B(new_n207), .C1(new_n351), .C2(new_n352), .ZN(new_n353));
  XOR2_X1   g152(.A(G127gat), .B(G155gat), .Z(new_n354));
  XNOR2_X1  g153(.A(new_n354), .B(KEYINPUT93), .ZN(new_n355));
  XNOR2_X1  g154(.A(new_n353), .B(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(G231gat), .A2(G233gat), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n351), .A2(new_n352), .A3(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n358), .ZN(new_n360));
  AOI22_X1  g159(.A1(new_n340), .A2(new_n344), .B1(new_n346), .B2(new_n349), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n360), .B1(new_n361), .B2(KEYINPUT21), .ZN(new_n362));
  XNOR2_X1  g161(.A(KEYINPUT92), .B(KEYINPUT19), .ZN(new_n363));
  XNOR2_X1  g162(.A(new_n363), .B(KEYINPUT20), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  AND3_X1   g164(.A1(new_n359), .A2(new_n362), .A3(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n365), .B1(new_n359), .B2(new_n362), .ZN(new_n367));
  XOR2_X1   g166(.A(G183gat), .B(G211gat), .Z(new_n368));
  NOR3_X1   g167(.A1(new_n366), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n368), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n359), .A2(new_n362), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(new_n364), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n359), .A2(new_n362), .A3(new_n365), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n370), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n357), .B1(new_n369), .B2(new_n374), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n368), .B1(new_n366), .B2(new_n367), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n372), .A2(new_n370), .A3(new_n373), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n376), .A2(new_n377), .A3(new_n356), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n375), .A2(new_n378), .ZN(new_n379));
  OAI21_X1  g178(.A(KEYINPUT99), .B1(new_n327), .B2(new_n379), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n315), .A2(new_n319), .A3(new_n323), .ZN(new_n381));
  AND2_X1   g180(.A1(new_n315), .A2(new_n323), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n381), .B1(new_n382), .B2(new_n325), .ZN(new_n383));
  AND3_X1   g182(.A1(new_n376), .A2(new_n377), .A3(new_n356), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n356), .B1(new_n376), .B2(new_n377), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT99), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n383), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(G230gat), .A2(G233gat), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n351), .A2(new_n308), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n292), .A2(new_n298), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(KEYINPUT100), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(new_n293), .ZN(new_n393));
  INV_X1    g192(.A(new_n293), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n391), .A2(KEYINPUT100), .A3(new_n394), .ZN(new_n395));
  NAND4_X1  g194(.A1(new_n345), .A2(new_n393), .A3(new_n350), .A4(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(KEYINPUT10), .B1(new_n390), .B2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT10), .ZN(new_n398));
  NOR3_X1   g197(.A1(new_n351), .A2(new_n398), .A3(new_n301), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n389), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  XOR2_X1   g199(.A(G120gat), .B(G148gat), .Z(new_n401));
  XNOR2_X1  g200(.A(G176gat), .B(G204gat), .ZN(new_n402));
  XNOR2_X1  g201(.A(new_n401), .B(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n390), .A2(new_n396), .ZN(new_n404));
  OR2_X1    g203(.A1(new_n404), .A2(new_n389), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n400), .A2(new_n403), .A3(new_n405), .ZN(new_n406));
  XOR2_X1   g205(.A(new_n403), .B(KEYINPUT101), .Z(new_n407));
  XOR2_X1   g206(.A(new_n389), .B(KEYINPUT102), .Z(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n409), .B1(new_n397), .B2(new_n399), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n407), .B1(new_n410), .B2(new_n405), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n411), .A2(KEYINPUT103), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT103), .ZN(new_n413));
  AOI211_X1 g212(.A(new_n413), .B(new_n407), .C1(new_n410), .C2(new_n405), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n406), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  AND3_X1   g215(.A1(new_n380), .A2(new_n388), .A3(new_n416), .ZN(new_n417));
  XNOR2_X1  g216(.A(KEYINPUT65), .B(G120gat), .ZN(new_n418));
  INV_X1    g217(.A(G113gat), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  XNOR2_X1  g219(.A(G127gat), .B(G134gat), .ZN(new_n421));
  INV_X1    g220(.A(G120gat), .ZN(new_n422));
  AOI21_X1  g221(.A(KEYINPUT1), .B1(new_n419), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT1), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n425), .B1(G113gat), .B2(G120gat), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n426), .B1(G113gat), .B2(G120gat), .ZN(new_n427));
  OAI22_X1  g226(.A1(new_n420), .A2(new_n424), .B1(new_n427), .B2(new_n421), .ZN(new_n428));
  AND2_X1   g227(.A1(G183gat), .A2(G190gat), .ZN(new_n429));
  INV_X1    g228(.A(G183gat), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(KEYINPUT27), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT27), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(G183gat), .ZN(new_n433));
  INV_X1    g232(.A(G190gat), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n431), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  AND2_X1   g234(.A1(KEYINPUT64), .A2(KEYINPUT28), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n429), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(G169gat), .A2(G176gat), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT26), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n440), .B1(G169gat), .B2(G176gat), .ZN(new_n441));
  NOR2_X1   g240(.A1(G169gat), .A2(G176gat), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(new_n439), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  NOR2_X1   g243(.A1(KEYINPUT64), .A2(KEYINPUT28), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n436), .A2(new_n445), .ZN(new_n446));
  XNOR2_X1  g245(.A(KEYINPUT27), .B(G183gat), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n446), .A2(new_n447), .A3(new_n434), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n437), .A2(new_n444), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(G183gat), .A2(G190gat), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n438), .B1(new_n450), .B2(KEYINPUT24), .ZN(new_n451));
  OAI21_X1  g250(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT23), .ZN(new_n453));
  INV_X1    g252(.A(G169gat), .ZN(new_n454));
  INV_X1    g253(.A(G176gat), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n453), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n451), .B1(new_n452), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n430), .A2(new_n434), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n458), .A2(KEYINPUT24), .A3(new_n450), .ZN(new_n459));
  AOI21_X1  g258(.A(KEYINPUT25), .B1(new_n457), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n451), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n456), .A2(new_n452), .ZN(new_n462));
  AND4_X1   g261(.A1(KEYINPUT25), .A2(new_n461), .A3(new_n462), .A4(new_n459), .ZN(new_n463));
  OAI211_X1 g262(.A(new_n428), .B(new_n449), .C1(new_n460), .C2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n457), .A2(KEYINPUT25), .A3(new_n459), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n461), .A2(new_n462), .A3(new_n459), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT25), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n428), .B1(new_n470), .B2(new_n449), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n465), .A2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(G227gat), .ZN(new_n473));
  INV_X1    g272(.A(G233gat), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  OAI21_X1  g274(.A(KEYINPUT34), .B1(new_n472), .B2(new_n475), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n449), .B1(new_n460), .B2(new_n463), .ZN(new_n477));
  INV_X1    g276(.A(G134gat), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(G127gat), .ZN(new_n479));
  INV_X1    g278(.A(G127gat), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(G134gat), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n482), .A2(new_n426), .ZN(new_n483));
  AND2_X1   g282(.A1(new_n422), .A2(KEYINPUT65), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n422), .A2(KEYINPUT65), .ZN(new_n485));
  OAI21_X1  g284(.A(G113gat), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n423), .B1(new_n419), .B2(new_n422), .ZN(new_n487));
  AOI22_X1  g286(.A1(new_n483), .A2(new_n486), .B1(new_n487), .B2(new_n482), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n477), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(new_n464), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT34), .ZN(new_n491));
  INV_X1    g290(.A(new_n475), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n490), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  AOI21_X1  g292(.A(KEYINPUT33), .B1(new_n472), .B2(new_n475), .ZN(new_n494));
  XNOR2_X1  g293(.A(G15gat), .B(G43gat), .ZN(new_n495));
  XNOR2_X1  g294(.A(G71gat), .B(G99gat), .ZN(new_n496));
  XNOR2_X1  g295(.A(new_n495), .B(new_n496), .ZN(new_n497));
  OAI211_X1 g296(.A(new_n476), .B(new_n493), .C1(new_n494), .C2(new_n497), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n489), .A2(new_n475), .A3(new_n464), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT33), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n497), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n491), .B1(new_n490), .B2(new_n492), .ZN(new_n502));
  AOI211_X1 g301(.A(KEYINPUT34), .B(new_n475), .C1(new_n489), .C2(new_n464), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n498), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n499), .A2(KEYINPUT32), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n506), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n498), .A2(new_n504), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  OR2_X1    g309(.A1(G141gat), .A2(G148gat), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT71), .ZN(new_n512));
  NAND2_X1  g311(.A1(G141gat), .A2(G148gat), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n511), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  AND2_X1   g313(.A1(G141gat), .A2(G148gat), .ZN(new_n515));
  NOR2_X1   g314(.A1(G141gat), .A2(G148gat), .ZN(new_n516));
  OAI21_X1  g315(.A(KEYINPUT71), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  OR2_X1    g316(.A1(KEYINPUT72), .A2(KEYINPUT2), .ZN(new_n518));
  NAND2_X1  g317(.A1(KEYINPUT72), .A2(KEYINPUT2), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n514), .A2(new_n517), .A3(new_n520), .ZN(new_n521));
  AND2_X1   g320(.A1(G155gat), .A2(G162gat), .ZN(new_n522));
  NOR2_X1   g321(.A1(G155gat), .A2(G162gat), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  XNOR2_X1  g323(.A(G141gat), .B(G148gat), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT2), .ZN(new_n527));
  OAI21_X1  g326(.A(KEYINPUT73), .B1(new_n522), .B2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT73), .ZN(new_n529));
  INV_X1    g328(.A(G155gat), .ZN(new_n530));
  INV_X1    g329(.A(G162gat), .ZN(new_n531));
  OAI211_X1 g330(.A(new_n529), .B(KEYINPUT2), .C1(new_n530), .C2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n528), .A2(new_n532), .ZN(new_n533));
  AOI22_X1  g332(.A1(new_n521), .A2(new_n524), .B1(new_n526), .B2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT67), .ZN(new_n535));
  NAND2_X1  g334(.A1(G211gat), .A2(G218gat), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  NOR2_X1   g336(.A1(G211gat), .A2(G218gat), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n535), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(G211gat), .ZN(new_n540));
  INV_X1    g339(.A(G218gat), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n542), .A2(KEYINPUT67), .A3(new_n536), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n539), .A2(new_n543), .ZN(new_n544));
  OR2_X1    g343(.A1(KEYINPUT66), .A2(KEYINPUT22), .ZN(new_n545));
  NAND2_X1  g344(.A1(KEYINPUT66), .A2(KEYINPUT22), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n545), .A2(new_n536), .A3(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(G197gat), .B(G204gat), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT68), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n544), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT29), .ZN(new_n552));
  AOI21_X1  g351(.A(KEYINPUT68), .B1(new_n547), .B2(new_n548), .ZN(new_n553));
  OAI211_X1 g352(.A(new_n551), .B(new_n552), .C1(new_n544), .C2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT3), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n534), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n521), .A2(new_n524), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n526), .A2(new_n533), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n557), .A2(new_n558), .A3(new_n555), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n549), .A2(new_n550), .ZN(new_n560));
  AND2_X1   g359(.A1(new_n539), .A2(new_n543), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AOI22_X1  g361(.A1(new_n559), .A2(new_n552), .B1(new_n562), .B2(new_n551), .ZN(new_n563));
  NAND2_X1  g362(.A1(G228gat), .A2(G233gat), .ZN(new_n564));
  NOR3_X1   g363(.A1(new_n556), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT80), .ZN(new_n567));
  AOI21_X1  g366(.A(KEYINPUT29), .B1(new_n544), .B2(new_n549), .ZN(new_n568));
  NAND4_X1  g367(.A1(new_n539), .A2(new_n547), .A3(new_n543), .A4(new_n548), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n534), .B1(new_n570), .B2(new_n555), .ZN(new_n571));
  OAI211_X1 g370(.A(new_n567), .B(new_n564), .C1(new_n563), .C2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  AOI21_X1  g372(.A(KEYINPUT29), .B1(new_n534), .B2(new_n555), .ZN(new_n574));
  AND2_X1   g373(.A1(new_n562), .A2(new_n551), .ZN(new_n575));
  AOI21_X1  g374(.A(KEYINPUT3), .B1(new_n568), .B2(new_n569), .ZN(new_n576));
  OAI22_X1  g375(.A1(new_n574), .A2(new_n575), .B1(new_n576), .B2(new_n534), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n567), .B1(new_n577), .B2(new_n564), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n566), .B1(new_n573), .B2(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(G78gat), .B(G106gat), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n580), .B(G50gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(KEYINPUT79), .B(KEYINPUT31), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n581), .B(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n579), .A2(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(KEYINPUT81), .B(G22gat), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n564), .B1(new_n563), .B2(new_n571), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n586), .A2(KEYINPUT80), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(new_n572), .ZN(new_n588));
  INV_X1    g387(.A(new_n583), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n588), .A2(new_n589), .A3(new_n566), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n584), .A2(new_n585), .A3(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n585), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n589), .B1(new_n588), .B2(new_n566), .ZN(new_n593));
  AOI211_X1 g392(.A(new_n583), .B(new_n565), .C1(new_n587), .C2(new_n572), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n592), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n510), .B1(new_n591), .B2(new_n595), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n488), .A2(new_n557), .A3(new_n558), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(KEYINPUT4), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT4), .ZN(new_n599));
  NAND4_X1  g398(.A1(new_n488), .A2(new_n557), .A3(new_n558), .A4(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n557), .A2(new_n558), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n602), .A2(KEYINPUT3), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n603), .A2(new_n559), .A3(new_n428), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT5), .ZN(new_n605));
  NAND2_X1  g404(.A1(G225gat), .A2(G233gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(KEYINPUT74), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  NAND4_X1  g407(.A1(new_n601), .A2(new_n604), .A3(new_n605), .A4(new_n608), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n428), .B1(new_n534), .B2(new_n555), .ZN(new_n610));
  INV_X1    g409(.A(new_n559), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n608), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT75), .ZN(new_n613));
  NAND4_X1  g412(.A1(new_n534), .A2(new_n613), .A3(new_n599), .A4(new_n488), .ZN(new_n614));
  AND2_X1   g413(.A1(new_n598), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n600), .A2(KEYINPUT75), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n612), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n524), .ZN(new_n618));
  AOI22_X1  g417(.A1(new_n525), .A2(KEYINPUT71), .B1(new_n518), .B2(new_n519), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n618), .B1(new_n619), .B2(new_n514), .ZN(new_n620));
  AND2_X1   g419(.A1(new_n526), .A2(new_n533), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n428), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT76), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n622), .A2(new_n623), .A3(new_n597), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n602), .A2(KEYINPUT76), .A3(new_n428), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n624), .A2(new_n607), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n626), .A2(KEYINPUT5), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n609), .B1(new_n617), .B2(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(G57gat), .B(G85gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(KEYINPUT78), .ZN(new_n630));
  XNOR2_X1  g429(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(G1gat), .B(G29gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n628), .A2(KEYINPUT6), .A3(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n635), .A2(KEYINPUT82), .ZN(new_n636));
  INV_X1    g435(.A(new_n634), .ZN(new_n637));
  AND3_X1   g436(.A1(new_n616), .A2(new_n614), .A3(new_n598), .ZN(new_n638));
  OAI211_X1 g437(.A(KEYINPUT5), .B(new_n626), .C1(new_n638), .C2(new_n612), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n637), .B1(new_n639), .B2(new_n609), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT82), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n640), .A2(new_n641), .A3(KEYINPUT6), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n636), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n628), .A2(new_n634), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT6), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n639), .A2(new_n637), .A3(new_n609), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n644), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  AOI21_X1  g446(.A(KEYINPUT35), .B1(new_n643), .B2(new_n647), .ZN(new_n648));
  AOI22_X1  g447(.A1(new_n477), .A2(new_n552), .B1(G226gat), .B2(G233gat), .ZN(new_n649));
  NAND2_X1  g448(.A1(G226gat), .A2(G233gat), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n650), .B1(new_n470), .B2(new_n449), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n575), .B1(new_n649), .B2(new_n651), .ZN(new_n652));
  AND3_X1   g451(.A1(new_n431), .A2(new_n433), .A3(new_n434), .ZN(new_n653));
  AOI22_X1  g452(.A1(new_n653), .A2(new_n446), .B1(new_n441), .B2(new_n443), .ZN(new_n654));
  AOI22_X1  g453(.A1(new_n469), .A2(new_n466), .B1(new_n654), .B2(new_n437), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n650), .B1(new_n655), .B2(KEYINPUT29), .ZN(new_n656));
  INV_X1    g455(.A(new_n575), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n477), .A2(G226gat), .A3(G233gat), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n656), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n652), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g459(.A(G8gat), .B(G36gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(G64gat), .B(G92gat), .ZN(new_n662));
  XOR2_X1   g461(.A(new_n661), .B(new_n662), .Z(new_n663));
  AOI21_X1  g462(.A(KEYINPUT70), .B1(new_n660), .B2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT70), .ZN(new_n665));
  INV_X1    g464(.A(new_n663), .ZN(new_n666));
  AOI211_X1 g465(.A(new_n665), .B(new_n666), .C1(new_n652), .C2(new_n659), .ZN(new_n667));
  NOR3_X1   g466(.A1(new_n664), .A2(new_n667), .A3(KEYINPUT30), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT69), .ZN(new_n669));
  NOR3_X1   g468(.A1(new_n649), .A2(new_n575), .A3(new_n651), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n657), .B1(new_n656), .B2(new_n658), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n669), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n652), .A2(new_n659), .A3(KEYINPUT69), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n672), .A2(new_n673), .A3(new_n666), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n660), .A2(KEYINPUT30), .A3(new_n663), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n668), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n596), .A2(new_n648), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n595), .A2(new_n591), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n647), .A2(new_n635), .ZN(new_n680));
  AND3_X1   g479(.A1(new_n498), .A2(new_n504), .A3(new_n508), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n508), .B1(new_n498), .B2(new_n504), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND4_X1  g482(.A1(new_n679), .A2(new_n677), .A3(new_n680), .A4(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(KEYINPUT35), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n678), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n677), .A2(new_n680), .ZN(new_n687));
  AND2_X1   g486(.A1(new_n595), .A2(new_n591), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n507), .A2(KEYINPUT36), .A3(new_n509), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT36), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n690), .B1(new_n681), .B2(new_n682), .ZN(new_n691));
  AOI22_X1  g490(.A1(new_n687), .A2(new_n688), .B1(new_n689), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n624), .A2(new_n625), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(new_n608), .ZN(new_n694));
  AND2_X1   g493(.A1(new_n601), .A2(new_n604), .ZN(new_n695));
  OAI211_X1 g494(.A(new_n694), .B(KEYINPUT39), .C1(new_n695), .C2(new_n608), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT39), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n608), .B1(new_n601), .B2(new_n604), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n634), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  AOI21_X1  g498(.A(KEYINPUT40), .B1(new_n696), .B2(new_n699), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n700), .A2(new_n640), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n696), .A2(new_n699), .A3(KEYINPUT40), .ZN(new_n702));
  OAI211_X1 g501(.A(new_n701), .B(new_n702), .C1(new_n668), .C2(new_n676), .ZN(new_n703));
  INV_X1    g502(.A(new_n642), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n641), .B1(new_n640), .B2(KEYINPUT6), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n647), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT37), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n707), .B1(new_n670), .B2(new_n671), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT38), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n652), .A2(new_n659), .A3(KEYINPUT37), .ZN(new_n710));
  NAND4_X1  g509(.A1(new_n708), .A2(new_n709), .A3(new_n666), .A4(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n660), .A2(new_n663), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(new_n665), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n660), .A2(KEYINPUT70), .A3(new_n663), .ZN(new_n714));
  AND3_X1   g513(.A1(new_n711), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n672), .A2(KEYINPUT37), .A3(new_n673), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n663), .B1(new_n660), .B2(new_n707), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(KEYINPUT38), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n715), .A2(new_n719), .ZN(new_n720));
  OAI211_X1 g519(.A(new_n679), .B(new_n703), .C1(new_n706), .C2(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n692), .A2(new_n721), .ZN(new_n722));
  AND3_X1   g521(.A1(new_n686), .A2(new_n722), .A3(KEYINPUT83), .ZN(new_n723));
  AOI21_X1  g522(.A(KEYINPUT83), .B1(new_n686), .B2(new_n722), .ZN(new_n724));
  OAI211_X1 g523(.A(new_n281), .B(new_n417), .C1(new_n723), .C2(new_n724), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n725), .A2(new_n680), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(new_n203), .ZN(G1324gat));
  INV_X1    g526(.A(KEYINPUT104), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT42), .ZN(new_n729));
  OAI21_X1  g528(.A(G8gat), .B1(new_n725), .B2(new_n677), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n686), .A2(new_n722), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT83), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n686), .A2(new_n722), .A3(KEYINPUT83), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n280), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n713), .A2(new_n714), .ZN(new_n736));
  OAI211_X1 g535(.A(new_n674), .B(new_n675), .C1(new_n736), .C2(KEYINPUT30), .ZN(new_n737));
  XOR2_X1   g536(.A(KEYINPUT16), .B(G8gat), .Z(new_n738));
  NAND4_X1  g537(.A1(new_n735), .A2(new_n737), .A3(new_n417), .A4(new_n738), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n729), .B1(new_n730), .B2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n739), .A2(new_n729), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n728), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  AND2_X1   g542(.A1(new_n739), .A2(new_n729), .ZN(new_n744));
  NOR3_X1   g543(.A1(new_n740), .A2(new_n744), .A3(KEYINPUT104), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n743), .A2(new_n745), .ZN(G1325gat));
  OAI21_X1  g545(.A(new_n208), .B1(new_n725), .B2(new_n510), .ZN(new_n747));
  OR2_X1    g546(.A1(new_n747), .A2(KEYINPUT105), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(KEYINPUT105), .ZN(new_n749));
  INV_X1    g548(.A(new_n725), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n691), .A2(new_n689), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n751), .A2(new_n208), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(KEYINPUT106), .ZN(new_n753));
  AOI22_X1  g552(.A1(new_n748), .A2(new_n749), .B1(new_n750), .B2(new_n753), .ZN(G1326gat));
  NOR2_X1   g553(.A1(new_n725), .A2(new_n679), .ZN(new_n755));
  XOR2_X1   g554(.A(KEYINPUT43), .B(G22gat), .Z(new_n756));
  XNOR2_X1  g555(.A(new_n755), .B(new_n756), .ZN(G1327gat));
  NOR2_X1   g556(.A1(new_n415), .A2(new_n386), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n735), .A2(new_n327), .A3(new_n758), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n680), .A2(G29gat), .ZN(new_n760));
  INV_X1    g559(.A(new_n760), .ZN(new_n761));
  OAI21_X1  g560(.A(KEYINPUT107), .B1(new_n759), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n758), .A2(new_n327), .ZN(new_n763));
  AOI211_X1 g562(.A(new_n280), .B(new_n763), .C1(new_n733), .C2(new_n734), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT107), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n764), .A2(new_n765), .A3(new_n760), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n762), .A2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT45), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n762), .A2(KEYINPUT45), .A3(new_n766), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT44), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n383), .A2(new_n771), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n772), .B1(new_n723), .B2(new_n724), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n731), .A2(new_n327), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(new_n771), .ZN(new_n775));
  AND2_X1   g574(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  AND2_X1   g575(.A1(new_n647), .A2(new_n635), .ZN(new_n777));
  NOR3_X1   g576(.A1(new_n280), .A2(new_n386), .A3(new_n415), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n776), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(KEYINPUT108), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(G29gat), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n779), .A2(KEYINPUT108), .ZN(new_n782));
  OAI211_X1 g581(.A(new_n769), .B(new_n770), .C1(new_n781), .C2(new_n782), .ZN(G1328gat));
  NOR3_X1   g582(.A1(new_n759), .A2(G36gat), .A3(new_n677), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n784), .B(KEYINPUT46), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n776), .A2(new_n737), .A3(new_n778), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(G36gat), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n785), .A2(new_n787), .ZN(G1329gat));
  INV_X1    g587(.A(KEYINPUT109), .ZN(new_n789));
  INV_X1    g588(.A(new_n751), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n773), .A2(new_n790), .A3(new_n775), .A4(new_n778), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(G43gat), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n510), .A2(G43gat), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n764), .A2(new_n793), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n789), .B1(new_n792), .B2(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT47), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n795), .B(new_n796), .ZN(G1330gat));
  NAND4_X1  g596(.A1(new_n773), .A2(new_n688), .A3(new_n775), .A4(new_n778), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(G50gat), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n688), .A2(new_n218), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n800), .B(KEYINPUT110), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n764), .A2(new_n801), .ZN(new_n802));
  OAI211_X1 g601(.A(new_n799), .B(new_n802), .C1(KEYINPUT111), .C2(KEYINPUT48), .ZN(new_n803));
  NAND2_X1  g602(.A1(KEYINPUT111), .A2(KEYINPUT48), .ZN(new_n804));
  XNOR2_X1  g603(.A(new_n803), .B(new_n804), .ZN(G1331gat));
  NAND4_X1  g604(.A1(new_n280), .A2(new_n380), .A3(new_n388), .A4(new_n415), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n806), .B1(new_n686), .B2(new_n722), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(new_n777), .ZN(new_n808));
  XNOR2_X1  g607(.A(new_n808), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g608(.A(new_n677), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n807), .A2(new_n810), .ZN(new_n811));
  XOR2_X1   g610(.A(new_n811), .B(KEYINPUT112), .Z(new_n812));
  NOR2_X1   g611(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n813));
  XNOR2_X1  g612(.A(new_n812), .B(new_n813), .ZN(G1333gat));
  INV_X1    g613(.A(G71gat), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n807), .A2(new_n815), .A3(new_n683), .ZN(new_n816));
  AND2_X1   g615(.A1(new_n807), .A2(new_n790), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n816), .B1(new_n817), .B2(new_n815), .ZN(new_n818));
  XOR2_X1   g617(.A(new_n818), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g618(.A1(new_n807), .A2(new_n688), .ZN(new_n820));
  XNOR2_X1  g619(.A(new_n820), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g620(.A1(new_n281), .A2(new_n386), .A3(new_n416), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n776), .A2(new_n777), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(G85gat), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n281), .A2(new_n386), .ZN(new_n825));
  AND2_X1   g624(.A1(new_n692), .A2(new_n721), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n679), .A2(new_n683), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n827), .A2(new_n737), .ZN(new_n828));
  AOI22_X1  g627(.A1(new_n828), .A2(new_n648), .B1(KEYINPUT35), .B2(new_n684), .ZN(new_n829));
  OAI211_X1 g628(.A(new_n327), .B(new_n825), .C1(new_n826), .C2(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT51), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT113), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n731), .A2(KEYINPUT51), .A3(new_n327), .A4(new_n825), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n832), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n830), .A2(KEYINPUT113), .A3(new_n831), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n416), .B1(new_n837), .B2(KEYINPUT114), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n838), .B1(KEYINPUT114), .B2(new_n837), .ZN(new_n839));
  OR2_X1    g638(.A1(new_n680), .A2(G85gat), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n824), .B1(new_n839), .B2(new_n840), .ZN(G1336gat));
  NAND3_X1  g640(.A1(new_n776), .A2(new_n737), .A3(new_n822), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(G92gat), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT52), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NOR3_X1   g644(.A1(new_n416), .A2(G92gat), .A3(new_n677), .ZN(new_n846));
  AND3_X1   g645(.A1(new_n835), .A2(new_n836), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n832), .A2(new_n834), .ZN(new_n848));
  AOI22_X1  g647(.A1(new_n842), .A2(G92gat), .B1(new_n848), .B2(new_n846), .ZN(new_n849));
  OAI22_X1  g648(.A1(new_n845), .A2(new_n847), .B1(new_n849), .B2(new_n844), .ZN(G1337gat));
  OR2_X1    g649(.A1(new_n510), .A2(G99gat), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n776), .A2(new_n790), .A3(new_n822), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(KEYINPUT115), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(G99gat), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n852), .A2(KEYINPUT115), .ZN(new_n855));
  OAI22_X1  g654(.A1(new_n839), .A2(new_n851), .B1(new_n854), .B2(new_n855), .ZN(G1338gat));
  INV_X1    g655(.A(KEYINPUT116), .ZN(new_n857));
  NAND4_X1  g656(.A1(new_n773), .A2(new_n688), .A3(new_n775), .A4(new_n822), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(G106gat), .ZN(new_n859));
  NOR3_X1   g658(.A1(new_n416), .A2(new_n679), .A3(G106gat), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n835), .A2(new_n836), .A3(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT53), .ZN(new_n862));
  AND3_X1   g661(.A1(new_n859), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n848), .A2(new_n860), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n862), .B1(new_n859), .B2(new_n864), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n857), .B1(new_n863), .B2(new_n865), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n859), .A2(new_n861), .A3(new_n862), .ZN(new_n867));
  AOI22_X1  g666(.A1(new_n858), .A2(G106gat), .B1(new_n848), .B2(new_n860), .ZN(new_n868));
  OAI211_X1 g667(.A(new_n867), .B(KEYINPUT116), .C1(new_n862), .C2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n866), .A2(new_n869), .ZN(G1339gat));
  AOI21_X1  g669(.A(new_n255), .B1(new_n262), .B2(new_n254), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n265), .A2(new_n266), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n272), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  AND2_X1   g672(.A1(new_n276), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n404), .A2(new_n398), .ZN(new_n875));
  INV_X1    g674(.A(new_n399), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n408), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT54), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n403), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NOR3_X1   g678(.A1(new_n397), .A2(new_n399), .A3(new_n409), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT117), .ZN(new_n881));
  OAI211_X1 g680(.A(KEYINPUT54), .B(new_n400), .C1(new_n880), .C2(new_n881), .ZN(new_n882));
  NOR4_X1   g681(.A1(new_n397), .A2(new_n399), .A3(KEYINPUT117), .A4(new_n409), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n879), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT55), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  OAI211_X1 g685(.A(new_n879), .B(KEYINPUT55), .C1(new_n882), .C2(new_n883), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n874), .A2(new_n886), .A3(new_n406), .A4(new_n887), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n386), .B1(new_n888), .B2(new_n327), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n327), .B1(new_n874), .B2(new_n415), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n886), .A2(new_n406), .A3(new_n887), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n890), .B1(new_n280), .B2(new_n891), .ZN(new_n892));
  AOI22_X1  g691(.A1(new_n889), .A2(new_n892), .B1(new_n417), .B2(new_n280), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n893), .A2(new_n680), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(new_n828), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n419), .B1(new_n895), .B2(new_n280), .ZN(new_n896));
  NOR4_X1   g695(.A1(new_n893), .A2(new_n680), .A3(new_n737), .A4(new_n827), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n897), .A2(G113gat), .A3(new_n281), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  XOR2_X1   g698(.A(new_n899), .B(KEYINPUT118), .Z(G1340gat));
  INV_X1    g699(.A(new_n895), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n901), .A2(new_n418), .A3(new_n415), .ZN(new_n902));
  AND2_X1   g701(.A1(new_n897), .A2(new_n415), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n902), .B1(new_n422), .B2(new_n903), .ZN(G1341gat));
  NOR3_X1   g703(.A1(new_n895), .A2(KEYINPUT119), .A3(new_n379), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n905), .A2(G127gat), .ZN(new_n906));
  OAI21_X1  g705(.A(KEYINPUT119), .B1(new_n895), .B2(new_n379), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n379), .A2(new_n480), .ZN(new_n908));
  AOI22_X1  g707(.A1(new_n906), .A2(new_n907), .B1(new_n897), .B2(new_n908), .ZN(G1342gat));
  AND2_X1   g708(.A1(new_n897), .A2(new_n327), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n910), .A2(new_n478), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n901), .A2(new_n478), .A3(new_n327), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n911), .B1(KEYINPUT56), .B2(new_n912), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n913), .B1(KEYINPUT56), .B2(new_n912), .ZN(G1343gat));
  INV_X1    g713(.A(KEYINPUT58), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n790), .A2(new_n679), .ZN(new_n916));
  INV_X1    g715(.A(new_n916), .ZN(new_n917));
  NOR3_X1   g716(.A1(new_n893), .A2(new_n680), .A3(new_n917), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n280), .A2(G141gat), .ZN(new_n919));
  AND3_X1   g718(.A1(new_n918), .A2(new_n677), .A3(new_n919), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n751), .A2(new_n777), .A3(new_n677), .ZN(new_n921));
  INV_X1    g720(.A(new_n921), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n889), .A2(new_n892), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n417), .A2(new_n280), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g724(.A(KEYINPUT57), .B1(new_n925), .B2(new_n688), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT57), .ZN(new_n927));
  NOR3_X1   g726(.A1(new_n893), .A2(new_n927), .A3(new_n679), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n922), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n929), .A2(KEYINPUT120), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n925), .A2(KEYINPUT57), .A3(new_n688), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n927), .B1(new_n893), .B2(new_n679), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT120), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n933), .A2(new_n934), .A3(new_n922), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n930), .A2(new_n281), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n920), .B1(new_n936), .B2(G141gat), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT122), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n933), .A2(new_n281), .A3(new_n922), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n939), .A2(G141gat), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n918), .A2(KEYINPUT121), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n925), .A2(new_n777), .A3(new_n916), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT121), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND4_X1  g743(.A1(new_n941), .A2(new_n944), .A3(new_n677), .A4(new_n919), .ZN(new_n945));
  AND4_X1   g744(.A1(new_n938), .A2(new_n940), .A3(new_n915), .A4(new_n945), .ZN(new_n946));
  AOI21_X1  g745(.A(KEYINPUT58), .B1(new_n939), .B2(G141gat), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n938), .B1(new_n947), .B2(new_n945), .ZN(new_n948));
  OAI22_X1  g747(.A1(new_n915), .A2(new_n937), .B1(new_n946), .B2(new_n948), .ZN(G1344gat));
  INV_X1    g748(.A(KEYINPUT59), .ZN(new_n950));
  AND3_X1   g749(.A1(new_n941), .A2(new_n944), .A3(new_n677), .ZN(new_n951));
  AOI211_X1 g750(.A(new_n950), .B(G148gat), .C1(new_n951), .C2(new_n415), .ZN(new_n952));
  NOR3_X1   g751(.A1(new_n921), .A2(new_n950), .A3(new_n416), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT123), .ZN(new_n954));
  XNOR2_X1  g753(.A(new_n924), .B(new_n954), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n955), .A2(new_n923), .ZN(new_n956));
  AOI21_X1  g755(.A(KEYINPUT57), .B1(new_n956), .B2(new_n688), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n953), .B1(new_n957), .B2(new_n928), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n934), .B1(new_n933), .B2(new_n922), .ZN(new_n959));
  AOI211_X1 g758(.A(KEYINPUT120), .B(new_n921), .C1(new_n931), .C2(new_n932), .ZN(new_n960));
  NOR3_X1   g759(.A1(new_n959), .A2(new_n960), .A3(new_n416), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n958), .B1(new_n961), .B2(KEYINPUT59), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n952), .B1(new_n962), .B2(G148gat), .ZN(G1345gat));
  NAND3_X1  g762(.A1(new_n951), .A2(new_n530), .A3(new_n386), .ZN(new_n964));
  NOR3_X1   g763(.A1(new_n959), .A2(new_n960), .A3(new_n379), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n964), .B1(new_n965), .B2(new_n530), .ZN(G1346gat));
  AOI21_X1  g765(.A(G162gat), .B1(new_n951), .B2(new_n327), .ZN(new_n967));
  NOR2_X1   g766(.A1(new_n959), .A2(new_n960), .ZN(new_n968));
  NOR2_X1   g767(.A1(new_n383), .A2(new_n531), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n967), .B1(new_n968), .B2(new_n969), .ZN(G1347gat));
  NAND2_X1  g769(.A1(new_n737), .A2(new_n680), .ZN(new_n971));
  XNOR2_X1  g770(.A(new_n971), .B(KEYINPUT124), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n972), .A2(new_n827), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n925), .A2(new_n973), .ZN(new_n974));
  NOR3_X1   g773(.A1(new_n974), .A2(new_n454), .A3(new_n280), .ZN(new_n975));
  NOR2_X1   g774(.A1(new_n893), .A2(new_n777), .ZN(new_n976));
  NOR2_X1   g775(.A1(new_n827), .A2(new_n677), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  INV_X1    g777(.A(new_n978), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n979), .A2(new_n281), .ZN(new_n980));
  AOI21_X1  g779(.A(new_n975), .B1(new_n980), .B2(new_n454), .ZN(G1348gat));
  OAI21_X1  g780(.A(G176gat), .B1(new_n974), .B2(new_n416), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n415), .A2(new_n455), .ZN(new_n983));
  OAI21_X1  g782(.A(new_n982), .B1(new_n978), .B2(new_n983), .ZN(G1349gat));
  OAI21_X1  g783(.A(G183gat), .B1(new_n974), .B2(new_n379), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n386), .A2(new_n447), .ZN(new_n986));
  OAI21_X1  g785(.A(new_n985), .B1(new_n978), .B2(new_n986), .ZN(new_n987));
  XNOR2_X1  g786(.A(new_n987), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g787(.A1(new_n979), .A2(new_n434), .A3(new_n327), .ZN(new_n989));
  NOR4_X1   g788(.A1(new_n893), .A2(new_n827), .A3(new_n383), .A4(new_n972), .ZN(new_n990));
  OAI21_X1  g789(.A(KEYINPUT125), .B1(new_n990), .B2(new_n434), .ZN(new_n991));
  INV_X1    g790(.A(KEYINPUT61), .ZN(new_n992));
  INV_X1    g791(.A(KEYINPUT125), .ZN(new_n993));
  OAI211_X1 g792(.A(new_n993), .B(G190gat), .C1(new_n974), .C2(new_n383), .ZN(new_n994));
  AND3_X1   g793(.A1(new_n991), .A2(new_n992), .A3(new_n994), .ZN(new_n995));
  AOI21_X1  g794(.A(new_n992), .B1(new_n991), .B2(new_n994), .ZN(new_n996));
  OAI21_X1  g795(.A(new_n989), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  INV_X1    g796(.A(KEYINPUT126), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  OAI211_X1 g798(.A(KEYINPUT126), .B(new_n989), .C1(new_n995), .C2(new_n996), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n999), .A2(new_n1000), .ZN(G1351gat));
  NOR2_X1   g800(.A1(new_n972), .A2(new_n790), .ZN(new_n1002));
  INV_X1    g801(.A(G197gat), .ZN(new_n1003));
  NOR2_X1   g802(.A1(new_n280), .A2(new_n1003), .ZN(new_n1004));
  OAI211_X1 g803(.A(new_n1002), .B(new_n1004), .C1(new_n957), .C2(new_n928), .ZN(new_n1005));
  NOR4_X1   g804(.A1(new_n893), .A2(new_n777), .A3(new_n677), .A4(new_n917), .ZN(new_n1006));
  NAND2_X1  g805(.A1(new_n1006), .A2(new_n281), .ZN(new_n1007));
  NAND2_X1  g806(.A1(new_n1007), .A2(new_n1003), .ZN(new_n1008));
  NAND2_X1  g807(.A1(new_n1005), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g808(.A1(new_n1009), .A2(KEYINPUT127), .ZN(new_n1010));
  INV_X1    g809(.A(KEYINPUT127), .ZN(new_n1011));
  NAND3_X1  g810(.A1(new_n1005), .A2(new_n1011), .A3(new_n1008), .ZN(new_n1012));
  NAND2_X1  g811(.A1(new_n1010), .A2(new_n1012), .ZN(G1352gat));
  OR2_X1    g812(.A1(new_n957), .A2(new_n928), .ZN(new_n1014));
  NAND3_X1  g813(.A1(new_n1014), .A2(new_n415), .A3(new_n1002), .ZN(new_n1015));
  NAND2_X1  g814(.A1(new_n1015), .A2(G204gat), .ZN(new_n1016));
  INV_X1    g815(.A(G204gat), .ZN(new_n1017));
  NAND3_X1  g816(.A1(new_n1006), .A2(new_n1017), .A3(new_n415), .ZN(new_n1018));
  XOR2_X1   g817(.A(new_n1018), .B(KEYINPUT62), .Z(new_n1019));
  NAND2_X1  g818(.A1(new_n1016), .A2(new_n1019), .ZN(G1353gat));
  NAND3_X1  g819(.A1(new_n1006), .A2(new_n540), .A3(new_n386), .ZN(new_n1021));
  OAI211_X1 g820(.A(new_n386), .B(new_n1002), .C1(new_n957), .C2(new_n928), .ZN(new_n1022));
  AND3_X1   g821(.A1(new_n1022), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1023));
  AOI21_X1  g822(.A(KEYINPUT63), .B1(new_n1022), .B2(G211gat), .ZN(new_n1024));
  OAI21_X1  g823(.A(new_n1021), .B1(new_n1023), .B2(new_n1024), .ZN(G1354gat));
  NAND3_X1  g824(.A1(new_n1014), .A2(new_n327), .A3(new_n1002), .ZN(new_n1026));
  NAND2_X1  g825(.A1(new_n1026), .A2(G218gat), .ZN(new_n1027));
  NAND3_X1  g826(.A1(new_n1006), .A2(new_n541), .A3(new_n327), .ZN(new_n1028));
  NAND2_X1  g827(.A1(new_n1027), .A2(new_n1028), .ZN(G1355gat));
endmodule


