//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 1 0 0 0 1 0 0 1 0 1 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 1 0 0 0 0 0 0 1 1 1 0 1 1 0 0 1 1 1 0 1 1 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:02 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n550, new_n551,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n624, new_n625, new_n628, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n855, new_n856, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1175;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT65), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT66), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(G2106), .ZN(new_n455));
  INV_X1    g030(.A(G567), .ZN(new_n456));
  OAI22_X1  g031(.A1(new_n451), .A2(new_n455), .B1(new_n456), .B2(new_n452), .ZN(new_n457));
  XNOR2_X1  g032(.A(new_n457), .B(KEYINPUT67), .ZN(G319));
  INV_X1    g033(.A(KEYINPUT68), .ZN(new_n459));
  AND2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  OAI211_X1 g036(.A(new_n459), .B(G125), .C1(new_n460), .C2(new_n461), .ZN(new_n462));
  NAND3_X1  g037(.A1(KEYINPUT69), .A2(G113), .A3(G2104), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT69), .ZN(new_n464));
  INV_X1    g039(.A(G113), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n462), .A2(new_n463), .A3(new_n467), .ZN(new_n468));
  OR2_X1    g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n459), .B1(new_n471), .B2(G125), .ZN(new_n472));
  OAI21_X1  g047(.A(G2105), .B1(new_n468), .B2(new_n472), .ZN(new_n473));
  AOI21_X1  g048(.A(G2105), .B1(new_n469), .B2(new_n470), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n466), .A2(G2105), .ZN(new_n475));
  AOI22_X1  g050(.A1(new_n474), .A2(G137), .B1(G101), .B2(new_n475), .ZN(new_n476));
  AND2_X1   g051(.A1(new_n473), .A2(new_n476), .ZN(G160));
  NAND2_X1  g052(.A1(new_n474), .A2(G136), .ZN(new_n478));
  INV_X1    g053(.A(G2105), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n479), .B1(new_n469), .B2(new_n470), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  OR2_X1    g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n482), .B(G2104), .C1(G112), .C2(new_n479), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n478), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  OAI211_X1 g060(.A(G126), .B(G2105), .C1(new_n460), .C2(new_n461), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n479), .A2(G114), .ZN(new_n487));
  OAI21_X1  g062(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n486), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  OAI211_X1 g064(.A(G138), .B(new_n479), .C1(new_n460), .C2(new_n461), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(KEYINPUT4), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n474), .A2(new_n492), .A3(G138), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n489), .B1(new_n491), .B2(new_n493), .ZN(G164));
  INV_X1    g069(.A(KEYINPUT70), .ZN(new_n495));
  INV_X1    g070(.A(G543), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n495), .B1(new_n496), .B2(KEYINPUT5), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT5), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n498), .A2(KEYINPUT70), .A3(G543), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n496), .A2(KEYINPUT5), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n500), .A2(G62), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(G75), .A2(G543), .ZN(new_n503));
  XOR2_X1   g078(.A(new_n503), .B(KEYINPUT71), .Z(new_n504));
  NAND2_X1  g079(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G651), .ZN(new_n506));
  XNOR2_X1  g081(.A(KEYINPUT6), .B(G651), .ZN(new_n507));
  NAND4_X1  g082(.A1(new_n500), .A2(G88), .A3(new_n501), .A4(new_n507), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n507), .A2(G50), .A3(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT72), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n506), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n514), .B1(new_n502), .B2(new_n504), .ZN(new_n515));
  OAI21_X1  g090(.A(KEYINPUT72), .B1(new_n515), .B2(new_n510), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n513), .A2(new_n516), .ZN(G166));
  NOR2_X1   g092(.A1(new_n498), .A2(G543), .ZN(new_n518));
  AOI21_X1  g093(.A(new_n518), .B1(new_n497), .B2(new_n499), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n519), .A2(G63), .A3(G651), .ZN(new_n520));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n521), .B(KEYINPUT7), .ZN(new_n522));
  INV_X1    g097(.A(G51), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n507), .A2(G543), .ZN(new_n524));
  OAI211_X1 g099(.A(new_n520), .B(new_n522), .C1(new_n523), .C2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n519), .A2(new_n507), .ZN(new_n526));
  XNOR2_X1  g101(.A(KEYINPUT73), .B(G89), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n525), .A2(new_n528), .ZN(G168));
  AND2_X1   g104(.A1(new_n519), .A2(new_n507), .ZN(new_n530));
  XNOR2_X1  g105(.A(KEYINPUT74), .B(G90), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(new_n524), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(G52), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n519), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  OAI211_X1 g110(.A(new_n532), .B(new_n534), .C1(new_n514), .C2(new_n535), .ZN(G301));
  INV_X1    g111(.A(G301), .ZN(G171));
  NAND3_X1  g112(.A1(new_n500), .A2(G56), .A3(new_n501), .ZN(new_n538));
  NAND2_X1  g113(.A1(G68), .A2(G543), .ZN(new_n539));
  AOI21_X1  g114(.A(new_n514), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  AND2_X1   g115(.A1(KEYINPUT75), .A2(G81), .ZN(new_n541));
  NOR2_X1   g116(.A1(KEYINPUT75), .A2(G81), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND4_X1  g118(.A1(new_n500), .A2(new_n501), .A3(new_n507), .A4(new_n543), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n507), .A2(G43), .A3(G543), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n540), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(G153));
  NAND4_X1  g123(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g124(.A1(G1), .A2(G3), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT8), .ZN(new_n551));
  NAND4_X1  g126(.A1(G319), .A2(G483), .A3(G661), .A4(new_n551), .ZN(G188));
  NAND3_X1  g127(.A1(new_n507), .A2(G53), .A3(G543), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(KEYINPUT9), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT9), .ZN(new_n555));
  NAND4_X1  g130(.A1(new_n507), .A2(new_n555), .A3(G53), .A4(G543), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n530), .A2(G91), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n500), .A2(G65), .A3(new_n501), .ZN(new_n558));
  NAND2_X1  g133(.A1(G78), .A2(G543), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  AOI21_X1  g135(.A(KEYINPUT76), .B1(new_n560), .B2(G651), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT76), .ZN(new_n562));
  AOI211_X1 g137(.A(new_n562), .B(new_n514), .C1(new_n558), .C2(new_n559), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n557), .B1(new_n561), .B2(new_n563), .ZN(G299));
  INV_X1    g139(.A(G168), .ZN(G286));
  INV_X1    g140(.A(G166), .ZN(G303));
  NAND3_X1  g141(.A1(new_n507), .A2(G49), .A3(G543), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT77), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n567), .B(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n530), .A2(G87), .ZN(new_n570));
  OAI21_X1  g145(.A(G651), .B1(new_n519), .B2(G74), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(G288));
  INV_X1    g147(.A(KEYINPUT78), .ZN(new_n573));
  NAND2_X1  g148(.A1(G73), .A2(G543), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n575), .B1(new_n519), .B2(G61), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n573), .B1(new_n576), .B2(new_n514), .ZN(new_n577));
  AND3_X1   g152(.A1(new_n498), .A2(KEYINPUT70), .A3(G543), .ZN(new_n578));
  AOI21_X1  g153(.A(KEYINPUT70), .B1(new_n498), .B2(G543), .ZN(new_n579));
  OAI211_X1 g154(.A(G61), .B(new_n501), .C1(new_n578), .C2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n580), .A2(new_n574), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n581), .A2(KEYINPUT78), .A3(G651), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n519), .A2(G86), .A3(new_n507), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n507), .A2(G48), .A3(G543), .ZN(new_n584));
  AND2_X1   g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n577), .A2(new_n582), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n586), .A2(KEYINPUT79), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT79), .ZN(new_n588));
  NAND4_X1  g163(.A1(new_n577), .A2(new_n582), .A3(new_n585), .A4(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(G305));
  INV_X1    g166(.A(KEYINPUT81), .ZN(new_n592));
  NAND2_X1  g167(.A1(G72), .A2(G543), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n594), .B1(new_n519), .B2(G60), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT80), .ZN(new_n596));
  OAI21_X1  g171(.A(G651), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  AOI211_X1 g172(.A(KEYINPUT80), .B(new_n594), .C1(new_n519), .C2(G60), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n592), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n500), .A2(G60), .A3(new_n501), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n600), .A2(new_n593), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n601), .A2(KEYINPUT80), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n595), .A2(new_n596), .ZN(new_n603));
  NAND4_X1  g178(.A1(new_n602), .A2(new_n603), .A3(KEYINPUT81), .A4(G651), .ZN(new_n604));
  INV_X1    g179(.A(G85), .ZN(new_n605));
  INV_X1    g180(.A(G47), .ZN(new_n606));
  OAI22_X1  g181(.A1(new_n526), .A2(new_n605), .B1(new_n606), .B2(new_n524), .ZN(new_n607));
  INV_X1    g182(.A(new_n607), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n599), .A2(new_n604), .A3(new_n608), .ZN(G290));
  NAND2_X1  g184(.A1(G301), .A2(G868), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n519), .A2(G66), .ZN(new_n611));
  NAND2_X1  g186(.A1(G79), .A2(G543), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  AOI22_X1  g188(.A1(new_n613), .A2(G651), .B1(G54), .B2(new_n533), .ZN(new_n614));
  INV_X1    g189(.A(KEYINPUT10), .ZN(new_n615));
  INV_X1    g190(.A(G92), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n526), .B2(new_n616), .ZN(new_n617));
  NAND4_X1  g192(.A1(new_n519), .A2(KEYINPUT10), .A3(G92), .A4(new_n507), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n614), .A2(new_n619), .ZN(new_n620));
  INV_X1    g195(.A(new_n620), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n610), .B1(new_n621), .B2(G868), .ZN(G284));
  OAI21_X1  g197(.A(new_n610), .B1(new_n621), .B2(G868), .ZN(G321));
  NAND2_X1  g198(.A1(G286), .A2(G868), .ZN(new_n624));
  INV_X1    g199(.A(G299), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n624), .B1(new_n625), .B2(G868), .ZN(G297));
  OAI21_X1  g201(.A(new_n624), .B1(new_n625), .B2(G868), .ZN(G280));
  INV_X1    g202(.A(G559), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n621), .B1(new_n628), .B2(G860), .ZN(G148));
  NOR2_X1   g204(.A1(new_n547), .A2(G868), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n621), .A2(KEYINPUT82), .A3(new_n628), .ZN(new_n631));
  INV_X1    g206(.A(KEYINPUT82), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n632), .B1(new_n620), .B2(G559), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  AOI21_X1  g209(.A(new_n630), .B1(new_n634), .B2(G868), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n635), .B(KEYINPUT83), .Z(G323));
  XNOR2_X1  g211(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g212(.A1(new_n471), .A2(new_n475), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n638), .B(KEYINPUT12), .Z(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(KEYINPUT13), .Z(new_n640));
  INV_X1    g215(.A(G2100), .ZN(new_n641));
  NOR2_X1   g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n642), .B(KEYINPUT84), .Z(new_n643));
  OR3_X1    g218(.A1(new_n479), .A2(KEYINPUT86), .A3(G111), .ZN(new_n644));
  OAI21_X1  g219(.A(KEYINPUT86), .B1(new_n479), .B2(G111), .ZN(new_n645));
  OR2_X1    g220(.A1(G99), .A2(G2105), .ZN(new_n646));
  AND4_X1   g221(.A1(G2104), .A2(new_n644), .A3(new_n645), .A4(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n474), .A2(G135), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(KEYINPUT85), .Z(new_n649));
  AOI211_X1 g224(.A(new_n647), .B(new_n649), .C1(G123), .C2(new_n480), .ZN(new_n650));
  INV_X1    g225(.A(G2096), .ZN(new_n651));
  AOI22_X1  g226(.A1(new_n650), .A2(new_n651), .B1(new_n640), .B2(new_n641), .ZN(new_n652));
  OAI211_X1 g227(.A(new_n643), .B(new_n652), .C1(new_n651), .C2(new_n650), .ZN(G156));
  XNOR2_X1  g228(.A(G2427), .B(G2438), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2430), .ZN(new_n655));
  XNOR2_X1  g230(.A(KEYINPUT15), .B(G2435), .ZN(new_n656));
  OR2_X1    g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n655), .A2(new_n656), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n657), .A2(KEYINPUT14), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT88), .ZN(new_n660));
  XOR2_X1   g235(.A(G1341), .B(G1348), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G2451), .B(G2454), .Z(new_n663));
  XNOR2_X1  g238(.A(G2443), .B(G2446), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n662), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(KEYINPUT87), .B(KEYINPUT16), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g243(.A(G14), .ZN(new_n669));
  AOI21_X1  g244(.A(new_n669), .B1(new_n666), .B2(new_n667), .ZN(new_n670));
  AND2_X1   g245(.A1(new_n668), .A2(new_n670), .ZN(G401));
  XOR2_X1   g246(.A(G2072), .B(G2078), .Z(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G2067), .B(G2678), .ZN(new_n674));
  XOR2_X1   g249(.A(G2084), .B(G2090), .Z(new_n675));
  NAND3_X1  g250(.A1(new_n673), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n676), .B(KEYINPUT18), .Z(new_n677));
  INV_X1    g252(.A(new_n674), .ZN(new_n678));
  AOI21_X1  g253(.A(new_n675), .B1(new_n678), .B2(new_n672), .ZN(new_n679));
  XOR2_X1   g254(.A(KEYINPUT89), .B(KEYINPUT17), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n672), .B(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n679), .B1(new_n682), .B2(new_n678), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n682), .A2(new_n678), .A3(new_n675), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n677), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(G2096), .B(G2100), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(G227));
  XNOR2_X1  g262(.A(G1971), .B(G1976), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT19), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(G1961), .B(G1966), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT90), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1956), .B(G2474), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n690), .A2(new_n692), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT20), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n690), .B1(new_n692), .B2(new_n694), .ZN(new_n697));
  OR2_X1    g272(.A1(new_n692), .A2(new_n694), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  OAI211_X1 g274(.A(new_n696), .B(new_n699), .C1(new_n689), .C2(new_n698), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT91), .ZN(new_n701));
  XNOR2_X1  g276(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  XOR2_X1   g278(.A(G1991), .B(G1996), .Z(new_n704));
  OR2_X1    g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n703), .A2(new_n704), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(G1981), .B(G1986), .ZN(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n705), .A2(new_n708), .A3(new_n706), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(G229));
  AND2_X1   g288(.A1(new_n475), .A2(G105), .ZN(new_n714));
  NAND3_X1  g289(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT26), .ZN(new_n716));
  AOI211_X1 g291(.A(new_n714), .B(new_n716), .C1(G141), .C2(new_n474), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n480), .A2(G129), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT97), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(G29), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(new_n722), .B2(G32), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT98), .ZN(new_n725));
  XNOR2_X1  g300(.A(KEYINPUT27), .B(G1996), .ZN(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  OR2_X1    g302(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n725), .A2(new_n727), .ZN(new_n729));
  INV_X1    g304(.A(G16), .ZN(new_n730));
  NOR2_X1   g305(.A1(G168), .A2(new_n730), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(new_n730), .B2(G21), .ZN(new_n732));
  INV_X1    g307(.A(G1966), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT99), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n728), .A2(new_n729), .A3(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(KEYINPUT30), .ZN(new_n737));
  AND2_X1   g312(.A1(new_n737), .A2(G28), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n722), .B1(new_n737), .B2(G28), .ZN(new_n739));
  AND2_X1   g314(.A1(KEYINPUT31), .A2(G11), .ZN(new_n740));
  NOR2_X1   g315(.A1(KEYINPUT31), .A2(G11), .ZN(new_n741));
  OAI22_X1  g316(.A1(new_n738), .A2(new_n739), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(new_n650), .B2(G29), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(new_n732), .B2(new_n733), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n730), .A2(G5), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(G171), .B2(new_n730), .ZN(new_n746));
  NAND2_X1  g321(.A1(G160), .A2(G29), .ZN(new_n747));
  INV_X1    g322(.A(G34), .ZN(new_n748));
  AOI21_X1  g323(.A(G29), .B1(new_n748), .B2(KEYINPUT24), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(KEYINPUT24), .B2(new_n748), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n747), .A2(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(G2084), .ZN(new_n752));
  AOI22_X1  g327(.A1(new_n746), .A2(G1961), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(G2072), .ZN(new_n754));
  AND2_X1   g329(.A1(new_n722), .A2(G33), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n471), .A2(G127), .ZN(new_n756));
  INV_X1    g331(.A(G115), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n756), .B1(new_n757), .B2(new_n466), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT95), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n479), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(new_n759), .B2(new_n758), .ZN(new_n761));
  INV_X1    g336(.A(KEYINPUT25), .ZN(new_n762));
  NAND2_X1  g337(.A1(G103), .A2(G2104), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n762), .B1(new_n763), .B2(G2105), .ZN(new_n764));
  NAND4_X1  g339(.A1(new_n479), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n765));
  AOI22_X1  g340(.A1(new_n474), .A2(G139), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n761), .A2(new_n766), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n755), .B1(new_n767), .B2(G29), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n753), .B1(new_n754), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n768), .A2(new_n754), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G1961), .B2(new_n746), .ZN(new_n771));
  NOR2_X1   g346(.A1(G27), .A2(G29), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(G164), .B2(G29), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(G2078), .ZN(new_n774));
  NOR4_X1   g349(.A1(new_n744), .A2(new_n769), .A3(new_n771), .A4(new_n774), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n751), .A2(new_n752), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT96), .Z(new_n777));
  NAND2_X1  g352(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(KEYINPUT100), .ZN(new_n779));
  OR3_X1    g354(.A1(new_n736), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  XOR2_X1   g355(.A(KEYINPUT102), .B(KEYINPUT23), .Z(new_n781));
  NAND2_X1  g356(.A1(new_n730), .A2(G20), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(new_n625), .B2(new_n730), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(G1956), .ZN(new_n785));
  NAND2_X1  g360(.A1(G162), .A2(G29), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(G29), .B2(G35), .ZN(new_n787));
  XNOR2_X1  g362(.A(KEYINPUT101), .B(KEYINPUT29), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(new_n789), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n785), .B1(G2090), .B2(new_n790), .ZN(new_n791));
  OR2_X1    g366(.A1(new_n791), .A2(KEYINPUT103), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n547), .A2(new_n730), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(new_n730), .B2(G19), .ZN(new_n794));
  INV_X1    g369(.A(new_n794), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n795), .A2(G1341), .ZN(new_n796));
  INV_X1    g371(.A(G1341), .ZN(new_n797));
  OAI22_X1  g372(.A1(new_n790), .A2(G2090), .B1(new_n797), .B2(new_n794), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n722), .A2(G26), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT28), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n474), .A2(G140), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n480), .A2(G128), .ZN(new_n802));
  OR2_X1    g377(.A1(G104), .A2(G2105), .ZN(new_n803));
  OAI211_X1 g378(.A(new_n803), .B(G2104), .C1(G116), .C2(new_n479), .ZN(new_n804));
  NAND3_X1  g379(.A1(new_n801), .A2(new_n802), .A3(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(new_n805), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n800), .B1(new_n806), .B2(new_n722), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(G2067), .ZN(new_n808));
  NOR2_X1   g383(.A1(G4), .A2(G16), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(new_n621), .B2(G16), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(G1348), .ZN(new_n811));
  OR4_X1    g386(.A1(new_n796), .A2(new_n798), .A3(new_n808), .A4(new_n811), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(new_n791), .B2(KEYINPUT103), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n779), .B1(new_n736), .B2(new_n778), .ZN(new_n814));
  NAND4_X1  g389(.A1(new_n780), .A2(new_n792), .A3(new_n813), .A4(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n730), .A2(G6), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(new_n590), .B2(new_n730), .ZN(new_n817));
  XNOR2_X1  g392(.A(KEYINPUT32), .B(G1981), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NOR2_X1   g394(.A1(G16), .A2(G23), .ZN(new_n820));
  XOR2_X1   g395(.A(new_n820), .B(KEYINPUT93), .Z(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(G288), .B2(new_n730), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT94), .ZN(new_n823));
  XNOR2_X1  g398(.A(KEYINPUT33), .B(G1976), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n823), .B(new_n824), .ZN(new_n825));
  OR2_X1    g400(.A1(new_n817), .A2(new_n818), .ZN(new_n826));
  NOR2_X1   g401(.A1(G16), .A2(G22), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n827), .B1(G166), .B2(G16), .ZN(new_n828));
  INV_X1    g403(.A(G1971), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n828), .B(new_n829), .ZN(new_n830));
  AND4_X1   g405(.A1(new_n819), .A2(new_n825), .A3(new_n826), .A4(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT34), .ZN(new_n832));
  OR2_X1    g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n831), .A2(new_n832), .ZN(new_n834));
  INV_X1    g409(.A(G290), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n835), .A2(G16), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n836), .B1(G16), .B2(G24), .ZN(new_n837));
  INV_X1    g412(.A(G1986), .ZN(new_n838));
  AND2_X1   g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n837), .A2(new_n838), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n474), .A2(G131), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n480), .A2(G119), .ZN(new_n842));
  OR2_X1    g417(.A1(G95), .A2(G2105), .ZN(new_n843));
  OAI211_X1 g418(.A(new_n843), .B(G2104), .C1(G107), .C2(new_n479), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n841), .A2(new_n842), .A3(new_n844), .ZN(new_n845));
  MUX2_X1   g420(.A(G25), .B(new_n845), .S(G29), .Z(new_n846));
  XOR2_X1   g421(.A(KEYINPUT35), .B(G1991), .Z(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT92), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n846), .B(new_n848), .ZN(new_n849));
  NOR3_X1   g424(.A1(new_n839), .A2(new_n840), .A3(new_n849), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n833), .A2(new_n834), .A3(new_n850), .ZN(new_n851));
  OR2_X1    g426(.A1(new_n851), .A2(KEYINPUT36), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(KEYINPUT36), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n815), .B1(new_n852), .B2(new_n853), .ZN(G311));
  NAND2_X1  g429(.A1(new_n852), .A2(new_n853), .ZN(new_n855));
  INV_X1    g430(.A(new_n815), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(G150));
  NAND2_X1  g432(.A1(new_n621), .A2(G559), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(KEYINPUT38), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n538), .A2(new_n539), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n860), .A2(G651), .ZN(new_n861));
  AND2_X1   g436(.A1(new_n544), .A2(new_n545), .ZN(new_n862));
  OAI211_X1 g437(.A(G67), .B(new_n501), .C1(new_n578), .C2(new_n579), .ZN(new_n863));
  NAND2_X1  g438(.A1(G80), .A2(G543), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n865), .A2(G651), .ZN(new_n866));
  NAND4_X1  g441(.A1(new_n500), .A2(G93), .A3(new_n501), .A4(new_n507), .ZN(new_n867));
  XOR2_X1   g442(.A(KEYINPUT104), .B(G55), .Z(new_n868));
  NAND3_X1  g443(.A1(new_n868), .A2(G543), .A3(new_n507), .ZN(new_n869));
  AND2_X1   g444(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  NAND4_X1  g445(.A1(new_n861), .A2(new_n862), .A3(new_n866), .A4(new_n870), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n514), .B1(new_n863), .B2(new_n864), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n867), .A2(new_n869), .ZN(new_n873));
  OAI22_X1  g448(.A1(new_n546), .A2(new_n540), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n871), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n859), .B(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT39), .ZN(new_n877));
  AOI21_X1  g452(.A(G860), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n878), .B1(new_n877), .B2(new_n876), .ZN(new_n879));
  OAI21_X1  g454(.A(G860), .B1(new_n872), .B2(new_n873), .ZN(new_n880));
  XOR2_X1   g455(.A(new_n880), .B(KEYINPUT37), .Z(new_n881));
  NAND2_X1  g456(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  XOR2_X1   g457(.A(new_n882), .B(KEYINPUT105), .Z(G145));
  XNOR2_X1  g458(.A(new_n767), .B(new_n720), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n639), .B(new_n845), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n884), .B(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(G164), .B(new_n805), .ZN(new_n887));
  AOI22_X1  g462(.A1(G130), .A2(new_n480), .B1(new_n474), .B2(G142), .ZN(new_n888));
  OAI21_X1  g463(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT106), .ZN(new_n890));
  INV_X1    g465(.A(G118), .ZN(new_n891));
  AOI22_X1  g466(.A1(new_n889), .A2(new_n890), .B1(new_n891), .B2(G2105), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n892), .B1(new_n890), .B2(new_n889), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n888), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n887), .B(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n886), .B(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(G160), .B(new_n484), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n650), .B(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(G37), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n899), .B1(new_n898), .B2(new_n896), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g476(.A(new_n634), .B(new_n875), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(G299), .A2(new_n620), .ZN(new_n904));
  AOI22_X1  g479(.A1(new_n519), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n562), .B1(new_n905), .B2(new_n514), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n560), .A2(KEYINPUT76), .A3(G651), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND4_X1  g483(.A1(new_n908), .A2(new_n557), .A3(new_n619), .A4(new_n614), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n904), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g485(.A(KEYINPUT107), .B1(new_n903), .B2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT41), .ZN(new_n912));
  AND3_X1   g487(.A1(new_n904), .A2(new_n912), .A3(new_n909), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n912), .B1(new_n904), .B2(new_n909), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n903), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT107), .ZN(new_n916));
  INV_X1    g491(.A(new_n910), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n902), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n911), .A2(new_n915), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(KEYINPUT42), .ZN(new_n920));
  AND3_X1   g495(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n602), .A2(G651), .A3(new_n603), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n607), .B1(new_n922), .B2(new_n592), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n921), .B1(new_n923), .B2(new_n604), .ZN(new_n924));
  AND4_X1   g499(.A1(new_n921), .A2(new_n599), .A3(new_n604), .A4(new_n608), .ZN(new_n925));
  OAI21_X1  g500(.A(KEYINPUT108), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  AND3_X1   g501(.A1(new_n587), .A2(G166), .A3(new_n589), .ZN(new_n927));
  AOI21_X1  g502(.A(G166), .B1(new_n587), .B2(new_n589), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(G290), .A2(G288), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT108), .ZN(new_n931));
  NAND4_X1  g506(.A1(new_n921), .A2(new_n599), .A3(new_n604), .A4(new_n608), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n926), .A2(new_n929), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n930), .A2(new_n932), .ZN(new_n935));
  OAI211_X1 g510(.A(new_n935), .B(KEYINPUT108), .C1(new_n928), .C2(new_n927), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT42), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n911), .A2(new_n915), .A3(new_n939), .A4(new_n918), .ZN(new_n940));
  AND3_X1   g515(.A1(new_n920), .A2(new_n938), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n938), .B1(new_n920), .B2(new_n940), .ZN(new_n942));
  OAI21_X1  g517(.A(G868), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n872), .A2(new_n873), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n943), .B1(G868), .B2(new_n944), .ZN(G295));
  OAI21_X1  g520(.A(new_n943), .B1(G868), .B2(new_n944), .ZN(G331));
  INV_X1    g521(.A(KEYINPUT111), .ZN(new_n947));
  AND3_X1   g522(.A1(new_n871), .A2(G301), .A3(new_n874), .ZN(new_n948));
  AOI21_X1  g523(.A(G301), .B1(new_n871), .B2(new_n874), .ZN(new_n949));
  NOR3_X1   g524(.A1(new_n948), .A2(new_n949), .A3(G286), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n875), .A2(G171), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n871), .A2(G301), .A3(new_n874), .ZN(new_n952));
  AOI21_X1  g527(.A(G168), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n917), .B1(new_n950), .B2(new_n953), .ZN(new_n954));
  OAI21_X1  g529(.A(G286), .B1(new_n948), .B2(new_n949), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n951), .A2(G168), .A3(new_n952), .ZN(new_n956));
  OAI211_X1 g531(.A(new_n955), .B(new_n956), .C1(new_n913), .C2(new_n914), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n934), .A2(new_n954), .A3(new_n936), .A4(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(G37), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  AOI22_X1  g535(.A1(new_n934), .A2(new_n936), .B1(new_n954), .B2(new_n957), .ZN(new_n961));
  OAI21_X1  g536(.A(KEYINPUT43), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT109), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  OAI211_X1 g539(.A(KEYINPUT109), .B(KEYINPUT43), .C1(new_n960), .C2(new_n961), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n955), .A2(new_n956), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT110), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n904), .A2(new_n909), .A3(new_n912), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n914), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n913), .A2(KEYINPUT110), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n966), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(new_n954), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n937), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT43), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n973), .A2(new_n974), .A3(new_n959), .A4(new_n958), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n964), .A2(new_n965), .A3(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT44), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n974), .B1(new_n960), .B2(new_n961), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n973), .A2(KEYINPUT43), .A3(new_n959), .A4(new_n958), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n977), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n947), .B1(new_n978), .B2(new_n982), .ZN(new_n983));
  AOI211_X1 g558(.A(KEYINPUT111), .B(new_n981), .C1(new_n976), .C2(new_n977), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n983), .A2(new_n984), .ZN(G397));
  XNOR2_X1  g560(.A(new_n805), .B(G2067), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n986), .B1(G1996), .B2(new_n720), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT45), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n988), .B1(G164), .B2(G1384), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n473), .A2(G40), .A3(new_n476), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(new_n991), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n987), .A2(new_n992), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n992), .A2(G1996), .ZN(new_n994));
  XNOR2_X1  g569(.A(new_n994), .B(KEYINPUT113), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n993), .B1(new_n995), .B2(new_n721), .ZN(new_n996));
  INV_X1    g571(.A(new_n847), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n845), .A2(new_n997), .ZN(new_n998));
  AND2_X1   g573(.A1(new_n845), .A2(new_n997), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n991), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  AND2_X1   g575(.A1(new_n996), .A2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n835), .A2(new_n991), .A3(new_n838), .ZN(new_n1002));
  XOR2_X1   g577(.A(new_n1002), .B(KEYINPUT127), .Z(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(KEYINPUT48), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1001), .A2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n1003), .A2(KEYINPUT48), .ZN(new_n1006));
  INV_X1    g581(.A(G2067), .ZN(new_n1007));
  AOI22_X1  g582(.A1(new_n996), .A2(new_n998), .B1(new_n1007), .B2(new_n806), .ZN(new_n1008));
  OAI22_X1  g583(.A1(new_n1005), .A2(new_n1006), .B1(new_n992), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT47), .ZN(new_n1010));
  XOR2_X1   g585(.A(new_n995), .B(KEYINPUT46), .Z(new_n1011));
  INV_X1    g586(.A(KEYINPUT126), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n991), .B1(new_n720), .B2(new_n986), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1011), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1012), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1010), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1016), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1018), .A2(KEYINPUT47), .A3(new_n1014), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1009), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT124), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n493), .A2(new_n491), .ZN(new_n1022));
  INV_X1    g597(.A(new_n489), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(G1384), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n990), .B1(new_n1026), .B2(new_n988), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1024), .A2(KEYINPUT45), .A3(new_n1025), .ZN(new_n1028));
  AOI21_X1  g603(.A(G1966), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g604(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1030));
  AND3_X1   g605(.A1(new_n473), .A2(G40), .A3(new_n476), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT50), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1024), .A2(new_n1032), .A3(new_n1025), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n1030), .A2(new_n1031), .A3(new_n1033), .A4(new_n752), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1034), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1021), .B1(new_n1029), .B2(new_n1035), .ZN(new_n1036));
  AND3_X1   g611(.A1(new_n989), .A2(new_n1031), .A3(new_n1028), .ZN(new_n1037));
  OAI211_X1 g612(.A(KEYINPUT124), .B(new_n1034), .C1(new_n1037), .C2(G1966), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1036), .A2(new_n1038), .A3(G168), .ZN(new_n1039));
  AND2_X1   g614(.A1(KEYINPUT51), .A2(G8), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g616(.A(G8), .B1(new_n1029), .B2(new_n1035), .ZN(new_n1042));
  INV_X1    g617(.A(G8), .ZN(new_n1043));
  NOR2_X1   g618(.A1(G168), .A2(new_n1043), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n1044), .A2(KEYINPUT51), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1042), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1041), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1044), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1048), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n989), .A2(new_n1031), .A3(new_n1028), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1051), .A2(G2078), .ZN(new_n1052));
  INV_X1    g627(.A(G1961), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1030), .A2(new_n1031), .A3(new_n1033), .ZN(new_n1054));
  AOI22_X1  g629(.A1(new_n1052), .A2(KEYINPUT53), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT53), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1056), .B1(new_n1051), .B2(G2078), .ZN(new_n1057));
  AOI21_X1  g632(.A(G301), .B1(new_n1055), .B2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(G2078), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1037), .A2(KEYINPUT53), .A3(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1054), .A2(new_n1053), .ZN(new_n1061));
  AND4_X1   g636(.A1(G301), .A2(new_n1060), .A3(new_n1057), .A4(new_n1061), .ZN(new_n1062));
  OAI21_X1  g637(.A(KEYINPUT54), .B1(new_n1058), .B2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1055), .A2(G301), .A3(new_n1057), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1060), .A2(new_n1057), .A3(new_n1061), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(G171), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT54), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1064), .A2(new_n1066), .A3(new_n1067), .ZN(new_n1068));
  AOI22_X1  g643(.A1(new_n1047), .A2(new_n1050), .B1(new_n1063), .B2(new_n1068), .ZN(new_n1069));
  XNOR2_X1  g644(.A(KEYINPUT56), .B(G2072), .ZN(new_n1070));
  INV_X1    g645(.A(G1956), .ZN(new_n1071));
  AOI22_X1  g646(.A1(new_n1037), .A2(new_n1070), .B1(new_n1054), .B2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n554), .A2(new_n556), .ZN(new_n1073));
  AOI21_X1  g648(.A(KEYINPUT57), .B1(new_n1073), .B2(KEYINPUT122), .ZN(new_n1074));
  XNOR2_X1  g649(.A(G299), .B(new_n1074), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1072), .A2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(G1348), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1026), .A2(new_n990), .ZN(new_n1078));
  AOI22_X1  g653(.A1(new_n1054), .A2(new_n1077), .B1(new_n1078), .B2(new_n1007), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1079), .A2(new_n620), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT123), .ZN(new_n1082));
  AOI22_X1  g657(.A1(new_n1081), .A2(new_n1082), .B1(new_n1075), .B2(new_n1072), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1080), .A2(KEYINPUT123), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1076), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1072), .A2(new_n1075), .ZN(new_n1086));
  OR2_X1    g661(.A1(new_n1086), .A2(KEYINPUT61), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n620), .A2(KEYINPUT60), .ZN(new_n1088));
  AOI22_X1  g663(.A1(new_n1086), .A2(KEYINPUT61), .B1(new_n1079), .B2(new_n1088), .ZN(new_n1089));
  AND2_X1   g664(.A1(new_n1079), .A2(new_n620), .ZN(new_n1090));
  OAI21_X1  g665(.A(KEYINPUT60), .B1(new_n1090), .B2(new_n1080), .ZN(new_n1091));
  XNOR2_X1  g666(.A(KEYINPUT58), .B(G1341), .ZN(new_n1092));
  OAI22_X1  g667(.A1(new_n1051), .A2(G1996), .B1(new_n1078), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(new_n547), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(KEYINPUT59), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT59), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1093), .A2(new_n1096), .A3(new_n547), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1087), .A2(new_n1089), .A3(new_n1091), .A4(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1085), .A2(new_n1099), .ZN(new_n1100));
  NOR2_X1   g675(.A1(G166), .A2(new_n1043), .ZN(new_n1101));
  XNOR2_X1  g676(.A(KEYINPUT114), .B(KEYINPUT55), .ZN(new_n1102));
  XNOR2_X1  g677(.A(new_n1101), .B(new_n1102), .ZN(new_n1103));
  OAI22_X1  g678(.A1(new_n1037), .A2(G1971), .B1(new_n1054), .B2(G2090), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(G8), .ZN(new_n1105));
  XNOR2_X1  g680(.A(new_n1103), .B(new_n1105), .ZN(new_n1106));
  XNOR2_X1  g681(.A(KEYINPUT116), .B(G86), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n519), .A2(new_n507), .A3(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(new_n584), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1109), .A2(KEYINPUT117), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT117), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1108), .A2(new_n1111), .A3(new_n584), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1110), .A2(new_n577), .A3(new_n1112), .A4(new_n582), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(G1981), .ZN(new_n1114));
  INV_X1    g689(.A(G1981), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n577), .A2(new_n582), .A3(new_n585), .A4(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1114), .A2(KEYINPUT49), .A3(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT118), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT49), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1114), .A2(KEYINPUT118), .A3(KEYINPUT49), .A4(new_n1116), .ZN(new_n1123));
  OAI21_X1  g698(.A(G8), .B1(new_n1026), .B2(new_n990), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(KEYINPUT115), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT115), .ZN(new_n1126));
  OAI211_X1 g701(.A(new_n1126), .B(G8), .C1(new_n1026), .C2(new_n990), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1125), .A2(new_n1127), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1119), .A2(new_n1122), .A3(new_n1123), .A4(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n921), .A2(G1976), .ZN(new_n1131));
  INV_X1    g706(.A(G1976), .ZN(new_n1132));
  AOI21_X1  g707(.A(KEYINPUT52), .B1(G288), .B2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1128), .A2(new_n1131), .A3(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT52), .ZN(new_n1135));
  AOI22_X1  g710(.A1(new_n1125), .A2(new_n1127), .B1(G1976), .B2(new_n921), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1134), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  OAI21_X1  g712(.A(KEYINPUT119), .B1(new_n1130), .B2(new_n1137), .ZN(new_n1138));
  OR2_X1    g713(.A1(new_n1136), .A2(new_n1135), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT119), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1139), .A2(new_n1140), .A3(new_n1129), .A4(new_n1134), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1106), .B1(new_n1138), .B2(new_n1141), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1069), .A2(new_n1100), .A3(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n921), .A2(new_n1132), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1116), .B1(new_n1130), .B2(new_n1144), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1130), .A2(new_n1137), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1147));
  AOI22_X1  g722(.A1(new_n1145), .A2(new_n1128), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1049), .B1(new_n1041), .B2(new_n1046), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT62), .ZN(new_n1150));
  OAI21_X1  g725(.A(KEYINPUT125), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT125), .ZN(new_n1152));
  AOI22_X1  g727(.A1(new_n1039), .A2(new_n1040), .B1(new_n1042), .B2(new_n1045), .ZN(new_n1153));
  OAI211_X1 g728(.A(new_n1152), .B(KEYINPUT62), .C1(new_n1153), .C2(new_n1049), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1151), .A2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1047), .A2(new_n1050), .A3(new_n1150), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1138), .A2(new_n1141), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1106), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1156), .A2(new_n1157), .A3(new_n1158), .A4(new_n1058), .ZN(new_n1159));
  OAI211_X1 g734(.A(new_n1143), .B(new_n1148), .C1(new_n1155), .C2(new_n1159), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n1042), .A2(G286), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1157), .A2(new_n1158), .A3(new_n1161), .ZN(new_n1162));
  XOR2_X1   g737(.A(KEYINPUT120), .B(KEYINPUT63), .Z(new_n1163));
  AOI21_X1  g738(.A(KEYINPUT121), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  AND4_X1   g739(.A1(KEYINPUT63), .A2(new_n1158), .A3(new_n1146), .A4(new_n1161), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1162), .A2(KEYINPUT121), .A3(new_n1163), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1160), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g743(.A1(G290), .A2(G1986), .A3(new_n991), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1002), .A2(new_n1169), .ZN(new_n1170));
  XOR2_X1   g745(.A(new_n1170), .B(KEYINPUT112), .Z(new_n1171));
  NAND2_X1  g746(.A1(new_n1001), .A2(new_n1171), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1020), .B1(new_n1168), .B2(new_n1172), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g748(.A1(G401), .A2(new_n457), .A3(G227), .ZN(new_n1175));
  AND4_X1   g749(.A1(new_n712), .A2(new_n900), .A3(new_n976), .A4(new_n1175), .ZN(G308));
  NAND4_X1  g750(.A1(new_n712), .A2(new_n900), .A3(new_n976), .A4(new_n1175), .ZN(G225));
endmodule


