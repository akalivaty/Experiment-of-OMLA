//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 1 1 0 0 1 1 1 0 0 0 0 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 1 1 1 0 0 1 1 0 1 1 1 0 1 0 0 0 0 1 1 1 1 0 1 0 1 0 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:11 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1206, new_n1207,
    new_n1208, new_n1209, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1284, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G250), .ZN(new_n206));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT64), .ZN(new_n208));
  INV_X1    g0008(.A(G13), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(G257), .ZN(new_n211));
  INV_X1    g0011(.A(G264), .ZN(new_n212));
  AOI211_X1 g0012(.A(new_n206), .B(new_n210), .C1(new_n211), .C2(new_n212), .ZN(new_n213));
  OR2_X1    g0013(.A1(new_n213), .A2(KEYINPUT0), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  INV_X1    g0015(.A(G20), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(new_n201), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n218), .A2(G50), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(new_n213), .A2(KEYINPUT0), .B1(new_n217), .B2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n225));
  AND4_X1   g0025(.A1(new_n222), .A2(new_n223), .A3(new_n224), .A4(new_n225), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n226), .A2(new_n208), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT1), .ZN(new_n228));
  AND3_X1   g0028(.A1(new_n214), .A2(new_n221), .A3(new_n228), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT2), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G226), .ZN(new_n232));
  INV_X1    g0032(.A(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G250), .B(G257), .Z(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n234), .B(new_n237), .Z(G358));
  XNOR2_X1  g0038(.A(G50), .B(G58), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT65), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G68), .B(G77), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XOR2_X1   g0043(.A(G107), .B(G116), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  INV_X1    g0045(.A(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n242), .B(new_n246), .ZN(G351));
  NOR2_X1   g0047(.A1(new_n209), .A2(G1), .ZN(new_n248));
  INV_X1    g0048(.A(G68), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n248), .A2(G20), .A3(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n250), .B(KEYINPUT12), .ZN(new_n251));
  NAND3_X1  g0051(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(new_n215), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n254), .B1(G1), .B2(new_n216), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n251), .B1(new_n249), .B2(new_n255), .ZN(new_n256));
  NOR2_X1   g0056(.A1(G20), .A2(G33), .ZN(new_n257));
  AOI22_X1  g0057(.A1(new_n257), .A2(G50), .B1(G20), .B2(new_n249), .ZN(new_n258));
  INV_X1    g0058(.A(G77), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n216), .A2(G33), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n258), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  AND3_X1   g0061(.A1(new_n261), .A2(KEYINPUT11), .A3(new_n253), .ZN(new_n262));
  AOI21_X1  g0062(.A(KEYINPUT11), .B1(new_n261), .B2(new_n253), .ZN(new_n263));
  NOR3_X1   g0063(.A1(new_n256), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT68), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT13), .ZN(new_n267));
  INV_X1    g0067(.A(G1698), .ZN(new_n268));
  AND2_X1   g0068(.A1(KEYINPUT3), .A2(G33), .ZN(new_n269));
  NOR2_X1   g0069(.A1(KEYINPUT3), .A2(G33), .ZN(new_n270));
  OAI211_X1 g0070(.A(G226), .B(new_n268), .C1(new_n269), .C2(new_n270), .ZN(new_n271));
  OAI211_X1 g0071(.A(G232), .B(G1698), .C1(new_n269), .C2(new_n270), .ZN(new_n272));
  NAND2_X1  g0072(.A1(G33), .A2(G97), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n271), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n215), .B1(G33), .B2(G41), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT67), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n274), .A2(KEYINPUT67), .A3(new_n275), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G1), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n281), .B1(G41), .B2(G45), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  AND2_X1   g0083(.A1(new_n283), .A2(G274), .ZN(new_n284));
  INV_X1    g0084(.A(G33), .ZN(new_n285));
  INV_X1    g0085(.A(G41), .ZN(new_n286));
  OAI211_X1 g0086(.A(G1), .B(G13), .C1(new_n285), .C2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(new_n282), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n284), .B1(new_n289), .B2(G238), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n267), .B1(new_n280), .B2(new_n290), .ZN(new_n291));
  AND3_X1   g0091(.A1(new_n274), .A2(KEYINPUT67), .A3(new_n275), .ZN(new_n292));
  AOI21_X1  g0092(.A(KEYINPUT67), .B1(new_n274), .B2(new_n275), .ZN(new_n293));
  OAI211_X1 g0093(.A(new_n267), .B(new_n290), .C1(new_n292), .C2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  OAI21_X1  g0095(.A(G169), .B1(new_n291), .B2(new_n295), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n291), .A2(new_n295), .ZN(new_n297));
  AOI22_X1  g0097(.A1(new_n296), .A2(KEYINPUT14), .B1(new_n297), .B2(G179), .ZN(new_n298));
  INV_X1    g0098(.A(G169), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n290), .B1(new_n292), .B2(new_n293), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(KEYINPUT13), .ZN(new_n301));
  AOI211_X1 g0101(.A(KEYINPUT14), .B(new_n299), .C1(new_n301), .C2(new_n294), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n266), .B1(new_n298), .B2(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n301), .A2(G179), .A3(new_n294), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n299), .B1(new_n301), .B2(new_n294), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT14), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n305), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NOR3_X1   g0108(.A1(new_n308), .A2(KEYINPUT68), .A3(new_n302), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n265), .B1(new_n304), .B2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(G190), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n297), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(G200), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n313), .B1(new_n291), .B2(new_n295), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n265), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n310), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT71), .ZN(new_n318));
  XNOR2_X1  g0118(.A(KEYINPUT8), .B(G58), .ZN(new_n319));
  INV_X1    g0119(.A(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n255), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n281), .A2(G13), .A3(G20), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n319), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(KEYINPUT70), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT70), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n321), .A2(new_n326), .A3(new_n323), .ZN(new_n327));
  AND2_X1   g0127(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT3), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(new_n285), .ZN(new_n330));
  NAND2_X1  g0130(.A1(KEYINPUT3), .A2(G33), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n332), .A2(G223), .A3(new_n268), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n332), .A2(G226), .A3(G1698), .ZN(new_n334));
  NAND2_X1  g0134(.A1(G33), .A2(G87), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n333), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(new_n275), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n283), .A2(G274), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n338), .B1(new_n288), .B2(new_n233), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n337), .A2(new_n311), .A3(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n339), .B1(new_n336), .B2(new_n275), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n341), .B1(G200), .B2(new_n342), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n269), .A2(new_n270), .ZN(new_n344));
  AOI21_X1  g0144(.A(KEYINPUT7), .B1(new_n344), .B2(new_n216), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n330), .A2(KEYINPUT7), .A3(new_n216), .A4(new_n331), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  OAI21_X1  g0147(.A(G68), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(G58), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n349), .A2(new_n249), .ZN(new_n350));
  OAI21_X1  g0150(.A(G20), .B1(new_n350), .B2(new_n201), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n257), .A2(G159), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  AOI21_X1  g0154(.A(KEYINPUT16), .B1(new_n348), .B2(new_n354), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n348), .A2(KEYINPUT16), .A3(new_n354), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n355), .B1(KEYINPUT69), .B2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT16), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n330), .A2(new_n216), .A3(new_n331), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT7), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n249), .B1(new_n361), .B2(new_n346), .ZN(new_n362));
  OAI211_X1 g0162(.A(KEYINPUT69), .B(new_n358), .C1(new_n362), .C2(new_n353), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(new_n253), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n328), .B(new_n343), .C1(new_n357), .C2(new_n364), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n318), .B1(new_n365), .B2(KEYINPUT17), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n325), .A2(new_n327), .ZN(new_n367));
  AND2_X1   g0167(.A1(new_n363), .A2(new_n253), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n358), .B1(new_n362), .B2(new_n353), .ZN(new_n369));
  NOR3_X1   g0169(.A1(new_n362), .A2(new_n358), .A3(new_n353), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT69), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n369), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n367), .B1(new_n368), .B2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT17), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n373), .A2(KEYINPUT71), .A3(new_n374), .A4(new_n343), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n366), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n365), .A2(KEYINPUT17), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n328), .B1(new_n357), .B2(new_n364), .ZN(new_n379));
  XNOR2_X1  g0179(.A(KEYINPUT66), .B(G179), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n342), .A2(new_n380), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n381), .B1(G169), .B2(new_n342), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n379), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(KEYINPUT18), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n368), .A2(new_n372), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n382), .B1(new_n386), .B2(new_n328), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT18), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  AND2_X1   g0189(.A1(new_n385), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n378), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n322), .A2(new_n202), .ZN(new_n392));
  INV_X1    g0192(.A(new_n255), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n392), .B1(new_n393), .B2(new_n202), .ZN(new_n394));
  AOI22_X1  g0194(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n257), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n395), .B1(new_n260), .B2(new_n319), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(new_n253), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n394), .A2(new_n397), .ZN(new_n398));
  XNOR2_X1  g0198(.A(new_n398), .B(KEYINPUT9), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n344), .A2(G1698), .ZN(new_n400));
  AOI22_X1  g0200(.A1(new_n400), .A2(G222), .B1(G77), .B2(new_n344), .ZN(new_n401));
  INV_X1    g0201(.A(G223), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n332), .A2(G1698), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n401), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(new_n275), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n284), .B1(new_n289), .B2(G226), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(G200), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n405), .A2(G190), .A3(new_n406), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n399), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  XNOR2_X1  g0210(.A(new_n410), .B(KEYINPUT10), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n407), .A2(G169), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n412), .B1(new_n380), .B2(new_n407), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(new_n398), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n411), .A2(new_n414), .ZN(new_n415));
  AOI22_X1  g0215(.A1(new_n400), .A2(G232), .B1(G107), .B2(new_n344), .ZN(new_n416));
  INV_X1    g0216(.A(G238), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n416), .B1(new_n417), .B2(new_n403), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(new_n275), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n284), .B1(new_n289), .B2(G244), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n421), .A2(new_n380), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n299), .B1(new_n419), .B2(new_n420), .ZN(new_n423));
  OR2_X1    g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n322), .A2(G77), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n425), .B1(new_n393), .B2(G77), .ZN(new_n426));
  NAND2_X1  g0226(.A1(G20), .A2(G77), .ZN(new_n427));
  INV_X1    g0227(.A(new_n257), .ZN(new_n428));
  XNOR2_X1  g0228(.A(KEYINPUT15), .B(G87), .ZN(new_n429));
  OAI221_X1 g0229(.A(new_n427), .B1(new_n319), .B2(new_n428), .C1(new_n260), .C2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(new_n253), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n426), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n424), .A2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n432), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n421), .A2(G190), .ZN(new_n435));
  AOI21_X1  g0235(.A(G200), .B1(new_n419), .B2(new_n420), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n434), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n433), .A2(new_n437), .ZN(new_n438));
  NOR4_X1   g0238(.A1(new_n317), .A2(new_n391), .A3(new_n415), .A4(new_n438), .ZN(new_n439));
  OAI211_X1 g0239(.A(G250), .B(new_n268), .C1(new_n269), .C2(new_n270), .ZN(new_n440));
  OAI211_X1 g0240(.A(G257), .B(G1698), .C1(new_n269), .C2(new_n270), .ZN(new_n441));
  NAND2_X1  g0241(.A1(G33), .A2(G294), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n440), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n281), .A2(G45), .ZN(new_n444));
  OR2_X1    g0244(.A1(KEYINPUT5), .A2(G41), .ZN(new_n445));
  NAND2_X1  g0245(.A1(KEYINPUT5), .A2(G41), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n444), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n447), .A2(new_n275), .ZN(new_n448));
  AOI22_X1  g0248(.A1(new_n275), .A2(new_n443), .B1(new_n448), .B2(G264), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n447), .A2(G274), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n449), .A2(KEYINPUT81), .A3(G179), .A4(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT81), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n443), .A2(new_n275), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n445), .A2(new_n446), .ZN(new_n454));
  INV_X1    g0254(.A(new_n444), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n456), .A2(G264), .A3(new_n287), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n453), .A2(new_n457), .A3(new_n450), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n452), .B1(new_n458), .B2(G169), .ZN(new_n459));
  INV_X1    g0259(.A(G179), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n451), .B1(new_n459), .B2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT74), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n463), .B1(new_n285), .B2(G1), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n281), .A2(KEYINPUT74), .A3(G33), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n464), .A2(new_n322), .A3(new_n465), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n466), .A2(new_n253), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(G107), .ZN(new_n468));
  INV_X1    g0268(.A(G107), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n248), .A2(G20), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(KEYINPUT25), .ZN(new_n471));
  OR2_X1    g0271(.A1(new_n470), .A2(KEYINPUT25), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n468), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT23), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n474), .B1(new_n216), .B2(G107), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n469), .A2(KEYINPUT23), .A3(G20), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n216), .A2(G33), .A3(G116), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n216), .B(G87), .C1(new_n269), .C2(new_n270), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(KEYINPUT22), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT22), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n332), .A2(new_n482), .A3(new_n216), .A4(G87), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n479), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n254), .B1(new_n484), .B2(KEYINPUT24), .ZN(new_n485));
  INV_X1    g0285(.A(new_n479), .ZN(new_n486));
  AOI21_X1  g0286(.A(G20), .B1(new_n330), .B2(new_n331), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n482), .B1(new_n487), .B2(G87), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n480), .A2(KEYINPUT22), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n486), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT24), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n473), .B1(new_n485), .B2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n462), .A2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n458), .A2(new_n313), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n449), .A2(new_n311), .A3(new_n450), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(new_n493), .ZN(new_n500));
  INV_X1    g0300(.A(new_n500), .ZN(new_n501));
  OAI21_X1  g0301(.A(KEYINPUT82), .B1(new_n496), .B2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT82), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n495), .A2(new_n503), .A3(new_n500), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT19), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n216), .B1(new_n273), .B2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(G87), .ZN(new_n508));
  INV_X1    g0308(.A(G97), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n508), .A2(new_n509), .A3(new_n469), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n216), .B(G68), .C1(new_n269), .C2(new_n270), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n506), .B1(new_n273), .B2(G20), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n511), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(new_n322), .ZN(new_n515));
  AOI22_X1  g0315(.A1(new_n514), .A2(new_n253), .B1(new_n515), .B2(new_n429), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n467), .A2(G87), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n444), .A2(G250), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n281), .A2(G45), .A3(G274), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n275), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  OAI211_X1 g0320(.A(G244), .B(G1698), .C1(new_n269), .C2(new_n270), .ZN(new_n521));
  OAI211_X1 g0321(.A(G238), .B(new_n268), .C1(new_n269), .C2(new_n270), .ZN(new_n522));
  NAND2_X1  g0322(.A1(G33), .A2(G116), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n520), .B1(new_n524), .B2(new_n275), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n516), .B(new_n517), .C1(new_n525), .C2(new_n313), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT78), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n524), .A2(new_n275), .ZN(new_n528));
  INV_X1    g0328(.A(new_n520), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n527), .B1(new_n530), .B2(new_n311), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n525), .A2(KEYINPUT78), .A3(G190), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n526), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(new_n467), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n516), .B1(new_n429), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n530), .A2(new_n299), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n525), .A2(new_n380), .ZN(new_n537));
  AND3_X1   g0337(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  OAI21_X1  g0338(.A(KEYINPUT79), .B1(new_n533), .B2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT20), .ZN(new_n540));
  INV_X1    g0340(.A(G116), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n216), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(G33), .A2(G283), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n543), .B1(new_n509), .B2(G33), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n542), .B1(new_n544), .B2(new_n216), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n540), .B1(new_n545), .B2(new_n254), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n285), .A2(G97), .ZN(new_n547));
  AOI21_X1  g0347(.A(G20), .B1(new_n547), .B2(new_n543), .ZN(new_n548));
  OAI211_X1 g0348(.A(KEYINPUT20), .B(new_n253), .C1(new_n548), .C2(new_n542), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n322), .A2(new_n541), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n551), .B1(new_n467), .B2(new_n541), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n299), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  AOI22_X1  g0353(.A1(new_n448), .A2(G270), .B1(G274), .B2(new_n447), .ZN(new_n554));
  OAI211_X1 g0354(.A(G264), .B(G1698), .C1(new_n269), .C2(new_n270), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n330), .A2(G303), .A3(new_n331), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  OAI211_X1 g0357(.A(G257), .B(new_n268), .C1(new_n269), .C2(new_n270), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT80), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n332), .A2(KEYINPUT80), .A3(G257), .A4(new_n268), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n557), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n554), .B1(new_n562), .B2(new_n287), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n553), .A2(KEYINPUT21), .A3(new_n563), .ZN(new_n564));
  AND2_X1   g0364(.A1(new_n560), .A2(new_n561), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n275), .B1(new_n565), .B2(new_n557), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n550), .A2(new_n552), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n566), .A2(new_n567), .A3(G179), .A4(new_n554), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n564), .A2(new_n568), .ZN(new_n569));
  AOI21_X1  g0369(.A(KEYINPUT21), .B1(new_n553), .B2(new_n563), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT79), .ZN(new_n573));
  AND3_X1   g0373(.A1(new_n525), .A2(KEYINPUT78), .A3(G190), .ZN(new_n574));
  AOI21_X1  g0374(.A(KEYINPUT78), .B1(new_n525), .B2(G190), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n572), .B(new_n573), .C1(new_n576), .C2(new_n526), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n563), .A2(new_n313), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n578), .B1(G190), .B2(new_n563), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n579), .A2(new_n550), .A3(new_n552), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n539), .A2(new_n571), .A3(new_n577), .A4(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT75), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT73), .ZN(new_n583));
  AOI211_X1 g0383(.A(new_n583), .B(new_n469), .C1(new_n361), .C2(new_n346), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT6), .ZN(new_n585));
  XNOR2_X1  g0385(.A(G97), .B(G107), .ZN(new_n586));
  NAND2_X1  g0386(.A1(KEYINPUT6), .A2(G97), .ZN(new_n587));
  OAI21_X1  g0387(.A(KEYINPUT72), .B1(new_n587), .B2(G107), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT72), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n589), .A2(new_n469), .A3(KEYINPUT6), .A4(G97), .ZN(new_n590));
  AOI22_X1  g0390(.A1(new_n585), .A2(new_n586), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  OAI22_X1  g0391(.A1(new_n591), .A2(new_n216), .B1(new_n259), .B2(new_n428), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n584), .A2(new_n592), .ZN(new_n593));
  OAI21_X1  g0393(.A(G107), .B1(new_n345), .B2(new_n347), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n583), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n254), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n515), .A2(G97), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n597), .B1(new_n534), .B2(G97), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n582), .B1(new_n596), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n456), .A2(new_n287), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n450), .B1(new_n600), .B2(new_n211), .ZN(new_n601));
  NOR2_X1   g0401(.A1(KEYINPUT76), .A2(KEYINPUT4), .ZN(new_n602));
  INV_X1    g0402(.A(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n400), .A2(G244), .A3(new_n603), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n332), .A2(G244), .A3(new_n268), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(new_n602), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n332), .A2(G250), .A3(G1698), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n604), .A2(new_n606), .A3(new_n543), .A4(new_n607), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n601), .B1(new_n608), .B2(new_n275), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n311), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n610), .B1(new_n609), .B2(G200), .ZN(new_n611));
  OAI211_X1 g0411(.A(KEYINPUT73), .B(G107), .C1(new_n345), .C2(new_n347), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n586), .A2(new_n585), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n588), .A2(new_n590), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  AOI22_X1  g0415(.A1(new_n615), .A2(G20), .B1(G77), .B2(new_n257), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n595), .A2(new_n612), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(new_n253), .ZN(new_n618));
  INV_X1    g0418(.A(new_n598), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n618), .A2(KEYINPUT75), .A3(new_n619), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n599), .A2(new_n611), .A3(new_n620), .ZN(new_n621));
  OAI21_X1  g0421(.A(KEYINPUT77), .B1(new_n596), .B2(new_n598), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT77), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n618), .A2(new_n623), .A3(new_n619), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n543), .B(new_n607), .C1(new_n605), .C2(new_n602), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n603), .B1(new_n400), .B2(G244), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n275), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n601), .ZN(new_n628));
  AND3_X1   g0428(.A1(new_n627), .A2(new_n380), .A3(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(G169), .B1(new_n627), .B2(new_n628), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n622), .A2(new_n624), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n621), .A2(new_n632), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n581), .A2(new_n633), .ZN(new_n634));
  AND3_X1   g0434(.A1(new_n439), .A2(new_n505), .A3(new_n634), .ZN(G372));
  NAND2_X1  g0435(.A1(new_n539), .A2(new_n577), .ZN(new_n636));
  OAI21_X1  g0436(.A(KEYINPUT26), .B1(new_n636), .B2(new_n632), .ZN(new_n637));
  INV_X1    g0437(.A(new_n570), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n564), .A2(new_n568), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n495), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT83), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n520), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n518), .A2(new_n519), .ZN(new_n643));
  AND3_X1   g0443(.A1(new_n643), .A2(new_n641), .A3(new_n287), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n528), .B1(new_n642), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(G200), .ZN(new_n646));
  AND2_X1   g0446(.A1(new_n516), .A2(new_n517), .ZN(new_n647));
  OAI211_X1 g0447(.A(new_n646), .B(new_n647), .C1(new_n574), .C2(new_n575), .ZN(new_n648));
  INV_X1    g0448(.A(new_n645), .ZN(new_n649));
  OAI211_X1 g0449(.A(new_n537), .B(new_n535), .C1(new_n649), .C2(G169), .ZN(new_n650));
  AND3_X1   g0450(.A1(new_n500), .A2(new_n648), .A3(new_n650), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n640), .A2(new_n621), .A3(new_n651), .A4(new_n632), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n599), .A2(new_n620), .ZN(new_n653));
  AND2_X1   g0453(.A1(new_n648), .A2(new_n650), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT26), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n653), .A2(new_n654), .A3(new_n655), .A4(new_n631), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n637), .A2(new_n652), .A3(new_n650), .A4(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n439), .A2(new_n657), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n315), .A2(new_n433), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n298), .A2(new_n266), .A3(new_n303), .ZN(new_n660));
  OAI21_X1  g0460(.A(KEYINPUT68), .B1(new_n308), .B2(new_n302), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n659), .B1(new_n662), .B2(new_n265), .ZN(new_n663));
  AOI22_X1  g0463(.A1(new_n366), .A2(new_n375), .B1(KEYINPUT17), .B2(new_n365), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n390), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  AOI22_X1  g0465(.A1(new_n665), .A2(new_n411), .B1(new_n398), .B2(new_n413), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n658), .A2(new_n666), .ZN(G369));
  INV_X1    g0467(.A(new_n248), .ZN(new_n668));
  OR3_X1    g0468(.A1(new_n668), .A2(KEYINPUT27), .A3(G20), .ZN(new_n669));
  OAI21_X1  g0469(.A(KEYINPUT27), .B1(new_n668), .B2(G20), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n669), .A2(G213), .A3(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n672), .A2(KEYINPUT84), .A3(G343), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT84), .ZN(new_n674));
  INV_X1    g0474(.A(G343), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n674), .B1(new_n671), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n494), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g0478(.A(new_n678), .B(KEYINPUT86), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n505), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n496), .A2(new_n677), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n571), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n677), .A2(new_n567), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n571), .A2(new_n580), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n686), .B1(new_n687), .B2(new_n685), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(G330), .ZN(new_n689));
  OR2_X1    g0489(.A1(new_n689), .A2(KEYINPUT85), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(KEYINPUT85), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n683), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n571), .A2(new_n677), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n505), .A2(new_n679), .A3(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n677), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n696), .B1(new_n496), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n693), .A2(new_n698), .ZN(new_n699));
  XOR2_X1   g0499(.A(new_n699), .B(KEYINPUT87), .Z(G399));
  NOR2_X1   g0500(.A1(new_n210), .A2(G41), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n701), .A2(new_n281), .ZN(new_n702));
  NOR4_X1   g0502(.A1(G87), .A2(G97), .A3(G107), .A4(G116), .ZN(new_n703));
  AOI22_X1  g0503(.A1(new_n702), .A2(new_n703), .B1(new_n220), .B2(new_n701), .ZN(new_n704));
  XOR2_X1   g0504(.A(new_n704), .B(KEYINPUT28), .Z(new_n705));
  NAND3_X1  g0505(.A1(new_n609), .A2(new_n449), .A3(new_n525), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n566), .A2(G179), .A3(new_n554), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT30), .ZN(new_n708));
  OR3_X1    g0508(.A1(new_n706), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n609), .B1(new_n566), .B2(new_n554), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n710), .A2(new_n380), .A3(new_n458), .A4(new_n645), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n708), .B1(new_n706), .B2(new_n707), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n709), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n713), .A2(KEYINPUT31), .A3(new_n677), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT88), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n713), .A2(KEYINPUT88), .A3(KEYINPUT31), .A4(new_n677), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  OR2_X1    g0518(.A1(new_n713), .A2(KEYINPUT31), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT31), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n720), .B1(new_n634), .B2(new_n505), .ZN(new_n721));
  OAI211_X1 g0521(.A(new_n718), .B(new_n719), .C1(new_n721), .C2(new_n677), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(G330), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n632), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n725), .A2(new_n655), .A3(new_n577), .A4(new_n539), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n653), .A2(new_n654), .A3(new_n631), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(KEYINPUT26), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n726), .A2(new_n728), .A3(new_n650), .A4(new_n652), .ZN(new_n729));
  AND2_X1   g0529(.A1(new_n729), .A2(new_n697), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(KEYINPUT29), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n657), .A2(new_n697), .ZN(new_n732));
  XOR2_X1   g0532(.A(KEYINPUT89), .B(KEYINPUT29), .Z(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n724), .B1(new_n731), .B2(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n705), .B1(new_n735), .B2(G1), .ZN(G364));
  NAND2_X1  g0536(.A1(new_n690), .A2(new_n691), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n209), .A2(G20), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(G45), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n702), .A2(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n740), .B1(new_n688), .B2(G330), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n737), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g0542(.A(new_n742), .B(KEYINPUT90), .ZN(new_n743));
  INV_X1    g0543(.A(new_n210), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n744), .A2(G355), .A3(new_n332), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n745), .B1(G116), .B2(new_n744), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n242), .A2(G45), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n747), .B1(G45), .B2(new_n220), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n210), .A2(new_n332), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n746), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(G13), .A2(G33), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(G20), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n215), .B1(G20), .B2(new_n299), .ZN(new_n754));
  NOR3_X1   g0554(.A1(new_n750), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(new_n740), .ZN(new_n756));
  INV_X1    g0556(.A(new_n754), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n216), .A2(G190), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n313), .A2(G179), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(G283), .ZN(new_n761));
  INV_X1    g0561(.A(G303), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n759), .A2(G20), .A3(G190), .ZN(new_n763));
  OAI221_X1 g0563(.A(new_n344), .B1(new_n760), .B2(new_n761), .C1(new_n762), .C2(new_n763), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n758), .A2(new_n460), .A3(new_n313), .ZN(new_n765));
  INV_X1    g0565(.A(KEYINPUT91), .ZN(new_n766));
  OR2_X1    g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n765), .A2(new_n766), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR4_X1   g0570(.A1(new_n380), .A2(new_n216), .A3(new_n311), .A4(new_n313), .ZN(new_n771));
  AOI22_X1  g0571(.A1(new_n770), .A2(G329), .B1(G326), .B2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(G311), .ZN(new_n773));
  INV_X1    g0573(.A(new_n380), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(new_n758), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(G200), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n772), .B1(new_n773), .B2(new_n777), .ZN(new_n778));
  NOR3_X1   g0578(.A1(new_n311), .A2(G179), .A3(G200), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(new_n216), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  AOI211_X1 g0581(.A(new_n764), .B(new_n778), .C1(G294), .C2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n775), .A2(new_n313), .ZN(new_n783));
  XNOR2_X1  g0583(.A(KEYINPUT33), .B(G317), .ZN(new_n784));
  NOR4_X1   g0584(.A1(new_n380), .A2(new_n216), .A3(new_n311), .A4(G200), .ZN(new_n785));
  AOI22_X1  g0585(.A1(new_n783), .A2(new_n784), .B1(G322), .B2(new_n785), .ZN(new_n786));
  XNOR2_X1  g0586(.A(new_n786), .B(KEYINPUT92), .ZN(new_n787));
  INV_X1    g0587(.A(G159), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n769), .A2(new_n788), .ZN(new_n789));
  XNOR2_X1  g0589(.A(new_n789), .B(KEYINPUT32), .ZN(new_n790));
  AOI22_X1  g0590(.A1(new_n776), .A2(G77), .B1(G58), .B2(new_n785), .ZN(new_n791));
  INV_X1    g0591(.A(new_n771), .ZN(new_n792));
  INV_X1    g0592(.A(new_n783), .ZN(new_n793));
  OAI221_X1 g0593(.A(new_n791), .B1(new_n202), .B2(new_n792), .C1(new_n249), .C2(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n780), .A2(new_n509), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n760), .A2(new_n469), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n332), .B1(new_n763), .B2(new_n508), .ZN(new_n797));
  NOR4_X1   g0597(.A1(new_n794), .A2(new_n795), .A3(new_n796), .A4(new_n797), .ZN(new_n798));
  AOI22_X1  g0598(.A1(new_n782), .A2(new_n787), .B1(new_n790), .B2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n753), .ZN(new_n800));
  OAI221_X1 g0600(.A(new_n756), .B1(new_n757), .B2(new_n799), .C1(new_n688), .C2(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n743), .A2(new_n801), .ZN(G396));
  INV_X1    g0602(.A(new_n740), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n757), .A2(new_n752), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n803), .B1(G77), .B2(new_n804), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n777), .A2(new_n541), .B1(new_n762), .B2(new_n792), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n806), .B1(G283), .B2(new_n783), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n344), .B1(new_n763), .B2(new_n469), .ZN(new_n808));
  INV_X1    g0608(.A(new_n760), .ZN(new_n809));
  AOI211_X1 g0609(.A(new_n808), .B(new_n795), .C1(G87), .C2(new_n809), .ZN(new_n810));
  AOI22_X1  g0610(.A1(new_n770), .A2(G311), .B1(G294), .B2(new_n785), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n807), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n332), .B1(new_n780), .B2(new_n349), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n813), .B1(new_n770), .B2(G132), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n760), .A2(new_n249), .ZN(new_n815));
  INV_X1    g0615(.A(new_n763), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n815), .B1(G50), .B2(new_n816), .ZN(new_n817));
  XNOR2_X1  g0617(.A(new_n817), .B(KEYINPUT93), .ZN(new_n818));
  AOI22_X1  g0618(.A1(new_n776), .A2(G159), .B1(G137), .B2(new_n771), .ZN(new_n819));
  INV_X1    g0619(.A(G143), .ZN(new_n820));
  INV_X1    g0620(.A(new_n785), .ZN(new_n821));
  INV_X1    g0621(.A(G150), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n819), .B1(new_n820), .B2(new_n821), .C1(new_n822), .C2(new_n793), .ZN(new_n823));
  INV_X1    g0623(.A(KEYINPUT34), .ZN(new_n824));
  OAI211_X1 g0624(.A(new_n814), .B(new_n818), .C1(new_n823), .C2(new_n824), .ZN(new_n825));
  AND2_X1   g0625(.A1(new_n823), .A2(new_n824), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n812), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n805), .B1(new_n827), .B2(new_n754), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n828), .B(KEYINPUT94), .ZN(new_n829));
  OAI211_X1 g0629(.A(new_n432), .B(new_n697), .C1(new_n422), .C2(new_n423), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n437), .B1(new_n434), .B2(new_n697), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n831), .B1(new_n832), .B2(new_n433), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n829), .B1(new_n752), .B2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n833), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n732), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n657), .A2(new_n697), .A3(new_n833), .ZN(new_n837));
  AND2_X1   g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n740), .B1(new_n839), .B2(new_n723), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n840), .A2(KEYINPUT95), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n841), .B1(new_n724), .B2(new_n838), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n840), .A2(KEYINPUT95), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n834), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  XOR2_X1   g0644(.A(new_n844), .B(KEYINPUT96), .Z(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(G384));
  NAND2_X1  g0646(.A1(new_n265), .A2(new_n677), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n310), .A2(new_n316), .A3(new_n847), .ZN(new_n848));
  OAI211_X1 g0648(.A(new_n265), .B(new_n677), .C1(new_n662), .C2(new_n315), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  XOR2_X1   g0650(.A(new_n830), .B(KEYINPUT98), .Z(new_n851));
  NAND2_X1  g0651(.A1(new_n837), .A2(new_n851), .ZN(new_n852));
  AND3_X1   g0652(.A1(new_n850), .A2(new_n852), .A3(KEYINPUT99), .ZN(new_n853));
  AOI21_X1  g0653(.A(KEYINPUT99), .B1(new_n850), .B2(new_n852), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n369), .A2(new_n356), .A3(new_n253), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(new_n324), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(new_n672), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n385), .A2(new_n389), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n858), .B1(new_n664), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n379), .A2(new_n672), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT37), .ZN(new_n862));
  NAND4_X1  g0662(.A1(new_n384), .A2(new_n861), .A3(new_n862), .A4(new_n365), .ZN(new_n863));
  INV_X1    g0663(.A(new_n365), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n382), .A2(new_n671), .B1(new_n324), .B2(new_n855), .ZN(new_n865));
  OAI21_X1  g0665(.A(KEYINPUT37), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n863), .A2(new_n866), .ZN(new_n867));
  AND3_X1   g0667(.A1(new_n860), .A2(KEYINPUT38), .A3(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(KEYINPUT38), .B1(new_n860), .B2(new_n867), .ZN(new_n869));
  OAI22_X1  g0669(.A1(new_n853), .A2(new_n854), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n859), .A2(new_n671), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(KEYINPUT100), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n864), .A2(new_n387), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT101), .ZN(new_n875));
  NAND4_X1  g0675(.A1(new_n874), .A2(new_n875), .A3(new_n862), .A4(new_n861), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n863), .A2(KEYINPUT101), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n384), .A2(new_n861), .A3(new_n365), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(KEYINPUT37), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n876), .A2(new_n877), .A3(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n861), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n881), .B1(new_n664), .B2(new_n859), .ZN(new_n882));
  AOI21_X1  g0682(.A(KEYINPUT38), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n867), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n884), .B1(new_n391), .B2(new_n858), .ZN(new_n885));
  AOI22_X1  g0685(.A1(new_n883), .A2(KEYINPUT102), .B1(new_n885), .B2(KEYINPUT38), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n880), .A2(new_n882), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT38), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT102), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT39), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n886), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(KEYINPUT39), .B1(new_n868), .B2(new_n869), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(KEYINPUT103), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  NAND4_X1  g0696(.A1(new_n886), .A2(new_n891), .A3(KEYINPUT103), .A4(new_n892), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n310), .A2(new_n677), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT100), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n870), .A2(new_n901), .A3(new_n871), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n873), .A2(new_n900), .A3(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n439), .A2(new_n731), .A3(new_n734), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n666), .ZN(new_n905));
  XOR2_X1   g0705(.A(new_n905), .B(KEYINPUT104), .Z(new_n906));
  XNOR2_X1  g0706(.A(new_n903), .B(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n886), .A2(new_n891), .ZN(new_n908));
  OAI211_X1 g0708(.A(new_n719), .B(new_n714), .C1(new_n721), .C2(new_n677), .ZN(new_n909));
  AND2_X1   g0709(.A1(new_n909), .A2(new_n833), .ZN(new_n910));
  NAND4_X1  g0710(.A1(new_n908), .A2(KEYINPUT40), .A3(new_n850), .A4(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT40), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n850), .A2(new_n909), .A3(new_n833), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n868), .A2(new_n869), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n912), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n911), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n439), .A2(new_n909), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n916), .B(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(G330), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  OAI22_X1  g0720(.A1(new_n907), .A2(new_n920), .B1(new_n281), .B2(new_n738), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n921), .B1(new_n907), .B2(new_n920), .ZN(new_n922));
  OAI211_X1 g0722(.A(G116), .B(new_n217), .C1(new_n615), .C2(KEYINPUT35), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n923), .B1(KEYINPUT35), .B2(new_n615), .ZN(new_n924));
  XOR2_X1   g0724(.A(KEYINPUT97), .B(KEYINPUT36), .Z(new_n925));
  XNOR2_X1  g0725(.A(new_n924), .B(new_n925), .ZN(new_n926));
  OR3_X1    g0726(.A1(new_n219), .A2(new_n259), .A3(new_n350), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n202), .A2(G68), .ZN(new_n928));
  AOI211_X1 g0728(.A(new_n281), .B(G13), .C1(new_n927), .C2(new_n928), .ZN(new_n929));
  OR3_X1    g0729(.A1(new_n922), .A2(new_n926), .A3(new_n929), .ZN(G367));
  NAND2_X1  g0730(.A1(new_n653), .A2(new_n677), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n931), .A2(new_n621), .A3(new_n632), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n653), .A2(new_n631), .A3(new_n677), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  AND3_X1   g0734(.A1(new_n692), .A2(KEYINPUT106), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(KEYINPUT106), .B1(new_n692), .B2(new_n934), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n697), .A2(new_n647), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n654), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n938), .B1(new_n650), .B2(new_n937), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n939), .A2(KEYINPUT43), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n940), .B(KEYINPUT105), .ZN(new_n941));
  OR3_X1    g0741(.A1(new_n935), .A2(new_n936), .A3(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n941), .B1(new_n935), .B2(new_n936), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n495), .B1(new_n932), .B2(new_n933), .ZN(new_n945));
  OR2_X1    g0745(.A1(new_n945), .A2(new_n725), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n695), .B1(new_n932), .B2(new_n933), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT42), .ZN(new_n948));
  AOI22_X1  g0748(.A1(new_n697), .A2(new_n946), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  OR2_X1    g0749(.A1(new_n947), .A2(new_n948), .ZN(new_n950));
  AOI22_X1  g0750(.A1(new_n949), .A2(new_n950), .B1(KEYINPUT43), .B2(new_n939), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n944), .B(new_n951), .ZN(new_n952));
  XOR2_X1   g0752(.A(new_n701), .B(KEYINPUT41), .Z(new_n953));
  NAND2_X1  g0753(.A1(new_n698), .A2(new_n934), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n954), .B(KEYINPUT45), .ZN(new_n955));
  OR3_X1    g0755(.A1(new_n698), .A2(KEYINPUT44), .A3(new_n934), .ZN(new_n956));
  OAI21_X1  g0756(.A(KEYINPUT44), .B1(new_n698), .B2(new_n934), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  OR3_X1    g0758(.A1(new_n955), .A2(new_n958), .A3(new_n692), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n692), .B1(new_n955), .B2(new_n958), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n695), .B1(new_n682), .B2(new_n694), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n737), .B(new_n961), .ZN(new_n962));
  NAND4_X1  g0762(.A1(new_n959), .A2(new_n735), .A3(new_n960), .A4(new_n962), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n953), .B1(new_n963), .B2(new_n735), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n739), .A2(G1), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n952), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(new_n749), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n967), .A2(new_n237), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n753), .A2(new_n754), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n969), .B1(new_n744), .B2(new_n429), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n803), .B1(new_n968), .B2(new_n970), .ZN(new_n971));
  XOR2_X1   g0771(.A(KEYINPUT108), .B(G317), .Z(new_n972));
  AOI22_X1  g0772(.A1(new_n770), .A2(new_n972), .B1(G311), .B2(new_n771), .ZN(new_n973));
  INV_X1    g0773(.A(G294), .ZN(new_n974));
  OAI221_X1 g0774(.A(new_n973), .B1(new_n974), .B2(new_n793), .C1(new_n762), .C2(new_n821), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT46), .ZN(new_n976));
  NOR3_X1   g0776(.A1(new_n763), .A2(new_n976), .A3(new_n541), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n809), .A2(G97), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n976), .B1(new_n763), .B2(new_n541), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n978), .A2(new_n979), .A3(new_n344), .ZN(new_n980));
  NOR3_X1   g0780(.A1(new_n975), .A2(new_n977), .A3(new_n980), .ZN(new_n981));
  AOI22_X1  g0781(.A1(new_n776), .A2(G283), .B1(G107), .B2(new_n781), .ZN(new_n982));
  XOR2_X1   g0782(.A(new_n982), .B(KEYINPUT107), .Z(new_n983));
  NAND2_X1  g0783(.A1(new_n781), .A2(G68), .ZN(new_n984));
  OAI221_X1 g0784(.A(new_n984), .B1(new_n821), .B2(new_n822), .C1(new_n820), .C2(new_n792), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT109), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  AOI22_X1  g0787(.A1(new_n770), .A2(G137), .B1(new_n776), .B2(G50), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n760), .A2(new_n259), .ZN(new_n989));
  AOI211_X1 g0789(.A(new_n344), .B(new_n989), .C1(G58), .C2(new_n816), .ZN(new_n990));
  OAI211_X1 g0790(.A(new_n988), .B(new_n990), .C1(new_n788), .C2(new_n793), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n985), .A2(new_n986), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  AOI22_X1  g0793(.A1(new_n981), .A2(new_n983), .B1(new_n987), .B2(new_n993), .ZN(new_n994));
  OR2_X1    g0794(.A1(new_n994), .A2(KEYINPUT47), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n757), .B1(new_n994), .B2(KEYINPUT47), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n971), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n997), .B1(new_n800), .B2(new_n939), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n966), .A2(new_n998), .ZN(G387));
  INV_X1    g0799(.A(new_n701), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n1000), .B1(new_n962), .B2(new_n735), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1001), .B1(new_n735), .B2(new_n962), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n344), .B1(new_n760), .B2(new_n541), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(new_n781), .A2(G283), .B1(new_n816), .B2(G294), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n783), .A2(G311), .B1(new_n785), .B2(new_n972), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(new_n776), .A2(G303), .B1(G322), .B2(new_n771), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT48), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1004), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1009), .B1(new_n1008), .B2(new_n1007), .ZN(new_n1010));
  XOR2_X1   g0810(.A(KEYINPUT110), .B(KEYINPUT49), .Z(new_n1011));
  XNOR2_X1  g0811(.A(new_n1010), .B(new_n1011), .ZN(new_n1012));
  AOI211_X1 g0812(.A(new_n1003), .B(new_n1012), .C1(G326), .C2(new_n770), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n770), .A2(G150), .B1(new_n776), .B2(G68), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(new_n202), .B2(new_n821), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n429), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n781), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n816), .A2(G77), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n1017), .A2(new_n332), .A3(new_n978), .A4(new_n1018), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n793), .A2(new_n319), .B1(new_n788), .B2(new_n792), .ZN(new_n1020));
  NOR3_X1   g0820(.A1(new_n1015), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n754), .B1(new_n1013), .B2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n234), .A2(G45), .A3(new_n344), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n249), .A2(new_n259), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n320), .A2(KEYINPUT50), .A3(new_n202), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT50), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1026), .B1(new_n319), .B2(G50), .ZN(new_n1027));
  AOI211_X1 g0827(.A(G45), .B(new_n1024), .C1(new_n1025), .C2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n703), .B1(new_n1028), .B2(new_n332), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n210), .B1(new_n1023), .B2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n969), .B1(new_n744), .B2(new_n469), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n1022), .B(new_n803), .C1(new_n1030), .C2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1032), .B1(new_n683), .B2(new_n753), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1033), .B1(new_n962), .B2(new_n965), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1002), .A2(new_n1034), .ZN(G393));
  NOR2_X1   g0835(.A1(new_n246), .A2(new_n967), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n969), .B1(new_n744), .B2(new_n509), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n344), .B1(new_n760), .B2(new_n469), .C1(new_n761), .C2(new_n763), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n770), .A2(G322), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n1039), .B1(new_n974), .B2(new_n777), .C1(new_n762), .C2(new_n793), .ZN(new_n1040));
  AOI211_X1 g0840(.A(new_n1038), .B(new_n1040), .C1(G116), .C2(new_n781), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(G311), .A2(new_n785), .B1(new_n771), .B2(G317), .ZN(new_n1042));
  XOR2_X1   g0842(.A(new_n1042), .B(KEYINPUT52), .Z(new_n1043));
  AOI22_X1  g0843(.A1(G150), .A2(new_n771), .B1(new_n785), .B2(G159), .ZN(new_n1044));
  XOR2_X1   g0844(.A(new_n1044), .B(KEYINPUT51), .Z(new_n1045));
  AOI22_X1  g0845(.A1(new_n770), .A2(G143), .B1(new_n776), .B2(new_n320), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1046), .B1(new_n202), .B2(new_n793), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n780), .A2(new_n259), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n763), .A2(new_n249), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n332), .B1(new_n760), .B2(new_n508), .ZN(new_n1050));
  NOR4_X1   g0850(.A1(new_n1047), .A2(new_n1048), .A3(new_n1049), .A4(new_n1050), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n1041), .A2(new_n1043), .B1(new_n1045), .B2(new_n1051), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n803), .B1(new_n1036), .B2(new_n1037), .C1(new_n1052), .C2(new_n757), .ZN(new_n1053));
  XOR2_X1   g0853(.A(new_n1053), .B(KEYINPUT111), .Z(new_n1054));
  OAI21_X1  g0854(.A(new_n1054), .B1(new_n800), .B2(new_n934), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n959), .A2(new_n960), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n965), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1055), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  AND2_X1   g0858(.A1(new_n963), .A2(new_n701), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n962), .A2(new_n735), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1056), .A2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1058), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n1062), .ZN(G390));
  AOI22_X1  g0863(.A1(new_n848), .A2(new_n849), .B1(new_n837), .B2(new_n851), .ZN(new_n1064));
  OAI21_X1  g0864(.A(KEYINPUT112), .B1(new_n1064), .B2(new_n899), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n850), .A2(new_n852), .ZN(new_n1066));
  INV_X1    g0866(.A(KEYINPUT112), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n899), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1066), .A2(new_n1067), .A3(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1065), .A2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1070), .A2(new_n896), .A3(new_n897), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n850), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n851), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1073), .B1(new_n730), .B2(new_n833), .ZN(new_n1074));
  OAI211_X1 g0874(.A(new_n908), .B(new_n1068), .C1(new_n1072), .C2(new_n1074), .ZN(new_n1075));
  NAND4_X1  g0875(.A1(new_n722), .A2(new_n850), .A3(G330), .A4(new_n833), .ZN(new_n1076));
  AND3_X1   g0876(.A1(new_n1071), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1077));
  NAND4_X1  g0877(.A1(new_n850), .A2(new_n909), .A3(G330), .A4(new_n833), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1078), .B1(new_n1071), .B2(new_n1075), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n896), .A2(new_n751), .A3(new_n897), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n803), .B1(new_n320), .B2(new_n804), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n816), .A2(G150), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(new_n1083), .B(KEYINPUT53), .ZN(new_n1084));
  XNOR2_X1  g0884(.A(KEYINPUT54), .B(G143), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n777), .A2(new_n1085), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n1084), .B(new_n1086), .C1(G125), .C2(new_n770), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(G128), .A2(new_n771), .B1(new_n785), .B2(G132), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(new_n1088), .B(KEYINPUT113), .ZN(new_n1089));
  OAI221_X1 g0889(.A(new_n332), .B1(new_n760), .B2(new_n202), .C1(new_n780), .C2(new_n788), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(G137), .B2(new_n783), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1087), .A2(new_n1089), .A3(new_n1091), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(G97), .A2(new_n776), .B1(new_n783), .B2(G107), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1093), .B(KEYINPUT114), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n344), .B1(new_n763), .B2(new_n508), .ZN(new_n1095));
  NOR3_X1   g0895(.A1(new_n1048), .A2(new_n1095), .A3(new_n815), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n769), .A2(new_n974), .B1(new_n821), .B2(new_n541), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1097), .B1(G283), .B2(new_n771), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1094), .A2(new_n1096), .A3(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1092), .A2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1082), .B1(new_n1100), .B2(new_n754), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n1080), .A2(new_n965), .B1(new_n1081), .B2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n439), .A2(G330), .A3(new_n909), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n904), .A2(new_n1103), .A3(new_n666), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n850), .B1(new_n910), .B2(G330), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1076), .A2(new_n1074), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1107), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1072), .B1(new_n723), .B2(new_n835), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1109), .A2(new_n1078), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(new_n852), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1104), .B1(new_n1108), .B2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n701), .B1(new_n1080), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1104), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n1109), .A2(new_n1078), .B1(new_n837), .B2(new_n851), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1114), .B1(new_n1115), .B2(new_n1107), .ZN(new_n1116));
  NOR3_X1   g0916(.A1(new_n1077), .A2(new_n1079), .A3(new_n1116), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1102), .B1(new_n1113), .B2(new_n1117), .ZN(G378));
  INV_X1    g0918(.A(new_n908), .ZN(new_n1119));
  NAND4_X1  g0919(.A1(new_n850), .A2(new_n909), .A3(KEYINPUT40), .A4(new_n833), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n915), .B(G330), .C1(new_n1119), .C2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n398), .A2(new_n672), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(new_n415), .B(new_n1122), .ZN(new_n1123));
  XOR2_X1   g0923(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1124));
  XNOR2_X1  g0924(.A(new_n1123), .B(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1121), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1125), .ZN(new_n1127));
  NAND4_X1  g0927(.A1(new_n911), .A2(new_n1127), .A3(G330), .A4(new_n915), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1129));
  OR2_X1    g0929(.A1(new_n903), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n903), .A2(new_n1129), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1071), .A2(new_n1075), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1078), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1071), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1135), .A2(new_n1136), .A3(new_n1112), .ZN(new_n1137));
  AND3_X1   g0937(.A1(new_n1137), .A2(KEYINPUT117), .A3(new_n1114), .ZN(new_n1138));
  AOI21_X1  g0938(.A(KEYINPUT117), .B1(new_n1137), .B2(new_n1114), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1132), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n1140), .A2(KEYINPUT57), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT57), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT117), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1143), .B1(new_n1117), .B2(new_n1104), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1137), .A2(KEYINPUT117), .A3(new_n1114), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1142), .B1(new_n1146), .B2(new_n1132), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n701), .B1(new_n1141), .B2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1125), .A2(new_n751), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n803), .B1(G50), .B2(new_n804), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n780), .A2(new_n822), .B1(new_n763), .B2(new_n1085), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(new_n776), .A2(G137), .B1(G128), .B2(new_n785), .ZN(new_n1152));
  INV_X1    g0952(.A(G132), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1152), .B1(new_n1153), .B2(new_n793), .ZN(new_n1154));
  AOI211_X1 g0954(.A(new_n1151), .B(new_n1154), .C1(G125), .C2(new_n771), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT59), .ZN(new_n1156));
  OR2_X1    g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n285), .B(new_n286), .C1(new_n760), .C2(new_n788), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1159), .B1(new_n770), .B2(G124), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1157), .A2(new_n1158), .A3(new_n1160), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n332), .A2(G41), .ZN(new_n1162));
  AOI211_X1 g0962(.A(G50), .B(new_n1162), .C1(new_n285), .C2(new_n286), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(G97), .A2(new_n783), .B1(new_n776), .B2(new_n1016), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n770), .A2(G283), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n760), .A2(new_n349), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1166), .ZN(new_n1167));
  AND4_X1   g0967(.A1(new_n984), .A2(new_n1018), .A3(new_n1167), .A4(new_n1162), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(G107), .A2(new_n785), .B1(new_n771), .B2(G116), .ZN(new_n1169));
  NAND4_X1  g0969(.A1(new_n1164), .A2(new_n1165), .A3(new_n1168), .A4(new_n1169), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(KEYINPUT115), .B(KEYINPUT58), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1163), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n1161), .B(new_n1172), .C1(new_n1171), .C2(new_n1170), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(new_n1174));
  OR2_X1    g0974(.A1(new_n1174), .A2(KEYINPUT116), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n757), .B1(new_n1174), .B2(KEYINPUT116), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1150), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n1132), .A2(new_n965), .B1(new_n1149), .B2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1148), .A2(new_n1178), .ZN(G375));
  NOR2_X1   g0979(.A1(new_n1115), .A2(new_n1107), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n1180), .A2(new_n1057), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1072), .A2(new_n751), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n803), .B1(G68), .B2(new_n804), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(new_n770), .A2(G128), .B1(G132), .B2(new_n771), .ZN(new_n1184));
  AOI211_X1 g0984(.A(new_n344), .B(new_n1166), .C1(G159), .C2(new_n816), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n1184), .B(new_n1185), .C1(new_n202), .C2(new_n780), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n785), .A2(G137), .ZN(new_n1187));
  OAI221_X1 g0987(.A(new_n1187), .B1(new_n793), .B2(new_n1085), .C1(new_n822), .C2(new_n777), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(new_n770), .A2(G303), .B1(G294), .B2(new_n771), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1189), .B1(new_n541), .B2(new_n793), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n776), .A2(G107), .B1(G283), .B2(new_n785), .ZN(new_n1191));
  AOI211_X1 g0991(.A(new_n332), .B(new_n989), .C1(G97), .C2(new_n816), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1191), .A2(new_n1192), .A3(new_n1017), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n1186), .A2(new_n1188), .B1(new_n1190), .B2(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1183), .B1(new_n1194), .B2(new_n754), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1181), .B1(new_n1182), .B2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1180), .A2(new_n1104), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n953), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1197), .A2(new_n1198), .A3(new_n1116), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1196), .A2(new_n1199), .ZN(G381));
  NOR2_X1   g1000(.A1(G375), .A2(G378), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1062), .A2(new_n966), .A3(new_n998), .ZN(new_n1202));
  OR2_X1    g1002(.A1(G393), .A2(G396), .ZN(new_n1203));
  NOR4_X1   g1003(.A1(new_n1202), .A2(G384), .A3(G381), .A4(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1201), .A2(new_n1204), .ZN(G407));
  NAND2_X1  g1005(.A1(new_n675), .A2(G213), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1201), .A2(new_n1207), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(G407), .A2(new_n1208), .A3(G213), .ZN(new_n1209));
  XNOR2_X1  g1009(.A(new_n1209), .B(KEYINPUT118), .ZN(G409));
  INV_X1    g1010(.A(KEYINPUT61), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1148), .A2(G378), .A3(new_n1178), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT119), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n953), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1214), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1215), .A2(new_n1178), .ZN(new_n1216));
  INV_X1    g1016(.A(G378), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1213), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  AOI211_X1 g1018(.A(KEYINPUT119), .B(G378), .C1(new_n1215), .C2(new_n1178), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1207), .B1(new_n1212), .B2(new_n1220), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1180), .A2(KEYINPUT60), .A3(new_n1104), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT120), .ZN(new_n1223));
  XNOR2_X1  g1023(.A(new_n1222), .B(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT60), .ZN(new_n1225));
  AOI211_X1 g1025(.A(new_n1000), .B(new_n1112), .C1(new_n1225), .C2(new_n1197), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT121), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1224), .A2(new_n1226), .A3(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1228), .A2(new_n1196), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1227), .B1(new_n1224), .B2(new_n1226), .ZN(new_n1230));
  OAI21_X1  g1030(.A(G384), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1230), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n1232), .A2(new_n845), .A3(new_n1196), .A4(new_n1228), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1207), .A2(G2897), .ZN(new_n1234));
  AND3_X1   g1034(.A1(new_n1231), .A2(new_n1233), .A3(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1234), .B1(new_n1231), .B2(new_n1233), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1211), .B1(new_n1221), .B2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT124), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1231), .A2(new_n1233), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1140), .A2(KEYINPUT57), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1146), .A2(new_n1142), .A3(new_n1132), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1000), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1132), .A2(new_n965), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1149), .A2(new_n1177), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  NOR3_X1   g1047(.A1(new_n1244), .A2(new_n1217), .A3(new_n1247), .ZN(new_n1248));
  AND3_X1   g1048(.A1(new_n870), .A2(new_n901), .A3(new_n871), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n901), .B1(new_n870), .B2(new_n871), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(new_n1251), .A2(new_n900), .B1(new_n1126), .B2(new_n1128), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n903), .A2(new_n1129), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1198), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1254), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1217), .B1(new_n1247), .B2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1256), .A2(KEYINPUT119), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1216), .A2(new_n1213), .A3(new_n1217), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  OAI211_X1 g1059(.A(new_n1206), .B(new_n1241), .C1(new_n1248), .C2(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT62), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1221), .A2(KEYINPUT62), .A3(new_n1241), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  OAI211_X1 g1064(.A(KEYINPUT124), .B(new_n1211), .C1(new_n1221), .C2(new_n1237), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1240), .A2(new_n1264), .A3(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(G393), .A2(G396), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT122), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1202), .A2(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1062), .B1(new_n966), .B2(new_n998), .ZN(new_n1270));
  OAI211_X1 g1070(.A(new_n1203), .B(new_n1267), .C1(new_n1269), .C2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1270), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1203), .A2(new_n1267), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1272), .A2(new_n1268), .A3(new_n1202), .A4(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1271), .A2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1266), .A2(new_n1275), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1275), .A2(KEYINPUT61), .ZN(new_n1277));
  XNOR2_X1  g1077(.A(new_n1277), .B(KEYINPUT123), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1221), .A2(new_n1237), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT63), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1260), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  OAI211_X1 g1081(.A(new_n1278), .B(new_n1281), .C1(new_n1280), .C2(new_n1260), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1276), .A2(new_n1282), .ZN(G405));
  AOI21_X1  g1083(.A(KEYINPUT125), .B1(new_n1271), .B2(new_n1274), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1241), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1217), .B1(new_n1148), .B2(new_n1178), .ZN(new_n1286));
  OR3_X1    g1086(.A1(new_n1201), .A2(new_n1285), .A3(new_n1286), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1285), .B1(new_n1201), .B2(new_n1286), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1284), .B1(new_n1287), .B2(new_n1288), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1271), .A2(new_n1274), .A3(KEYINPUT125), .ZN(new_n1290));
  XOR2_X1   g1090(.A(new_n1290), .B(KEYINPUT126), .Z(new_n1291));
  XNOR2_X1  g1091(.A(new_n1289), .B(new_n1291), .ZN(G402));
endmodule


