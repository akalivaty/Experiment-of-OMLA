

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781;

  XNOR2_X1 U375 ( .A(n663), .B(n662), .ZN(n664) );
  XNOR2_X1 U376 ( .A(n670), .B(n669), .ZN(n671) );
  XNOR2_X1 U377 ( .A(n658), .B(KEYINPUT59), .ZN(n659) );
  AND2_X1 U378 ( .A1(n396), .A2(n393), .ZN(n364) );
  INV_X1 U379 ( .A(KEYINPUT32), .ZN(n355) );
  OR2_X1 U380 ( .A1(n585), .A2(n422), .ZN(n421) );
  XNOR2_X1 U381 ( .A(n354), .B(KEYINPUT107), .ZN(n704) );
  AND2_X1 U382 ( .A1(n701), .A2(n700), .ZN(n354) );
  XNOR2_X1 U383 ( .A(n443), .B(G116), .ZN(n403) );
  NAND2_X2 U384 ( .A1(n605), .A2(n700), .ZN(n514) );
  XNOR2_X1 U385 ( .A(n352), .B(n495), .ZN(n589) );
  NOR2_X2 U386 ( .A1(n585), .A2(n733), .ZN(n352) );
  NAND2_X1 U387 ( .A1(n353), .A2(n621), .ZN(n373) );
  NAND2_X1 U388 ( .A1(n679), .A2(n694), .ZN(n353) );
  AND2_X2 U389 ( .A1(n455), .A2(n453), .ZN(n452) );
  NAND2_X2 U390 ( .A1(n452), .A2(n449), .ZN(n774) );
  BUF_X2 U391 ( .A(n605), .Z(n643) );
  NAND2_X1 U392 ( .A1(n757), .A2(n767), .ZN(n738) );
  XNOR2_X2 U393 ( .A(n598), .B(KEYINPUT45), .ZN(n757) );
  NAND2_X1 U394 ( .A1(n778), .A2(n397), .ZN(n395) );
  XNOR2_X2 U395 ( .A(n356), .B(n355), .ZN(n778) );
  AND2_X4 U396 ( .A1(n438), .A2(n387), .ZN(n742) );
  NOR2_X2 U397 ( .A1(n774), .A2(n780), .ZN(n618) );
  NAND2_X1 U398 ( .A1(n594), .A2(n400), .ZN(n356) );
  XOR2_X1 U399 ( .A(G143), .B(G128), .Z(n501) );
  NAND2_X1 U400 ( .A1(n738), .A2(n737), .ZN(n739) );
  XOR2_X1 U401 ( .A(KEYINPUT38), .B(n643), .Z(n701) );
  XNOR2_X1 U402 ( .A(n470), .B(n522), .ZN(n670) );
  XNOR2_X1 U403 ( .A(n375), .B(KEYINPUT8), .ZN(n569) );
  XNOR2_X1 U404 ( .A(n501), .B(G134), .ZN(n573) );
  NOR2_X1 U405 ( .A1(G953), .A2(G237), .ZN(n549) );
  XNOR2_X1 U406 ( .A(KEYINPUT16), .B(G122), .ZN(n507) );
  XNOR2_X1 U407 ( .A(n632), .B(n515), .ZN(n357) );
  XNOR2_X1 U408 ( .A(n632), .B(n515), .ZN(n619) );
  AND2_X1 U409 ( .A1(n475), .A2(n473), .ZN(n472) );
  BUF_X2 U410 ( .A(n579), .Z(n585) );
  XNOR2_X1 U411 ( .A(G146), .B(G125), .ZN(n527) );
  OR2_X1 U412 ( .A1(G237), .A2(G902), .ZN(n511) );
  NOR2_X1 U413 ( .A1(n670), .A2(n414), .ZN(n413) );
  NAND2_X1 U414 ( .A1(n500), .A2(n415), .ZN(n414) );
  INV_X1 U415 ( .A(G902), .ZN(n415) );
  NAND2_X1 U416 ( .A1(n418), .A2(n417), .ZN(n416) );
  NAND2_X1 U417 ( .A1(G472), .A2(G902), .ZN(n417) );
  NAND2_X1 U418 ( .A1(n670), .A2(G472), .ZN(n418) );
  XNOR2_X1 U419 ( .A(n573), .B(n496), .ZN(n763) );
  XNOR2_X1 U420 ( .A(G131), .B(KEYINPUT4), .ZN(n496) );
  XNOR2_X1 U421 ( .A(n369), .B(n368), .ZN(n611) );
  INV_X1 U422 ( .A(G469), .ZN(n368) );
  OR2_X1 U423 ( .A1(n651), .A2(G902), .ZN(n369) );
  XNOR2_X1 U424 ( .A(n542), .B(n484), .ZN(n483) );
  NOR2_X1 U425 ( .A1(G902), .A2(n747), .ZN(n543) );
  INV_X1 U426 ( .A(KEYINPUT91), .ZN(n484) );
  OR2_X1 U427 ( .A1(n716), .A2(n611), .ZN(n604) );
  XNOR2_X1 U428 ( .A(n763), .B(G146), .ZN(n522) );
  XNOR2_X1 U429 ( .A(G119), .B(G113), .ZN(n493) );
  XOR2_X1 U430 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n506) );
  NOR2_X1 U431 ( .A1(n380), .A2(n378), .ZN(n447) );
  XNOR2_X1 U432 ( .A(n627), .B(n379), .ZN(n378) );
  NAND2_X1 U433 ( .A1(n637), .A2(n628), .ZN(n380) );
  INV_X1 U434 ( .A(KEYINPUT79), .ZN(n379) );
  AND2_X1 U435 ( .A1(n402), .A2(n676), .ZN(n401) );
  AND2_X1 U436 ( .A1(n395), .A2(n394), .ZN(n393) );
  NAND2_X1 U437 ( .A1(n392), .A2(n391), .ZN(n390) );
  XNOR2_X1 U438 ( .A(KEYINPUT15), .B(G902), .ZN(n647) );
  NAND2_X1 U439 ( .A1(G234), .A2(G237), .ZN(n516) );
  NOR2_X1 U440 ( .A1(n458), .A2(n620), .ZN(n457) );
  XNOR2_X1 U441 ( .A(KEYINPUT88), .B(n512), .ZN(n700) );
  XNOR2_X1 U442 ( .A(n383), .B(n382), .ZN(n716) );
  INV_X1 U443 ( .A(KEYINPUT67), .ZN(n382) );
  INV_X1 U444 ( .A(n577), .ZN(n482) );
  NAND2_X1 U445 ( .A1(n360), .A2(n609), .ZN(n377) );
  OR2_X1 U446 ( .A1(n410), .A2(n407), .ZN(n630) );
  NAND2_X1 U447 ( .A1(n409), .A2(n408), .ZN(n407) );
  NOR2_X1 U448 ( .A1(n416), .A2(n411), .ZN(n410) );
  XNOR2_X1 U449 ( .A(KEYINPUT64), .B(G953), .ZN(n504) );
  XNOR2_X1 U450 ( .A(n522), .B(n370), .ZN(n651) );
  XNOR2_X1 U451 ( .A(n526), .B(n359), .ZN(n370) );
  XNOR2_X1 U452 ( .A(n442), .B(n441), .ZN(n661) );
  XNOR2_X1 U453 ( .A(n750), .B(n362), .ZN(n442) );
  XNOR2_X1 U454 ( .A(n505), .B(n477), .ZN(n476) );
  NOR2_X1 U455 ( .A1(n463), .A2(KEYINPUT42), .ZN(n454) );
  XNOR2_X1 U456 ( .A(n606), .B(n494), .ZN(n466) );
  XNOR2_X1 U457 ( .A(n611), .B(n405), .ZN(n406) );
  INV_X1 U458 ( .A(KEYINPUT1), .ZN(n405) );
  INV_X1 U459 ( .A(n604), .ZN(n424) );
  XNOR2_X1 U460 ( .A(n762), .B(n538), .ZN(n747) );
  NAND2_X1 U461 ( .A1(n569), .A2(G221), .ZN(n536) );
  NAND2_X1 U462 ( .A1(n777), .A2(KEYINPUT44), .ZN(n402) );
  NOR2_X1 U463 ( .A1(n492), .A2(n596), .ZN(n397) );
  INV_X1 U464 ( .A(KEYINPUT0), .ZN(n474) );
  OR2_X1 U465 ( .A1(n521), .A2(n474), .ZN(n473) );
  NAND2_X1 U466 ( .A1(n412), .A2(KEYINPUT6), .ZN(n411) );
  INV_X1 U467 ( .A(n413), .ZN(n412) );
  NAND2_X1 U468 ( .A1(n416), .A2(n419), .ZN(n409) );
  XOR2_X1 U469 ( .A(G137), .B(G140), .Z(n530) );
  XOR2_X1 U470 ( .A(KEYINPUT12), .B(KEYINPUT96), .Z(n551) );
  XNOR2_X1 U471 ( .A(n553), .B(n552), .ZN(n554) );
  INV_X1 U472 ( .A(KEYINPUT11), .ZN(n552) );
  XNOR2_X1 U473 ( .A(G113), .B(G131), .ZN(n553) );
  XOR2_X1 U474 ( .A(G140), .B(G104), .Z(n548) );
  XNOR2_X1 U475 ( .A(G143), .B(G122), .ZN(n547) );
  XNOR2_X1 U476 ( .A(KEYINPUT10), .B(KEYINPUT68), .ZN(n529) );
  XNOR2_X1 U477 ( .A(n527), .B(KEYINPUT4), .ZN(n477) );
  XNOR2_X1 U478 ( .A(n501), .B(n506), .ZN(n425) );
  XOR2_X1 U479 ( .A(KEYINPUT74), .B(KEYINPUT75), .Z(n502) );
  XNOR2_X1 U480 ( .A(n446), .B(n445), .ZN(n444) );
  INV_X1 U481 ( .A(KEYINPUT48), .ZN(n445) );
  NAND2_X1 U482 ( .A1(n448), .A2(n447), .ZN(n446) );
  OR2_X1 U483 ( .A1(n704), .A2(n460), .ZN(n459) );
  NAND2_X1 U484 ( .A1(n461), .A2(n615), .ZN(n460) );
  INV_X1 U485 ( .A(n703), .ZN(n461) );
  XNOR2_X1 U486 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U487 ( .A(n562), .B(n437), .ZN(n588) );
  INV_X1 U488 ( .A(G475), .ZN(n437) );
  XNOR2_X1 U489 ( .A(G110), .B(KEYINPUT90), .ZN(n532) );
  XNOR2_X1 U490 ( .A(G119), .B(G128), .ZN(n531) );
  XNOR2_X1 U491 ( .A(KEYINPUT101), .B(KEYINPUT100), .ZN(n565) );
  XOR2_X1 U492 ( .A(KEYINPUT7), .B(KEYINPUT99), .Z(n566) );
  XNOR2_X1 U493 ( .A(G116), .B(G122), .ZN(n563) );
  XOR2_X1 U494 ( .A(KEYINPUT9), .B(G107), .Z(n564) );
  NOR2_X1 U495 ( .A1(n504), .A2(n376), .ZN(n375) );
  INV_X1 U496 ( .A(n647), .ZN(n433) );
  XNOR2_X1 U497 ( .A(n436), .B(n435), .ZN(n732) );
  INV_X1 U498 ( .A(KEYINPUT89), .ZN(n435) );
  NAND2_X1 U499 ( .A1(n363), .A2(n371), .ZN(n724) );
  INV_X1 U500 ( .A(n716), .ZN(n371) );
  NOR2_X1 U501 ( .A1(n604), .A2(n603), .ZN(n624) );
  XNOR2_X1 U502 ( .A(n469), .B(n468), .ZN(n467) );
  INV_X1 U503 ( .A(KEYINPUT30), .ZN(n468) );
  INV_X1 U504 ( .A(KEYINPUT19), .ZN(n515) );
  AND2_X1 U505 ( .A1(n714), .A2(n629), .ZN(n610) );
  XNOR2_X1 U506 ( .A(n499), .B(G137), .ZN(n404) );
  XNOR2_X1 U507 ( .A(n372), .B(G107), .ZN(n749) );
  XNOR2_X1 U508 ( .A(G104), .B(G110), .ZN(n372) );
  XNOR2_X1 U509 ( .A(n651), .B(n650), .ZN(n652) );
  NAND2_X1 U510 ( .A1(n451), .A2(n450), .ZN(n449) );
  AND2_X1 U511 ( .A1(n463), .A2(KEYINPUT42), .ZN(n450) );
  INV_X1 U512 ( .A(KEYINPUT40), .ZN(n616) );
  AND2_X1 U513 ( .A1(n593), .A2(n406), .ZN(n400) );
  NAND2_X1 U514 ( .A1(n426), .A2(n427), .ZN(n684) );
  AND2_X1 U515 ( .A1(n429), .A2(n608), .ZN(n428) );
  INV_X1 U516 ( .A(KEYINPUT95), .ZN(n420) );
  NAND2_X1 U517 ( .A1(n424), .A2(n423), .ZN(n422) );
  INV_X1 U518 ( .A(n710), .ZN(n389) );
  XNOR2_X1 U519 ( .A(n746), .B(n747), .ZN(n398) );
  INV_X1 U520 ( .A(KEYINPUT60), .ZN(n485) );
  AND2_X1 U521 ( .A1(n384), .A2(n399), .ZN(n741) );
  AND2_X1 U522 ( .A1(n740), .A2(n756), .ZN(n399) );
  OR2_X1 U523 ( .A1(n413), .A2(n416), .ZN(n714) );
  OR2_X1 U524 ( .A1(n423), .A2(KEYINPUT66), .ZN(n358) );
  XOR2_X1 U525 ( .A(n524), .B(n523), .Z(n359) );
  OR2_X1 U526 ( .A1(n602), .A2(n601), .ZN(n360) );
  XNOR2_X1 U527 ( .A(n543), .B(n483), .ZN(n591) );
  INV_X1 U528 ( .A(n591), .ZN(n608) );
  XNOR2_X1 U529 ( .A(KEYINPUT78), .B(n607), .ZN(n361) );
  XOR2_X1 U530 ( .A(n425), .B(n503), .Z(n362) );
  AND2_X1 U531 ( .A1(n406), .A2(n714), .ZN(n363) );
  NAND2_X1 U532 ( .A1(n521), .A2(n474), .ZN(n365) );
  INV_X1 U533 ( .A(n406), .ZN(n717) );
  AND2_X1 U534 ( .A1(n459), .A2(n462), .ZN(n366) );
  INV_X1 U535 ( .A(KEYINPUT6), .ZN(n419) );
  XNOR2_X1 U536 ( .A(KEYINPUT108), .B(KEYINPUT41), .ZN(n615) );
  OR2_X1 U537 ( .A1(n737), .A2(n645), .ZN(n367) );
  INV_X1 U538 ( .A(KEYINPUT42), .ZN(n464) );
  INV_X1 U539 ( .A(KEYINPUT65), .ZN(n492) );
  XNOR2_X1 U540 ( .A(n373), .B(KEYINPUT102), .ZN(n583) );
  XNOR2_X2 U541 ( .A(n421), .B(n420), .ZN(n679) );
  XNOR2_X1 U542 ( .A(n546), .B(KEYINPUT31), .ZN(n694) );
  INV_X1 U543 ( .A(n504), .ZN(n768) );
  INV_X1 U544 ( .A(G234), .ZN(n376) );
  NOR2_X1 U545 ( .A1(n591), .A2(n377), .ZN(n629) );
  NOR2_X2 U546 ( .A1(n381), .A2(n699), .ZN(n767) );
  NOR2_X1 U547 ( .A1(n381), .A2(n361), .ZN(n479) );
  NAND2_X1 U548 ( .A1(n444), .A2(n775), .ZN(n381) );
  NAND2_X1 U549 ( .A1(n591), .A2(n482), .ZN(n383) );
  XNOR2_X1 U550 ( .A(n385), .B(KEYINPUT80), .ZN(n384) );
  NAND2_X1 U551 ( .A1(n739), .A2(n387), .ZN(n385) );
  XNOR2_X2 U552 ( .A(n386), .B(n507), .ZN(n750) );
  XNOR2_X1 U553 ( .A(n386), .B(n404), .ZN(n470) );
  XNOR2_X2 U554 ( .A(n403), .B(n493), .ZN(n386) );
  XNOR2_X2 U555 ( .A(n478), .B(KEYINPUT72), .ZN(n387) );
  INV_X1 U556 ( .A(n388), .ZN(n430) );
  NAND2_X1 U557 ( .A1(n594), .A2(n717), .ZN(n388) );
  NAND2_X1 U558 ( .A1(n388), .A2(n590), .ZN(n432) );
  AND2_X1 U559 ( .A1(n430), .A2(n389), .ZN(n582) );
  NAND2_X1 U560 ( .A1(n684), .A2(n397), .ZN(n396) );
  NOR2_X1 U561 ( .A1(n684), .A2(n778), .ZN(n597) );
  NAND2_X1 U562 ( .A1(n364), .A2(n390), .ZN(n491) );
  NOR2_X1 U563 ( .A1(n778), .A2(KEYINPUT65), .ZN(n391) );
  INV_X1 U564 ( .A(n684), .ZN(n392) );
  NAND2_X1 U565 ( .A1(n492), .A2(n596), .ZN(n394) );
  NOR2_X1 U566 ( .A1(n398), .A2(n748), .ZN(G66) );
  NAND2_X1 U567 ( .A1(n439), .A2(n367), .ZN(n438) );
  NAND2_X1 U568 ( .A1(n430), .A2(n428), .ZN(n427) );
  NAND2_X1 U569 ( .A1(n401), .A2(n583), .ZN(n489) );
  NAND2_X1 U570 ( .A1(n406), .A2(n630), .ZN(n481) );
  NAND2_X1 U571 ( .A1(n413), .A2(n419), .ZN(n408) );
  INV_X1 U572 ( .A(n714), .ZN(n423) );
  NAND2_X1 U573 ( .A1(n431), .A2(n608), .ZN(n426) );
  NOR2_X1 U574 ( .A1(n714), .A2(n590), .ZN(n429) );
  NAND2_X1 U575 ( .A1(n432), .A2(n358), .ZN(n431) );
  NAND2_X1 U576 ( .A1(n434), .A2(n433), .ZN(n439) );
  INV_X1 U577 ( .A(n738), .ZN(n434) );
  NAND2_X1 U578 ( .A1(n518), .A2(G952), .ZN(n436) );
  NAND2_X1 U579 ( .A1(n661), .A2(n647), .ZN(n440) );
  NAND2_X1 U580 ( .A1(n742), .A2(G210), .ZN(n665) );
  NOR2_X1 U581 ( .A1(n658), .A2(G902), .ZN(n561) );
  NOR2_X1 U582 ( .A1(n588), .A2(n587), .ZN(n576) );
  XNOR2_X2 U583 ( .A(n440), .B(n510), .ZN(n605) );
  XNOR2_X1 U584 ( .A(n525), .B(n476), .ZN(n441) );
  XNOR2_X2 U585 ( .A(G101), .B(KEYINPUT3), .ZN(n443) );
  XNOR2_X1 U586 ( .A(n618), .B(KEYINPUT46), .ZN(n448) );
  NAND2_X1 U587 ( .A1(n704), .A2(n465), .ZN(n463) );
  INV_X1 U588 ( .A(n456), .ZN(n451) );
  INV_X1 U589 ( .A(n454), .ZN(n453) );
  NAND2_X1 U590 ( .A1(n456), .A2(n464), .ZN(n455) );
  NAND2_X1 U591 ( .A1(n366), .A2(n463), .ZN(n734) );
  NAND2_X1 U592 ( .A1(n459), .A2(n457), .ZN(n456) );
  INV_X1 U593 ( .A(n462), .ZN(n458) );
  NAND2_X1 U594 ( .A1(n703), .A2(n465), .ZN(n462) );
  INV_X1 U595 ( .A(n615), .ZN(n465) );
  NAND2_X1 U596 ( .A1(n466), .A2(n690), .ZN(n617) );
  NAND2_X1 U597 ( .A1(n466), .A2(n685), .ZN(n646) );
  NAND2_X1 U598 ( .A1(n467), .A2(n360), .ZN(n603) );
  NAND2_X1 U599 ( .A1(n714), .A2(n700), .ZN(n469) );
  NAND2_X1 U600 ( .A1(n472), .A2(n471), .ZN(n579) );
  OR2_X1 U601 ( .A1(n357), .A2(n365), .ZN(n471) );
  NAND2_X1 U602 ( .A1(n619), .A2(KEYINPUT0), .ZN(n475) );
  NAND2_X1 U603 ( .A1(n757), .A2(n479), .ZN(n478) );
  XNOR2_X2 U604 ( .A(n480), .B(KEYINPUT35), .ZN(n777) );
  NAND2_X1 U605 ( .A1(n589), .A2(n623), .ZN(n480) );
  NOR2_X1 U606 ( .A1(n716), .A2(n481), .ZN(n584) );
  XNOR2_X1 U607 ( .A(n486), .B(n485), .ZN(G60) );
  NAND2_X1 U608 ( .A1(n487), .A2(n673), .ZN(n486) );
  XNOR2_X1 U609 ( .A(n660), .B(n659), .ZN(n487) );
  NAND2_X1 U610 ( .A1(n491), .A2(n488), .ZN(n598) );
  NOR2_X1 U611 ( .A1(n490), .A2(n489), .ZN(n488) );
  AND2_X1 U612 ( .A1(n597), .A2(n595), .ZN(n490) );
  XNOR2_X1 U613 ( .A(KEYINPUT82), .B(KEYINPUT39), .ZN(n494) );
  XNOR2_X1 U614 ( .A(KEYINPUT34), .B(KEYINPUT76), .ZN(n495) );
  INV_X1 U615 ( .A(n697), .ZN(n637) );
  XNOR2_X1 U616 ( .A(n502), .B(KEYINPUT86), .ZN(n503) );
  XNOR2_X1 U617 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U618 ( .A(n498), .B(n497), .ZN(n499) );
  OR2_X1 U619 ( .A1(n703), .A2(n577), .ZN(n578) );
  XNOR2_X1 U620 ( .A(n541), .B(n540), .ZN(n542) );
  INV_X1 U621 ( .A(KEYINPUT66), .ZN(n590) );
  XNOR2_X1 U622 ( .A(n672), .B(n671), .ZN(n674) );
  XNOR2_X1 U623 ( .A(n665), .B(n664), .ZN(n666) );
  INV_X1 U624 ( .A(KEYINPUT122), .ZN(n656) );
  XNOR2_X1 U625 ( .A(n617), .B(n616), .ZN(n780) );
  XNOR2_X1 U626 ( .A(n657), .B(n656), .ZN(G54) );
  XOR2_X1 U627 ( .A(KEYINPUT94), .B(KEYINPUT5), .Z(n498) );
  NAND2_X1 U628 ( .A1(n549), .A2(G210), .ZN(n497) );
  INV_X1 U629 ( .A(G472), .ZN(n500) );
  NAND2_X1 U630 ( .A1(G224), .A2(n768), .ZN(n505) );
  XOR2_X1 U631 ( .A(KEYINPUT69), .B(n749), .Z(n525) );
  XOR2_X1 U632 ( .A(KEYINPUT77), .B(KEYINPUT87), .Z(n509) );
  NAND2_X1 U633 ( .A1(G210), .A2(n511), .ZN(n508) );
  NAND2_X1 U634 ( .A1(n511), .A2(G214), .ZN(n512) );
  INV_X1 U635 ( .A(KEYINPUT83), .ZN(n513) );
  XNOR2_X2 U636 ( .A(n514), .B(n513), .ZN(n632) );
  INV_X1 U637 ( .A(G953), .ZN(n756) );
  NOR2_X1 U638 ( .A1(G898), .A2(n756), .ZN(n752) );
  XOR2_X1 U639 ( .A(KEYINPUT71), .B(KEYINPUT14), .Z(n517) );
  XNOR2_X1 U640 ( .A(n517), .B(n516), .ZN(n518) );
  AND2_X1 U641 ( .A1(G902), .A2(n518), .ZN(n599) );
  NAND2_X1 U642 ( .A1(n752), .A2(n599), .ZN(n520) );
  NOR2_X1 U643 ( .A1(G953), .A2(n732), .ZN(n602) );
  INV_X1 U644 ( .A(n602), .ZN(n519) );
  NAND2_X1 U645 ( .A1(n520), .A2(n519), .ZN(n521) );
  XOR2_X1 U646 ( .A(G101), .B(n530), .Z(n524) );
  NAND2_X1 U647 ( .A1(G227), .A2(n768), .ZN(n523) );
  INV_X1 U648 ( .A(n525), .ZN(n526) );
  INV_X1 U649 ( .A(n527), .ZN(n528) );
  XOR2_X1 U650 ( .A(n529), .B(n528), .Z(n558) );
  XNOR2_X1 U651 ( .A(n530), .B(n558), .ZN(n762) );
  XNOR2_X1 U652 ( .A(n531), .B(KEYINPUT23), .ZN(n535) );
  XOR2_X1 U653 ( .A(KEYINPUT73), .B(KEYINPUT24), .Z(n533) );
  XNOR2_X1 U654 ( .A(n533), .B(n532), .ZN(n534) );
  XOR2_X1 U655 ( .A(n535), .B(n534), .Z(n537) );
  XNOR2_X1 U656 ( .A(n537), .B(n536), .ZN(n538) );
  NAND2_X1 U657 ( .A1(G234), .A2(n647), .ZN(n539) );
  XNOR2_X1 U658 ( .A(KEYINPUT20), .B(n539), .ZN(n544) );
  NAND2_X1 U659 ( .A1(G217), .A2(n544), .ZN(n541) );
  XNOR2_X1 U660 ( .A(KEYINPUT92), .B(KEYINPUT25), .ZN(n540) );
  NAND2_X1 U661 ( .A1(G221), .A2(n544), .ZN(n545) );
  XNOR2_X1 U662 ( .A(KEYINPUT21), .B(n545), .ZN(n709) );
  INV_X1 U663 ( .A(n709), .ZN(n609) );
  XNOR2_X1 U664 ( .A(KEYINPUT93), .B(n609), .ZN(n577) );
  NOR2_X1 U665 ( .A1(n585), .A2(n724), .ZN(n546) );
  XNOR2_X1 U666 ( .A(n548), .B(n547), .ZN(n557) );
  NAND2_X1 U667 ( .A1(G214), .A2(n549), .ZN(n550) );
  XNOR2_X1 U668 ( .A(n551), .B(n550), .ZN(n555) );
  XNOR2_X1 U669 ( .A(n557), .B(n556), .ZN(n559) );
  XNOR2_X1 U670 ( .A(n559), .B(n558), .ZN(n658) );
  XNOR2_X1 U671 ( .A(KEYINPUT97), .B(KEYINPUT13), .ZN(n560) );
  XNOR2_X1 U672 ( .A(n561), .B(n560), .ZN(n562) );
  XOR2_X1 U673 ( .A(KEYINPUT98), .B(n588), .Z(n575) );
  XNOR2_X1 U674 ( .A(n564), .B(n563), .ZN(n568) );
  XNOR2_X1 U675 ( .A(n566), .B(n565), .ZN(n567) );
  XOR2_X1 U676 ( .A(n568), .B(n567), .Z(n571) );
  NAND2_X1 U677 ( .A1(G217), .A2(n569), .ZN(n570) );
  XNOR2_X1 U678 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U679 ( .A(n573), .B(n572), .ZN(n744) );
  NOR2_X1 U680 ( .A1(n744), .A2(G902), .ZN(n574) );
  XOR2_X1 U681 ( .A(n574), .B(G478), .Z(n587) );
  NAND2_X1 U682 ( .A1(n575), .A2(n587), .ZN(n695) );
  INV_X1 U683 ( .A(n695), .ZN(n685) );
  NOR2_X1 U684 ( .A1(n575), .A2(n587), .ZN(n690) );
  NOR2_X1 U685 ( .A1(n685), .A2(n690), .ZN(n705) );
  INV_X1 U686 ( .A(n705), .ZN(n621) );
  XNOR2_X1 U687 ( .A(n608), .B(KEYINPUT104), .ZN(n710) );
  XNOR2_X1 U688 ( .A(n576), .B(KEYINPUT103), .ZN(n703) );
  NOR2_X1 U689 ( .A1(n579), .A2(n578), .ZN(n581) );
  XNOR2_X1 U690 ( .A(KEYINPUT22), .B(KEYINPUT70), .ZN(n580) );
  XNOR2_X1 U691 ( .A(n581), .B(n580), .ZN(n594) );
  INV_X1 U692 ( .A(n630), .ZN(n592) );
  NAND2_X1 U693 ( .A1(n582), .A2(n592), .ZN(n676) );
  XNOR2_X1 U694 ( .A(n584), .B(KEYINPUT33), .ZN(n733) );
  AND2_X1 U695 ( .A1(n588), .A2(n587), .ZN(n623) );
  NOR2_X1 U696 ( .A1(n777), .A2(KEYINPUT44), .ZN(n595) );
  AND2_X1 U697 ( .A1(n592), .A2(n710), .ZN(n593) );
  INV_X1 U698 ( .A(KEYINPUT44), .ZN(n596) );
  NAND2_X1 U699 ( .A1(n599), .A2(n504), .ZN(n600) );
  NOR2_X1 U700 ( .A1(G900), .A2(n600), .ZN(n601) );
  NAND2_X1 U701 ( .A1(n624), .A2(n701), .ZN(n606) );
  NAND2_X1 U702 ( .A1(KEYINPUT2), .A2(n646), .ZN(n607) );
  XNOR2_X1 U703 ( .A(KEYINPUT28), .B(n610), .ZN(n613) );
  INV_X1 U704 ( .A(n611), .ZN(n612) );
  NAND2_X1 U705 ( .A1(n613), .A2(n612), .ZN(n620) );
  NOR2_X1 U706 ( .A1(n620), .A2(n357), .ZN(n689) );
  NAND2_X1 U707 ( .A1(n689), .A2(n621), .ZN(n622) );
  OR2_X1 U708 ( .A1(KEYINPUT47), .A2(n622), .ZN(n628) );
  NAND2_X1 U709 ( .A1(n622), .A2(KEYINPUT47), .ZN(n626) );
  AND2_X1 U710 ( .A1(n624), .A2(n623), .ZN(n625) );
  NAND2_X1 U711 ( .A1(n643), .A2(n625), .ZN(n688) );
  NAND2_X1 U712 ( .A1(n626), .A2(n688), .ZN(n627) );
  XNOR2_X1 U713 ( .A(KEYINPUT109), .B(KEYINPUT36), .ZN(n635) );
  INV_X1 U714 ( .A(n690), .ZN(n692) );
  NAND2_X1 U715 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U716 ( .A1(n692), .A2(n631), .ZN(n639) );
  INV_X1 U717 ( .A(n639), .ZN(n633) );
  NOR2_X1 U718 ( .A1(n633), .A2(n632), .ZN(n634) );
  XNOR2_X1 U719 ( .A(n635), .B(n634), .ZN(n636) );
  NOR2_X1 U720 ( .A1(n717), .A2(n636), .ZN(n697) );
  AND2_X1 U721 ( .A1(n700), .A2(n717), .ZN(n638) );
  NAND2_X1 U722 ( .A1(n639), .A2(n638), .ZN(n640) );
  XNOR2_X1 U723 ( .A(KEYINPUT105), .B(n640), .ZN(n641) );
  XNOR2_X1 U724 ( .A(n641), .B(KEYINPUT43), .ZN(n642) );
  NOR2_X1 U725 ( .A1(n643), .A2(n642), .ZN(n644) );
  XOR2_X1 U726 ( .A(KEYINPUT106), .B(n644), .Z(n775) );
  INV_X1 U727 ( .A(KEYINPUT2), .ZN(n737) );
  XOR2_X1 U728 ( .A(KEYINPUT81), .B(n647), .Z(n645) );
  INV_X1 U729 ( .A(n646), .ZN(n699) );
  NAND2_X1 U730 ( .A1(n742), .A2(G469), .ZN(n653) );
  XOR2_X1 U731 ( .A(KEYINPUT121), .B(KEYINPUT120), .Z(n649) );
  XNOR2_X1 U732 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n648) );
  XNOR2_X1 U733 ( .A(n649), .B(n648), .ZN(n650) );
  XNOR2_X1 U734 ( .A(n653), .B(n652), .ZN(n655) );
  NOR2_X1 U735 ( .A1(n768), .A2(G952), .ZN(n654) );
  XOR2_X1 U736 ( .A(KEYINPUT85), .B(n654), .Z(n748) );
  INV_X1 U737 ( .A(n748), .ZN(n673) );
  NAND2_X1 U738 ( .A1(n655), .A2(n673), .ZN(n657) );
  NAND2_X1 U739 ( .A1(n742), .A2(G475), .ZN(n660) );
  XNOR2_X1 U740 ( .A(n661), .B(KEYINPUT55), .ZN(n663) );
  XOR2_X1 U741 ( .A(KEYINPUT118), .B(KEYINPUT54), .Z(n662) );
  NAND2_X1 U742 ( .A1(n666), .A2(n673), .ZN(n668) );
  XNOR2_X1 U743 ( .A(KEYINPUT119), .B(KEYINPUT56), .ZN(n667) );
  XNOR2_X1 U744 ( .A(n668), .B(n667), .ZN(G51) );
  NAND2_X1 U745 ( .A1(n742), .A2(G472), .ZN(n672) );
  XOR2_X1 U746 ( .A(KEYINPUT62), .B(KEYINPUT84), .Z(n669) );
  NAND2_X1 U747 ( .A1(n674), .A2(n673), .ZN(n675) );
  XNOR2_X1 U748 ( .A(n675), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U749 ( .A(G101), .B(n676), .ZN(G3) );
  NOR2_X1 U750 ( .A1(n692), .A2(n679), .ZN(n677) );
  XOR2_X1 U751 ( .A(KEYINPUT110), .B(n677), .Z(n678) );
  XNOR2_X1 U752 ( .A(G104), .B(n678), .ZN(G6) );
  NOR2_X1 U753 ( .A1(n679), .A2(n695), .ZN(n683) );
  XOR2_X1 U754 ( .A(KEYINPUT111), .B(KEYINPUT26), .Z(n681) );
  XNOR2_X1 U755 ( .A(G107), .B(KEYINPUT27), .ZN(n680) );
  XNOR2_X1 U756 ( .A(n681), .B(n680), .ZN(n682) );
  XNOR2_X1 U757 ( .A(n683), .B(n682), .ZN(G9) );
  XOR2_X1 U758 ( .A(n684), .B(G110), .Z(G12) );
  XOR2_X1 U759 ( .A(G128), .B(KEYINPUT29), .Z(n687) );
  NAND2_X1 U760 ( .A1(n689), .A2(n685), .ZN(n686) );
  XNOR2_X1 U761 ( .A(n687), .B(n686), .ZN(G30) );
  XNOR2_X1 U762 ( .A(G143), .B(n688), .ZN(G45) );
  NAND2_X1 U763 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U764 ( .A(G146), .B(n691), .ZN(G48) );
  NOR2_X1 U765 ( .A1(n692), .A2(n694), .ZN(n693) );
  XOR2_X1 U766 ( .A(G113), .B(n693), .Z(G15) );
  NOR2_X1 U767 ( .A1(n695), .A2(n694), .ZN(n696) );
  XOR2_X1 U768 ( .A(G116), .B(n696), .Z(G18) );
  XNOR2_X1 U769 ( .A(G125), .B(n697), .ZN(n698) );
  XNOR2_X1 U770 ( .A(n698), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U771 ( .A(G134), .B(n699), .Z(G36) );
  NOR2_X1 U772 ( .A1(n701), .A2(n700), .ZN(n702) );
  NOR2_X1 U773 ( .A1(n703), .A2(n702), .ZN(n707) );
  NOR2_X1 U774 ( .A1(n705), .A2(n704), .ZN(n706) );
  NOR2_X1 U775 ( .A1(n707), .A2(n706), .ZN(n708) );
  NOR2_X1 U776 ( .A1(n708), .A2(n733), .ZN(n729) );
  NAND2_X1 U777 ( .A1(n710), .A2(n709), .ZN(n713) );
  XNOR2_X1 U778 ( .A(KEYINPUT114), .B(KEYINPUT49), .ZN(n711) );
  XNOR2_X1 U779 ( .A(n711), .B(KEYINPUT113), .ZN(n712) );
  XNOR2_X1 U780 ( .A(n713), .B(n712), .ZN(n715) );
  NAND2_X1 U781 ( .A1(n715), .A2(n423), .ZN(n722) );
  XOR2_X1 U782 ( .A(KEYINPUT116), .B(KEYINPUT50), .Z(n719) );
  NAND2_X1 U783 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U784 ( .A(n719), .B(n718), .ZN(n720) );
  XOR2_X1 U785 ( .A(KEYINPUT115), .B(n720), .Z(n721) );
  NOR2_X1 U786 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U787 ( .A(n723), .B(KEYINPUT117), .ZN(n725) );
  NAND2_X1 U788 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U789 ( .A(KEYINPUT51), .B(n726), .ZN(n727) );
  NOR2_X1 U790 ( .A1(n734), .A2(n727), .ZN(n728) );
  NOR2_X1 U791 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U792 ( .A(n730), .B(KEYINPUT52), .ZN(n731) );
  NOR2_X1 U793 ( .A1(n732), .A2(n731), .ZN(n736) );
  NOR2_X1 U794 ( .A1(n734), .A2(n733), .ZN(n735) );
  NOR2_X1 U795 ( .A1(n736), .A2(n735), .ZN(n740) );
  XNOR2_X1 U796 ( .A(n741), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U797 ( .A1(G478), .A2(n742), .ZN(n743) );
  XNOR2_X1 U798 ( .A(n743), .B(n744), .ZN(n745) );
  NOR2_X1 U799 ( .A1(n748), .A2(n745), .ZN(G63) );
  NAND2_X1 U800 ( .A1(G217), .A2(n742), .ZN(n746) );
  XNOR2_X1 U801 ( .A(n750), .B(n749), .ZN(n751) );
  NOR2_X1 U802 ( .A1(n752), .A2(n751), .ZN(n761) );
  XOR2_X1 U803 ( .A(KEYINPUT61), .B(KEYINPUT123), .Z(n754) );
  NAND2_X1 U804 ( .A1(G224), .A2(G953), .ZN(n753) );
  XNOR2_X1 U805 ( .A(n754), .B(n753), .ZN(n755) );
  NAND2_X1 U806 ( .A1(n755), .A2(G898), .ZN(n759) );
  NAND2_X1 U807 ( .A1(n757), .A2(n756), .ZN(n758) );
  NAND2_X1 U808 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U809 ( .A(n761), .B(n760), .ZN(G69) );
  XNOR2_X1 U810 ( .A(n763), .B(n762), .ZN(n766) );
  XOR2_X1 U811 ( .A(G227), .B(n766), .Z(n764) );
  NAND2_X1 U812 ( .A1(n764), .A2(G900), .ZN(n765) );
  NAND2_X1 U813 ( .A1(n765), .A2(G953), .ZN(n771) );
  XNOR2_X1 U814 ( .A(n767), .B(n766), .ZN(n769) );
  NAND2_X1 U815 ( .A1(n769), .A2(n768), .ZN(n770) );
  NAND2_X1 U816 ( .A1(n771), .A2(n770), .ZN(n772) );
  XNOR2_X1 U817 ( .A(n772), .B(KEYINPUT124), .ZN(G72) );
  XOR2_X1 U818 ( .A(G137), .B(KEYINPUT126), .Z(n773) );
  XNOR2_X1 U819 ( .A(n774), .B(n773), .ZN(G39) );
  XNOR2_X1 U820 ( .A(G140), .B(n775), .ZN(n776) );
  XNOR2_X1 U821 ( .A(n776), .B(KEYINPUT112), .ZN(G42) );
  XOR2_X1 U822 ( .A(n777), .B(G122), .Z(G24) );
  XNOR2_X1 U823 ( .A(G119), .B(KEYINPUT125), .ZN(n779) );
  XNOR2_X1 U824 ( .A(n779), .B(n778), .ZN(G21) );
  XNOR2_X1 U825 ( .A(G131), .B(KEYINPUT127), .ZN(n781) );
  XNOR2_X1 U826 ( .A(n781), .B(n780), .ZN(G33) );
endmodule

