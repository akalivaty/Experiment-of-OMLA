//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 1 1 0 0 1 0 0 1 0 1 1 0 1 1 1 1 0 0 1 1 1 0 1 1 0 1 0 1 0 0 1 1 1 0 1 1 1 0 1 0 0 0 0 1 1 0 1 0 0 0 1 0 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:03 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1222, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1277, new_n1278, new_n1279, new_n1280, new_n1281,
    new_n1282, new_n1283, new_n1284;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  OAI21_X1  g0012(.A(G50), .B1(G58), .B2(G68), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n207), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  XNOR2_X1  g0017(.A(KEYINPUT64), .B(G238), .ZN(new_n218));
  INV_X1    g0018(.A(G68), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G107), .A2(G264), .ZN(new_n224));
  NAND4_X1  g0024(.A1(new_n221), .A2(new_n222), .A3(new_n223), .A4(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n209), .B1(new_n220), .B2(new_n225), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n212), .B(new_n217), .C1(KEYINPUT1), .C2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XOR2_X1   g0028(.A(G250), .B(G257), .Z(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT65), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G264), .B(G270), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  INV_X1    g0033(.A(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n232), .B(new_n237), .ZN(G358));
  XNOR2_X1  g0038(.A(G50), .B(G68), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G58), .B(G77), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n239), .B(new_n240), .Z(new_n241));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G351));
  INV_X1    g0045(.A(G274), .ZN(new_n246));
  INV_X1    g0046(.A(new_n215), .ZN(new_n247));
  NAND2_X1  g0047(.A1(G33), .A2(G41), .ZN(new_n248));
  AOI21_X1  g0048(.A(new_n246), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NOR2_X1   g0049(.A1(G41), .A2(G45), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n250), .A2(G1), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  OAI21_X1  g0052(.A(KEYINPUT66), .B1(new_n250), .B2(G1), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT66), .ZN(new_n254));
  OAI211_X1 g0054(.A(new_n254), .B(new_n206), .C1(G41), .C2(G45), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n248), .A2(G1), .A3(G13), .ZN(new_n256));
  AND3_X1   g0056(.A1(new_n253), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G226), .ZN(new_n258));
  OR2_X1    g0058(.A1(KEYINPUT3), .A2(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(KEYINPUT3), .A2(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n261), .A2(G223), .A3(G1698), .ZN(new_n262));
  INV_X1    g0062(.A(G77), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n262), .B1(new_n263), .B2(new_n261), .ZN(new_n264));
  AOI21_X1  g0064(.A(G1698), .B1(new_n259), .B2(new_n260), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n264), .B1(G222), .B2(new_n265), .ZN(new_n266));
  OAI211_X1 g0066(.A(new_n252), .B(new_n258), .C1(new_n266), .C2(new_n256), .ZN(new_n267));
  XNOR2_X1  g0067(.A(new_n267), .B(KEYINPUT67), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(G200), .ZN(new_n269));
  NAND3_X1  g0069(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(new_n215), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n271), .B1(new_n206), .B2(G20), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G50), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n203), .A2(G20), .ZN(new_n275));
  INV_X1    g0075(.A(G150), .ZN(new_n276));
  NOR2_X1   g0076(.A1(G20), .A2(G33), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n275), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  XNOR2_X1  g0079(.A(KEYINPUT8), .B(G58), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(KEYINPUT68), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT8), .ZN(new_n282));
  OR3_X1    g0082(.A1(new_n282), .A2(KEYINPUT68), .A3(G58), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n207), .A2(G33), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n279), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(new_n271), .ZN(new_n289));
  OAI221_X1 g0089(.A(new_n273), .B1(G50), .B2(new_n274), .C1(new_n288), .C2(new_n289), .ZN(new_n290));
  XNOR2_X1  g0090(.A(new_n290), .B(KEYINPUT9), .ZN(new_n291));
  INV_X1    g0091(.A(G190), .ZN(new_n292));
  OAI211_X1 g0092(.A(new_n269), .B(new_n291), .C1(new_n292), .C2(new_n268), .ZN(new_n293));
  XNOR2_X1  g0093(.A(new_n293), .B(KEYINPUT10), .ZN(new_n294));
  OR2_X1    g0094(.A1(new_n268), .A2(G179), .ZN(new_n295));
  INV_X1    g0095(.A(G169), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n268), .A2(new_n296), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n295), .A2(new_n290), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n294), .A2(new_n298), .ZN(new_n299));
  AND3_X1   g0099(.A1(KEYINPUT73), .A2(G58), .A3(G68), .ZN(new_n300));
  AOI21_X1  g0100(.A(KEYINPUT73), .B1(G58), .B2(G68), .ZN(new_n301));
  NOR3_X1   g0101(.A1(new_n300), .A2(new_n301), .A3(new_n201), .ZN(new_n302));
  INV_X1    g0102(.A(G159), .ZN(new_n303));
  OAI22_X1  g0103(.A1(new_n302), .A2(new_n207), .B1(new_n303), .B2(new_n278), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT74), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  OAI221_X1 g0106(.A(KEYINPUT74), .B1(new_n303), .B2(new_n278), .C1(new_n302), .C2(new_n207), .ZN(new_n307));
  AND2_X1   g0107(.A1(KEYINPUT3), .A2(G33), .ZN(new_n308));
  NOR2_X1   g0108(.A1(KEYINPUT3), .A2(G33), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  AOI21_X1  g0110(.A(KEYINPUT7), .B1(new_n310), .B2(new_n207), .ZN(new_n311));
  AND4_X1   g0111(.A1(KEYINPUT7), .A2(new_n259), .A3(new_n207), .A4(new_n260), .ZN(new_n312));
  OAI21_X1  g0112(.A(G68), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n306), .A2(new_n307), .A3(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT16), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND4_X1  g0116(.A1(new_n306), .A2(KEYINPUT16), .A3(new_n307), .A4(new_n313), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n316), .A2(new_n317), .A3(new_n271), .ZN(new_n318));
  NAND4_X1  g0118(.A1(new_n253), .A2(G232), .A3(new_n255), .A4(new_n256), .ZN(new_n319));
  NOR2_X1   g0119(.A1(G223), .A2(G1698), .ZN(new_n320));
  INV_X1    g0120(.A(G226), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n320), .B1(new_n321), .B2(G1698), .ZN(new_n322));
  AOI22_X1  g0122(.A1(new_n322), .A2(new_n261), .B1(G33), .B2(G87), .ZN(new_n323));
  OAI211_X1 g0123(.A(new_n319), .B(new_n252), .C1(new_n323), .C2(new_n256), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(G200), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n321), .A2(G1698), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n326), .B1(G223), .B2(G1698), .ZN(new_n327));
  INV_X1    g0127(.A(G33), .ZN(new_n328));
  INV_X1    g0128(.A(G87), .ZN(new_n329));
  OAI22_X1  g0129(.A1(new_n327), .A2(new_n310), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n256), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND4_X1  g0132(.A1(new_n332), .A2(G190), .A3(new_n319), .A4(new_n252), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n325), .A2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n284), .A2(new_n272), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n336), .B1(new_n284), .B2(new_n274), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n318), .A2(new_n335), .A3(new_n338), .ZN(new_n339));
  XNOR2_X1  g0139(.A(new_n339), .B(KEYINPUT17), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n324), .A2(new_n296), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n341), .B1(G179), .B2(new_n324), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n342), .B1(new_n318), .B2(new_n338), .ZN(new_n343));
  NOR2_X1   g0143(.A1(KEYINPUT75), .A2(KEYINPUT18), .ZN(new_n344));
  INV_X1    g0144(.A(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(KEYINPUT75), .A2(KEYINPUT18), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n289), .B1(new_n314), .B2(new_n315), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n337), .B1(new_n348), .B2(new_n317), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n344), .B1(new_n349), .B2(new_n342), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n346), .A2(new_n347), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n340), .A2(new_n351), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n277), .A2(G50), .B1(G20), .B2(new_n219), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n353), .B1(new_n263), .B2(new_n286), .ZN(new_n354));
  AND2_X1   g0154(.A1(new_n354), .A2(new_n271), .ZN(new_n355));
  OR2_X1    g0155(.A1(new_n355), .A2(KEYINPUT11), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(KEYINPUT11), .ZN(new_n357));
  OR3_X1    g0157(.A1(new_n274), .A2(KEYINPUT12), .A3(G68), .ZN(new_n358));
  OAI21_X1  g0158(.A(KEYINPUT12), .B1(new_n274), .B2(G68), .ZN(new_n359));
  AOI22_X1  g0159(.A1(G68), .A2(new_n272), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n356), .A2(new_n357), .A3(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT14), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n253), .A2(G238), .A3(new_n255), .A4(new_n256), .ZN(new_n363));
  NAND2_X1  g0163(.A1(G33), .A2(G97), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  NOR2_X1   g0165(.A1(G226), .A2(G1698), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n366), .B1(new_n234), .B2(G1698), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n365), .B1(new_n367), .B2(new_n261), .ZN(new_n368));
  OAI211_X1 g0168(.A(new_n252), .B(new_n363), .C1(new_n368), .C2(new_n256), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(KEYINPUT13), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n234), .A2(G1698), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n371), .B1(G226), .B2(G1698), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n364), .B1(new_n372), .B2(new_n310), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(new_n331), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT13), .ZN(new_n375));
  NAND4_X1  g0175(.A1(new_n374), .A2(new_n375), .A3(new_n252), .A4(new_n363), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n370), .A2(new_n376), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n362), .B1(new_n377), .B2(G169), .ZN(new_n378));
  AOI211_X1 g0178(.A(KEYINPUT14), .B(new_n296), .C1(new_n370), .C2(new_n376), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n370), .A2(G179), .A3(new_n376), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT71), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n370), .A2(new_n376), .A3(KEYINPUT71), .A4(G179), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  AND3_X1   g0185(.A1(new_n380), .A2(KEYINPUT72), .A3(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(KEYINPUT72), .B1(new_n380), .B2(new_n385), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n361), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  OR3_X1    g0188(.A1(new_n377), .A2(KEYINPUT70), .A3(new_n292), .ZN(new_n389));
  OAI21_X1  g0189(.A(KEYINPUT70), .B1(new_n377), .B2(new_n292), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n361), .B1(G200), .B2(new_n377), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n388), .A2(new_n393), .ZN(new_n394));
  XNOR2_X1  g0194(.A(KEYINPUT15), .B(G87), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n396), .A2(KEYINPUT69), .A3(new_n287), .ZN(new_n397));
  OAI221_X1 g0197(.A(new_n397), .B1(new_n207), .B2(new_n263), .C1(new_n278), .C2(new_n280), .ZN(new_n398));
  AOI21_X1  g0198(.A(KEYINPUT69), .B1(new_n396), .B2(new_n287), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n271), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n274), .A2(G77), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n401), .B1(new_n272), .B2(G77), .ZN(new_n402));
  AND2_X1   g0202(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n257), .A2(G244), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(new_n252), .ZN(new_n405));
  AOI22_X1  g0205(.A1(new_n265), .A2(G232), .B1(new_n310), .B2(G107), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n261), .A2(G1698), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n406), .B1(new_n218), .B2(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n405), .B1(new_n331), .B2(new_n408), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n409), .A2(G169), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n403), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(G179), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n409), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n409), .A2(G190), .ZN(new_n415));
  INV_X1    g0215(.A(G200), .ZN(new_n416));
  OAI211_X1 g0216(.A(new_n403), .B(new_n415), .C1(new_n416), .C2(new_n409), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n414), .A2(new_n417), .ZN(new_n418));
  NOR4_X1   g0218(.A1(new_n299), .A2(new_n352), .A3(new_n394), .A4(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(new_n274), .ZN(new_n421));
  INV_X1    g0221(.A(G107), .ZN(new_n422));
  AOI21_X1  g0222(.A(KEYINPUT25), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n421), .A2(KEYINPUT25), .A3(new_n422), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n274), .B1(G1), .B2(new_n328), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n426), .A2(new_n271), .ZN(new_n427));
  AOI22_X1  g0227(.A1(new_n424), .A2(new_n425), .B1(new_n427), .B2(G107), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT22), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT83), .ZN(new_n430));
  AOI21_X1  g0230(.A(G20), .B1(new_n259), .B2(new_n260), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n430), .B1(new_n431), .B2(G87), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n207), .B(G87), .C1(new_n308), .C2(new_n309), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n433), .A2(KEYINPUT83), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n429), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n431), .A2(new_n430), .A3(G87), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n433), .A2(KEYINPUT83), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n436), .A2(KEYINPUT22), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n287), .A2(G116), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT23), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n440), .A2(new_n422), .A3(G20), .ZN(new_n441));
  OAI21_X1  g0241(.A(KEYINPUT23), .B1(new_n207), .B2(G107), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n439), .A2(KEYINPUT84), .A3(new_n441), .A4(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(G116), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n442), .B(new_n441), .C1(new_n444), .C2(new_n286), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT84), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n443), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n435), .A2(new_n438), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(KEYINPUT24), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT24), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n435), .A2(new_n451), .A3(new_n438), .A4(new_n448), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(KEYINPUT85), .B1(new_n453), .B2(new_n271), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT85), .ZN(new_n455));
  AOI211_X1 g0255(.A(new_n455), .B(new_n289), .C1(new_n450), .C2(new_n452), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n428), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n261), .A2(G257), .A3(G1698), .ZN(new_n458));
  INV_X1    g0258(.A(G1698), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n261), .A2(G250), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(G33), .A2(G294), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n458), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(G45), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n463), .A2(G1), .ZN(new_n464));
  NOR2_X1   g0264(.A1(KEYINPUT5), .A2(G41), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(KEYINPUT5), .A2(G41), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n331), .B1(new_n464), .B2(new_n468), .ZN(new_n469));
  AOI22_X1  g0269(.A1(new_n462), .A2(new_n331), .B1(G264), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n256), .A2(G274), .ZN(new_n471));
  INV_X1    g0271(.A(new_n467), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n464), .B1(new_n472), .B2(new_n465), .ZN(new_n473));
  OAI21_X1  g0273(.A(KEYINPUT78), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT78), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n249), .A2(new_n468), .A3(new_n475), .A4(new_n464), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n470), .A2(new_n477), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n478), .A2(G179), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n479), .B1(new_n296), .B2(new_n478), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n457), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n478), .A2(new_n416), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n482), .B1(G190), .B2(new_n478), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n428), .B(new_n483), .C1(new_n454), .C2(new_n456), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT21), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n310), .A2(G303), .ZN(new_n486));
  OAI211_X1 g0286(.A(G264), .B(G1698), .C1(new_n308), .C2(new_n309), .ZN(new_n487));
  OAI211_X1 g0287(.A(G257), .B(new_n459), .C1(new_n308), .C2(new_n309), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n486), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT80), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n486), .A2(KEYINPUT80), .A3(new_n487), .A4(new_n488), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n256), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n469), .A2(G270), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n477), .A2(new_n494), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(G33), .A2(G283), .ZN(new_n497));
  INV_X1    g0297(.A(G97), .ZN(new_n498));
  OAI211_X1 g0298(.A(new_n497), .B(new_n207), .C1(G33), .C2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n444), .A2(G20), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n499), .A2(new_n271), .A3(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT20), .ZN(new_n502));
  XNOR2_X1  g0302(.A(new_n501), .B(new_n502), .ZN(new_n503));
  OR3_X1    g0303(.A1(new_n274), .A2(KEYINPUT81), .A3(G116), .ZN(new_n504));
  OAI21_X1  g0304(.A(KEYINPUT81), .B1(new_n274), .B2(G116), .ZN(new_n505));
  AOI22_X1  g0305(.A1(new_n427), .A2(G116), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(G169), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n485), .B1(new_n496), .B2(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n296), .B1(new_n503), .B2(new_n506), .ZN(new_n510));
  OAI211_X1 g0310(.A(new_n510), .B(KEYINPUT21), .C1(new_n493), .C2(new_n495), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n496), .A2(G179), .A3(new_n507), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n509), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(new_n507), .ZN(new_n514));
  OAI21_X1  g0314(.A(G200), .B1(new_n493), .B2(new_n495), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n491), .A2(new_n492), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(new_n331), .ZN(new_n517));
  INV_X1    g0317(.A(new_n495), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n514), .B(new_n515), .C1(new_n519), .C2(new_n292), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(KEYINPUT82), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n507), .B1(new_n496), .B2(G190), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT82), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n522), .A2(new_n523), .A3(new_n515), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n513), .B1(new_n521), .B2(new_n524), .ZN(new_n525));
  OAI211_X1 g0325(.A(G238), .B(new_n459), .C1(new_n308), .C2(new_n309), .ZN(new_n526));
  OAI211_X1 g0326(.A(G244), .B(G1698), .C1(new_n308), .C2(new_n309), .ZN(new_n527));
  NAND2_X1  g0327(.A1(G33), .A2(G116), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n331), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n256), .A2(G274), .A3(new_n464), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n206), .A2(G45), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n256), .A2(G250), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n530), .A2(new_n535), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n536), .A2(new_n292), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT19), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n207), .B1(new_n364), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g0339(.A1(G97), .A2(G107), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n329), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n207), .B(G68), .C1(new_n308), .C2(new_n309), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n538), .B1(new_n286), .B2(new_n498), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  AOI22_X1  g0345(.A1(new_n545), .A2(new_n271), .B1(new_n421), .B2(new_n395), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n427), .A2(G87), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n534), .B1(new_n331), .B2(new_n529), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n546), .B(new_n547), .C1(new_n548), .C2(new_n416), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n537), .B1(new_n549), .B2(KEYINPUT79), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n536), .A2(G200), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT79), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n551), .A2(new_n552), .A3(new_n546), .A4(new_n547), .ZN(new_n553));
  INV_X1    g0353(.A(new_n427), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n546), .B1(new_n395), .B2(new_n554), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n548), .A2(G169), .ZN(new_n556));
  AND3_X1   g0356(.A1(new_n530), .A2(new_n412), .A3(new_n535), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  AOI22_X1  g0358(.A1(new_n550), .A2(new_n553), .B1(new_n555), .B2(new_n558), .ZN(new_n559));
  AND2_X1   g0359(.A1(G97), .A2(G107), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT76), .ZN(new_n561));
  OAI22_X1  g0361(.A1(new_n560), .A2(new_n540), .B1(new_n561), .B2(KEYINPUT6), .ZN(new_n562));
  MUX2_X1   g0362(.A(new_n561), .B(G97), .S(KEYINPUT6), .Z(new_n563));
  XNOR2_X1  g0363(.A(G97), .B(G107), .ZN(new_n564));
  OAI211_X1 g0364(.A(G20), .B(new_n562), .C1(new_n563), .C2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n277), .A2(G77), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n565), .A2(KEYINPUT77), .A3(new_n566), .ZN(new_n567));
  OAI21_X1  g0367(.A(G107), .B1(new_n311), .B2(new_n312), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  AOI21_X1  g0369(.A(KEYINPUT77), .B1(new_n565), .B2(new_n566), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n271), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n274), .A2(G97), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n572), .B1(new_n427), .B2(G97), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  AOI22_X1  g0374(.A1(new_n474), .A2(new_n476), .B1(new_n469), .B2(G257), .ZN(new_n575));
  OAI211_X1 g0375(.A(G250), .B(G1698), .C1(new_n308), .C2(new_n309), .ZN(new_n576));
  OAI211_X1 g0376(.A(G244), .B(new_n459), .C1(new_n308), .C2(new_n309), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT4), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n497), .B(new_n576), .C1(new_n577), .C2(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(KEYINPUT4), .B1(new_n265), .B2(G244), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n331), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n575), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n296), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n575), .A2(new_n412), .A3(new_n581), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n574), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(new_n573), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n565), .A2(new_n566), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT77), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n589), .A2(new_n568), .A3(new_n567), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n586), .B1(new_n590), .B2(new_n271), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n582), .A2(G200), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n575), .A2(G190), .A3(new_n581), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  AND3_X1   g0394(.A1(new_n559), .A2(new_n585), .A3(new_n594), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n481), .A2(new_n484), .A3(new_n525), .A4(new_n595), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n420), .A2(new_n596), .ZN(G372));
  INV_X1    g0397(.A(new_n294), .ZN(new_n598));
  AOI211_X1 g0398(.A(new_n337), .B(new_n334), .C1(new_n348), .C2(new_n317), .ZN(new_n599));
  XNOR2_X1  g0399(.A(new_n599), .B(KEYINPUT17), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n393), .A2(new_n413), .A3(new_n411), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n600), .B1(new_n388), .B2(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT18), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT88), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n318), .A2(new_n338), .ZN(new_n605));
  INV_X1    g0405(.A(new_n342), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n604), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NOR3_X1   g0407(.A1(new_n349), .A2(KEYINPUT88), .A3(new_n342), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n603), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n343), .A2(new_n604), .ZN(new_n610));
  OAI21_X1  g0410(.A(KEYINPUT88), .B1(new_n349), .B2(new_n342), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n610), .A2(KEYINPUT18), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n609), .A2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(new_n613), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n602), .A2(new_n614), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n298), .B1(new_n598), .B2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT89), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  OAI211_X1 g0418(.A(KEYINPUT89), .B(new_n298), .C1(new_n598), .C2(new_n615), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n536), .A2(new_n296), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n548), .A2(new_n412), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n555), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n583), .A2(new_n584), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n625), .A2(new_n591), .ZN(new_n626));
  XNOR2_X1  g0426(.A(KEYINPUT86), .B(KEYINPUT26), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n559), .A2(new_n626), .A3(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT26), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n623), .B1(new_n549), .B2(new_n537), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n630), .B1(new_n585), .B2(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n624), .B1(new_n629), .B2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT87), .ZN(new_n634));
  OR2_X1    g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(new_n513), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n481), .A2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n549), .ZN(new_n638));
  INV_X1    g0438(.A(new_n537), .ZN(new_n639));
  AOI22_X1  g0439(.A1(new_n555), .A2(new_n558), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  AND3_X1   g0440(.A1(new_n640), .A2(new_n585), .A3(new_n594), .ZN(new_n641));
  AND2_X1   g0441(.A1(new_n484), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n637), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n633), .A2(new_n634), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n635), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n419), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n620), .A2(new_n646), .ZN(G369));
  INV_X1    g0447(.A(G13), .ZN(new_n648));
  NOR3_X1   g0448(.A1(new_n648), .A2(G1), .A3(G20), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  AND3_X1   g0450(.A1(new_n650), .A2(KEYINPUT90), .A3(KEYINPUT27), .ZN(new_n651));
  AOI21_X1  g0451(.A(KEYINPUT90), .B1(new_n650), .B2(KEYINPUT27), .ZN(new_n652));
  OAI221_X1 g0452(.A(G213), .B1(KEYINPUT27), .B2(new_n650), .C1(new_n651), .C2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(G343), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(new_n507), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n525), .A2(new_n656), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n657), .B1(new_n636), .B2(new_n656), .ZN(new_n658));
  XOR2_X1   g0458(.A(KEYINPUT91), .B(G330), .Z(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n481), .A2(new_n484), .ZN(new_n663));
  AND2_X1   g0463(.A1(new_n457), .A2(new_n655), .ZN(new_n664));
  INV_X1    g0464(.A(new_n655), .ZN(new_n665));
  OAI22_X1  g0465(.A1(new_n663), .A2(new_n664), .B1(new_n481), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n662), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n457), .A2(new_n480), .A3(new_n665), .ZN(new_n668));
  INV_X1    g0468(.A(new_n663), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n636), .A2(new_n655), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n667), .A2(new_n668), .A3(new_n671), .ZN(G399));
  INV_X1    g0472(.A(new_n210), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n673), .A2(G41), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n541), .A2(G116), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n675), .A2(G1), .A3(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n677), .B1(new_n213), .B2(new_n675), .ZN(new_n678));
  XNOR2_X1  g0478(.A(new_n678), .B(KEYINPUT28), .ZN(new_n679));
  AOI211_X1 g0479(.A(KEYINPUT92), .B(KEYINPUT29), .C1(new_n645), .C2(new_n665), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT94), .ZN(new_n681));
  XNOR2_X1  g0481(.A(new_n623), .B(KEYINPUT93), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n628), .B1(new_n559), .B2(new_n626), .ZN(new_n684));
  NOR3_X1   g0484(.A1(new_n585), .A2(new_n631), .A3(new_n630), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n683), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n686), .B1(new_n637), .B2(new_n642), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n681), .B1(new_n687), .B2(new_n655), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n513), .B1(new_n457), .B2(new_n480), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n484), .A2(new_n641), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  OAI211_X1 g0491(.A(KEYINPUT94), .B(new_n665), .C1(new_n691), .C2(new_n686), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n688), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(KEYINPUT29), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT92), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n645), .A2(new_n665), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT29), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n695), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n680), .B1(new_n694), .B2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT30), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n517), .A2(G179), .A3(new_n518), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n470), .A2(new_n575), .A3(new_n548), .A4(new_n581), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n700), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  AND4_X1   g0503(.A1(new_n470), .A2(new_n548), .A3(new_n575), .A4(new_n581), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n704), .A2(KEYINPUT30), .A3(G179), .A4(new_n496), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n548), .A2(G179), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n519), .A2(new_n478), .A3(new_n582), .A4(new_n706), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n703), .A2(new_n705), .A3(new_n707), .ZN(new_n708));
  AND3_X1   g0508(.A1(new_n708), .A2(KEYINPUT31), .A3(new_n655), .ZN(new_n709));
  AOI21_X1  g0509(.A(KEYINPUT31), .B1(new_n708), .B2(new_n655), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n711), .B1(new_n596), .B2(new_n655), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(new_n660), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n699), .A2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n679), .B1(new_n715), .B2(G1), .ZN(G364));
  NOR2_X1   g0516(.A1(new_n658), .A2(new_n660), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n648), .A2(G20), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n206), .B1(new_n718), .B2(G45), .ZN(new_n719));
  AOI211_X1 g0519(.A(new_n717), .B(new_n662), .C1(new_n675), .C2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n719), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n674), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n210), .A2(new_n261), .ZN(new_n723));
  INV_X1    g0523(.A(G355), .ZN(new_n724));
  OAI22_X1  g0524(.A1(new_n723), .A2(new_n724), .B1(G116), .B2(new_n210), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n673), .A2(new_n261), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n727), .B1(new_n463), .B2(new_n214), .ZN(new_n728));
  OR2_X1    g0528(.A1(new_n241), .A2(new_n463), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n725), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n215), .B1(G20), .B2(new_n296), .ZN(new_n731));
  NOR3_X1   g0531(.A1(G13), .A2(G20), .A3(G33), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n722), .B1(new_n730), .B2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n207), .A2(G190), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT96), .ZN(new_n737));
  XNOR2_X1  g0537(.A(new_n736), .B(new_n737), .ZN(new_n738));
  NOR3_X1   g0538(.A1(new_n738), .A2(G179), .A3(G200), .ZN(new_n739));
  XOR2_X1   g0539(.A(new_n739), .B(KEYINPUT98), .Z(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(G329), .ZN(new_n741));
  NOR2_X1   g0541(.A1(G179), .A2(G200), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n207), .B1(new_n742), .B2(G190), .ZN(new_n743));
  INV_X1    g0543(.A(G294), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g0545(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(G190), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  OR2_X1    g0548(.A1(KEYINPUT33), .A2(G317), .ZN(new_n749));
  NAND2_X1  g0549(.A1(KEYINPUT33), .A2(G317), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n748), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n746), .A2(new_n292), .ZN(new_n752));
  AOI211_X1 g0552(.A(new_n745), .B(new_n751), .C1(G326), .C2(new_n752), .ZN(new_n753));
  NOR3_X1   g0553(.A1(new_n738), .A2(G179), .A3(new_n416), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(G283), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n207), .A2(new_n292), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n756), .A2(new_n412), .A3(G200), .ZN(new_n757));
  INV_X1    g0557(.A(G303), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n412), .A2(G200), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n756), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(G322), .ZN(new_n761));
  OAI22_X1  g0561(.A1(new_n757), .A2(new_n758), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n736), .A2(new_n759), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  AOI211_X1 g0564(.A(new_n261), .B(new_n762), .C1(G311), .C2(new_n764), .ZN(new_n765));
  NAND4_X1  g0565(.A1(new_n741), .A2(new_n753), .A3(new_n755), .A4(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n739), .A2(G159), .ZN(new_n767));
  XNOR2_X1  g0567(.A(KEYINPUT97), .B(KEYINPUT32), .ZN(new_n768));
  XNOR2_X1  g0568(.A(new_n767), .B(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n743), .A2(new_n498), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n261), .B1(new_n757), .B2(new_n329), .ZN(new_n771));
  AOI211_X1 g0571(.A(new_n770), .B(new_n771), .C1(G68), .C2(new_n747), .ZN(new_n772));
  INV_X1    g0572(.A(new_n754), .ZN(new_n773));
  OAI211_X1 g0573(.A(new_n769), .B(new_n772), .C1(new_n422), .C2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n760), .ZN(new_n775));
  AOI22_X1  g0575(.A1(G58), .A2(new_n775), .B1(new_n764), .B2(G77), .ZN(new_n776));
  INV_X1    g0576(.A(new_n752), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n776), .B1(new_n202), .B2(new_n777), .ZN(new_n778));
  XOR2_X1   g0578(.A(new_n778), .B(KEYINPUT95), .Z(new_n779));
  OAI21_X1  g0579(.A(new_n766), .B1(new_n774), .B2(new_n779), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n735), .B1(new_n780), .B2(new_n731), .ZN(new_n781));
  XOR2_X1   g0581(.A(new_n732), .B(KEYINPUT99), .Z(new_n782));
  OAI21_X1  g0582(.A(new_n781), .B1(new_n658), .B2(new_n782), .ZN(new_n783));
  XOR2_X1   g0583(.A(new_n783), .B(KEYINPUT100), .Z(new_n784));
  NOR2_X1   g0584(.A1(new_n720), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(G396));
  NOR2_X1   g0586(.A1(G13), .A2(G33), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n731), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n722), .B1(G77), .B2(new_n789), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT101), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n740), .A2(G311), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n777), .A2(new_n758), .ZN(new_n793));
  AOI211_X1 g0593(.A(new_n770), .B(new_n793), .C1(G283), .C2(new_n747), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n754), .A2(G87), .ZN(new_n795));
  OAI22_X1  g0595(.A1(new_n757), .A2(new_n422), .B1(new_n760), .B2(new_n744), .ZN(new_n796));
  AOI211_X1 g0596(.A(new_n261), .B(new_n796), .C1(G116), .C2(new_n764), .ZN(new_n797));
  NAND4_X1  g0597(.A1(new_n792), .A2(new_n794), .A3(new_n795), .A4(new_n797), .ZN(new_n798));
  AOI22_X1  g0598(.A1(G143), .A2(new_n775), .B1(new_n764), .B2(G159), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n799), .B1(new_n276), .B2(new_n748), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n800), .B1(G137), .B2(new_n752), .ZN(new_n801));
  XNOR2_X1  g0601(.A(KEYINPUT102), .B(KEYINPUT34), .ZN(new_n802));
  XNOR2_X1  g0602(.A(new_n801), .B(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n743), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n310), .B1(new_n804), .B2(G58), .ZN(new_n805));
  INV_X1    g0605(.A(G132), .ZN(new_n806));
  INV_X1    g0606(.A(new_n740), .ZN(new_n807));
  OAI211_X1 g0607(.A(new_n803), .B(new_n805), .C1(new_n806), .C2(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n754), .A2(G68), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n809), .B1(new_n202), .B2(new_n757), .ZN(new_n810));
  XNOR2_X1  g0610(.A(new_n810), .B(KEYINPUT103), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n798), .B1(new_n808), .B2(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n791), .B1(new_n812), .B2(new_n731), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n414), .A2(new_n655), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n417), .B1(new_n403), .B2(new_n665), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(new_n414), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n787), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n813), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n418), .A2(new_n655), .ZN(new_n822));
  AOI22_X1  g0622(.A1(new_n696), .A2(new_n818), .B1(new_n645), .B2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n713), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n722), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT104), .ZN(new_n826));
  OAI22_X1  g0626(.A1(new_n825), .A2(new_n826), .B1(new_n824), .B2(new_n823), .ZN(new_n827));
  AND2_X1   g0627(.A1(new_n825), .A2(new_n826), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n821), .B1(new_n827), .B2(new_n828), .ZN(G384));
  NOR2_X1   g0629(.A1(new_n718), .A2(new_n206), .ZN(new_n830));
  INV_X1    g0630(.A(new_n699), .ZN(new_n831));
  AOI22_X1  g0631(.A1(new_n831), .A2(new_n419), .B1(new_n618), .B2(new_n619), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n599), .A2(new_n343), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n653), .B1(new_n318), .B2(new_n338), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT105), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NOR3_X1   g0636(.A1(new_n349), .A2(KEYINPUT105), .A3(new_n653), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n833), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n838), .A2(KEYINPUT37), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT37), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n840), .B1(new_n349), .B2(new_n342), .ZN(new_n841));
  NOR3_X1   g0641(.A1(new_n841), .A2(new_n599), .A3(new_n834), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n839), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n834), .A2(new_n835), .ZN(new_n845));
  OAI21_X1  g0645(.A(KEYINPUT105), .B1(new_n349), .B2(new_n653), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n847), .B1(new_n340), .B2(new_n351), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n844), .A2(new_n849), .A3(KEYINPUT38), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT38), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n842), .B1(new_n838), .B2(KEYINPUT37), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n851), .B1(new_n852), .B2(new_n848), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n850), .A2(new_n853), .A3(KEYINPUT39), .ZN(new_n854));
  NOR3_X1   g0654(.A1(new_n852), .A2(new_n848), .A3(new_n851), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n600), .B1(new_n609), .B2(new_n612), .ZN(new_n856));
  INV_X1    g0656(.A(new_n834), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n610), .A2(new_n611), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n599), .A2(new_n834), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n840), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  OAI22_X1  g0660(.A1(new_n856), .A2(new_n857), .B1(new_n842), .B2(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n855), .B1(new_n861), .B2(new_n851), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n854), .B1(new_n862), .B2(KEYINPUT39), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n388), .A2(new_n655), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n361), .A2(new_n655), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n388), .A2(new_n393), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n377), .A2(G169), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n869), .A2(KEYINPUT14), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n377), .A2(new_n362), .A3(G169), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n385), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT72), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n380), .A2(KEYINPUT72), .A3(new_n385), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n393), .ZN(new_n877));
  OAI211_X1 g0677(.A(new_n361), .B(new_n655), .C1(new_n876), .C2(new_n877), .ZN(new_n878));
  AND2_X1   g0678(.A1(new_n868), .A2(new_n878), .ZN(new_n879));
  OAI22_X1  g0679(.A1(new_n689), .A2(new_n690), .B1(new_n633), .B2(new_n634), .ZN(new_n880));
  INV_X1    g0680(.A(new_n644), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n822), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n879), .B1(new_n882), .B2(new_n815), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n850), .A2(new_n853), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n653), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n885), .B1(new_n613), .B2(new_n886), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n866), .A2(new_n887), .ZN(new_n888));
  XNOR2_X1  g0688(.A(new_n832), .B(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n868), .A2(new_n878), .ZN(new_n890));
  AND3_X1   g0690(.A1(new_n890), .A2(new_n712), .A3(new_n819), .ZN(new_n891));
  AOI21_X1  g0691(.A(KEYINPUT40), .B1(new_n891), .B2(new_n884), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT106), .ZN(new_n893));
  NAND4_X1  g0693(.A1(new_n890), .A2(new_n712), .A3(KEYINPUT40), .A4(new_n819), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n893), .B1(new_n862), .B2(new_n894), .ZN(new_n895));
  AND4_X1   g0695(.A1(KEYINPUT40), .A2(new_n890), .A3(new_n712), .A4(new_n819), .ZN(new_n896));
  AND3_X1   g0696(.A1(new_n610), .A2(KEYINPUT18), .A3(new_n611), .ZN(new_n897));
  AOI21_X1  g0697(.A(KEYINPUT18), .B1(new_n610), .B2(new_n611), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n340), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n859), .B1(new_n607), .B2(new_n608), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(KEYINPUT37), .ZN(new_n901));
  AOI22_X1  g0701(.A1(new_n899), .A2(new_n834), .B1(new_n901), .B2(new_n843), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n850), .B1(new_n902), .B2(KEYINPUT38), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n896), .A2(new_n903), .A3(KEYINPUT106), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n892), .B1(new_n895), .B2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n419), .A2(new_n712), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n659), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n908), .B1(new_n907), .B2(new_n906), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n830), .B1(new_n889), .B2(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n910), .B1(new_n889), .B2(new_n909), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n562), .B1(new_n563), .B2(new_n564), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT35), .ZN(new_n913));
  OAI211_X1 g0713(.A(G116), .B(new_n216), .C1(new_n912), .C2(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n914), .B1(new_n913), .B2(new_n912), .ZN(new_n915));
  XOR2_X1   g0715(.A(new_n915), .B(KEYINPUT36), .Z(new_n916));
  NOR4_X1   g0716(.A1(new_n301), .A2(new_n300), .A3(new_n213), .A4(new_n263), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n219), .A2(G50), .ZN(new_n918));
  OAI211_X1 g0718(.A(G1), .B(new_n648), .C1(new_n917), .C2(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n911), .A2(new_n916), .A3(new_n919), .ZN(G367));
  NAND2_X1  g0720(.A1(new_n671), .A2(new_n668), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n585), .B(new_n594), .C1(new_n591), .C2(new_n665), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n626), .A2(new_n655), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(new_n924), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n921), .A2(new_n925), .ZN(new_n926));
  AND2_X1   g0726(.A1(new_n926), .A2(KEYINPUT45), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n926), .A2(KEYINPUT45), .ZN(new_n928));
  AOI21_X1  g0728(.A(KEYINPUT44), .B1(new_n921), .B2(new_n925), .ZN(new_n929));
  AND3_X1   g0729(.A1(new_n921), .A2(KEYINPUT44), .A3(new_n925), .ZN(new_n930));
  OAI22_X1  g0730(.A1(new_n927), .A2(new_n928), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(new_n667), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n931), .B(new_n932), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n671), .A2(KEYINPUT109), .ZN(new_n934));
  OR2_X1    g0734(.A1(new_n666), .A2(new_n670), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT109), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n934), .B1(new_n937), .B2(new_n671), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n938), .B(new_n661), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(new_n715), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n715), .B1(new_n933), .B2(new_n940), .ZN(new_n941));
  XOR2_X1   g0741(.A(new_n674), .B(KEYINPUT41), .Z(new_n942));
  INV_X1    g0742(.A(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n721), .B1(new_n941), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n546), .A2(new_n547), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n655), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n640), .A2(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(new_n623), .B2(new_n946), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(KEYINPUT43), .ZN(new_n949));
  XOR2_X1   g0749(.A(new_n949), .B(KEYINPUT108), .Z(new_n950));
  NAND3_X1  g0750(.A1(new_n669), .A2(new_n670), .A3(new_n924), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(KEYINPUT42), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n585), .B1(new_n481), .B2(new_n922), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(new_n665), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n951), .A2(KEYINPUT42), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n950), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n948), .A2(KEYINPUT43), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n958), .B(KEYINPUT107), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n957), .B(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n932), .A2(new_n924), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n960), .B(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(G283), .ZN(new_n963));
  OAI22_X1  g0763(.A1(new_n760), .A2(new_n758), .B1(new_n763), .B2(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(new_n757), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(G116), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT46), .ZN(new_n967));
  INV_X1    g0767(.A(G311), .ZN(new_n968));
  OAI221_X1 g0768(.A(new_n967), .B1(new_n744), .B2(new_n748), .C1(new_n968), .C2(new_n777), .ZN(new_n969));
  AOI211_X1 g0769(.A(new_n964), .B(new_n969), .C1(G107), .C2(new_n804), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT110), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n754), .A2(G97), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n739), .A2(G317), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n972), .A2(new_n973), .A3(new_n310), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n970), .B1(new_n971), .B2(new_n974), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n975), .B1(new_n971), .B2(new_n974), .ZN(new_n976));
  XOR2_X1   g0776(.A(new_n976), .B(KEYINPUT111), .Z(new_n977));
  NAND2_X1  g0777(.A1(new_n804), .A2(G68), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n752), .A2(G143), .ZN(new_n979));
  OAI211_X1 g0779(.A(new_n978), .B(new_n979), .C1(new_n303), .C2(new_n748), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n754), .A2(G77), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n310), .B1(new_n965), .B2(G58), .ZN(new_n982));
  AOI22_X1  g0782(.A1(G150), .A2(new_n775), .B1(new_n764), .B2(G50), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n981), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  AOI211_X1 g0784(.A(new_n980), .B(new_n984), .C1(G137), .C2(new_n739), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n977), .A2(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n731), .B1(new_n986), .B2(KEYINPUT47), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n987), .B1(KEYINPUT47), .B2(new_n986), .ZN(new_n988));
  AND2_X1   g0788(.A1(new_n232), .A2(new_n726), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n733), .B1(new_n210), .B2(new_n395), .ZN(new_n990));
  OAI221_X1 g0790(.A(new_n722), .B1(new_n989), .B2(new_n990), .C1(new_n948), .C2(new_n782), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n944), .A2(new_n962), .B1(new_n988), .B2(new_n991), .ZN(G387));
  OR2_X1    g0792(.A1(new_n666), .A2(new_n782), .ZN(new_n993));
  OAI22_X1  g0793(.A1(new_n723), .A2(new_n676), .B1(G107), .B2(new_n210), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n237), .A2(G45), .ZN(new_n995));
  INV_X1    g0795(.A(new_n676), .ZN(new_n996));
  AOI211_X1 g0796(.A(G45), .B(new_n996), .C1(G68), .C2(G77), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n280), .A2(G50), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n998), .B(KEYINPUT50), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n727), .B1(new_n997), .B2(new_n999), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n994), .B1(new_n995), .B2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n722), .B1(new_n1001), .B2(new_n734), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n743), .A2(new_n395), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n310), .B1(new_n764), .B2(G68), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n1004), .B1(new_n202), .B2(new_n760), .C1(new_n263), .C2(new_n757), .ZN(new_n1005));
  AOI211_X1 g0805(.A(new_n1003), .B(new_n1005), .C1(G159), .C2(new_n752), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n739), .A2(G150), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n285), .A2(new_n747), .ZN(new_n1008));
  NAND4_X1  g0808(.A1(new_n1006), .A2(new_n972), .A3(new_n1007), .A4(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n261), .B1(new_n739), .B2(G326), .ZN(new_n1010));
  OAI22_X1  g0810(.A1(new_n757), .A2(new_n744), .B1(new_n743), .B2(new_n963), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(G317), .A2(new_n775), .B1(new_n764), .B2(G303), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n1012), .B1(new_n777), .B2(new_n761), .C1(new_n968), .C2(new_n748), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT48), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1011), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1015), .B1(new_n1014), .B2(new_n1013), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT49), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n1010), .B1(new_n444), .B2(new_n773), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1018));
  AND2_X1   g0818(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1009), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1002), .B1(new_n1020), .B2(new_n731), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n939), .A2(new_n721), .B1(new_n993), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n940), .A2(new_n674), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n939), .A2(new_n715), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1022), .B1(new_n1023), .B2(new_n1024), .ZN(G393));
  OR2_X1    g0825(.A1(new_n933), .A2(KEYINPUT112), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n719), .B1(new_n933), .B2(KEYINPUT112), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n925), .A2(new_n732), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n733), .B1(new_n498), .B2(new_n210), .C1(new_n727), .C2(new_n244), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1029), .A2(new_n722), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n775), .A2(G311), .B1(G317), .B2(new_n752), .ZN(new_n1031));
  XOR2_X1   g0831(.A(new_n1031), .B(KEYINPUT52), .Z(new_n1032));
  OAI21_X1  g0832(.A(new_n310), .B1(new_n763), .B2(new_n744), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1033), .B1(G283), .B2(new_n965), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n804), .A2(G116), .B1(G303), .B2(new_n747), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(G107), .A2(new_n754), .B1(new_n739), .B2(G322), .ZN(new_n1036));
  NAND4_X1  g0836(.A1(new_n1032), .A2(new_n1034), .A3(new_n1035), .A4(new_n1036), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n743), .A2(new_n263), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n261), .B1(new_n763), .B2(new_n280), .C1(new_n757), .C2(new_n219), .ZN(new_n1039));
  AOI211_X1 g0839(.A(new_n1038), .B(new_n1039), .C1(G50), .C2(new_n747), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n739), .A2(G143), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1040), .A2(new_n795), .A3(new_n1041), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n777), .A2(new_n276), .B1(new_n760), .B2(new_n303), .ZN(new_n1043));
  XOR2_X1   g0843(.A(new_n1043), .B(KEYINPUT51), .Z(new_n1044));
  OAI21_X1  g0844(.A(new_n1037), .B1(new_n1042), .B2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1030), .B1(new_n1045), .B2(new_n731), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n1026), .A2(new_n1027), .B1(new_n1028), .B2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n674), .B1(new_n933), .B2(new_n940), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT113), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n933), .A2(new_n940), .ZN(new_n1051));
  AND3_X1   g0851(.A1(new_n1049), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1050), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1047), .B1(new_n1052), .B2(new_n1053), .ZN(G390));
  INV_X1    g0854(.A(KEYINPUT114), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n814), .B1(new_n645), .B2(new_n822), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n865), .B1(new_n1056), .B2(new_n879), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n688), .A2(new_n692), .A3(new_n815), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1058), .A2(new_n817), .A3(new_n890), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n857), .B1(new_n613), .B2(new_n340), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n860), .A2(new_n842), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n851), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n864), .B1(new_n1062), .B2(new_n850), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n863), .A2(new_n1057), .B1(new_n1059), .B2(new_n1063), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n879), .A2(new_n818), .ZN(new_n1065));
  AND2_X1   g0865(.A1(new_n712), .A2(G330), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1055), .B1(new_n1064), .B2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1059), .A2(new_n1063), .ZN(new_n1069));
  AOI21_X1  g0869(.A(KEYINPUT39), .B1(new_n1062), .B2(new_n850), .ZN(new_n1070));
  AND3_X1   g0870(.A1(new_n850), .A2(new_n853), .A3(KEYINPUT39), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n1070), .A2(new_n1071), .B1(new_n883), .B2(new_n864), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1069), .A2(new_n1072), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1067), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1073), .A2(KEYINPUT114), .A3(new_n1074), .ZN(new_n1075));
  NOR3_X1   g0875(.A1(new_n713), .A2(new_n879), .A3(new_n818), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n1076), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1069), .A2(new_n1072), .A3(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1078), .A2(KEYINPUT115), .ZN(new_n1079));
  INV_X1    g0879(.A(KEYINPUT115), .ZN(new_n1080));
  NAND4_X1  g0880(.A1(new_n1069), .A2(new_n1072), .A3(new_n1080), .A4(new_n1077), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n1068), .A2(new_n1075), .B1(new_n1079), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n721), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n863), .A2(new_n787), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n722), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n285), .A2(new_n789), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n740), .A2(G294), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n777), .A2(new_n963), .ZN(new_n1088));
  AOI211_X1 g0888(.A(new_n1038), .B(new_n1088), .C1(G107), .C2(new_n747), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n760), .A2(new_n444), .B1(new_n763), .B2(new_n498), .ZN(new_n1090));
  AOI211_X1 g0890(.A(new_n261), .B(new_n1090), .C1(G87), .C2(new_n965), .ZN(new_n1091));
  NAND4_X1  g0891(.A1(new_n1087), .A2(new_n809), .A3(new_n1089), .A4(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(G125), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n310), .B1(new_n754), .B2(G50), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n807), .A2(new_n1093), .B1(new_n1094), .B2(KEYINPUT116), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1094), .A2(KEYINPUT116), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n752), .A2(G128), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(KEYINPUT54), .B(G143), .ZN(new_n1098));
  OAI221_X1 g0898(.A(new_n1097), .B1(new_n763), .B2(new_n1098), .C1(new_n806), .C2(new_n760), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(new_n804), .A2(G159), .B1(G137), .B2(new_n747), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n757), .A2(new_n276), .ZN(new_n1102));
  XOR2_X1   g0902(.A(KEYINPUT117), .B(KEYINPUT53), .Z(new_n1103));
  XNOR2_X1  g0903(.A(new_n1102), .B(new_n1103), .ZN(new_n1104));
  NAND4_X1  g0904(.A1(new_n1096), .A2(new_n1100), .A3(new_n1101), .A4(new_n1104), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1092), .B1(new_n1095), .B2(new_n1105), .ZN(new_n1106));
  AOI211_X1 g0906(.A(new_n1085), .B(new_n1086), .C1(new_n1106), .C2(new_n731), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1084), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n419), .A2(new_n1066), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n620), .B(new_n1109), .C1(new_n699), .C2(new_n420), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n890), .B1(new_n1066), .B2(new_n819), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n1111), .A2(new_n1076), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1058), .A2(new_n817), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n879), .B1(new_n713), .B2(new_n818), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1067), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1056), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n1112), .A2(new_n1113), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n1110), .A2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n674), .B1(new_n1082), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1068), .A2(new_n1075), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1120), .A2(new_n1121), .A3(new_n1118), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n1083), .B(new_n1108), .C1(new_n1119), .C2(new_n1123), .ZN(G378));
  AOI21_X1  g0924(.A(new_n1110), .B1(new_n1082), .B2(new_n1118), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n891), .A2(new_n884), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT40), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NOR3_X1   g0928(.A1(new_n862), .A2(new_n893), .A3(new_n894), .ZN(new_n1129));
  AOI21_X1  g0929(.A(KEYINPUT106), .B1(new_n896), .B2(new_n903), .ZN(new_n1130));
  OAI211_X1 g0930(.A(G330), .B(new_n1128), .C1(new_n1129), .C2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n290), .A2(new_n886), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n299), .A2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n294), .A2(new_n298), .A3(new_n1132), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1134), .A2(new_n1135), .A3(new_n1137), .ZN(new_n1140));
  AND2_X1   g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1131), .A2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n905), .A2(G330), .A3(new_n1143), .ZN(new_n1144));
  AND3_X1   g0944(.A1(new_n1142), .A2(new_n888), .A3(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n888), .B1(new_n1142), .B2(new_n1144), .ZN(new_n1146));
  OAI21_X1  g0946(.A(KEYINPUT57), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n674), .B1(new_n1125), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1110), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1122), .A2(new_n1149), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n1131), .A2(new_n1141), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1143), .B1(new_n905), .B2(G330), .ZN(new_n1152));
  OAI22_X1  g0952(.A1(new_n1151), .A2(new_n1152), .B1(new_n866), .B2(new_n887), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1142), .A2(new_n1144), .A3(new_n888), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(KEYINPUT57), .B1(new_n1150), .B2(new_n1155), .ZN(new_n1156));
  OR2_X1    g0956(.A1(new_n1148), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1141), .A2(new_n787), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n722), .B1(G50), .B2(new_n789), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n754), .A2(G58), .ZN(new_n1160));
  XOR2_X1   g0960(.A(new_n1160), .B(KEYINPUT118), .Z(new_n1161));
  OAI221_X1 g0961(.A(new_n978), .B1(new_n777), .B2(new_n444), .C1(new_n498), .C2(new_n748), .ZN(new_n1162));
  OAI22_X1  g0962(.A1(new_n757), .A2(new_n263), .B1(new_n763), .B2(new_n395), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n760), .A2(new_n422), .ZN(new_n1164));
  OR2_X1    g0964(.A1(new_n261), .A2(G41), .ZN(new_n1165));
  NOR4_X1   g0965(.A1(new_n1162), .A2(new_n1163), .A3(new_n1164), .A4(new_n1165), .ZN(new_n1166));
  OAI211_X1 g0966(.A(new_n1161), .B(new_n1166), .C1(new_n807), .C2(new_n963), .ZN(new_n1167));
  INV_X1    g0967(.A(KEYINPUT58), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  OAI211_X1 g0969(.A(new_n1165), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1170));
  AND2_X1   g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n748), .A2(new_n806), .B1(new_n276), .B2(new_n743), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n764), .A2(G137), .ZN(new_n1173));
  INV_X1    g0973(.A(G128), .ZN(new_n1174));
  OAI221_X1 g0974(.A(new_n1173), .B1(new_n1174), .B2(new_n760), .C1(new_n757), .C2(new_n1098), .ZN(new_n1175));
  AOI211_X1 g0975(.A(new_n1172), .B(new_n1175), .C1(G125), .C2(new_n752), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1176), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n1177), .A2(KEYINPUT59), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1177), .A2(KEYINPUT59), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n754), .A2(G159), .ZN(new_n1180));
  AOI211_X1 g0980(.A(G33), .B(G41), .C1(new_n739), .C2(G124), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1179), .A2(new_n1180), .A3(new_n1181), .ZN(new_n1182));
  OAI221_X1 g0982(.A(new_n1171), .B1(new_n1168), .B2(new_n1167), .C1(new_n1178), .C2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1159), .B1(new_n1183), .B2(new_n731), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(new_n1155), .A2(new_n721), .B1(new_n1158), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1157), .A2(new_n1185), .ZN(G375));
  INV_X1    g0986(.A(new_n1118), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1110), .A2(new_n1117), .ZN(new_n1188));
  XOR2_X1   g0988(.A(new_n942), .B(KEYINPUT119), .Z(new_n1189));
  NAND3_X1  g0989(.A1(new_n1187), .A2(new_n1188), .A3(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1117), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n879), .A2(new_n787), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n722), .B1(G68), .B2(new_n789), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n981), .A2(new_n310), .ZN(new_n1194));
  XNOR2_X1  g0994(.A(new_n1194), .B(KEYINPUT120), .ZN(new_n1195));
  OAI22_X1  g0995(.A1(new_n757), .A2(new_n498), .B1(new_n760), .B2(new_n963), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1003), .B1(new_n747), .B2(G116), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1197), .B1(new_n744), .B2(new_n777), .ZN(new_n1198));
  AOI211_X1 g0998(.A(new_n1196), .B(new_n1198), .C1(G107), .C2(new_n764), .ZN(new_n1199));
  OAI211_X1 g0999(.A(new_n1195), .B(new_n1199), .C1(new_n758), .C2(new_n807), .ZN(new_n1200));
  XOR2_X1   g1000(.A(new_n1200), .B(KEYINPUT121), .Z(new_n1201));
  OAI221_X1 g1001(.A(new_n261), .B1(new_n763), .B2(new_n276), .C1(new_n757), .C2(new_n303), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(G50), .B2(new_n804), .ZN(new_n1203));
  OAI211_X1 g1003(.A(new_n1161), .B(new_n1203), .C1(new_n807), .C2(new_n1174), .ZN(new_n1204));
  INV_X1    g1004(.A(KEYINPUT122), .ZN(new_n1205));
  AND2_X1   g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n748), .A2(new_n1098), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1207), .B1(G137), .B2(new_n775), .ZN(new_n1208));
  OAI221_X1 g1008(.A(new_n1208), .B1(new_n806), .B2(new_n777), .C1(new_n1204), .C2(new_n1205), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1201), .B1(new_n1206), .B2(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1193), .B1(new_n1210), .B2(new_n731), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n1191), .A2(new_n721), .B1(new_n1192), .B2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1190), .A2(new_n1212), .ZN(G381));
  INV_X1    g1013(.A(G375), .ZN(new_n1214));
  OR4_X1    g1014(.A1(G396), .A2(G381), .A3(G393), .A4(G384), .ZN(new_n1215));
  NOR3_X1   g1015(.A1(new_n1215), .A2(G390), .A3(G387), .ZN(new_n1216));
  INV_X1    g1016(.A(G378), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1214), .A2(new_n1216), .A3(new_n1217), .ZN(new_n1218));
  AND2_X1   g1018(.A1(new_n1218), .A2(KEYINPUT123), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n1218), .A2(KEYINPUT123), .ZN(new_n1220));
  OR2_X1    g1020(.A1(new_n1219), .A2(new_n1220), .ZN(G407));
  NAND2_X1  g1021(.A1(new_n1217), .A2(new_n654), .ZN(new_n1222));
  OAI221_X1 g1022(.A(G213), .B1(G375), .B2(new_n1222), .C1(new_n1219), .C2(new_n1220), .ZN(G409));
  INV_X1    g1023(.A(KEYINPUT63), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1189), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1225));
  OAI21_X1  g1025(.A(KEYINPUT124), .B1(new_n1125), .B2(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1189), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1227), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT124), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1150), .A2(new_n1228), .A3(new_n1229), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1226), .A2(new_n1185), .A3(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1231), .A2(new_n1217), .ZN(new_n1232));
  OAI211_X1 g1032(.A(G378), .B(new_n1185), .C1(new_n1148), .C2(new_n1156), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(G213), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n1235), .A2(G343), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1234), .A2(new_n1237), .ZN(new_n1238));
  XNOR2_X1  g1038(.A(KEYINPUT125), .B(KEYINPUT60), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1188), .B1(new_n1118), .B2(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT60), .ZN(new_n1242));
  OAI211_X1 g1042(.A(new_n1241), .B(new_n674), .C1(new_n1242), .C2(new_n1188), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1243), .A2(G384), .A3(new_n1212), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(G384), .B1(new_n1243), .B2(new_n1212), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1247), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1224), .B1(new_n1238), .B2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1236), .A2(G2897), .ZN(new_n1250));
  XOR2_X1   g1050(.A(new_n1250), .B(KEYINPUT126), .Z(new_n1251));
  OAI21_X1  g1051(.A(new_n1251), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1246), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1251), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1253), .A2(new_n1244), .A3(new_n1254), .ZN(new_n1255));
  AND2_X1   g1055(.A1(new_n1252), .A2(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(KEYINPUT61), .B1(new_n1238), .B2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(G387), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(G390), .A2(new_n1258), .ZN(new_n1259));
  OAI211_X1 g1059(.A(G387), .B(new_n1047), .C1(new_n1052), .C2(new_n1053), .ZN(new_n1260));
  XNOR2_X1  g1060(.A(G393), .B(new_n785), .ZN(new_n1261));
  AND3_X1   g1061(.A1(new_n1259), .A2(new_n1260), .A3(new_n1261), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1261), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1236), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1265), .A2(KEYINPUT63), .A3(new_n1247), .ZN(new_n1266));
  NAND4_X1  g1066(.A1(new_n1249), .A2(new_n1257), .A3(new_n1264), .A4(new_n1266), .ZN(new_n1267));
  XOR2_X1   g1067(.A(KEYINPUT127), .B(KEYINPUT62), .Z(new_n1268));
  AND3_X1   g1068(.A1(new_n1265), .A2(new_n1247), .A3(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT61), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1252), .A2(new_n1255), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1270), .B1(new_n1265), .B2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1273), .B1(new_n1265), .B2(new_n1247), .ZN(new_n1274));
  NOR3_X1   g1074(.A1(new_n1269), .A2(new_n1272), .A3(new_n1274), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1267), .B1(new_n1275), .B2(new_n1264), .ZN(G405));
  NAND2_X1  g1076(.A1(G375), .A2(new_n1217), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1277), .A2(new_n1233), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1278), .A2(new_n1247), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1277), .A2(new_n1248), .A3(new_n1233), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1264), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1279), .A2(new_n1264), .A3(new_n1280), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1283), .A2(new_n1284), .ZN(G402));
endmodule


