

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U554 ( .A1(n522), .A2(G2104), .ZN(n879) );
  NOR2_X2 U555 ( .A1(G2104), .A2(G2105), .ZN(n526) );
  XNOR2_X1 U556 ( .A(KEYINPUT29), .B(KEYINPUT95), .ZN(n710) );
  NAND2_X1 U557 ( .A1(n756), .A2(n755), .ZN(n757) );
  AND2_X1 U558 ( .A1(n520), .A2(n769), .ZN(n770) );
  NAND2_X1 U559 ( .A1(G40), .A2(G160), .ZN(n788) );
  NOR2_X1 U560 ( .A1(n813), .A2(n803), .ZN(n804) );
  NAND2_X1 U561 ( .A1(n771), .A2(n770), .ZN(n805) );
  XNOR2_X1 U562 ( .A(KEYINPUT100), .B(n765), .ZN(n520) );
  NOR2_X1 U563 ( .A1(n687), .A2(n1013), .ZN(n695) );
  INV_X1 U564 ( .A(n686), .ZN(n712) );
  BUF_X1 U565 ( .A(n686), .Z(n689) );
  XNOR2_X1 U566 ( .A(n711), .B(n710), .ZN(n716) );
  OR2_X1 U567 ( .A1(n729), .A2(n728), .ZN(n747) );
  INV_X1 U568 ( .A(n1021), .ZN(n755) );
  INV_X1 U569 ( .A(n817), .ZN(n803) );
  NOR2_X1 U570 ( .A1(G1384), .A2(G164), .ZN(n681) );
  NOR2_X1 U571 ( .A1(G651), .A2(n646), .ZN(n650) );
  NOR2_X1 U572 ( .A1(n531), .A2(n530), .ZN(G160) );
  INV_X1 U573 ( .A(G2105), .ZN(n522) );
  NAND2_X1 U574 ( .A1(G101), .A2(n879), .ZN(n521) );
  XOR2_X1 U575 ( .A(KEYINPUT23), .B(n521), .Z(n525) );
  NOR2_X1 U576 ( .A1(G2104), .A2(n522), .ZN(n547) );
  NAND2_X1 U577 ( .A1(G125), .A2(n547), .ZN(n523) );
  XOR2_X1 U578 ( .A(KEYINPUT65), .B(n523), .Z(n524) );
  NAND2_X1 U579 ( .A1(n525), .A2(n524), .ZN(n531) );
  XOR2_X2 U580 ( .A(KEYINPUT17), .B(n526), .Z(n876) );
  NAND2_X1 U581 ( .A1(G137), .A2(n876), .ZN(n529) );
  NAND2_X1 U582 ( .A1(G2105), .A2(G2104), .ZN(n527) );
  XOR2_X1 U583 ( .A(KEYINPUT66), .B(n527), .Z(n549) );
  NAND2_X1 U584 ( .A1(G113), .A2(n549), .ZN(n528) );
  NAND2_X1 U585 ( .A1(n529), .A2(n528), .ZN(n530) );
  NAND2_X1 U586 ( .A1(G138), .A2(n876), .ZN(n533) );
  NAND2_X1 U587 ( .A1(G102), .A2(n879), .ZN(n532) );
  NAND2_X1 U588 ( .A1(n533), .A2(n532), .ZN(n537) );
  BUF_X1 U589 ( .A(n547), .Z(n854) );
  NAND2_X1 U590 ( .A1(G126), .A2(n854), .ZN(n535) );
  NAND2_X1 U591 ( .A1(G114), .A2(n549), .ZN(n534) );
  NAND2_X1 U592 ( .A1(n535), .A2(n534), .ZN(n536) );
  NOR2_X1 U593 ( .A1(n537), .A2(n536), .ZN(G164) );
  NOR2_X1 U594 ( .A1(G651), .A2(G543), .ZN(n637) );
  NAND2_X1 U595 ( .A1(G85), .A2(n637), .ZN(n539) );
  XOR2_X1 U596 ( .A(G543), .B(KEYINPUT0), .Z(n646) );
  INV_X1 U597 ( .A(G651), .ZN(n540) );
  NOR2_X1 U598 ( .A1(n646), .A2(n540), .ZN(n635) );
  NAND2_X1 U599 ( .A1(G72), .A2(n635), .ZN(n538) );
  NAND2_X1 U600 ( .A1(n539), .A2(n538), .ZN(n545) );
  NOR2_X1 U601 ( .A1(G543), .A2(n540), .ZN(n541) );
  XOR2_X1 U602 ( .A(KEYINPUT1), .B(n541), .Z(n589) );
  NAND2_X1 U603 ( .A1(G60), .A2(n589), .ZN(n543) );
  NAND2_X1 U604 ( .A1(G47), .A2(n650), .ZN(n542) );
  NAND2_X1 U605 ( .A1(n543), .A2(n542), .ZN(n544) );
  OR2_X1 U606 ( .A1(n545), .A2(n544), .ZN(G290) );
  AND2_X1 U607 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U608 ( .A1(G135), .A2(n876), .ZN(n546) );
  XNOR2_X1 U609 ( .A(n546), .B(KEYINPUT76), .ZN(n556) );
  NAND2_X1 U610 ( .A1(n854), .A2(G123), .ZN(n548) );
  XNOR2_X1 U611 ( .A(n548), .B(KEYINPUT18), .ZN(n551) );
  BUF_X1 U612 ( .A(n549), .Z(n872) );
  NAND2_X1 U613 ( .A1(G111), .A2(n872), .ZN(n550) );
  NAND2_X1 U614 ( .A1(n551), .A2(n550), .ZN(n554) );
  NAND2_X1 U615 ( .A1(G99), .A2(n879), .ZN(n552) );
  XNOR2_X1 U616 ( .A(KEYINPUT77), .B(n552), .ZN(n553) );
  NOR2_X1 U617 ( .A1(n554), .A2(n553), .ZN(n555) );
  NAND2_X1 U618 ( .A1(n556), .A2(n555), .ZN(n972) );
  XNOR2_X1 U619 ( .A(G2096), .B(n972), .ZN(n557) );
  OR2_X1 U620 ( .A1(G2100), .A2(n557), .ZN(G156) );
  INV_X1 U621 ( .A(G57), .ZN(G237) );
  NAND2_X1 U622 ( .A1(G88), .A2(n637), .ZN(n559) );
  NAND2_X1 U623 ( .A1(G75), .A2(n635), .ZN(n558) );
  NAND2_X1 U624 ( .A1(n559), .A2(n558), .ZN(n563) );
  NAND2_X1 U625 ( .A1(G62), .A2(n589), .ZN(n561) );
  NAND2_X1 U626 ( .A1(G50), .A2(n650), .ZN(n560) );
  NAND2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n562) );
  NOR2_X1 U628 ( .A1(n563), .A2(n562), .ZN(G166) );
  NAND2_X1 U629 ( .A1(G64), .A2(n589), .ZN(n565) );
  NAND2_X1 U630 ( .A1(G52), .A2(n650), .ZN(n564) );
  NAND2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n570) );
  NAND2_X1 U632 ( .A1(G90), .A2(n637), .ZN(n567) );
  NAND2_X1 U633 ( .A1(G77), .A2(n635), .ZN(n566) );
  NAND2_X1 U634 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U635 ( .A(KEYINPUT9), .B(n568), .Z(n569) );
  NOR2_X1 U636 ( .A1(n570), .A2(n569), .ZN(G171) );
  NAND2_X1 U637 ( .A1(n637), .A2(G89), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n571), .B(KEYINPUT4), .ZN(n573) );
  NAND2_X1 U639 ( .A1(G76), .A2(n635), .ZN(n572) );
  NAND2_X1 U640 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n574), .B(KEYINPUT5), .ZN(n580) );
  NAND2_X1 U642 ( .A1(n650), .A2(G51), .ZN(n575) );
  XNOR2_X1 U643 ( .A(n575), .B(KEYINPUT72), .ZN(n577) );
  NAND2_X1 U644 ( .A1(G63), .A2(n589), .ZN(n576) );
  NAND2_X1 U645 ( .A1(n577), .A2(n576), .ZN(n578) );
  XOR2_X1 U646 ( .A(KEYINPUT6), .B(n578), .Z(n579) );
  NAND2_X1 U647 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U648 ( .A(n581), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U649 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U650 ( .A1(G7), .A2(G661), .ZN(n582) );
  XNOR2_X1 U651 ( .A(n582), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U652 ( .A(KEYINPUT11), .B(KEYINPUT68), .Z(n584) );
  INV_X1 U653 ( .A(G223), .ZN(n826) );
  NAND2_X1 U654 ( .A1(G567), .A2(n826), .ZN(n583) );
  XNOR2_X1 U655 ( .A(n584), .B(n583), .ZN(G234) );
  NAND2_X1 U656 ( .A1(n637), .A2(G81), .ZN(n585) );
  XNOR2_X1 U657 ( .A(n585), .B(KEYINPUT12), .ZN(n587) );
  NAND2_X1 U658 ( .A1(G68), .A2(n635), .ZN(n586) );
  NAND2_X1 U659 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U660 ( .A(KEYINPUT13), .B(n588), .Z(n593) );
  NAND2_X1 U661 ( .A1(G56), .A2(n589), .ZN(n590) );
  XNOR2_X1 U662 ( .A(n590), .B(KEYINPUT14), .ZN(n591) );
  XNOR2_X1 U663 ( .A(n591), .B(KEYINPUT69), .ZN(n592) );
  NOR2_X1 U664 ( .A1(n593), .A2(n592), .ZN(n595) );
  NAND2_X1 U665 ( .A1(n650), .A2(G43), .ZN(n594) );
  NAND2_X1 U666 ( .A1(n595), .A2(n594), .ZN(n1013) );
  INV_X1 U667 ( .A(n1013), .ZN(n596) );
  NAND2_X1 U668 ( .A1(n596), .A2(G860), .ZN(n597) );
  XNOR2_X1 U669 ( .A(KEYINPUT70), .B(n597), .ZN(G153) );
  INV_X1 U670 ( .A(G171), .ZN(G301) );
  NAND2_X1 U671 ( .A1(G868), .A2(G301), .ZN(n607) );
  NAND2_X1 U672 ( .A1(G54), .A2(n650), .ZN(n604) );
  NAND2_X1 U673 ( .A1(G79), .A2(n635), .ZN(n599) );
  NAND2_X1 U674 ( .A1(G66), .A2(n589), .ZN(n598) );
  NAND2_X1 U675 ( .A1(n599), .A2(n598), .ZN(n602) );
  NAND2_X1 U676 ( .A1(G92), .A2(n637), .ZN(n600) );
  XNOR2_X1 U677 ( .A(KEYINPUT71), .B(n600), .ZN(n601) );
  NOR2_X1 U678 ( .A1(n602), .A2(n601), .ZN(n603) );
  NAND2_X1 U679 ( .A1(n604), .A2(n603), .ZN(n605) );
  XNOR2_X1 U680 ( .A(n605), .B(KEYINPUT15), .ZN(n1000) );
  OR2_X1 U681 ( .A1(n1000), .A2(G868), .ZN(n606) );
  NAND2_X1 U682 ( .A1(n607), .A2(n606), .ZN(G284) );
  NAND2_X1 U683 ( .A1(G65), .A2(n589), .ZN(n609) );
  NAND2_X1 U684 ( .A1(G53), .A2(n650), .ZN(n608) );
  NAND2_X1 U685 ( .A1(n609), .A2(n608), .ZN(n613) );
  NAND2_X1 U686 ( .A1(G91), .A2(n637), .ZN(n611) );
  NAND2_X1 U687 ( .A1(G78), .A2(n635), .ZN(n610) );
  NAND2_X1 U688 ( .A1(n611), .A2(n610), .ZN(n612) );
  NOR2_X1 U689 ( .A1(n613), .A2(n612), .ZN(n1007) );
  XNOR2_X1 U690 ( .A(n1007), .B(KEYINPUT67), .ZN(G299) );
  NAND2_X1 U691 ( .A1(G286), .A2(G868), .ZN(n616) );
  INV_X1 U692 ( .A(G868), .ZN(n614) );
  NAND2_X1 U693 ( .A1(G299), .A2(n614), .ZN(n615) );
  NAND2_X1 U694 ( .A1(n616), .A2(n615), .ZN(G297) );
  INV_X1 U695 ( .A(G559), .ZN(n617) );
  NOR2_X1 U696 ( .A1(G860), .A2(n617), .ZN(n618) );
  XNOR2_X1 U697 ( .A(KEYINPUT73), .B(n618), .ZN(n619) );
  NAND2_X1 U698 ( .A1(n619), .A2(n1000), .ZN(n620) );
  XNOR2_X1 U699 ( .A(n620), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U700 ( .A1(n1000), .A2(G868), .ZN(n621) );
  NOR2_X1 U701 ( .A1(G559), .A2(n621), .ZN(n622) );
  XNOR2_X1 U702 ( .A(n622), .B(KEYINPUT74), .ZN(n624) );
  NOR2_X1 U703 ( .A1(n1013), .A2(G868), .ZN(n623) );
  NOR2_X1 U704 ( .A1(n624), .A2(n623), .ZN(n625) );
  XOR2_X1 U705 ( .A(KEYINPUT75), .B(n625), .Z(G282) );
  XNOR2_X1 U706 ( .A(n1013), .B(KEYINPUT78), .ZN(n627) );
  NAND2_X1 U707 ( .A1(n1000), .A2(G559), .ZN(n626) );
  XNOR2_X1 U708 ( .A(n627), .B(n626), .ZN(n661) );
  NOR2_X1 U709 ( .A1(G860), .A2(n661), .ZN(n634) );
  NAND2_X1 U710 ( .A1(G67), .A2(n589), .ZN(n629) );
  NAND2_X1 U711 ( .A1(G55), .A2(n650), .ZN(n628) );
  NAND2_X1 U712 ( .A1(n629), .A2(n628), .ZN(n633) );
  NAND2_X1 U713 ( .A1(G93), .A2(n637), .ZN(n631) );
  NAND2_X1 U714 ( .A1(G80), .A2(n635), .ZN(n630) );
  NAND2_X1 U715 ( .A1(n631), .A2(n630), .ZN(n632) );
  NOR2_X1 U716 ( .A1(n633), .A2(n632), .ZN(n657) );
  XNOR2_X1 U717 ( .A(n634), .B(n657), .ZN(G145) );
  NAND2_X1 U718 ( .A1(G73), .A2(n635), .ZN(n636) );
  XOR2_X1 U719 ( .A(KEYINPUT2), .B(n636), .Z(n642) );
  NAND2_X1 U720 ( .A1(G86), .A2(n637), .ZN(n639) );
  NAND2_X1 U721 ( .A1(G61), .A2(n589), .ZN(n638) );
  NAND2_X1 U722 ( .A1(n639), .A2(n638), .ZN(n640) );
  XOR2_X1 U723 ( .A(KEYINPUT81), .B(n640), .Z(n641) );
  NOR2_X1 U724 ( .A1(n642), .A2(n641), .ZN(n644) );
  NAND2_X1 U725 ( .A1(n650), .A2(G48), .ZN(n643) );
  NAND2_X1 U726 ( .A1(n644), .A2(n643), .ZN(G305) );
  NAND2_X1 U727 ( .A1(G74), .A2(G651), .ZN(n645) );
  XNOR2_X1 U728 ( .A(n645), .B(KEYINPUT80), .ZN(n648) );
  NAND2_X1 U729 ( .A1(n646), .A2(G87), .ZN(n647) );
  NAND2_X1 U730 ( .A1(n648), .A2(n647), .ZN(n649) );
  NOR2_X1 U731 ( .A1(n589), .A2(n649), .ZN(n653) );
  NAND2_X1 U732 ( .A1(G49), .A2(n650), .ZN(n651) );
  XOR2_X1 U733 ( .A(KEYINPUT79), .B(n651), .Z(n652) );
  NAND2_X1 U734 ( .A1(n653), .A2(n652), .ZN(G288) );
  NOR2_X1 U735 ( .A1(G868), .A2(n657), .ZN(n654) );
  XOR2_X1 U736 ( .A(n654), .B(KEYINPUT82), .Z(n664) );
  XNOR2_X1 U737 ( .A(G166), .B(KEYINPUT19), .ZN(n660) );
  XOR2_X1 U738 ( .A(G305), .B(G288), .Z(n655) );
  XNOR2_X1 U739 ( .A(G299), .B(n655), .ZN(n656) );
  XNOR2_X1 U740 ( .A(n657), .B(n656), .ZN(n658) );
  XNOR2_X1 U741 ( .A(n658), .B(G290), .ZN(n659) );
  XNOR2_X1 U742 ( .A(n660), .B(n659), .ZN(n900) );
  XNOR2_X1 U743 ( .A(n661), .B(n900), .ZN(n662) );
  NAND2_X1 U744 ( .A1(G868), .A2(n662), .ZN(n663) );
  NAND2_X1 U745 ( .A1(n664), .A2(n663), .ZN(G295) );
  NAND2_X1 U746 ( .A1(G2084), .A2(G2078), .ZN(n665) );
  XNOR2_X1 U747 ( .A(n665), .B(KEYINPUT83), .ZN(n666) );
  XNOR2_X1 U748 ( .A(KEYINPUT20), .B(n666), .ZN(n667) );
  NAND2_X1 U749 ( .A1(n667), .A2(G2090), .ZN(n668) );
  XNOR2_X1 U750 ( .A(n668), .B(KEYINPUT21), .ZN(n669) );
  XNOR2_X1 U751 ( .A(KEYINPUT84), .B(n669), .ZN(n670) );
  NAND2_X1 U752 ( .A1(n670), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U753 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U754 ( .A1(G69), .A2(G120), .ZN(n671) );
  NOR2_X1 U755 ( .A1(G237), .A2(n671), .ZN(n672) );
  NAND2_X1 U756 ( .A1(G108), .A2(n672), .ZN(n830) );
  NAND2_X1 U757 ( .A1(n830), .A2(G567), .ZN(n679) );
  XOR2_X1 U758 ( .A(KEYINPUT22), .B(KEYINPUT85), .Z(n674) );
  NAND2_X1 U759 ( .A1(G132), .A2(G82), .ZN(n673) );
  XNOR2_X1 U760 ( .A(n674), .B(n673), .ZN(n675) );
  NOR2_X1 U761 ( .A1(G218), .A2(n675), .ZN(n676) );
  NAND2_X1 U762 ( .A1(G96), .A2(n676), .ZN(n677) );
  XNOR2_X1 U763 ( .A(KEYINPUT86), .B(n677), .ZN(n831) );
  NAND2_X1 U764 ( .A1(G2106), .A2(n831), .ZN(n678) );
  NAND2_X1 U765 ( .A1(n679), .A2(n678), .ZN(n832) );
  NAND2_X1 U766 ( .A1(G661), .A2(G483), .ZN(n680) );
  NOR2_X1 U767 ( .A1(n832), .A2(n680), .ZN(n829) );
  NAND2_X1 U768 ( .A1(n829), .A2(G36), .ZN(G176) );
  INV_X1 U769 ( .A(G166), .ZN(G303) );
  INV_X1 U770 ( .A(KEYINPUT92), .ZN(n684) );
  XNOR2_X1 U771 ( .A(n788), .B(KEYINPUT87), .ZN(n682) );
  XNOR2_X1 U772 ( .A(n681), .B(KEYINPUT64), .ZN(n789) );
  NAND2_X1 U773 ( .A1(n682), .A2(n789), .ZN(n686) );
  AND2_X1 U774 ( .A1(G8), .A2(n686), .ZN(n683) );
  XNOR2_X2 U775 ( .A(n684), .B(n683), .ZN(n763) );
  AND2_X1 U776 ( .A1(n712), .A2(G1996), .ZN(n685) );
  XOR2_X1 U777 ( .A(n685), .B(KEYINPUT26), .Z(n696) );
  AND2_X1 U778 ( .A1(n689), .A2(G1341), .ZN(n687) );
  AND2_X1 U779 ( .A1(n695), .A2(n1000), .ZN(n688) );
  NAND2_X1 U780 ( .A1(n696), .A2(n688), .ZN(n693) );
  NOR2_X1 U781 ( .A1(n712), .A2(G1348), .ZN(n691) );
  NOR2_X1 U782 ( .A1(G2067), .A2(n689), .ZN(n690) );
  NOR2_X1 U783 ( .A1(n691), .A2(n690), .ZN(n692) );
  NAND2_X1 U784 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U785 ( .A(n694), .B(KEYINPUT94), .ZN(n699) );
  AND2_X1 U786 ( .A1(n696), .A2(n695), .ZN(n697) );
  OR2_X1 U787 ( .A1(n697), .A2(n1000), .ZN(n698) );
  NAND2_X1 U788 ( .A1(n699), .A2(n698), .ZN(n705) );
  XOR2_X1 U789 ( .A(KEYINPUT93), .B(KEYINPUT27), .Z(n701) );
  NAND2_X1 U790 ( .A1(G2072), .A2(n712), .ZN(n700) );
  XNOR2_X1 U791 ( .A(n701), .B(n700), .ZN(n703) );
  AND2_X1 U792 ( .A1(n689), .A2(G1956), .ZN(n702) );
  NOR2_X1 U793 ( .A1(n703), .A2(n702), .ZN(n706) );
  NAND2_X1 U794 ( .A1(n1007), .A2(n706), .ZN(n704) );
  NAND2_X1 U795 ( .A1(n705), .A2(n704), .ZN(n709) );
  NOR2_X1 U796 ( .A1(n1007), .A2(n706), .ZN(n707) );
  XOR2_X1 U797 ( .A(n707), .B(KEYINPUT28), .Z(n708) );
  NAND2_X1 U798 ( .A1(n709), .A2(n708), .ZN(n711) );
  NOR2_X1 U799 ( .A1(n712), .A2(G1961), .ZN(n714) );
  XOR2_X1 U800 ( .A(G2078), .B(KEYINPUT25), .Z(n956) );
  NOR2_X1 U801 ( .A1(n956), .A2(n689), .ZN(n713) );
  NOR2_X1 U802 ( .A1(n714), .A2(n713), .ZN(n721) );
  OR2_X1 U803 ( .A1(G301), .A2(n721), .ZN(n715) );
  NAND2_X1 U804 ( .A1(n716), .A2(n715), .ZN(n738) );
  NOR2_X1 U805 ( .A1(n763), .A2(G1966), .ZN(n726) );
  NOR2_X1 U806 ( .A1(G2084), .A2(n689), .ZN(n725) );
  NOR2_X1 U807 ( .A1(n726), .A2(n725), .ZN(n717) );
  AND2_X1 U808 ( .A1(n717), .A2(G8), .ZN(n718) );
  XNOR2_X1 U809 ( .A(n718), .B(KEYINPUT30), .ZN(n720) );
  INV_X1 U810 ( .A(G168), .ZN(n719) );
  NAND2_X1 U811 ( .A1(n720), .A2(n719), .ZN(n723) );
  NAND2_X1 U812 ( .A1(n721), .A2(G301), .ZN(n722) );
  NAND2_X1 U813 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U814 ( .A(n724), .B(KEYINPUT31), .ZN(n736) );
  AND2_X1 U815 ( .A1(n738), .A2(n736), .ZN(n729) );
  AND2_X1 U816 ( .A1(G8), .A2(n725), .ZN(n727) );
  OR2_X1 U817 ( .A1(n727), .A2(n726), .ZN(n728) );
  INV_X1 U818 ( .A(G8), .ZN(n735) );
  NOR2_X1 U819 ( .A1(n763), .A2(G1971), .ZN(n730) );
  XNOR2_X1 U820 ( .A(n730), .B(KEYINPUT96), .ZN(n732) );
  NOR2_X1 U821 ( .A1(n689), .A2(G2090), .ZN(n731) );
  NOR2_X1 U822 ( .A1(n732), .A2(n731), .ZN(n733) );
  NAND2_X1 U823 ( .A1(n733), .A2(G303), .ZN(n734) );
  OR2_X1 U824 ( .A1(n735), .A2(n734), .ZN(n739) );
  AND2_X1 U825 ( .A1(n736), .A2(n739), .ZN(n737) );
  NAND2_X1 U826 ( .A1(n738), .A2(n737), .ZN(n743) );
  INV_X1 U827 ( .A(n739), .ZN(n741) );
  AND2_X1 U828 ( .A1(G286), .A2(G8), .ZN(n740) );
  OR2_X1 U829 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U830 ( .A1(n743), .A2(n742), .ZN(n745) );
  XOR2_X1 U831 ( .A(KEYINPUT32), .B(KEYINPUT97), .Z(n744) );
  XNOR2_X1 U832 ( .A(n745), .B(n744), .ZN(n746) );
  NAND2_X1 U833 ( .A1(n747), .A2(n746), .ZN(n761) );
  NOR2_X1 U834 ( .A1(G1971), .A2(G303), .ZN(n748) );
  NOR2_X1 U835 ( .A1(G1976), .A2(G288), .ZN(n1003) );
  NOR2_X1 U836 ( .A1(n748), .A2(n1003), .ZN(n749) );
  NAND2_X1 U837 ( .A1(n761), .A2(n749), .ZN(n750) );
  NAND2_X1 U838 ( .A1(G1976), .A2(G288), .ZN(n1005) );
  NAND2_X1 U839 ( .A1(n750), .A2(n1005), .ZN(n751) );
  XNOR2_X1 U840 ( .A(KEYINPUT98), .B(n751), .ZN(n752) );
  NOR2_X1 U841 ( .A1(n763), .A2(n752), .ZN(n753) );
  NOR2_X1 U842 ( .A1(KEYINPUT33), .A2(n753), .ZN(n758) );
  AND2_X1 U843 ( .A1(n1003), .A2(KEYINPUT33), .ZN(n754) );
  INV_X1 U844 ( .A(n763), .ZN(n767) );
  NAND2_X1 U845 ( .A1(n754), .A2(n767), .ZN(n756) );
  XNOR2_X1 U846 ( .A(G1981), .B(G305), .ZN(n1021) );
  OR2_X1 U847 ( .A1(n758), .A2(n757), .ZN(n771) );
  NAND2_X1 U848 ( .A1(G8), .A2(G166), .ZN(n759) );
  NOR2_X1 U849 ( .A1(G2090), .A2(n759), .ZN(n760) );
  XNOR2_X1 U850 ( .A(KEYINPUT99), .B(n760), .ZN(n762) );
  NAND2_X1 U851 ( .A1(n762), .A2(n761), .ZN(n764) );
  NAND2_X1 U852 ( .A1(n764), .A2(n763), .ZN(n765) );
  NOR2_X1 U853 ( .A1(G1981), .A2(G305), .ZN(n766) );
  XNOR2_X1 U854 ( .A(n766), .B(KEYINPUT24), .ZN(n768) );
  NAND2_X1 U855 ( .A1(n768), .A2(n767), .ZN(n769) );
  NAND2_X1 U856 ( .A1(G119), .A2(n854), .ZN(n773) );
  NAND2_X1 U857 ( .A1(G107), .A2(n872), .ZN(n772) );
  NAND2_X1 U858 ( .A1(n773), .A2(n772), .ZN(n774) );
  XOR2_X1 U859 ( .A(KEYINPUT90), .B(n774), .Z(n778) );
  NAND2_X1 U860 ( .A1(G131), .A2(n876), .ZN(n776) );
  NAND2_X1 U861 ( .A1(G95), .A2(n879), .ZN(n775) );
  AND2_X1 U862 ( .A1(n776), .A2(n775), .ZN(n777) );
  NAND2_X1 U863 ( .A1(n778), .A2(n777), .ZN(n894) );
  NAND2_X1 U864 ( .A1(G1991), .A2(n894), .ZN(n787) );
  NAND2_X1 U865 ( .A1(G141), .A2(n876), .ZN(n780) );
  NAND2_X1 U866 ( .A1(G129), .A2(n854), .ZN(n779) );
  NAND2_X1 U867 ( .A1(n780), .A2(n779), .ZN(n783) );
  NAND2_X1 U868 ( .A1(n879), .A2(G105), .ZN(n781) );
  XOR2_X1 U869 ( .A(KEYINPUT38), .B(n781), .Z(n782) );
  NOR2_X1 U870 ( .A1(n783), .A2(n782), .ZN(n785) );
  NAND2_X1 U871 ( .A1(G117), .A2(n872), .ZN(n784) );
  NAND2_X1 U872 ( .A1(n785), .A2(n784), .ZN(n885) );
  NAND2_X1 U873 ( .A1(G1996), .A2(n885), .ZN(n786) );
  NAND2_X1 U874 ( .A1(n787), .A2(n786), .ZN(n975) );
  XOR2_X1 U875 ( .A(n788), .B(KEYINPUT87), .Z(n790) );
  NOR2_X1 U876 ( .A1(n790), .A2(n789), .ZN(n821) );
  NAND2_X1 U877 ( .A1(n975), .A2(n821), .ZN(n791) );
  XNOR2_X1 U878 ( .A(n791), .B(KEYINPUT91), .ZN(n813) );
  XNOR2_X1 U879 ( .A(G2067), .B(KEYINPUT37), .ZN(n792) );
  XNOR2_X1 U880 ( .A(n792), .B(KEYINPUT88), .ZN(n809) );
  NAND2_X1 U881 ( .A1(G140), .A2(n876), .ZN(n794) );
  NAND2_X1 U882 ( .A1(G104), .A2(n879), .ZN(n793) );
  NAND2_X1 U883 ( .A1(n794), .A2(n793), .ZN(n795) );
  XNOR2_X1 U884 ( .A(KEYINPUT34), .B(n795), .ZN(n801) );
  NAND2_X1 U885 ( .A1(G128), .A2(n854), .ZN(n797) );
  NAND2_X1 U886 ( .A1(G116), .A2(n872), .ZN(n796) );
  NAND2_X1 U887 ( .A1(n797), .A2(n796), .ZN(n798) );
  XNOR2_X1 U888 ( .A(KEYINPUT35), .B(n798), .ZN(n799) );
  XNOR2_X1 U889 ( .A(KEYINPUT89), .B(n799), .ZN(n800) );
  NOR2_X1 U890 ( .A1(n801), .A2(n800), .ZN(n802) );
  XNOR2_X1 U891 ( .A(KEYINPUT36), .B(n802), .ZN(n897) );
  NOR2_X1 U892 ( .A1(n809), .A2(n897), .ZN(n991) );
  NAND2_X1 U893 ( .A1(n821), .A2(n991), .ZN(n817) );
  NAND2_X1 U894 ( .A1(n805), .A2(n804), .ZN(n806) );
  XNOR2_X1 U895 ( .A(KEYINPUT101), .B(n806), .ZN(n808) );
  XNOR2_X1 U896 ( .A(G1986), .B(G290), .ZN(n1010) );
  NAND2_X1 U897 ( .A1(n1010), .A2(n821), .ZN(n807) );
  NAND2_X1 U898 ( .A1(n808), .A2(n807), .ZN(n824) );
  NAND2_X1 U899 ( .A1(n809), .A2(n897), .ZN(n980) );
  NOR2_X1 U900 ( .A1(G1996), .A2(n885), .ZN(n978) );
  NOR2_X1 U901 ( .A1(G1991), .A2(n894), .ZN(n971) );
  NOR2_X1 U902 ( .A1(G1986), .A2(G290), .ZN(n810) );
  XNOR2_X1 U903 ( .A(KEYINPUT102), .B(n810), .ZN(n811) );
  NOR2_X1 U904 ( .A1(n971), .A2(n811), .ZN(n812) );
  NOR2_X1 U905 ( .A1(n813), .A2(n812), .ZN(n814) );
  XOR2_X1 U906 ( .A(KEYINPUT103), .B(n814), .Z(n815) );
  NOR2_X1 U907 ( .A1(n978), .A2(n815), .ZN(n816) );
  XNOR2_X1 U908 ( .A(n816), .B(KEYINPUT39), .ZN(n818) );
  NAND2_X1 U909 ( .A1(n818), .A2(n817), .ZN(n819) );
  NAND2_X1 U910 ( .A1(n980), .A2(n819), .ZN(n820) );
  XNOR2_X1 U911 ( .A(KEYINPUT104), .B(n820), .ZN(n822) );
  NAND2_X1 U912 ( .A1(n822), .A2(n821), .ZN(n823) );
  NAND2_X1 U913 ( .A1(n824), .A2(n823), .ZN(n825) );
  XNOR2_X1 U914 ( .A(n825), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U915 ( .A1(G2106), .A2(n826), .ZN(G217) );
  AND2_X1 U916 ( .A1(G15), .A2(G2), .ZN(n827) );
  NAND2_X1 U917 ( .A1(G661), .A2(n827), .ZN(G259) );
  NAND2_X1 U918 ( .A1(G3), .A2(G1), .ZN(n828) );
  NAND2_X1 U919 ( .A1(n829), .A2(n828), .ZN(G188) );
  INV_X1 U921 ( .A(G132), .ZN(G219) );
  INV_X1 U922 ( .A(G120), .ZN(G236) );
  INV_X1 U923 ( .A(G96), .ZN(G221) );
  INV_X1 U924 ( .A(G82), .ZN(G220) );
  INV_X1 U925 ( .A(G69), .ZN(G235) );
  NOR2_X1 U926 ( .A1(n831), .A2(n830), .ZN(G325) );
  INV_X1 U927 ( .A(G325), .ZN(G261) );
  INV_X1 U928 ( .A(n832), .ZN(G319) );
  XOR2_X1 U929 ( .A(KEYINPUT42), .B(KEYINPUT108), .Z(n834) );
  XNOR2_X1 U930 ( .A(KEYINPUT106), .B(G2096), .ZN(n833) );
  XNOR2_X1 U931 ( .A(n834), .B(n833), .ZN(n835) );
  XOR2_X1 U932 ( .A(n835), .B(KEYINPUT107), .Z(n837) );
  XNOR2_X1 U933 ( .A(G2067), .B(G2072), .ZN(n836) );
  XNOR2_X1 U934 ( .A(n837), .B(n836), .ZN(n841) );
  XOR2_X1 U935 ( .A(G2100), .B(G2090), .Z(n839) );
  XNOR2_X1 U936 ( .A(G2078), .B(G2084), .ZN(n838) );
  XNOR2_X1 U937 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U938 ( .A(n841), .B(n840), .Z(n843) );
  XNOR2_X1 U939 ( .A(G2678), .B(KEYINPUT43), .ZN(n842) );
  XNOR2_X1 U940 ( .A(n843), .B(n842), .ZN(G227) );
  XOR2_X1 U941 ( .A(G1961), .B(G1956), .Z(n845) );
  XNOR2_X1 U942 ( .A(G1976), .B(G1971), .ZN(n844) );
  XNOR2_X1 U943 ( .A(n845), .B(n844), .ZN(n849) );
  XOR2_X1 U944 ( .A(G1966), .B(G1981), .Z(n847) );
  XNOR2_X1 U945 ( .A(G1996), .B(G1991), .ZN(n846) );
  XNOR2_X1 U946 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U947 ( .A(n849), .B(n848), .Z(n851) );
  XNOR2_X1 U948 ( .A(KEYINPUT109), .B(KEYINPUT41), .ZN(n850) );
  XNOR2_X1 U949 ( .A(n851), .B(n850), .ZN(n853) );
  XOR2_X1 U950 ( .A(G1986), .B(G2474), .Z(n852) );
  XNOR2_X1 U951 ( .A(n853), .B(n852), .ZN(G229) );
  NAND2_X1 U952 ( .A1(n854), .A2(G124), .ZN(n855) );
  XNOR2_X1 U953 ( .A(n855), .B(KEYINPUT44), .ZN(n857) );
  NAND2_X1 U954 ( .A1(G112), .A2(n872), .ZN(n856) );
  NAND2_X1 U955 ( .A1(n857), .A2(n856), .ZN(n861) );
  NAND2_X1 U956 ( .A1(G136), .A2(n876), .ZN(n859) );
  NAND2_X1 U957 ( .A1(G100), .A2(n879), .ZN(n858) );
  NAND2_X1 U958 ( .A1(n859), .A2(n858), .ZN(n860) );
  NOR2_X1 U959 ( .A1(n861), .A2(n860), .ZN(G162) );
  NAND2_X1 U960 ( .A1(G118), .A2(n872), .ZN(n862) );
  XNOR2_X1 U961 ( .A(n862), .B(KEYINPUT110), .ZN(n864) );
  NAND2_X1 U962 ( .A1(G130), .A2(n854), .ZN(n863) );
  NAND2_X1 U963 ( .A1(n864), .A2(n863), .ZN(n870) );
  XNOR2_X1 U964 ( .A(KEYINPUT45), .B(KEYINPUT111), .ZN(n868) );
  NAND2_X1 U965 ( .A1(G142), .A2(n876), .ZN(n866) );
  NAND2_X1 U966 ( .A1(G106), .A2(n879), .ZN(n865) );
  NAND2_X1 U967 ( .A1(n866), .A2(n865), .ZN(n867) );
  XNOR2_X1 U968 ( .A(n868), .B(n867), .ZN(n869) );
  NOR2_X1 U969 ( .A1(n870), .A2(n869), .ZN(n896) );
  NAND2_X1 U970 ( .A1(n854), .A2(G127), .ZN(n871) );
  XNOR2_X1 U971 ( .A(n871), .B(KEYINPUT114), .ZN(n874) );
  NAND2_X1 U972 ( .A1(G115), .A2(n872), .ZN(n873) );
  NAND2_X1 U973 ( .A1(n874), .A2(n873), .ZN(n875) );
  XNOR2_X1 U974 ( .A(n875), .B(KEYINPUT47), .ZN(n878) );
  NAND2_X1 U975 ( .A1(G139), .A2(n876), .ZN(n877) );
  NAND2_X1 U976 ( .A1(n878), .A2(n877), .ZN(n882) );
  NAND2_X1 U977 ( .A1(G103), .A2(n879), .ZN(n880) );
  XNOR2_X1 U978 ( .A(KEYINPUT113), .B(n880), .ZN(n881) );
  NOR2_X1 U979 ( .A1(n882), .A2(n881), .ZN(n982) );
  XOR2_X1 U980 ( .A(n982), .B(G162), .Z(n883) );
  XNOR2_X1 U981 ( .A(n972), .B(n883), .ZN(n887) );
  XOR2_X1 U982 ( .A(G164), .B(G160), .Z(n884) );
  XNOR2_X1 U983 ( .A(n885), .B(n884), .ZN(n886) );
  XOR2_X1 U984 ( .A(n887), .B(n886), .Z(n892) );
  XOR2_X1 U985 ( .A(KEYINPUT112), .B(KEYINPUT48), .Z(n889) );
  XNOR2_X1 U986 ( .A(KEYINPUT46), .B(KEYINPUT116), .ZN(n888) );
  XNOR2_X1 U987 ( .A(n889), .B(n888), .ZN(n890) );
  XNOR2_X1 U988 ( .A(KEYINPUT115), .B(n890), .ZN(n891) );
  XNOR2_X1 U989 ( .A(n892), .B(n891), .ZN(n893) );
  XOR2_X1 U990 ( .A(n894), .B(n893), .Z(n895) );
  XNOR2_X1 U991 ( .A(n896), .B(n895), .ZN(n898) );
  XOR2_X1 U992 ( .A(n898), .B(n897), .Z(n899) );
  NOR2_X1 U993 ( .A1(G37), .A2(n899), .ZN(G395) );
  XNOR2_X1 U994 ( .A(G286), .B(n1013), .ZN(n901) );
  XNOR2_X1 U995 ( .A(n901), .B(n900), .ZN(n903) );
  XOR2_X1 U996 ( .A(G171), .B(n1000), .Z(n902) );
  XNOR2_X1 U997 ( .A(n903), .B(n902), .ZN(n904) );
  NOR2_X1 U998 ( .A1(G37), .A2(n904), .ZN(G397) );
  XOR2_X1 U999 ( .A(KEYINPUT105), .B(G2427), .Z(n906) );
  XNOR2_X1 U1000 ( .A(G2435), .B(G2438), .ZN(n905) );
  XNOR2_X1 U1001 ( .A(n906), .B(n905), .ZN(n913) );
  XOR2_X1 U1002 ( .A(G2443), .B(G2430), .Z(n908) );
  XNOR2_X1 U1003 ( .A(G2454), .B(G2446), .ZN(n907) );
  XNOR2_X1 U1004 ( .A(n908), .B(n907), .ZN(n909) );
  XOR2_X1 U1005 ( .A(n909), .B(G2451), .Z(n911) );
  XNOR2_X1 U1006 ( .A(G1341), .B(G1348), .ZN(n910) );
  XNOR2_X1 U1007 ( .A(n911), .B(n910), .ZN(n912) );
  XNOR2_X1 U1008 ( .A(n913), .B(n912), .ZN(n914) );
  NAND2_X1 U1009 ( .A1(n914), .A2(G14), .ZN(n920) );
  NAND2_X1 U1010 ( .A1(G319), .A2(n920), .ZN(n917) );
  NOR2_X1 U1011 ( .A1(G227), .A2(G229), .ZN(n915) );
  XNOR2_X1 U1012 ( .A(KEYINPUT49), .B(n915), .ZN(n916) );
  NOR2_X1 U1013 ( .A1(n917), .A2(n916), .ZN(n919) );
  NOR2_X1 U1014 ( .A1(G395), .A2(G397), .ZN(n918) );
  NAND2_X1 U1015 ( .A1(n919), .A2(n918), .ZN(G225) );
  INV_X1 U1016 ( .A(G225), .ZN(G308) );
  INV_X1 U1017 ( .A(G108), .ZN(G238) );
  INV_X1 U1018 ( .A(n920), .ZN(G401) );
  XOR2_X1 U1019 ( .A(KEYINPUT60), .B(KEYINPUT126), .Z(n931) );
  XNOR2_X1 U1020 ( .A(KEYINPUT59), .B(G1348), .ZN(n921) );
  XNOR2_X1 U1021 ( .A(n921), .B(G4), .ZN(n929) );
  XNOR2_X1 U1022 ( .A(G1956), .B(G20), .ZN(n927) );
  XNOR2_X1 U1023 ( .A(G1981), .B(G6), .ZN(n922) );
  XNOR2_X1 U1024 ( .A(n922), .B(KEYINPUT124), .ZN(n924) );
  XNOR2_X1 U1025 ( .A(G19), .B(G1341), .ZN(n923) );
  NOR2_X1 U1026 ( .A1(n924), .A2(n923), .ZN(n925) );
  XNOR2_X1 U1027 ( .A(KEYINPUT125), .B(n925), .ZN(n926) );
  NOR2_X1 U1028 ( .A1(n927), .A2(n926), .ZN(n928) );
  NAND2_X1 U1029 ( .A1(n929), .A2(n928), .ZN(n930) );
  XNOR2_X1 U1030 ( .A(n931), .B(n930), .ZN(n935) );
  XNOR2_X1 U1031 ( .A(G1966), .B(G21), .ZN(n933) );
  XNOR2_X1 U1032 ( .A(G1961), .B(G5), .ZN(n932) );
  NOR2_X1 U1033 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1034 ( .A1(n935), .A2(n934), .ZN(n943) );
  XNOR2_X1 U1035 ( .A(G1986), .B(G24), .ZN(n937) );
  XNOR2_X1 U1036 ( .A(G22), .B(G1971), .ZN(n936) );
  NOR2_X1 U1037 ( .A1(n937), .A2(n936), .ZN(n940) );
  XNOR2_X1 U1038 ( .A(G1976), .B(KEYINPUT127), .ZN(n938) );
  XNOR2_X1 U1039 ( .A(n938), .B(G23), .ZN(n939) );
  NAND2_X1 U1040 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1041 ( .A(KEYINPUT58), .B(n941), .ZN(n942) );
  NOR2_X1 U1042 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1043 ( .A(KEYINPUT61), .B(n944), .ZN(n946) );
  INV_X1 U1044 ( .A(G16), .ZN(n945) );
  NAND2_X1 U1045 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1046 ( .A1(n947), .A2(G11), .ZN(n999) );
  XOR2_X1 U1047 ( .A(KEYINPUT120), .B(G34), .Z(n949) );
  XNOR2_X1 U1048 ( .A(G2084), .B(KEYINPUT54), .ZN(n948) );
  XNOR2_X1 U1049 ( .A(n949), .B(n948), .ZN(n966) );
  XNOR2_X1 U1050 ( .A(G2090), .B(G35), .ZN(n964) );
  XOR2_X1 U1051 ( .A(G2067), .B(G26), .Z(n955) );
  XOR2_X1 U1052 ( .A(G2072), .B(G33), .Z(n950) );
  NAND2_X1 U1053 ( .A1(n950), .A2(G28), .ZN(n953) );
  XNOR2_X1 U1054 ( .A(G25), .B(G1991), .ZN(n951) );
  XNOR2_X1 U1055 ( .A(KEYINPUT118), .B(n951), .ZN(n952) );
  NOR2_X1 U1056 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1057 ( .A1(n955), .A2(n954), .ZN(n961) );
  XNOR2_X1 U1058 ( .A(G1996), .B(G32), .ZN(n958) );
  XNOR2_X1 U1059 ( .A(n956), .B(G27), .ZN(n957) );
  NOR2_X1 U1060 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1061 ( .A(n959), .B(KEYINPUT119), .ZN(n960) );
  NOR2_X1 U1062 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1063 ( .A(KEYINPUT53), .B(n962), .ZN(n963) );
  NOR2_X1 U1064 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1065 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1066 ( .A(KEYINPUT55), .B(n967), .ZN(n968) );
  NOR2_X1 U1067 ( .A1(G29), .A2(n968), .ZN(n969) );
  XNOR2_X1 U1068 ( .A(n969), .B(KEYINPUT121), .ZN(n997) );
  XOR2_X1 U1069 ( .A(G160), .B(G2084), .Z(n970) );
  NOR2_X1 U1070 ( .A1(n971), .A2(n970), .ZN(n973) );
  NAND2_X1 U1071 ( .A1(n973), .A2(n972), .ZN(n974) );
  NOR2_X1 U1072 ( .A1(n975), .A2(n974), .ZN(n989) );
  XNOR2_X1 U1073 ( .A(G2090), .B(G162), .ZN(n976) );
  XNOR2_X1 U1074 ( .A(n976), .B(KEYINPUT117), .ZN(n977) );
  NOR2_X1 U1075 ( .A1(n978), .A2(n977), .ZN(n979) );
  XOR2_X1 U1076 ( .A(KEYINPUT51), .B(n979), .Z(n981) );
  NAND2_X1 U1077 ( .A1(n981), .A2(n980), .ZN(n987) );
  XOR2_X1 U1078 ( .A(G2072), .B(n982), .Z(n984) );
  XOR2_X1 U1079 ( .A(G164), .B(G2078), .Z(n983) );
  NOR2_X1 U1080 ( .A1(n984), .A2(n983), .ZN(n985) );
  XOR2_X1 U1081 ( .A(KEYINPUT50), .B(n985), .Z(n986) );
  NOR2_X1 U1082 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1083 ( .A1(n989), .A2(n988), .ZN(n990) );
  NOR2_X1 U1084 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1085 ( .A(n992), .B(KEYINPUT52), .ZN(n994) );
  INV_X1 U1086 ( .A(KEYINPUT55), .ZN(n993) );
  NAND2_X1 U1087 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1088 ( .A1(G29), .A2(n995), .ZN(n996) );
  NAND2_X1 U1089 ( .A1(n997), .A2(n996), .ZN(n998) );
  NOR2_X1 U1090 ( .A1(n999), .A2(n998), .ZN(n1028) );
  XNOR2_X1 U1091 ( .A(KEYINPUT56), .B(G16), .ZN(n1026) );
  XNOR2_X1 U1092 ( .A(G171), .B(G1961), .ZN(n1002) );
  XNOR2_X1 U1093 ( .A(n1000), .B(G1348), .ZN(n1001) );
  NAND2_X1 U1094 ( .A1(n1002), .A2(n1001), .ZN(n1019) );
  INV_X1 U1095 ( .A(n1003), .ZN(n1004) );
  NAND2_X1 U1096 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1097 ( .A(n1006), .B(KEYINPUT123), .ZN(n1017) );
  XNOR2_X1 U1098 ( .A(G1956), .B(n1007), .ZN(n1008) );
  XNOR2_X1 U1099 ( .A(n1008), .B(KEYINPUT122), .ZN(n1012) );
  XOR2_X1 U1100 ( .A(G1971), .B(G166), .Z(n1009) );
  NOR2_X1 U1101 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1102 ( .A1(n1012), .A2(n1011), .ZN(n1015) );
  XNOR2_X1 U1103 ( .A(G1341), .B(n1013), .ZN(n1014) );
  NOR2_X1 U1104 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1105 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NOR2_X1 U1106 ( .A1(n1019), .A2(n1018), .ZN(n1024) );
  XOR2_X1 U1107 ( .A(G1966), .B(G168), .Z(n1020) );
  NOR2_X1 U1108 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XOR2_X1 U1109 ( .A(KEYINPUT57), .B(n1022), .Z(n1023) );
  NAND2_X1 U1110 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1111 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1112 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XOR2_X1 U1113 ( .A(KEYINPUT62), .B(n1029), .Z(G311) );
  INV_X1 U1114 ( .A(G311), .ZN(G150) );
endmodule

