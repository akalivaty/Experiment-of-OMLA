//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 1 0 1 1 0 1 1 1 0 0 1 1 0 1 0 1 1 1 0 0 1 0 0 1 1 0 1 0 0 0 0 1 0 1 1 0 1 0 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:21 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1230,
    new_n1231, new_n1232, new_n1234, new_n1235, new_n1236, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT64), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n210), .B1(new_n216), .B2(new_n219), .ZN(new_n220));
  OR2_X1    g0020(.A1(new_n220), .A2(KEYINPUT1), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n203), .A2(G50), .ZN(new_n222));
  XOR2_X1   g0022(.A(new_n222), .B(KEYINPUT65), .Z(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G13), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n224), .A2(new_n208), .ZN(new_n225));
  INV_X1    g0025(.A(new_n225), .ZN(new_n226));
  OR2_X1    g0026(.A1(new_n223), .A2(new_n226), .ZN(new_n227));
  NAND3_X1  g0027(.A1(new_n213), .A2(new_n221), .A3(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n220), .ZN(G361));
  XNOR2_X1  g0029(.A(G250), .B(G257), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT66), .ZN(new_n231));
  XOR2_X1   g0031(.A(G264), .B(G270), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  INV_X1    g0034(.A(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n233), .B(new_n238), .ZN(G358));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XOR2_X1   g0040(.A(G107), .B(G116), .Z(new_n241));
  XOR2_X1   g0041(.A(new_n240), .B(new_n241), .Z(new_n242));
  XOR2_X1   g0042(.A(new_n242), .B(KEYINPUT67), .Z(new_n243));
  INV_X1    g0043(.A(G50), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n244), .A2(G68), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n202), .A2(G50), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G58), .B(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n243), .B(new_n249), .ZN(G351));
  INV_X1    g0050(.A(KEYINPUT74), .ZN(new_n251));
  NAND3_X1  g0051(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(new_n224), .ZN(new_n253));
  AND3_X1   g0053(.A1(KEYINPUT68), .A2(KEYINPUT8), .A3(G58), .ZN(new_n254));
  AOI21_X1  g0054(.A(KEYINPUT8), .B1(KEYINPUT68), .B2(G58), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n208), .A2(G33), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  OAI21_X1  g0059(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n260));
  INV_X1    g0060(.A(G150), .ZN(new_n261));
  NOR2_X1   g0061(.A1(G20), .A2(G33), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n260), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n253), .B1(new_n259), .B2(new_n264), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n207), .A2(G13), .A3(G20), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n266), .A2(G50), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n253), .B1(new_n207), .B2(G20), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n267), .B1(new_n268), .B2(G50), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n265), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT9), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n265), .A2(KEYINPUT9), .A3(new_n269), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT69), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(KEYINPUT10), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n272), .A2(new_n273), .A3(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n274), .A2(KEYINPUT10), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G41), .ZN(new_n280));
  INV_X1    g0080(.A(G45), .ZN(new_n281));
  AOI21_X1  g0081(.A(G1), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(G33), .A2(G41), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n283), .A2(G1), .A3(G13), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n282), .A2(new_n284), .A3(G274), .ZN(new_n285));
  INV_X1    g0085(.A(G226), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n284), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n285), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  XNOR2_X1  g0089(.A(KEYINPUT3), .B(G33), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n290), .A2(G223), .A3(G1698), .ZN(new_n291));
  INV_X1    g0091(.A(G77), .ZN(new_n292));
  INV_X1    g0092(.A(G1698), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n290), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G222), .ZN(new_n295));
  OAI221_X1 g0095(.A(new_n291), .B1(new_n292), .B2(new_n290), .C1(new_n294), .C2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n284), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n289), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(G190), .ZN(new_n299));
  INV_X1    g0099(.A(new_n298), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(G200), .ZN(new_n301));
  NAND4_X1  g0101(.A1(new_n277), .A2(new_n279), .A3(new_n299), .A4(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n299), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n278), .B1(new_n303), .B2(new_n276), .ZN(new_n304));
  AND2_X1   g0104(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n286), .A2(new_n293), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n235), .A2(G1698), .ZN(new_n307));
  AND2_X1   g0107(.A1(KEYINPUT3), .A2(G33), .ZN(new_n308));
  NOR2_X1   g0108(.A1(KEYINPUT3), .A2(G33), .ZN(new_n309));
  OAI211_X1 g0109(.A(new_n306), .B(new_n307), .C1(new_n308), .C2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(G33), .A2(G97), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(new_n297), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n284), .A2(G238), .A3(new_n287), .ZN(new_n314));
  AND2_X1   g0114(.A1(new_n285), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT13), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n313), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT70), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n284), .B1(new_n310), .B2(new_n311), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n285), .A2(new_n314), .ZN(new_n320));
  OAI21_X1  g0120(.A(KEYINPUT13), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n317), .A2(new_n318), .A3(new_n321), .ZN(new_n322));
  OAI211_X1 g0122(.A(KEYINPUT70), .B(KEYINPUT13), .C1(new_n319), .C2(new_n320), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n322), .A2(G169), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(KEYINPUT14), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT14), .ZN(new_n326));
  NAND4_X1  g0126(.A1(new_n322), .A2(new_n326), .A3(G169), .A4(new_n323), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n317), .A2(G179), .A3(new_n321), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n325), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n266), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(new_n202), .ZN(new_n331));
  OAI21_X1  g0131(.A(KEYINPUT12), .B1(new_n331), .B2(KEYINPUT71), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(KEYINPUT71), .ZN(new_n333));
  XNOR2_X1  g0133(.A(new_n332), .B(new_n333), .ZN(new_n334));
  AOI22_X1  g0134(.A1(new_n262), .A2(G50), .B1(G20), .B2(new_n202), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n335), .B1(new_n292), .B2(new_n258), .ZN(new_n336));
  AOI21_X1  g0136(.A(KEYINPUT11), .B1(new_n336), .B2(new_n253), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n337), .B1(G68), .B2(new_n268), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n336), .A2(KEYINPUT11), .A3(new_n253), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n334), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n329), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(G169), .ZN(new_n342));
  AOI22_X1  g0142(.A1(new_n300), .A2(new_n342), .B1(new_n265), .B2(new_n269), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n343), .B1(G179), .B2(new_n300), .ZN(new_n344));
  INV_X1    g0144(.A(new_n340), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n317), .A2(G190), .A3(new_n321), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n322), .A2(G200), .A3(new_n323), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n290), .A2(G238), .A3(G1698), .ZN(new_n351));
  INV_X1    g0151(.A(G107), .ZN(new_n352));
  OAI221_X1 g0152(.A(new_n351), .B1(new_n352), .B2(new_n290), .C1(new_n294), .C2(new_n235), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(new_n297), .ZN(new_n354));
  INV_X1    g0154(.A(G244), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n285), .B1(new_n355), .B2(new_n288), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n354), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(new_n342), .ZN(new_n359));
  XNOR2_X1  g0159(.A(KEYINPUT8), .B(G58), .ZN(new_n360));
  OAI22_X1  g0160(.A1(new_n360), .A2(new_n263), .B1(new_n208), .B2(new_n292), .ZN(new_n361));
  XNOR2_X1  g0161(.A(KEYINPUT15), .B(G87), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n362), .A2(new_n258), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n253), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n268), .A2(G77), .ZN(new_n365));
  OAI211_X1 g0165(.A(new_n364), .B(new_n365), .C1(G77), .C2(new_n266), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n356), .B1(new_n353), .B2(new_n297), .ZN(new_n367));
  INV_X1    g0167(.A(G179), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n359), .A2(new_n366), .A3(new_n369), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n366), .B1(new_n367), .B2(G190), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n358), .A2(G200), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n370), .A2(new_n373), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n350), .A2(new_n374), .ZN(new_n375));
  NAND4_X1  g0175(.A1(new_n305), .A2(new_n341), .A3(new_n344), .A4(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT16), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT72), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n262), .A2(G159), .ZN(new_n379));
  NAND2_X1  g0179(.A1(G58), .A2(G68), .ZN(new_n380));
  AND2_X1   g0180(.A1(new_n203), .A2(new_n380), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n378), .B(new_n379), .C1(new_n381), .C2(new_n208), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n208), .B1(new_n203), .B2(new_n380), .ZN(new_n383));
  INV_X1    g0183(.A(new_n379), .ZN(new_n384));
  OAI21_X1  g0184(.A(KEYINPUT72), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n382), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT7), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n387), .B1(new_n290), .B2(G20), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n308), .A2(new_n309), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n389), .A2(KEYINPUT7), .A3(new_n208), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n202), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n377), .B1(new_n386), .B2(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(KEYINPUT7), .B1(new_n389), .B2(new_n208), .ZN(new_n393));
  NOR4_X1   g0193(.A1(new_n308), .A2(new_n309), .A3(new_n387), .A4(G20), .ZN(new_n394));
  OAI21_X1  g0194(.A(G68), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n395), .A2(KEYINPUT16), .A3(new_n382), .A4(new_n385), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n392), .A2(new_n396), .A3(new_n253), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n256), .A2(new_n266), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n398), .B1(new_n256), .B2(new_n268), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  OAI211_X1 g0200(.A(G223), .B(new_n293), .C1(new_n308), .C2(new_n309), .ZN(new_n401));
  OAI211_X1 g0201(.A(G226), .B(G1698), .C1(new_n308), .C2(new_n309), .ZN(new_n402));
  INV_X1    g0202(.A(G33), .ZN(new_n403));
  INV_X1    g0203(.A(G87), .ZN(new_n404));
  OAI211_X1 g0204(.A(new_n401), .B(new_n402), .C1(new_n403), .C2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(new_n297), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(new_n368), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n284), .A2(G232), .A3(new_n287), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n285), .A2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT73), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n285), .A2(new_n408), .A3(KEYINPUT73), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n409), .B1(new_n405), .B2(new_n297), .ZN(new_n414));
  OAI22_X1  g0214(.A1(new_n407), .A2(new_n413), .B1(new_n414), .B2(G169), .ZN(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n400), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(KEYINPUT18), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n415), .B1(new_n397), .B2(new_n399), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT18), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(G190), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n406), .A2(new_n422), .ZN(new_n423));
  OAI22_X1  g0223(.A1(new_n423), .A2(new_n413), .B1(new_n414), .B2(G200), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n397), .A2(new_n424), .A3(new_n399), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT17), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n397), .A2(new_n424), .A3(KEYINPUT17), .A4(new_n399), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n418), .A2(new_n421), .A3(new_n427), .A4(new_n428), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n251), .B1(new_n376), .B2(new_n429), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n302), .A2(new_n304), .A3(new_n344), .ZN(new_n431));
  NOR3_X1   g0231(.A1(new_n431), .A2(new_n350), .A3(new_n374), .ZN(new_n432));
  INV_X1    g0232(.A(new_n429), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n432), .A2(new_n433), .A3(KEYINPUT74), .A4(new_n341), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n430), .A2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT6), .ZN(new_n436));
  INV_X1    g0236(.A(G97), .ZN(new_n437));
  NOR3_X1   g0237(.A1(new_n436), .A2(new_n437), .A3(G107), .ZN(new_n438));
  XNOR2_X1  g0238(.A(G97), .B(G107), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n438), .B1(new_n436), .B2(new_n439), .ZN(new_n440));
  OAI22_X1  g0240(.A1(new_n440), .A2(new_n208), .B1(new_n292), .B2(new_n263), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n352), .B1(new_n388), .B2(new_n390), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n253), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT75), .ZN(new_n444));
  NOR3_X1   g0244(.A1(new_n266), .A2(new_n444), .A3(G97), .ZN(new_n445));
  AOI21_X1  g0245(.A(KEYINPUT75), .B1(new_n330), .B2(new_n437), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n207), .A2(G33), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n266), .A2(new_n447), .A3(new_n224), .A4(new_n252), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  AOI211_X1 g0249(.A(new_n445), .B(new_n446), .C1(G97), .C2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT76), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n443), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n451), .B1(new_n443), .B2(new_n450), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  XNOR2_X1  g0255(.A(KEYINPUT5), .B(G41), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n207), .A2(G45), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n224), .ZN(new_n459));
  AOI22_X1  g0259(.A1(new_n456), .A2(new_n458), .B1(new_n459), .B2(new_n283), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(G257), .ZN(new_n461));
  OR2_X1    g0261(.A1(KEYINPUT5), .A2(G41), .ZN(new_n462));
  NAND2_X1  g0262(.A1(KEYINPUT5), .A2(G41), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n457), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(G274), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n465), .B1(new_n459), .B2(new_n283), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n461), .A2(new_n467), .ZN(new_n468));
  OAI211_X1 g0268(.A(G250), .B(G1698), .C1(new_n308), .C2(new_n309), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT77), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n290), .A2(KEYINPUT77), .A3(G250), .A4(G1698), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n290), .A2(KEYINPUT4), .A3(G244), .A4(new_n293), .ZN(new_n474));
  NAND2_X1  g0274(.A1(G33), .A2(G283), .ZN(new_n475));
  OAI211_X1 g0275(.A(G244), .B(new_n293), .C1(new_n308), .C2(new_n309), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT4), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n473), .A2(new_n474), .A3(new_n475), .A4(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n468), .B1(new_n479), .B2(new_n297), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(new_n422), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n481), .B1(G200), .B2(new_n480), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n443), .A2(new_n450), .ZN(new_n483));
  AND2_X1   g0283(.A1(new_n471), .A2(new_n472), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n478), .A2(new_n474), .A3(new_n475), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n297), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(new_n468), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n486), .A2(G179), .A3(new_n487), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n488), .B1(new_n480), .B2(new_n342), .ZN(new_n489));
  AOI22_X1  g0289(.A1(new_n455), .A2(new_n482), .B1(new_n483), .B2(new_n489), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n208), .B(G68), .C1(new_n308), .C2(new_n309), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT19), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n492), .B1(new_n258), .B2(new_n437), .ZN(new_n493));
  NAND3_X1  g0293(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n494));
  NOR2_X1   g0294(.A1(G97), .A2(G107), .ZN(new_n495));
  AOI22_X1  g0295(.A1(new_n208), .A2(new_n494), .B1(new_n495), .B2(new_n404), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT78), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n491), .B(new_n493), .C1(new_n496), .C2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n494), .A2(new_n208), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n495), .A2(new_n404), .ZN(new_n500));
  AND3_X1   g0300(.A1(new_n499), .A2(new_n500), .A3(new_n497), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n253), .B1(new_n498), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n362), .A2(new_n330), .ZN(new_n503));
  AND3_X1   g0303(.A1(new_n502), .A2(KEYINPUT79), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g0304(.A(KEYINPUT79), .B1(new_n502), .B2(new_n503), .ZN(new_n505));
  OAI22_X1  g0305(.A1(new_n504), .A2(new_n505), .B1(new_n404), .B2(new_n448), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n466), .A2(new_n458), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n284), .A2(G250), .A3(new_n457), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  OAI211_X1 g0309(.A(G238), .B(new_n293), .C1(new_n308), .C2(new_n309), .ZN(new_n510));
  OAI211_X1 g0310(.A(G244), .B(G1698), .C1(new_n308), .C2(new_n309), .ZN(new_n511));
  NAND2_X1  g0311(.A1(G33), .A2(G116), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n509), .B1(new_n297), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(G190), .ZN(new_n515));
  INV_X1    g0315(.A(G200), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n515), .B1(new_n516), .B2(new_n514), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n506), .A2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(new_n362), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n449), .A2(new_n519), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n520), .B1(new_n504), .B2(new_n505), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(KEYINPUT80), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT80), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n523), .B(new_n520), .C1(new_n504), .C2(new_n505), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n514), .A2(G169), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n526), .B1(new_n368), .B2(new_n514), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n518), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  OAI211_X1 g0328(.A(G257), .B(G1698), .C1(new_n308), .C2(new_n309), .ZN(new_n529));
  OAI211_X1 g0329(.A(G250), .B(new_n293), .C1(new_n308), .C2(new_n309), .ZN(new_n530));
  NAND2_X1  g0330(.A1(G33), .A2(G294), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n529), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  AOI22_X1  g0332(.A1(new_n532), .A2(new_n297), .B1(new_n460), .B2(G264), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n533), .A2(new_n368), .A3(new_n467), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n467), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n342), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n208), .B(G87), .C1(new_n308), .C2(new_n309), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(KEYINPUT22), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT22), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n290), .A2(new_n539), .A3(new_n208), .A4(G87), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n512), .A2(G20), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT23), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n543), .B1(new_n208), .B2(G107), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n352), .A2(KEYINPUT23), .A3(G20), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n542), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n541), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(KEYINPUT24), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT24), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n541), .A2(new_n549), .A3(new_n546), .ZN(new_n550));
  AOI22_X1  g0350(.A1(new_n548), .A2(new_n550), .B1(new_n224), .B2(new_n252), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n330), .A2(KEYINPUT25), .A3(new_n352), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(KEYINPUT82), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT25), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n554), .B1(new_n266), .B2(G107), .ZN(new_n555));
  OR2_X1    g0355(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n553), .A2(new_n555), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n449), .A2(G107), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n534), .B(new_n536), .C1(new_n551), .C2(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT81), .ZN(new_n562));
  INV_X1    g0362(.A(G116), .ZN(new_n563));
  AOI22_X1  g0363(.A1(new_n252), .A2(new_n224), .B1(G20), .B2(new_n563), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n475), .B(new_n208), .C1(G33), .C2(new_n437), .ZN(new_n565));
  AND3_X1   g0365(.A1(new_n564), .A2(KEYINPUT20), .A3(new_n565), .ZN(new_n566));
  AOI21_X1  g0366(.A(KEYINPUT20), .B1(new_n564), .B2(new_n565), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n330), .A2(new_n563), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n569), .B1(new_n448), .B2(new_n563), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  AOI22_X1  g0371(.A1(new_n460), .A2(G270), .B1(new_n466), .B2(new_n464), .ZN(new_n572));
  OAI211_X1 g0372(.A(G264), .B(G1698), .C1(new_n308), .C2(new_n309), .ZN(new_n573));
  INV_X1    g0373(.A(new_n309), .ZN(new_n574));
  NAND2_X1  g0374(.A1(KEYINPUT3), .A2(G33), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n574), .A2(G303), .A3(new_n575), .ZN(new_n576));
  OAI211_X1 g0376(.A(G257), .B(new_n293), .C1(new_n308), .C2(new_n309), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n573), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(new_n297), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n572), .A2(new_n579), .A3(G190), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n571), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n516), .B1(new_n572), .B2(new_n579), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n562), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(new_n582), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n584), .A2(KEYINPUT81), .A3(new_n571), .A4(new_n580), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n572), .A2(new_n579), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n449), .A2(G116), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n588), .B(new_n569), .C1(new_n566), .C2(new_n567), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n587), .A2(new_n589), .A3(KEYINPUT21), .A4(G169), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n589), .A2(G179), .A3(new_n579), .A4(new_n572), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n342), .B1(new_n572), .B2(new_n579), .ZN(new_n593));
  AOI21_X1  g0393(.A(KEYINPUT21), .B1(new_n593), .B2(new_n589), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(new_n550), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n549), .B1(new_n541), .B2(new_n546), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n253), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  AOI22_X1  g0398(.A1(new_n556), .A2(new_n557), .B1(G107), .B2(new_n449), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n535), .A2(G190), .ZN(new_n600));
  AOI21_X1  g0400(.A(G200), .B1(new_n533), .B2(new_n467), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n598), .B(new_n599), .C1(new_n600), .C2(new_n601), .ZN(new_n602));
  AND4_X1   g0402(.A1(new_n561), .A2(new_n586), .A3(new_n595), .A4(new_n602), .ZN(new_n603));
  AND4_X1   g0403(.A1(new_n435), .A2(new_n490), .A3(new_n528), .A4(new_n603), .ZN(G372));
  INV_X1    g0404(.A(new_n344), .ZN(new_n605));
  AND2_X1   g0405(.A1(new_n418), .A2(new_n421), .ZN(new_n606));
  INV_X1    g0406(.A(new_n350), .ZN(new_n607));
  INV_X1    g0407(.A(new_n370), .ZN(new_n608));
  AOI22_X1  g0408(.A1(new_n607), .A2(new_n608), .B1(new_n340), .B2(new_n329), .ZN(new_n609));
  AND2_X1   g0409(.A1(new_n609), .A2(KEYINPUT84), .ZN(new_n610));
  AND2_X1   g0410(.A1(new_n427), .A2(new_n428), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n611), .B1(new_n609), .B2(KEYINPUT84), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n606), .B1(new_n610), .B2(new_n612), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n605), .B1(new_n613), .B2(new_n305), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n502), .A2(new_n503), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT79), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n502), .A2(KEYINPUT79), .A3(new_n503), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n523), .B1(new_n619), .B2(new_n520), .ZN(new_n620));
  INV_X1    g0420(.A(new_n524), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n527), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n489), .A2(new_n483), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n518), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n622), .A2(KEYINPUT26), .A3(new_n624), .A4(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n514), .A2(new_n368), .ZN(new_n627));
  AOI21_X1  g0427(.A(KEYINPUT83), .B1(new_n513), .B2(new_n297), .ZN(new_n628));
  INV_X1    g0428(.A(new_n628), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n513), .A2(KEYINPUT83), .A3(new_n297), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n509), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n627), .B1(new_n631), .B2(G169), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n632), .B1(new_n522), .B2(new_n524), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n515), .B1(new_n631), .B2(new_n516), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n506), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n483), .A2(KEYINPUT76), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(new_n452), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(new_n489), .ZN(new_n638));
  NOR3_X1   g0438(.A1(new_n633), .A2(new_n635), .A3(new_n638), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n626), .B1(new_n639), .B2(KEYINPUT26), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n486), .A2(new_n487), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(new_n516), .ZN(new_n642));
  AND2_X1   g0442(.A1(new_n642), .A2(new_n481), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n623), .B1(new_n643), .B2(new_n637), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n602), .B1(new_n506), .B2(new_n634), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n595), .A2(new_n561), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n633), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n640), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n435), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n614), .A2(new_n650), .ZN(G369));
  AND2_X1   g0451(.A1(new_n561), .A2(new_n602), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n207), .A2(new_n208), .A3(G13), .ZN(new_n654));
  OR2_X1    g0454(.A1(new_n654), .A2(KEYINPUT27), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(KEYINPUT27), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n655), .A2(G213), .A3(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(G343), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n660), .B1(new_n598), .B2(new_n599), .ZN(new_n661));
  OAI22_X1  g0461(.A1(new_n653), .A2(new_n661), .B1(new_n561), .B2(new_n660), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n571), .A2(new_n660), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n663), .B1(new_n592), .B2(new_n594), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n586), .A2(new_n595), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n664), .B1(new_n665), .B2(new_n663), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n662), .A2(new_n666), .A3(G330), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n561), .A2(new_n659), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n595), .A2(new_n659), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n668), .B1(new_n652), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n667), .A2(new_n670), .ZN(G399));
  INV_X1    g0471(.A(new_n211), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n672), .A2(G41), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n673), .A2(new_n207), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n500), .A2(G116), .ZN(new_n675));
  INV_X1    g0475(.A(new_n222), .ZN(new_n676));
  AOI22_X1  g0476(.A1(new_n674), .A2(new_n675), .B1(new_n676), .B2(new_n673), .ZN(new_n677));
  XOR2_X1   g0477(.A(new_n677), .B(KEYINPUT28), .Z(new_n678));
  INV_X1    g0478(.A(KEYINPUT87), .ZN(new_n679));
  AOI21_X1  g0479(.A(KEYINPUT26), .B1(new_n528), .B2(new_n624), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT26), .ZN(new_n681));
  NOR4_X1   g0481(.A1(new_n633), .A2(new_n638), .A3(new_n681), .A4(new_n635), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n648), .B1(new_n680), .B2(new_n682), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n683), .A2(KEYINPUT29), .A3(new_n660), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n659), .B1(new_n640), .B2(new_n648), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n684), .B1(KEYINPUT29), .B2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(G330), .ZN(new_n687));
  AND4_X1   g0487(.A1(new_n486), .A2(new_n487), .A3(new_n514), .A4(new_n533), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n572), .A2(new_n579), .A3(G179), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(KEYINPUT85), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT85), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n572), .A2(new_n579), .A3(new_n691), .A4(G179), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n688), .A2(KEYINPUT30), .A3(new_n690), .A4(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n509), .ZN(new_n694));
  AND3_X1   g0494(.A1(new_n513), .A2(KEYINPUT83), .A3(new_n297), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n694), .B1(new_n695), .B2(new_n628), .ZN(new_n696));
  AOI21_X1  g0496(.A(G179), .B1(new_n572), .B2(new_n579), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n641), .A2(new_n535), .A3(new_n696), .A4(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT86), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT30), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n690), .A2(new_n692), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n486), .A2(new_n487), .A3(new_n514), .A4(new_n533), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n701), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  AND2_X1   g0504(.A1(new_n697), .A2(new_n535), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n705), .A2(KEYINPUT86), .A3(new_n641), .A4(new_n696), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n693), .A2(new_n700), .A3(new_n704), .A4(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(new_n659), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT31), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n693), .A2(new_n704), .A3(new_n698), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n660), .A2(new_n709), .ZN(new_n711));
  AOI22_X1  g0511(.A1(new_n708), .A2(new_n709), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n528), .A2(new_n490), .A3(new_n603), .A4(new_n660), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n687), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n679), .B1(new_n686), .B2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n686), .A2(new_n679), .A3(new_n715), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n678), .B1(new_n719), .B2(G1), .ZN(G364));
  NAND2_X1  g0520(.A1(new_n666), .A2(G330), .ZN(new_n721));
  OR2_X1    g0521(.A1(new_n721), .A2(KEYINPUT88), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(KEYINPUT88), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(G13), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n725), .A2(G20), .ZN(new_n726));
  XNOR2_X1  g0526(.A(new_n726), .B(KEYINPUT89), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(G45), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n674), .A2(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n729), .B1(new_n666), .B2(G330), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n724), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(G13), .A2(G33), .ZN(new_n732));
  XNOR2_X1  g0532(.A(new_n732), .B(KEYINPUT90), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(new_n208), .ZN(new_n735));
  XOR2_X1   g0535(.A(new_n735), .B(KEYINPUT91), .Z(new_n736));
  OR2_X1    g0536(.A1(new_n666), .A2(new_n736), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n224), .B1(G20), .B2(new_n342), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n208), .A2(G190), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n516), .A2(G179), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n290), .B1(new_n742), .B2(new_n352), .ZN(new_n743));
  NOR2_X1   g0543(.A1(G179), .A2(G200), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n208), .B1(new_n744), .B2(G190), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(new_n437), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n740), .A2(new_n744), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(G159), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n746), .B1(new_n749), .B2(KEYINPUT32), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n750), .B1(KEYINPUT32), .B2(new_n749), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n208), .A2(new_n422), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(new_n741), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  AOI211_X1 g0554(.A(new_n743), .B(new_n751), .C1(G87), .C2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n368), .A2(G200), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n752), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n756), .A2(new_n740), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  AOI22_X1  g0560(.A1(G58), .A2(new_n758), .B1(new_n760), .B2(G77), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n208), .A2(new_n368), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(G200), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(new_n422), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n761), .B1(new_n244), .B2(new_n765), .ZN(new_n766));
  XOR2_X1   g0566(.A(new_n766), .B(KEYINPUT92), .Z(new_n767));
  INV_X1    g0567(.A(new_n763), .ZN(new_n768));
  AND3_X1   g0568(.A1(new_n768), .A2(KEYINPUT93), .A3(new_n422), .ZN(new_n769));
  AOI21_X1  g0569(.A(KEYINPUT93), .B1(new_n768), .B2(new_n422), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  OAI211_X1 g0571(.A(new_n755), .B(new_n767), .C1(new_n202), .C2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n771), .ZN(new_n773));
  XNOR2_X1  g0573(.A(KEYINPUT33), .B(G317), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(G294), .ZN(new_n776));
  INV_X1    g0576(.A(G311), .ZN(new_n777));
  OAI221_X1 g0577(.A(new_n389), .B1(new_n745), .B2(new_n776), .C1(new_n777), .C2(new_n759), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n778), .B1(G326), .B2(new_n764), .ZN(new_n779));
  XNOR2_X1  g0579(.A(new_n753), .B(KEYINPUT94), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(G303), .ZN(new_n781));
  INV_X1    g0581(.A(G322), .ZN(new_n782));
  INV_X1    g0582(.A(G329), .ZN(new_n783));
  OAI22_X1  g0583(.A1(new_n757), .A2(new_n782), .B1(new_n747), .B2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n742), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n784), .B1(G283), .B2(new_n785), .ZN(new_n786));
  NAND4_X1  g0586(.A1(new_n775), .A2(new_n779), .A3(new_n781), .A4(new_n786), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n739), .B1(new_n772), .B2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n736), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(new_n738), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n672), .A2(new_n389), .ZN(new_n791));
  AOI22_X1  g0591(.A1(new_n791), .A2(G355), .B1(new_n563), .B2(new_n672), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n672), .A2(new_n290), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n793), .B1(new_n223), .B2(G45), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n249), .A2(new_n281), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n792), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  AOI211_X1 g0596(.A(new_n729), .B(new_n788), .C1(new_n790), .C2(new_n796), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n731), .B1(new_n737), .B2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(G396));
  INV_X1    g0599(.A(new_n729), .ZN(new_n800));
  INV_X1    g0600(.A(new_n369), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n366), .B1(new_n367), .B2(G169), .ZN(new_n802));
  OAI21_X1  g0602(.A(KEYINPUT96), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(KEYINPUT96), .ZN(new_n804));
  NAND4_X1  g0604(.A1(new_n359), .A2(new_n804), .A3(new_n366), .A4(new_n369), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n366), .A2(new_n659), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n373), .A2(new_n807), .ZN(new_n808));
  OAI21_X1  g0608(.A(KEYINPUT97), .B1(new_n806), .B2(new_n808), .ZN(new_n809));
  AND2_X1   g0609(.A1(new_n373), .A2(new_n807), .ZN(new_n810));
  INV_X1    g0610(.A(KEYINPUT97), .ZN(new_n811));
  NAND4_X1  g0611(.A1(new_n810), .A2(new_n803), .A3(new_n811), .A4(new_n805), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n809), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n649), .A2(new_n660), .A3(new_n813), .ZN(new_n814));
  OAI211_X1 g0614(.A(new_n809), .B(new_n812), .C1(new_n370), .C2(new_n660), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n814), .B1(new_n685), .B2(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n800), .B1(new_n816), .B2(new_n715), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n817), .B1(new_n715), .B2(new_n816), .ZN(new_n818));
  OR2_X1    g0618(.A1(new_n738), .A2(new_n732), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n800), .B1(G77), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n773), .A2(G283), .ZN(new_n821));
  INV_X1    g0621(.A(G303), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n765), .A2(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n742), .A2(new_n404), .ZN(new_n824));
  NOR4_X1   g0624(.A1(new_n823), .A2(new_n290), .A3(new_n746), .A4(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n780), .A2(G107), .ZN(new_n826));
  OAI22_X1  g0626(.A1(new_n757), .A2(new_n776), .B1(new_n747), .B2(new_n777), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n827), .B1(G116), .B2(new_n760), .ZN(new_n828));
  NAND4_X1  g0628(.A1(new_n821), .A2(new_n825), .A3(new_n826), .A4(new_n828), .ZN(new_n829));
  AOI22_X1  g0629(.A1(G143), .A2(new_n758), .B1(new_n760), .B2(G159), .ZN(new_n830));
  INV_X1    g0630(.A(G137), .ZN(new_n831));
  OAI221_X1 g0631(.A(new_n830), .B1(new_n831), .B2(new_n765), .C1(new_n771), .C2(new_n261), .ZN(new_n832));
  XOR2_X1   g0632(.A(new_n832), .B(KEYINPUT95), .Z(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(KEYINPUT34), .ZN(new_n834));
  INV_X1    g0634(.A(G132), .ZN(new_n835));
  OAI221_X1 g0635(.A(new_n290), .B1(new_n747), .B2(new_n835), .C1(new_n202), .C2(new_n742), .ZN(new_n836));
  INV_X1    g0636(.A(new_n745), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n836), .B1(G58), .B2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n780), .ZN(new_n839));
  OAI211_X1 g0639(.A(new_n834), .B(new_n838), .C1(new_n244), .C2(new_n839), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n833), .A2(KEYINPUT34), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n829), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n820), .B1(new_n842), .B2(new_n738), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n843), .B1(new_n733), .B2(new_n815), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n818), .A2(new_n844), .ZN(G384));
  NOR2_X1   g0645(.A1(new_n727), .A2(new_n207), .ZN(new_n846));
  INV_X1    g0646(.A(new_n657), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n400), .A2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n429), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n417), .A2(new_n848), .A3(new_n425), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(KEYINPUT37), .ZN(new_n852));
  XNOR2_X1  g0652(.A(KEYINPUT101), .B(KEYINPUT37), .ZN(new_n853));
  NAND4_X1  g0653(.A1(new_n417), .A2(new_n848), .A3(new_n425), .A4(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n850), .A2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT38), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n850), .A2(new_n855), .A3(KEYINPUT38), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  AND3_X1   g0660(.A1(new_n329), .A2(KEYINPUT100), .A3(new_n340), .ZN(new_n861));
  AOI21_X1  g0661(.A(KEYINPUT100), .B1(new_n329), .B2(new_n340), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n340), .A2(new_n659), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n863), .B1(new_n347), .B2(new_n349), .ZN(new_n864));
  NOR3_X1   g0664(.A1(new_n861), .A2(new_n862), .A3(new_n864), .ZN(new_n865));
  OAI211_X1 g0665(.A(new_n340), .B(new_n659), .C1(new_n350), .C2(new_n329), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n815), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n708), .A2(new_n709), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n707), .A2(KEYINPUT31), .A3(new_n659), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n622), .A2(new_n490), .A3(new_n625), .ZN(new_n873));
  NAND4_X1  g0673(.A1(new_n652), .A2(new_n595), .A3(new_n586), .A4(new_n660), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NOR3_X1   g0675(.A1(new_n872), .A2(new_n875), .A3(KEYINPUT102), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT102), .ZN(new_n877));
  AND3_X1   g0677(.A1(new_n707), .A2(KEYINPUT31), .A3(new_n659), .ZN(new_n878));
  AOI21_X1  g0678(.A(KEYINPUT31), .B1(new_n707), .B2(new_n659), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n877), .B1(new_n880), .B2(new_n713), .ZN(new_n881));
  OAI211_X1 g0681(.A(new_n860), .B(new_n869), .C1(new_n876), .C2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT40), .ZN(new_n883));
  OAI21_X1  g0683(.A(KEYINPUT102), .B1(new_n872), .B2(new_n875), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n880), .A2(new_n877), .A3(new_n713), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n868), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n853), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n851), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(new_n854), .ZN(new_n889));
  AOI21_X1  g0689(.A(KEYINPUT38), .B1(new_n850), .B2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n883), .B1(new_n891), .B2(new_n859), .ZN(new_n892));
  AOI22_X1  g0692(.A1(new_n882), .A2(new_n883), .B1(new_n886), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n884), .A2(new_n885), .ZN(new_n894));
  AND3_X1   g0694(.A1(new_n893), .A2(new_n435), .A3(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n893), .B1(new_n435), .B2(new_n894), .ZN(new_n896));
  NOR3_X1   g0696(.A1(new_n895), .A2(new_n896), .A3(new_n687), .ZN(new_n897));
  XNOR2_X1  g0697(.A(new_n897), .B(KEYINPUT103), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT100), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n341), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n329), .A2(KEYINPUT100), .A3(new_n340), .ZN(new_n902));
  INV_X1    g0702(.A(new_n864), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n866), .ZN(new_n905));
  AND2_X1   g0705(.A1(new_n809), .A2(new_n812), .ZN(new_n906));
  AOI211_X1 g0706(.A(new_n659), .B(new_n906), .C1(new_n640), .C2(new_n648), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n806), .A2(new_n660), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n860), .B(new_n905), .C1(new_n907), .C2(new_n909), .ZN(new_n910));
  OR2_X1    g0710(.A1(new_n606), .A2(new_n847), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT39), .ZN(new_n912));
  INV_X1    g0712(.A(new_n859), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n912), .B1(new_n913), .B2(new_n890), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n858), .A2(KEYINPUT39), .A3(new_n859), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n659), .B1(new_n901), .B2(new_n902), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n914), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n910), .A2(new_n911), .A3(new_n917), .ZN(new_n918));
  OAI211_X1 g0718(.A(new_n684), .B(new_n435), .C1(KEYINPUT29), .C2(new_n685), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(new_n614), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n918), .B(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n846), .B1(new_n899), .B2(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n922), .B1(new_n899), .B2(new_n921), .ZN(new_n923));
  INV_X1    g0723(.A(new_n440), .ZN(new_n924));
  AOI211_X1 g0724(.A(new_n563), .B(new_n226), .C1(new_n924), .C2(KEYINPUT35), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n925), .B1(KEYINPUT35), .B2(new_n924), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n926), .B(KEYINPUT36), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n676), .A2(G77), .A3(new_n380), .ZN(new_n928));
  AND2_X1   g0728(.A1(new_n928), .A2(KEYINPUT98), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n928), .A2(KEYINPUT98), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n245), .B(KEYINPUT99), .ZN(new_n931));
  NOR3_X1   g0731(.A1(new_n929), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n725), .A2(G1), .ZN(new_n933));
  OAI211_X1 g0733(.A(new_n923), .B(new_n927), .C1(new_n932), .C2(new_n933), .ZN(G367));
  NAND2_X1  g0734(.A1(new_n728), .A2(G1), .ZN(new_n935));
  INV_X1    g0735(.A(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(new_n718), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n937), .A2(new_n716), .ZN(new_n938));
  INV_X1    g0738(.A(new_n667), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n455), .A2(new_n660), .ZN(new_n940));
  OAI22_X1  g0740(.A1(new_n644), .A2(new_n940), .B1(new_n638), .B2(new_n660), .ZN(new_n941));
  OR3_X1    g0741(.A1(new_n941), .A2(new_n670), .A3(KEYINPUT104), .ZN(new_n942));
  OAI21_X1  g0742(.A(KEYINPUT104), .B1(new_n941), .B2(new_n670), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n942), .A2(KEYINPUT44), .A3(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT45), .ZN(new_n945));
  INV_X1    g0745(.A(new_n941), .ZN(new_n946));
  INV_X1    g0746(.A(new_n670), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n945), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n941), .A2(new_n670), .A3(KEYINPUT45), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n944), .A2(new_n950), .ZN(new_n951));
  AOI21_X1  g0751(.A(KEYINPUT44), .B1(new_n942), .B2(new_n943), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n939), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(new_n952), .ZN(new_n954));
  NAND4_X1  g0754(.A1(new_n954), .A2(new_n667), .A3(new_n950), .A4(new_n944), .ZN(new_n955));
  AND2_X1   g0755(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n652), .A2(new_n669), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(new_n662), .B2(new_n669), .ZN(new_n958));
  OR2_X1    g0758(.A1(new_n958), .A2(new_n721), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n958), .A2(new_n722), .A3(new_n723), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  OAI211_X1 g0762(.A(new_n956), .B(new_n962), .C1(new_n937), .C2(new_n716), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(KEYINPUT105), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT105), .ZN(new_n965));
  NAND4_X1  g0765(.A1(new_n719), .A2(new_n965), .A3(new_n962), .A4(new_n956), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n938), .B1(new_n964), .B2(new_n966), .ZN(new_n967));
  XOR2_X1   g0767(.A(new_n673), .B(KEYINPUT41), .Z(new_n968));
  OAI21_X1  g0768(.A(new_n936), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n946), .A2(new_n957), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n970), .B(KEYINPUT42), .Z(new_n971));
  OAI21_X1  g0771(.A(new_n623), .B1(new_n946), .B2(new_n561), .ZN(new_n972));
  AND2_X1   g0772(.A1(new_n972), .A2(new_n660), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT43), .ZN(new_n974));
  AOI211_X1 g0774(.A(new_n635), .B(new_n633), .C1(new_n506), .C2(new_n659), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n633), .A2(new_n506), .A3(new_n659), .ZN(new_n976));
  INV_X1    g0776(.A(new_n976), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  OAI22_X1  g0778(.A1(new_n971), .A2(new_n973), .B1(new_n974), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n974), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n979), .B(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n939), .A2(new_n941), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n981), .B(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n969), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n978), .A2(new_n789), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n790), .B1(new_n211), .B2(new_n362), .ZN(new_n986));
  AND2_X1   g0786(.A1(new_n233), .A2(new_n793), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n800), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n785), .A2(G77), .ZN(new_n989));
  INV_X1    g0789(.A(G143), .ZN(new_n990));
  OAI211_X1 g0790(.A(new_n290), .B(new_n989), .C1(new_n765), .C2(new_n990), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n745), .A2(new_n202), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  OAI22_X1  g0793(.A1(new_n201), .A2(new_n753), .B1(new_n757), .B2(new_n261), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n759), .A2(new_n244), .B1(new_n747), .B2(new_n831), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(G159), .ZN(new_n997));
  OAI211_X1 g0797(.A(new_n993), .B(new_n996), .C1(new_n997), .C2(new_n771), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n742), .A2(new_n437), .ZN(new_n999));
  AOI211_X1 g0799(.A(new_n290), .B(new_n999), .C1(G317), .C2(new_n748), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n773), .A2(G294), .B1(new_n1000), .B2(KEYINPUT106), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1001), .B1(KEYINPUT106), .B2(new_n1000), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n780), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT46), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1004), .B1(new_n753), .B2(new_n563), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(G303), .A2(new_n758), .B1(new_n760), .B2(G283), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(new_n764), .A2(G311), .B1(G107), .B2(new_n837), .ZN(new_n1007));
  NAND4_X1  g0807(.A1(new_n1003), .A2(new_n1005), .A3(new_n1006), .A4(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n998), .B1(new_n1002), .B2(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(KEYINPUT47), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n988), .B1(new_n1010), .B2(new_n738), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n985), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n984), .A2(new_n1012), .ZN(G387));
  NAND2_X1  g0813(.A1(new_n938), .A2(new_n961), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n719), .A2(new_n962), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1014), .A2(new_n1015), .A3(new_n673), .ZN(new_n1016));
  OR2_X1    g0816(.A1(new_n662), .A2(new_n736), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n790), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n791), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n1019), .A2(new_n675), .B1(G107), .B2(new_n211), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n793), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1021), .B1(new_n238), .B2(G45), .ZN(new_n1022));
  OAI211_X1 g0822(.A(new_n675), .B(new_n281), .C1(new_n202), .C2(new_n292), .ZN(new_n1023));
  INV_X1    g0823(.A(KEYINPUT107), .ZN(new_n1024));
  OR2_X1    g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n360), .A2(G50), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT50), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1025), .A2(new_n1026), .A3(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1020), .B1(new_n1022), .B2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n800), .B1(new_n1018), .B2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n754), .A2(G77), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(new_n261), .B2(new_n747), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT108), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n837), .A2(new_n519), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1035), .B1(new_n765), .B2(new_n997), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n757), .A2(new_n244), .B1(new_n759), .B2(new_n202), .ZN(new_n1037));
  NOR4_X1   g0837(.A1(new_n1036), .A2(new_n1037), .A3(new_n389), .A4(new_n999), .ZN(new_n1038));
  OAI211_X1 g0838(.A(new_n1034), .B(new_n1038), .C1(new_n257), .C2(new_n771), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n290), .B1(new_n748), .B2(G326), .ZN(new_n1040));
  INV_X1    g0840(.A(G283), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n753), .A2(new_n776), .B1(new_n745), .B2(new_n1041), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(G317), .A2(new_n758), .B1(new_n760), .B2(G303), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n1043), .B1(new_n782), .B2(new_n765), .C1(new_n771), .C2(new_n777), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT48), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1042), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1046), .B1(new_n1045), .B2(new_n1044), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT49), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n1040), .B1(new_n563), .B2(new_n742), .C1(new_n1047), .C2(new_n1048), .ZN(new_n1049));
  AND2_X1   g0849(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1039), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1031), .B1(new_n1051), .B2(new_n738), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n962), .A2(new_n935), .B1(new_n1017), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1016), .A2(new_n1053), .ZN(G393));
  OAI22_X1  g0854(.A1(new_n1021), .A2(new_n242), .B1(new_n437), .B2(new_n211), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n800), .B1(new_n1018), .B2(new_n1055), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n764), .A2(G317), .B1(new_n758), .B2(G311), .ZN(new_n1057));
  XOR2_X1   g0857(.A(new_n1057), .B(KEYINPUT52), .Z(new_n1058));
  OAI22_X1  g0858(.A1(new_n759), .A2(new_n776), .B1(new_n747), .B2(new_n782), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n389), .B1(new_n745), .B2(new_n563), .C1(new_n352), .C2(new_n742), .ZN(new_n1060));
  AOI211_X1 g0860(.A(new_n1059), .B(new_n1060), .C1(G283), .C2(new_n754), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n1058), .B(new_n1061), .C1(new_n822), .C2(new_n771), .ZN(new_n1062));
  XOR2_X1   g0862(.A(new_n1062), .B(KEYINPUT110), .Z(new_n1063));
  OAI22_X1  g0863(.A1(new_n771), .A2(new_n244), .B1(new_n360), .B2(new_n759), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n1064), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n1065), .A2(KEYINPUT109), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n764), .A2(G150), .B1(new_n758), .B2(G159), .ZN(new_n1067));
  XOR2_X1   g0867(.A(new_n1067), .B(KEYINPUT51), .Z(new_n1068));
  OAI22_X1  g0868(.A1(new_n753), .A2(new_n202), .B1(new_n747), .B2(new_n990), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n745), .A2(new_n292), .ZN(new_n1070));
  NOR4_X1   g0870(.A1(new_n1069), .A2(new_n824), .A3(new_n1070), .A4(new_n389), .ZN(new_n1071));
  INV_X1    g0871(.A(KEYINPUT109), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n1068), .B(new_n1071), .C1(new_n1064), .C2(new_n1072), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1063), .B1(new_n1066), .B2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1056), .B1(new_n1074), .B2(new_n738), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1075), .B1(new_n736), .B2(new_n941), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n956), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1076), .B1(new_n1077), .B2(new_n936), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n964), .A2(new_n966), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n673), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1080), .B1(new_n1015), .B2(new_n1077), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1078), .B1(new_n1079), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1082), .ZN(G390));
  NAND2_X1  g0883(.A1(new_n914), .A2(new_n915), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1084), .A2(new_n734), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n800), .B1(new_n256), .B2(new_n819), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n389), .B1(new_n742), .B2(new_n202), .ZN(new_n1087));
  AOI211_X1 g0887(.A(new_n1070), .B(new_n1087), .C1(G283), .C2(new_n764), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n757), .A2(new_n563), .B1(new_n759), .B2(new_n437), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1089), .B1(G294), .B2(new_n748), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n1088), .B(new_n1090), .C1(new_n404), .C2(new_n839), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n771), .A2(new_n352), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n290), .B1(new_n742), .B2(new_n244), .ZN(new_n1093));
  XOR2_X1   g0893(.A(new_n1093), .B(KEYINPUT111), .Z(new_n1094));
  OAI21_X1  g0894(.A(new_n1094), .B1(new_n831), .B2(new_n771), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n753), .A2(new_n261), .ZN(new_n1096));
  XOR2_X1   g0896(.A(KEYINPUT112), .B(KEYINPUT53), .Z(new_n1097));
  XNOR2_X1  g0897(.A(new_n1096), .B(new_n1097), .ZN(new_n1098));
  XNOR2_X1  g0898(.A(KEYINPUT54), .B(G143), .ZN(new_n1099));
  INV_X1    g0899(.A(G125), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n759), .A2(new_n1099), .B1(new_n747), .B2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(G132), .B2(new_n758), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n764), .A2(G128), .B1(G159), .B2(new_n837), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1098), .A2(new_n1102), .A3(new_n1103), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n1091), .A2(new_n1092), .B1(new_n1095), .B2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1086), .B1(new_n1105), .B2(new_n738), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1085), .A2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n916), .B1(new_n891), .B2(new_n859), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n683), .A2(new_n660), .A3(new_n813), .ZN(new_n1109));
  AND2_X1   g0909(.A1(new_n1109), .A2(new_n908), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n905), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1108), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1111), .B1(new_n814), .B2(new_n908), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1084), .B1(new_n1113), .B2(new_n916), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1115));
  AOI211_X1 g0915(.A(new_n687), .B(new_n868), .C1(new_n884), .C2(new_n885), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n710), .A2(new_n711), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n713), .A2(new_n870), .A3(new_n1118), .ZN(new_n1119));
  NAND4_X1  g0919(.A1(new_n1119), .A2(G330), .A3(new_n815), .A4(new_n905), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1112), .A2(new_n1114), .A3(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1117), .A2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1107), .B1(new_n1122), .B2(new_n936), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n894), .A2(G330), .A3(new_n435), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n919), .A2(new_n1124), .A3(new_n614), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n905), .B1(new_n714), .B2(new_n815), .ZN(new_n1126));
  OAI22_X1  g0926(.A1(new_n1116), .A2(new_n1126), .B1(new_n907), .B2(new_n909), .ZN(new_n1127));
  AND3_X1   g0927(.A1(new_n1109), .A2(new_n1120), .A3(new_n908), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n815), .ZN(new_n1129));
  AOI211_X1 g0929(.A(new_n687), .B(new_n1129), .C1(new_n884), .C2(new_n885), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1128), .B1(new_n1130), .B2(new_n905), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1125), .B1(new_n1127), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1080), .B1(new_n1122), .B2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1117), .A2(new_n1121), .A3(new_n1132), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1123), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(G378));
  AND3_X1   g0937(.A1(new_n910), .A2(new_n911), .A3(new_n917), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n882), .A2(new_n883), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n886), .A2(new_n892), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1139), .A2(new_n1140), .A3(G330), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1138), .A2(new_n1141), .ZN(new_n1142));
  XNOR2_X1  g0942(.A(KEYINPUT117), .B(KEYINPUT56), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(new_n1143), .B(KEYINPUT118), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(new_n431), .B(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n270), .A2(new_n847), .ZN(new_n1146));
  XOR2_X1   g0946(.A(new_n1146), .B(KEYINPUT55), .Z(new_n1147));
  XNOR2_X1  g0947(.A(new_n1147), .B(KEYINPUT116), .ZN(new_n1148));
  XNOR2_X1  g0948(.A(new_n1145), .B(new_n1148), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n1149), .A2(KEYINPUT120), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n918), .A2(G330), .A3(new_n893), .ZN(new_n1151));
  AND3_X1   g0951(.A1(new_n1142), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1150), .B1(new_n1142), .B2(new_n1151), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n935), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n800), .B1(G50), .B2(new_n819), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n290), .A2(G41), .ZN(new_n1156));
  AOI211_X1 g0956(.A(G50), .B(new_n1156), .C1(new_n403), .C2(new_n280), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(new_n1157), .B(KEYINPUT113), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n773), .A2(G97), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n757), .A2(new_n352), .B1(new_n759), .B2(new_n362), .ZN(new_n1160));
  OAI22_X1  g0960(.A1(new_n742), .A2(new_n201), .B1(new_n747), .B2(new_n1041), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n764), .A2(G116), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1032), .A2(new_n1156), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n1164), .A2(new_n992), .ZN(new_n1165));
  NAND4_X1  g0965(.A1(new_n1159), .A2(new_n1162), .A3(new_n1163), .A4(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1158), .B1(new_n1167), .B2(KEYINPUT58), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n745), .A2(new_n261), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n753), .A2(new_n1099), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT114), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  AOI211_X1 g0972(.A(new_n1169), .B(new_n1172), .C1(G125), .C2(new_n764), .ZN(new_n1173));
  INV_X1    g0973(.A(G128), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n757), .A2(new_n1174), .B1(new_n759), .B2(new_n831), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1175), .B1(new_n1171), .B2(new_n1170), .ZN(new_n1176));
  OAI211_X1 g0976(.A(new_n1173), .B(new_n1176), .C1(new_n835), .C2(new_n771), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1177), .A2(KEYINPUT59), .ZN(new_n1178));
  XOR2_X1   g0978(.A(KEYINPUT115), .B(G124), .Z(new_n1179));
  AOI211_X1 g0979(.A(G33), .B(G41), .C1(new_n748), .C2(new_n1179), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1178), .B(new_n1180), .C1(new_n997), .C2(new_n742), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n1177), .A2(KEYINPUT59), .ZN(new_n1182));
  OAI221_X1 g0982(.A(new_n1168), .B1(KEYINPUT58), .B2(new_n1167), .C1(new_n1181), .C2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1155), .B1(new_n1183), .B2(new_n738), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1184), .B1(new_n1149), .B2(new_n733), .ZN(new_n1185));
  XNOR2_X1  g0985(.A(new_n1185), .B(KEYINPUT119), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1154), .A2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1142), .A2(new_n1151), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1150), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1142), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1125), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n1192), .A2(new_n1193), .B1(new_n1135), .B2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1195), .A2(KEYINPUT57), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1196), .A2(new_n673), .ZN(new_n1197));
  INV_X1    g0997(.A(KEYINPUT57), .ZN(new_n1198));
  AND2_X1   g0998(.A1(new_n1135), .A2(new_n1194), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1198), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1189), .B1(new_n1197), .B2(new_n1202), .ZN(G375));
  INV_X1    g1003(.A(new_n968), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1127), .A2(new_n1131), .A3(new_n1125), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1133), .A2(new_n1204), .A3(new_n1205), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(new_n1206), .B(KEYINPUT121), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n764), .A2(G294), .ZN(new_n1208));
  NAND4_X1  g1008(.A1(new_n1208), .A2(new_n389), .A3(new_n989), .A4(new_n1035), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(G283), .A2(new_n758), .B1(new_n760), .B2(G107), .ZN(new_n1210));
  OAI221_X1 g1010(.A(new_n1210), .B1(new_n822), .B2(new_n747), .C1(new_n839), .C2(new_n437), .ZN(new_n1211));
  AOI211_X1 g1011(.A(new_n1209), .B(new_n1211), .C1(G116), .C2(new_n773), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(G137), .A2(new_n758), .B1(new_n760), .B2(G150), .ZN(new_n1213));
  OAI221_X1 g1013(.A(new_n1213), .B1(new_n1174), .B2(new_n747), .C1(new_n839), .C2(new_n997), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n771), .A2(new_n1099), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n389), .B1(new_n785), .B2(G58), .ZN(new_n1216));
  OAI221_X1 g1016(.A(new_n1216), .B1(new_n244), .B2(new_n745), .C1(new_n765), .C2(new_n835), .ZN(new_n1217));
  NOR3_X1   g1017(.A1(new_n1214), .A2(new_n1215), .A3(new_n1217), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n738), .B1(new_n1212), .B2(new_n1218), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1219), .B(new_n800), .C1(G68), .C2(new_n819), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1220), .B1(new_n1111), .B2(new_n732), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n909), .B1(new_n685), .B2(new_n813), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n687), .B1(new_n884), .B2(new_n885), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1126), .B1(new_n1223), .B2(new_n869), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n905), .B1(new_n1223), .B2(new_n815), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1109), .A2(new_n1120), .A3(new_n908), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n1222), .A2(new_n1224), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1221), .B1(new_n1227), .B2(new_n935), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1207), .A2(new_n1228), .ZN(G381));
  NOR3_X1   g1029(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1230));
  XOR2_X1   g1030(.A(new_n1230), .B(KEYINPUT122), .Z(new_n1231));
  NAND4_X1  g1031(.A1(new_n1136), .A2(new_n1207), .A3(new_n1082), .A4(new_n1228), .ZN(new_n1232));
  OR4_X1    g1032(.A1(G387), .A2(new_n1231), .A3(new_n1232), .A4(G375), .ZN(G407));
  NAND2_X1  g1033(.A1(new_n658), .A2(G213), .ZN(new_n1234));
  XOR2_X1   g1034(.A(new_n1234), .B(KEYINPUT123), .Z(new_n1235));
  NAND2_X1  g1035(.A1(new_n1136), .A2(new_n1235), .ZN(new_n1236));
  OAI211_X1 g1036(.A(G407), .B(G213), .C1(G375), .C2(new_n1236), .ZN(G409));
  NAND2_X1  g1037(.A1(G387), .A2(new_n1082), .ZN(new_n1238));
  XNOR2_X1  g1038(.A(G393), .B(new_n798), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n984), .A2(new_n1012), .A3(G390), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1238), .A2(new_n1239), .A3(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1239), .ZN(new_n1242));
  AOI21_X1  g1042(.A(G390), .B1(new_n984), .B2(new_n1012), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1012), .ZN(new_n1244));
  AOI211_X1 g1044(.A(new_n1244), .B(new_n1082), .C1(new_n969), .C2(new_n983), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1242), .B1(new_n1243), .B2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1241), .A2(new_n1246), .ZN(new_n1247));
  AND2_X1   g1047(.A1(new_n1235), .A2(G2897), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1127), .A2(new_n1131), .A3(KEYINPUT60), .A4(new_n1125), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT125), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  OAI211_X1 g1051(.A(G330), .B(new_n815), .C1(new_n876), .C2(new_n881), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1226), .B1(new_n1111), .B2(new_n1252), .ZN(new_n1253));
  OAI211_X1 g1053(.A(G330), .B(new_n869), .C1(new_n876), .C2(new_n881), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1126), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1222), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1253), .A2(new_n1256), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1257), .A2(KEYINPUT125), .A3(KEYINPUT60), .A4(new_n1125), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1080), .B1(new_n1227), .B2(new_n1194), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT60), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1205), .A2(new_n1260), .ZN(new_n1261));
  NAND4_X1  g1061(.A1(new_n1251), .A2(new_n1258), .A3(new_n1259), .A4(new_n1261), .ZN(new_n1262));
  AND3_X1   g1062(.A1(new_n1262), .A2(G384), .A3(new_n1228), .ZN(new_n1263));
  AOI21_X1  g1063(.A(G384), .B1(new_n1262), .B2(new_n1228), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1248), .B1(new_n1263), .B2(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1262), .A2(new_n1228), .ZN(new_n1266));
  INV_X1    g1066(.A(G384), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1262), .A2(G384), .A3(new_n1228), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n658), .A2(G213), .A3(G2897), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1268), .A2(new_n1269), .A3(new_n1270), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1265), .A2(new_n1271), .A3(KEYINPUT126), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT126), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1273), .A2(new_n1274), .A3(new_n1248), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1272), .A2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(KEYINPUT127), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1235), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1080), .B1(new_n1195), .B2(KEYINPUT57), .ZN(new_n1279));
  AOI211_X1 g1079(.A(new_n1188), .B(new_n1136), .C1(new_n1279), .C2(new_n1201), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT124), .ZN(new_n1281));
  AOI22_X1  g1081(.A1(new_n1188), .A2(new_n1281), .B1(new_n1195), .B2(new_n1204), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1154), .A2(KEYINPUT124), .A3(new_n1187), .ZN(new_n1283));
  AOI21_X1  g1083(.A(G378), .B1(new_n1282), .B2(new_n1283), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1278), .B1(new_n1280), .B2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT127), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1272), .A2(new_n1286), .A3(new_n1275), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1277), .A2(new_n1285), .A3(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT61), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1273), .ZN(new_n1291));
  OAI211_X1 g1091(.A(new_n1234), .B(new_n1291), .C1(new_n1280), .C2(new_n1284), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT62), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1188), .A2(new_n1281), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1195), .A2(new_n1204), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1294), .A2(new_n1283), .A3(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1296), .A2(new_n1136), .ZN(new_n1297));
  OAI211_X1 g1097(.A(G378), .B(new_n1189), .C1(new_n1197), .C2(new_n1202), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1235), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1299));
  NOR2_X1   g1099(.A1(new_n1273), .A2(new_n1293), .ZN(new_n1300));
  AOI22_X1  g1100(.A1(new_n1292), .A2(new_n1293), .B1(new_n1299), .B2(new_n1300), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1247), .B1(new_n1290), .B2(new_n1301), .ZN(new_n1302));
  NOR2_X1   g1102(.A1(new_n1247), .A2(KEYINPUT61), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT63), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1292), .A2(new_n1304), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1234), .B1(new_n1280), .B2(new_n1284), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1277), .A2(new_n1306), .A3(new_n1287), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1299), .A2(KEYINPUT63), .A3(new_n1291), .ZN(new_n1308));
  NAND4_X1  g1108(.A1(new_n1303), .A2(new_n1305), .A3(new_n1307), .A4(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1302), .A2(new_n1309), .ZN(G405));
  XNOR2_X1  g1110(.A(G375), .B(G378), .ZN(new_n1311));
  OR2_X1    g1111(.A1(new_n1311), .A2(new_n1273), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1311), .A2(new_n1273), .ZN(new_n1313));
  NAND4_X1  g1113(.A1(new_n1312), .A2(new_n1241), .A3(new_n1246), .A4(new_n1313), .ZN(new_n1314));
  AND2_X1   g1114(.A1(new_n1311), .A2(new_n1273), .ZN(new_n1315));
  NOR2_X1   g1115(.A1(new_n1311), .A2(new_n1273), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1247), .B1(new_n1315), .B2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1314), .A2(new_n1317), .ZN(G402));
endmodule


