//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 1 0 1 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 1 0 0 0 0 1 1 0 1 0 1 0 1 1 1 1 0 1 1 1 0 1 0 0 0 1 0 0 1 1 1 1 1 1 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n585, new_n586, new_n587, new_n588,
    new_n590, new_n591, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n663, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n690, new_n691,
    new_n692, new_n693, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n753, new_n754, new_n755, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n812, new_n813, new_n815, new_n816, new_n817, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n831, new_n832, new_n833, new_n834, new_n836,
    new_n837, new_n838, new_n840, new_n841, new_n842, new_n843, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n876,
    new_n877, new_n878, new_n879, new_n880;
  INV_X1    g000(.A(G8gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G15gat), .B(G22gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT16), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n203), .B1(new_n204), .B2(G1gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT86), .ZN(new_n206));
  AOI21_X1  g005(.A(new_n202), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n205), .B1(G1gat), .B2(new_n203), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  OAI221_X1 g008(.A(new_n205), .B1(new_n206), .B2(new_n202), .C1(G1gat), .C2(new_n203), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT88), .ZN(new_n212));
  XNOR2_X1  g011(.A(new_n211), .B(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(G71gat), .A2(G78gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT9), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  OR2_X1    g015(.A1(G57gat), .A2(G64gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(G57gat), .A2(G64gat), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT92), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n217), .A2(new_n220), .A3(new_n218), .ZN(new_n221));
  XNOR2_X1  g020(.A(G71gat), .B(G78gat), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n219), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  AND2_X1   g022(.A1(G57gat), .A2(G64gat), .ZN(new_n224));
  NOR2_X1   g023(.A1(G57gat), .A2(G64gat), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  AND2_X1   g025(.A1(G71gat), .A2(G78gat), .ZN(new_n227));
  NOR2_X1   g026(.A1(G71gat), .A2(G78gat), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OAI211_X1 g028(.A(new_n216), .B(new_n226), .C1(new_n229), .C2(new_n220), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n223), .A2(new_n230), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n213), .B1(KEYINPUT21), .B2(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n232), .B(KEYINPUT94), .ZN(new_n233));
  XOR2_X1   g032(.A(KEYINPUT93), .B(KEYINPUT19), .Z(new_n234));
  XNOR2_X1  g033(.A(new_n233), .B(new_n234), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n231), .A2(KEYINPUT21), .ZN(new_n236));
  NAND2_X1  g035(.A1(G231gat), .A2(G233gat), .ZN(new_n237));
  XNOR2_X1  g036(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(G127gat), .B(G155gat), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n239), .B(KEYINPUT20), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n238), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(G183gat), .B(G211gat), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n241), .B(new_n242), .ZN(new_n243));
  OR2_X1    g042(.A1(new_n235), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n235), .A2(new_n243), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(G99gat), .A2(G106gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(KEYINPUT8), .ZN(new_n248));
  NAND2_X1  g047(.A1(G85gat), .A2(G92gat), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT7), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(G85gat), .ZN(new_n252));
  INV_X1    g051(.A(G92gat), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g053(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n255));
  NAND4_X1  g054(.A1(new_n248), .A2(new_n251), .A3(new_n254), .A4(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(G99gat), .B(G106gat), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  AND3_X1   g058(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n260));
  AOI21_X1  g059(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  AOI22_X1  g061(.A1(KEYINPUT8), .A2(new_n247), .B1(new_n252), .B2(new_n253), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n262), .A2(new_n257), .A3(new_n263), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n259), .A2(KEYINPUT95), .A3(new_n264), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n257), .B1(new_n262), .B2(new_n263), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT95), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  AND2_X1   g067(.A1(new_n265), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  XOR2_X1   g069(.A(G43gat), .B(G50gat), .Z(new_n271));
  INV_X1    g070(.A(KEYINPUT15), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(G43gat), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n275), .A2(KEYINPUT85), .A3(G50gat), .ZN(new_n276));
  XNOR2_X1  g075(.A(KEYINPUT84), .B(KEYINPUT15), .ZN(new_n277));
  OAI211_X1 g076(.A(new_n276), .B(new_n277), .C1(new_n271), .C2(KEYINPUT85), .ZN(new_n278));
  NAND2_X1  g077(.A1(G29gat), .A2(G36gat), .ZN(new_n279));
  OR3_X1    g078(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n280));
  OAI21_X1  g079(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND4_X1  g081(.A1(new_n274), .A2(new_n278), .A3(new_n279), .A4(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT83), .ZN(new_n284));
  OR2_X1    g083(.A1(new_n281), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n281), .A2(new_n284), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n285), .A2(new_n280), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(new_n279), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(new_n273), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n283), .A2(new_n289), .ZN(new_n290));
  AND2_X1   g089(.A1(G232gat), .A2(G233gat), .ZN(new_n291));
  AOI22_X1  g090(.A1(new_n270), .A2(new_n290), .B1(KEYINPUT41), .B2(new_n291), .ZN(new_n292));
  AOI21_X1  g091(.A(KEYINPUT17), .B1(new_n283), .B2(new_n289), .ZN(new_n293));
  OR2_X1    g092(.A1(new_n293), .A2(new_n270), .ZN(new_n294));
  AND3_X1   g093(.A1(new_n289), .A2(new_n283), .A3(KEYINPUT17), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n292), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  XNOR2_X1  g095(.A(G190gat), .B(G218gat), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n296), .B(new_n297), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n291), .A2(KEYINPUT41), .ZN(new_n299));
  XNOR2_X1  g098(.A(G134gat), .B(G162gat), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n299), .B(new_n300), .ZN(new_n301));
  XNOR2_X1  g100(.A(new_n298), .B(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n246), .A2(new_n303), .ZN(new_n304));
  XNOR2_X1  g103(.A(G120gat), .B(G148gat), .ZN(new_n305));
  XNOR2_X1  g104(.A(G176gat), .B(G204gat), .ZN(new_n306));
  XOR2_X1   g105(.A(new_n305), .B(new_n306), .Z(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT10), .ZN(new_n309));
  AND2_X1   g108(.A1(new_n223), .A2(new_n230), .ZN(new_n310));
  NOR3_X1   g109(.A1(new_n269), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT97), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT96), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n259), .A2(new_n264), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n314), .B1(new_n310), .B2(new_n315), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n256), .A2(new_n258), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n317), .A2(new_n266), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n318), .A2(KEYINPUT96), .A3(new_n231), .ZN(new_n319));
  AOI22_X1  g118(.A1(new_n316), .A2(new_n319), .B1(new_n269), .B2(new_n310), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n313), .B1(new_n320), .B2(new_n309), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n316), .A2(new_n319), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n310), .A2(new_n265), .A3(new_n268), .ZN(new_n323));
  AND4_X1   g122(.A1(new_n313), .A2(new_n322), .A3(new_n309), .A4(new_n323), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n312), .B1(new_n321), .B2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT99), .ZN(new_n326));
  NAND2_X1  g125(.A1(G230gat), .A2(G233gat), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n325), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  NOR3_X1   g127(.A1(new_n310), .A2(new_n315), .A3(new_n314), .ZN(new_n329));
  AOI21_X1  g128(.A(KEYINPUT96), .B1(new_n318), .B2(new_n231), .ZN(new_n330));
  OAI211_X1 g129(.A(new_n309), .B(new_n323), .C1(new_n329), .C2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(KEYINPUT97), .ZN(new_n332));
  NAND4_X1  g131(.A1(new_n322), .A2(new_n313), .A3(new_n309), .A4(new_n323), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n311), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(new_n327), .ZN(new_n335));
  OAI21_X1  g134(.A(KEYINPUT99), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  AND2_X1   g135(.A1(new_n328), .A2(new_n336), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n320), .A2(new_n327), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n308), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT98), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n325), .A2(new_n340), .A3(new_n327), .ZN(new_n341));
  OAI21_X1  g140(.A(KEYINPUT98), .B1(new_n334), .B2(new_n335), .ZN(new_n342));
  AND2_X1   g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n338), .A2(new_n308), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n339), .A2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n304), .A2(new_n347), .ZN(new_n348));
  XNOR2_X1  g147(.A(G15gat), .B(G43gat), .ZN(new_n349));
  XNOR2_X1  g148(.A(G71gat), .B(G99gat), .ZN(new_n350));
  XNOR2_X1  g149(.A(new_n349), .B(new_n350), .ZN(new_n351));
  NOR2_X1   g150(.A1(G169gat), .A2(G176gat), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT26), .ZN(new_n354));
  NAND2_X1  g153(.A1(G169gat), .A2(G176gat), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(G183gat), .A2(G190gat), .ZN(new_n357));
  OAI211_X1 g156(.A(new_n356), .B(new_n357), .C1(new_n354), .C2(new_n353), .ZN(new_n358));
  OR2_X1    g157(.A1(new_n358), .A2(KEYINPUT66), .ZN(new_n359));
  XNOR2_X1  g158(.A(KEYINPUT27), .B(G183gat), .ZN(new_n360));
  INV_X1    g159(.A(G190gat), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT28), .ZN(new_n363));
  XNOR2_X1  g162(.A(new_n362), .B(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n358), .A2(KEYINPUT66), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n359), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT23), .ZN(new_n367));
  XNOR2_X1  g166(.A(new_n352), .B(new_n367), .ZN(new_n368));
  OR2_X1    g167(.A1(G183gat), .A2(G190gat), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n369), .A2(KEYINPUT24), .A3(new_n357), .ZN(new_n370));
  OR2_X1    g169(.A1(new_n357), .A2(KEYINPUT24), .ZN(new_n371));
  NOR2_X1   g170(.A1(KEYINPUT65), .A2(KEYINPUT25), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n372), .B1(G169gat), .B2(G176gat), .ZN(new_n373));
  NAND4_X1  g172(.A1(new_n368), .A2(new_n370), .A3(new_n371), .A4(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(KEYINPUT65), .A2(KEYINPUT25), .ZN(new_n375));
  XNOR2_X1  g174(.A(new_n374), .B(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n366), .A2(new_n376), .ZN(new_n377));
  XOR2_X1   g176(.A(G127gat), .B(G134gat), .Z(new_n378));
  INV_X1    g177(.A(KEYINPUT67), .ZN(new_n379));
  XOR2_X1   g178(.A(G113gat), .B(G120gat), .Z(new_n380));
  AOI21_X1  g179(.A(new_n378), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT1), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  XNOR2_X1  g182(.A(new_n381), .B(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  XNOR2_X1  g184(.A(new_n377), .B(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(G227gat), .A2(G233gat), .ZN(new_n387));
  XOR2_X1   g186(.A(new_n387), .B(KEYINPUT64), .Z(new_n388));
  NAND2_X1  g187(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT33), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n351), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n389), .A2(KEYINPUT32), .ZN(new_n392));
  XNOR2_X1  g191(.A(new_n391), .B(new_n392), .ZN(new_n393));
  NOR3_X1   g192(.A1(new_n386), .A2(KEYINPUT34), .A3(new_n388), .ZN(new_n394));
  INV_X1    g193(.A(new_n386), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(new_n387), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n394), .B1(KEYINPUT34), .B2(new_n396), .ZN(new_n397));
  XNOR2_X1  g196(.A(new_n393), .B(new_n397), .ZN(new_n398));
  XOR2_X1   g197(.A(new_n398), .B(KEYINPUT36), .Z(new_n399));
  INV_X1    g198(.A(KEYINPUT69), .ZN(new_n400));
  XNOR2_X1  g199(.A(new_n377), .B(new_n400), .ZN(new_n401));
  AND2_X1   g200(.A1(G226gat), .A2(G233gat), .ZN(new_n402));
  NOR3_X1   g201(.A1(new_n401), .A2(KEYINPUT29), .A3(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n377), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n403), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  XNOR2_X1  g204(.A(G197gat), .B(G204gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(KEYINPUT68), .B(G218gat), .ZN(new_n407));
  AND2_X1   g206(.A1(new_n407), .A2(G211gat), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n406), .B1(new_n408), .B2(KEYINPUT22), .ZN(new_n409));
  XNOR2_X1  g208(.A(G211gat), .B(G218gat), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n409), .B(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n405), .A2(new_n411), .ZN(new_n412));
  XOR2_X1   g211(.A(G8gat), .B(G36gat), .Z(new_n413));
  XNOR2_X1  g212(.A(new_n413), .B(KEYINPUT70), .ZN(new_n414));
  XNOR2_X1  g213(.A(G64gat), .B(G92gat), .ZN(new_n415));
  XOR2_X1   g214(.A(new_n414), .B(new_n415), .Z(new_n416));
  NOR3_X1   g215(.A1(new_n404), .A2(KEYINPUT29), .A3(new_n402), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n417), .B1(new_n401), .B2(new_n402), .ZN(new_n418));
  OR2_X1    g217(.A1(new_n418), .A2(new_n411), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n412), .A2(new_n416), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(KEYINPUT71), .ZN(new_n421));
  OR2_X1    g220(.A1(new_n421), .A2(KEYINPUT30), .ZN(new_n422));
  INV_X1    g221(.A(new_n416), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n412), .A2(new_n419), .ZN(new_n424));
  AOI22_X1  g223(.A1(new_n421), .A2(KEYINPUT30), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n422), .A2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  XNOR2_X1  g226(.A(G141gat), .B(G148gat), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT2), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n429), .B1(G155gat), .B2(G162gat), .ZN(new_n430));
  INV_X1    g229(.A(G155gat), .ZN(new_n431));
  INV_X1    g230(.A(G162gat), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  OAI22_X1  g232(.A1(new_n428), .A2(new_n430), .B1(KEYINPUT72), .B2(new_n433), .ZN(new_n434));
  XOR2_X1   g233(.A(G155gat), .B(G162gat), .Z(new_n435));
  OR2_X1    g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n434), .A2(new_n435), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT73), .ZN(new_n439));
  XNOR2_X1  g238(.A(new_n438), .B(new_n439), .ZN(new_n440));
  AND2_X1   g239(.A1(new_n440), .A2(new_n384), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(KEYINPUT4), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT3), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n438), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n436), .A2(KEYINPUT3), .A3(new_n437), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n385), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(G225gat), .A2(G233gat), .ZN(new_n447));
  AND2_X1   g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n384), .A2(new_n438), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT4), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n442), .A2(new_n448), .A3(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT5), .ZN(new_n453));
  XNOR2_X1  g252(.A(new_n384), .B(new_n438), .ZN(new_n454));
  INV_X1    g253(.A(new_n447), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n453), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n441), .A2(new_n450), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n449), .A2(KEYINPUT4), .ZN(new_n458));
  XNOR2_X1  g257(.A(new_n458), .B(KEYINPUT74), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  AND2_X1   g259(.A1(new_n448), .A2(new_n453), .ZN(new_n461));
  AOI22_X1  g260(.A1(new_n452), .A2(new_n456), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  XOR2_X1   g261(.A(G1gat), .B(G29gat), .Z(new_n463));
  XNOR2_X1  g262(.A(new_n463), .B(KEYINPUT0), .ZN(new_n464));
  XNOR2_X1  g263(.A(G57gat), .B(G85gat), .ZN(new_n465));
  XNOR2_X1  g264(.A(new_n464), .B(new_n465), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n462), .A2(new_n466), .ZN(new_n467));
  OR2_X1    g266(.A1(new_n467), .A2(KEYINPUT75), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT6), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n467), .A2(KEYINPUT75), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n462), .A2(new_n466), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n468), .A2(new_n469), .A3(new_n470), .A4(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n467), .A2(KEYINPUT6), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n427), .A2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT29), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n444), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(new_n411), .ZN(new_n478));
  XOR2_X1   g277(.A(new_n409), .B(new_n410), .Z(new_n479));
  AOI21_X1  g278(.A(KEYINPUT3), .B1(new_n479), .B2(new_n476), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n478), .B1(new_n480), .B2(new_n438), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n481), .A2(G228gat), .A3(G233gat), .ZN(new_n482));
  NAND2_X1  g281(.A1(G228gat), .A2(G233gat), .ZN(new_n483));
  OAI211_X1 g282(.A(new_n483), .B(new_n478), .C1(new_n480), .C2(new_n440), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  XNOR2_X1  g284(.A(new_n485), .B(KEYINPUT77), .ZN(new_n486));
  XOR2_X1   g285(.A(KEYINPUT31), .B(G50gat), .Z(new_n487));
  XNOR2_X1  g286(.A(new_n486), .B(new_n487), .ZN(new_n488));
  XOR2_X1   g287(.A(G78gat), .B(G106gat), .Z(new_n489));
  XNOR2_X1  g288(.A(new_n489), .B(KEYINPUT76), .ZN(new_n490));
  XNOR2_X1  g289(.A(new_n490), .B(G22gat), .ZN(new_n491));
  AND2_X1   g290(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n488), .A2(new_n491), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n399), .B1(new_n475), .B2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(new_n494), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n447), .B1(new_n460), .B2(new_n446), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT39), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  OR2_X1    g298(.A1(new_n454), .A2(new_n455), .ZN(new_n500));
  OR2_X1    g299(.A1(new_n500), .A2(KEYINPUT78), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(KEYINPUT78), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n501), .A2(KEYINPUT39), .A3(new_n502), .ZN(new_n503));
  OAI211_X1 g302(.A(new_n499), .B(new_n466), .C1(new_n497), .C2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT40), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n467), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  OAI211_X1 g305(.A(new_n426), .B(new_n506), .C1(new_n505), .C2(new_n504), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT37), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n418), .A2(new_n479), .ZN(new_n509));
  AOI211_X1 g308(.A(new_n508), .B(new_n509), .C1(new_n405), .C2(new_n479), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n510), .B(KEYINPUT79), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n423), .B1(new_n424), .B2(KEYINPUT37), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n512), .A2(KEYINPUT38), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  OR2_X1    g313(.A1(new_n473), .A2(KEYINPUT80), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n471), .A2(new_n469), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n516), .A2(new_n467), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n473), .A2(KEYINPUT80), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n515), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n508), .B1(new_n412), .B2(new_n419), .ZN(new_n520));
  OAI21_X1  g319(.A(KEYINPUT38), .B1(new_n512), .B2(new_n520), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n514), .A2(new_n420), .A3(new_n519), .A4(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n496), .A2(new_n507), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n495), .A2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(new_n398), .ZN(new_n525));
  OAI21_X1  g324(.A(KEYINPUT81), .B1(new_n494), .B2(new_n525), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n426), .B1(new_n473), .B2(new_n472), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT81), .ZN(new_n528));
  OAI211_X1 g327(.A(new_n528), .B(new_n398), .C1(new_n492), .C2(new_n493), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n526), .A2(new_n527), .A3(new_n529), .ZN(new_n530));
  AND2_X1   g329(.A1(new_n530), .A2(KEYINPUT35), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n422), .A2(new_n425), .A3(new_n398), .ZN(new_n532));
  NOR4_X1   g331(.A1(new_n494), .A2(new_n532), .A3(KEYINPUT35), .A4(new_n519), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n524), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT91), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n213), .B(new_n290), .ZN(new_n536));
  NAND2_X1  g335(.A1(G229gat), .A2(G233gat), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n537), .B(KEYINPUT87), .ZN(new_n538));
  XOR2_X1   g337(.A(new_n538), .B(KEYINPUT13), .Z(new_n539));
  NAND2_X1  g338(.A1(new_n536), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n213), .A2(new_n290), .ZN(new_n541));
  OR3_X1    g340(.A1(new_n295), .A2(new_n293), .A3(new_n211), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n541), .A2(new_n538), .A3(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT89), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT18), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n544), .A2(new_n545), .ZN(new_n547));
  NAND4_X1  g346(.A1(new_n541), .A2(new_n542), .A3(new_n538), .A4(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n540), .A2(new_n546), .A3(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT90), .ZN(new_n550));
  XNOR2_X1  g349(.A(G113gat), .B(G141gat), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n551), .B(G197gat), .ZN(new_n552));
  XOR2_X1   g351(.A(KEYINPUT11), .B(G169gat), .Z(new_n553));
  XNOR2_X1  g352(.A(new_n552), .B(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n554), .B(KEYINPUT12), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n555), .B(KEYINPUT82), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n549), .A2(new_n550), .A3(new_n556), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n540), .A2(new_n546), .A3(new_n548), .A4(new_n555), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n550), .B1(new_n549), .B2(new_n556), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n534), .A2(new_n535), .A3(new_n562), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n533), .B1(new_n530), .B2(KEYINPUT35), .ZN(new_n564));
  INV_X1    g363(.A(new_n524), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  OAI21_X1  g365(.A(KEYINPUT91), .B1(new_n566), .B2(new_n561), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n348), .B1(new_n563), .B2(new_n567), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n474), .A2(KEYINPUT100), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT100), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n570), .B1(new_n472), .B2(new_n473), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n568), .A2(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n573), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g373(.A1(new_n563), .A2(new_n567), .ZN(new_n575));
  INV_X1    g374(.A(new_n348), .ZN(new_n576));
  XOR2_X1   g375(.A(KEYINPUT16), .B(G8gat), .Z(new_n577));
  AND4_X1   g376(.A1(new_n426), .A2(new_n575), .A3(new_n576), .A4(new_n577), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n202), .B1(new_n568), .B2(new_n426), .ZN(new_n579));
  OAI21_X1  g378(.A(KEYINPUT42), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n568), .A2(new_n426), .A3(new_n577), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT42), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n580), .A2(new_n583), .ZN(G1325gat));
  INV_X1    g383(.A(new_n568), .ZN(new_n585));
  OR3_X1    g384(.A1(new_n585), .A2(G15gat), .A3(new_n525), .ZN(new_n586));
  INV_X1    g385(.A(new_n399), .ZN(new_n587));
  OAI21_X1  g386(.A(G15gat), .B1(new_n585), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n586), .A2(new_n588), .ZN(G1326gat));
  NAND2_X1  g388(.A1(new_n568), .A2(new_n494), .ZN(new_n590));
  XNOR2_X1  g389(.A(KEYINPUT43), .B(G22gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n590), .B(new_n591), .ZN(G1327gat));
  NAND3_X1  g391(.A1(new_n246), .A2(new_n303), .A3(new_n347), .ZN(new_n593));
  XOR2_X1   g392(.A(new_n593), .B(KEYINPUT101), .Z(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n595), .B1(new_n563), .B2(new_n567), .ZN(new_n596));
  INV_X1    g395(.A(G29gat), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n596), .A2(new_n597), .A3(new_n572), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT45), .ZN(new_n599));
  OR2_X1    g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n534), .A2(KEYINPUT44), .A3(new_n303), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT44), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n602), .B1(new_n566), .B2(new_n302), .ZN(new_n603));
  AND2_X1   g402(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n246), .B(KEYINPUT102), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n605), .A2(new_n562), .A3(new_n347), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(KEYINPUT103), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n604), .A2(new_n572), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(G29gat), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n598), .A2(new_n599), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n600), .A2(new_n609), .A3(new_n610), .ZN(G1328gat));
  INV_X1    g410(.A(G36gat), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n596), .A2(new_n612), .A3(new_n426), .ZN(new_n613));
  OR2_X1    g412(.A1(new_n613), .A2(KEYINPUT46), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n604), .A2(new_n426), .A3(new_n607), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n615), .A2(G36gat), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n613), .A2(KEYINPUT46), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n614), .A2(new_n616), .A3(new_n617), .ZN(G1329gat));
  NOR2_X1   g417(.A1(new_n587), .A2(new_n275), .ZN(new_n619));
  AND4_X1   g418(.A1(new_n603), .A2(new_n601), .A3(new_n607), .A4(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT47), .ZN(new_n622));
  AOI211_X1 g421(.A(new_n525), .B(new_n595), .C1(new_n563), .C2(new_n567), .ZN(new_n623));
  OAI211_X1 g422(.A(new_n621), .B(new_n622), .C1(new_n623), .C2(G43gat), .ZN(new_n624));
  AOI21_X1  g423(.A(G43gat), .B1(new_n596), .B2(new_n398), .ZN(new_n625));
  OAI21_X1  g424(.A(KEYINPUT47), .B1(new_n625), .B2(new_n620), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n624), .A2(new_n626), .ZN(G1330gat));
  AND2_X1   g426(.A1(new_n494), .A2(G50gat), .ZN(new_n628));
  AND4_X1   g427(.A1(new_n603), .A2(new_n601), .A3(new_n607), .A4(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT48), .ZN(new_n631));
  AOI211_X1 g430(.A(new_n496), .B(new_n595), .C1(new_n563), .C2(new_n567), .ZN(new_n632));
  OAI211_X1 g431(.A(new_n630), .B(new_n631), .C1(new_n632), .C2(G50gat), .ZN(new_n633));
  AOI21_X1  g432(.A(G50gat), .B1(new_n596), .B2(new_n494), .ZN(new_n634));
  OAI21_X1  g433(.A(KEYINPUT48), .B1(new_n634), .B2(new_n629), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n633), .A2(new_n635), .ZN(G1331gat));
  NOR4_X1   g435(.A1(new_n246), .A2(new_n562), .A3(new_n347), .A4(new_n303), .ZN(new_n637));
  AND2_X1   g436(.A1(new_n534), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n638), .A2(new_n572), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g439(.A(new_n427), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n638), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(KEYINPUT104), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n642), .A2(KEYINPUT104), .ZN(new_n645));
  OAI22_X1  g444(.A1(new_n644), .A2(new_n645), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n646));
  INV_X1    g445(.A(new_n645), .ZN(new_n647));
  NOR2_X1   g446(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n647), .A2(new_n648), .A3(new_n643), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n646), .A2(new_n649), .ZN(G1333gat));
  NAND3_X1  g449(.A1(new_n638), .A2(G71gat), .A3(new_n399), .ZN(new_n651));
  INV_X1    g450(.A(G71gat), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n534), .A2(new_n398), .A3(new_n637), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n652), .B1(new_n654), .B2(KEYINPUT105), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT105), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n651), .B1(new_n655), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n658), .A2(KEYINPUT50), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT50), .ZN(new_n660));
  OAI211_X1 g459(.A(new_n660), .B(new_n651), .C1(new_n655), .C2(new_n657), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n659), .A2(new_n661), .ZN(G1334gat));
  NAND2_X1  g461(.A1(new_n638), .A2(new_n494), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(G78gat), .ZN(G1335gat));
  INV_X1    g463(.A(new_n246), .ZN(new_n665));
  NOR3_X1   g464(.A1(new_n665), .A2(new_n562), .A3(new_n347), .ZN(new_n666));
  AND3_X1   g465(.A1(new_n604), .A2(new_n572), .A3(new_n666), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n665), .A2(new_n562), .ZN(new_n668));
  NAND4_X1  g467(.A1(new_n534), .A2(KEYINPUT51), .A3(new_n303), .A4(new_n668), .ZN(new_n669));
  OAI211_X1 g468(.A(new_n303), .B(new_n668), .C1(new_n564), .C2(new_n565), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT51), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n572), .A2(new_n252), .A3(new_n346), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(KEYINPUT106), .ZN(new_n676));
  OAI22_X1  g475(.A1(new_n667), .A2(new_n252), .B1(new_n674), .B2(new_n676), .ZN(G1336gat));
  INV_X1    g476(.A(KEYINPUT107), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n669), .A2(new_n672), .A3(new_n678), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n670), .A2(KEYINPUT107), .A3(new_n671), .ZN(new_n680));
  NOR3_X1   g479(.A1(new_n427), .A2(G92gat), .A3(new_n347), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n679), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  NAND4_X1  g481(.A1(new_n601), .A2(new_n603), .A3(new_n426), .A4(new_n666), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(G92gat), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n685), .A2(KEYINPUT52), .ZN(new_n686));
  AOI21_X1  g485(.A(KEYINPUT52), .B1(new_n673), .B2(new_n681), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(new_n684), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n686), .A2(new_n688), .ZN(G1337gat));
  NAND3_X1  g488(.A1(new_n604), .A2(new_n399), .A3(new_n666), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n690), .A2(G99gat), .ZN(new_n691));
  NOR3_X1   g490(.A1(new_n525), .A2(G99gat), .A3(new_n347), .ZN(new_n692));
  XOR2_X1   g491(.A(new_n692), .B(KEYINPUT108), .Z(new_n693));
  OAI21_X1  g492(.A(new_n691), .B1(new_n674), .B2(new_n693), .ZN(G1338gat));
  NOR3_X1   g493(.A1(new_n496), .A2(G106gat), .A3(new_n347), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n679), .A2(new_n680), .A3(new_n695), .ZN(new_n696));
  NAND4_X1  g495(.A1(new_n601), .A2(new_n603), .A3(new_n494), .A4(new_n666), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n697), .A2(G106gat), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(KEYINPUT53), .ZN(new_n700));
  AOI21_X1  g499(.A(KEYINPUT53), .B1(new_n673), .B2(new_n695), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(new_n698), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n700), .A2(new_n702), .ZN(G1339gat));
  INV_X1    g502(.A(new_n572), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT54), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n705), .B1(new_n334), .B2(new_n335), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n341), .A2(new_n342), .A3(new_n706), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n328), .A2(new_n705), .A3(new_n336), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT109), .ZN(new_n709));
  AND3_X1   g508(.A1(new_n708), .A2(new_n709), .A3(new_n308), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n709), .B1(new_n708), .B2(new_n308), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n707), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT55), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n707), .A2(KEYINPUT55), .ZN(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n716), .B1(new_n710), .B2(new_n711), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT110), .ZN(new_n718));
  AND3_X1   g517(.A1(new_n717), .A2(new_n718), .A3(new_n345), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n718), .B1(new_n717), .B2(new_n345), .ZN(new_n720));
  OAI211_X1 g519(.A(new_n562), .B(new_n714), .C1(new_n719), .C2(new_n720), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n536), .A2(new_n539), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n538), .B1(new_n541), .B2(new_n542), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n554), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  OR2_X1    g523(.A1(new_n724), .A2(KEYINPUT111), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(KEYINPUT111), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n725), .A2(new_n558), .A3(new_n726), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n347), .A2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n303), .B1(new_n721), .B2(new_n729), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n727), .A2(new_n302), .ZN(new_n731));
  OAI211_X1 g530(.A(new_n714), .B(new_n731), .C1(new_n719), .C2(new_n720), .ZN(new_n732));
  INV_X1    g531(.A(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n605), .B1(new_n730), .B2(new_n733), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n348), .A2(new_n562), .ZN(new_n735));
  INV_X1    g534(.A(new_n735), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n704), .B1(new_n734), .B2(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n526), .A2(new_n529), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n738), .A2(new_n426), .ZN(new_n739));
  AND2_X1   g538(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n561), .A2(G113gat), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n494), .B1(new_n734), .B2(new_n736), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n704), .A2(new_n532), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n742), .A2(new_n562), .A3(new_n743), .ZN(new_n744));
  AOI22_X1  g543(.A1(new_n740), .A2(new_n741), .B1(new_n744), .B2(G113gat), .ZN(new_n745));
  XOR2_X1   g544(.A(new_n745), .B(KEYINPUT112), .Z(G1340gat));
  NOR2_X1   g545(.A1(new_n347), .A2(G120gat), .ZN(new_n747));
  XOR2_X1   g546(.A(new_n747), .B(KEYINPUT113), .Z(new_n748));
  NAND2_X1  g547(.A1(new_n740), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n742), .A2(new_n743), .ZN(new_n750));
  OAI21_X1  g549(.A(G120gat), .B1(new_n750), .B2(new_n347), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n749), .A2(new_n751), .ZN(G1341gat));
  INV_X1    g551(.A(G127gat), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n740), .A2(new_n753), .A3(new_n665), .ZN(new_n754));
  OAI21_X1  g553(.A(G127gat), .B1(new_n750), .B2(new_n605), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(G1342gat));
  INV_X1    g555(.A(G134gat), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n740), .A2(new_n757), .A3(new_n303), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT56), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n758), .B(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT115), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n742), .A2(new_n303), .A3(new_n743), .ZN(new_n762));
  AOI21_X1  g561(.A(KEYINPUT114), .B1(new_n762), .B2(G134gat), .ZN(new_n763));
  AND3_X1   g562(.A1(new_n762), .A2(KEYINPUT114), .A3(G134gat), .ZN(new_n764));
  OAI211_X1 g563(.A(new_n760), .B(new_n761), .C1(new_n763), .C2(new_n764), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n758), .B(KEYINPUT56), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n764), .A2(new_n763), .ZN(new_n767));
  OAI21_X1  g566(.A(KEYINPUT115), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n765), .A2(new_n768), .ZN(G1343gat));
  NOR3_X1   g568(.A1(new_n496), .A2(new_n399), .A3(new_n426), .ZN(new_n770));
  AND2_X1   g569(.A1(new_n737), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n561), .A2(G141gat), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT58), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n773), .B1(KEYINPUT117), .B2(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n734), .A2(new_n736), .ZN(new_n776));
  AOI21_X1  g575(.A(KEYINPUT57), .B1(new_n776), .B2(new_n494), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n494), .A2(KEYINPUT57), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT116), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n561), .B1(new_n713), .B2(new_n712), .ZN(new_n780));
  AND2_X1   g579(.A1(new_n717), .A2(new_n345), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n728), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n779), .B1(new_n782), .B2(new_n303), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(new_n732), .ZN(new_n784));
  NOR3_X1   g583(.A1(new_n782), .A2(new_n779), .A3(new_n303), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n246), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n778), .B1(new_n786), .B2(new_n736), .ZN(new_n787));
  OR2_X1    g586(.A1(new_n777), .A2(new_n787), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n704), .A2(new_n426), .A3(new_n399), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n788), .A2(new_n562), .A3(new_n789), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n775), .B1(new_n790), .B2(G141gat), .ZN(new_n791));
  AND2_X1   g590(.A1(new_n774), .A2(KEYINPUT117), .ZN(new_n792));
  XNOR2_X1  g591(.A(new_n791), .B(new_n792), .ZN(G1344gat));
  INV_X1    g592(.A(G148gat), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n771), .A2(new_n794), .A3(new_n346), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n788), .A2(new_n789), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n796), .A2(new_n347), .ZN(new_n797));
  NOR3_X1   g596(.A1(new_n797), .A2(KEYINPUT59), .A3(new_n794), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT59), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT57), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n732), .B1(new_n782), .B2(new_n303), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n735), .B1(new_n801), .B2(new_n246), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n800), .B1(new_n802), .B2(new_n496), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n778), .B1(new_n734), .B2(new_n736), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n803), .B1(new_n804), .B2(KEYINPUT118), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT118), .ZN(new_n806));
  AOI211_X1 g605(.A(new_n806), .B(new_n778), .C1(new_n734), .C2(new_n736), .ZN(new_n807));
  OR2_X1    g606(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n808), .A2(new_n346), .A3(new_n789), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n799), .B1(new_n809), .B2(G148gat), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n795), .B1(new_n798), .B2(new_n810), .ZN(G1345gat));
  OAI21_X1  g610(.A(G155gat), .B1(new_n796), .B2(new_n605), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n771), .A2(new_n431), .A3(new_n665), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(G1346gat));
  NAND3_X1  g613(.A1(new_n771), .A2(new_n432), .A3(new_n303), .ZN(new_n815));
  XNOR2_X1  g614(.A(new_n815), .B(KEYINPUT119), .ZN(new_n816));
  OAI21_X1  g615(.A(G162gat), .B1(new_n796), .B2(new_n302), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(G1347gat));
  OAI21_X1  g617(.A(KEYINPUT120), .B1(new_n572), .B2(new_n427), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT120), .ZN(new_n820));
  OAI211_X1 g619(.A(new_n820), .B(new_n426), .C1(new_n569), .C2(new_n571), .ZN(new_n821));
  AND3_X1   g620(.A1(new_n819), .A2(new_n398), .A3(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(new_n742), .ZN(new_n823));
  INV_X1    g622(.A(G169gat), .ZN(new_n824));
  NOR3_X1   g623(.A1(new_n823), .A2(new_n824), .A3(new_n561), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n572), .B1(new_n734), .B2(new_n736), .ZN(new_n826));
  NAND4_X1  g625(.A1(new_n826), .A2(new_n426), .A3(new_n526), .A4(new_n529), .ZN(new_n827));
  INV_X1    g626(.A(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(new_n562), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n825), .B1(new_n824), .B2(new_n829), .ZN(G1348gat));
  AOI21_X1  g629(.A(G176gat), .B1(new_n828), .B2(new_n346), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n822), .A2(new_n742), .A3(G176gat), .A4(new_n346), .ZN(new_n832));
  AND2_X1   g631(.A1(new_n832), .A2(KEYINPUT121), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n832), .A2(KEYINPUT121), .ZN(new_n834));
  NOR3_X1   g633(.A1(new_n831), .A2(new_n833), .A3(new_n834), .ZN(G1349gat));
  OAI21_X1  g634(.A(G183gat), .B1(new_n823), .B2(new_n605), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n665), .A2(new_n360), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n836), .B1(new_n827), .B2(new_n837), .ZN(new_n838));
  XNOR2_X1  g637(.A(new_n838), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g638(.A1(new_n828), .A2(new_n361), .A3(new_n303), .ZN(new_n840));
  OAI21_X1  g639(.A(G190gat), .B1(new_n823), .B2(new_n302), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n841), .A2(KEYINPUT61), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n841), .A2(KEYINPUT61), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n840), .B1(new_n842), .B2(new_n843), .ZN(G1351gat));
  AND4_X1   g643(.A1(new_n426), .A2(new_n826), .A3(new_n494), .A4(new_n587), .ZN(new_n845));
  XNOR2_X1  g644(.A(KEYINPUT122), .B(G197gat), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n845), .A2(new_n562), .A3(new_n846), .ZN(new_n847));
  XOR2_X1   g646(.A(new_n847), .B(KEYINPUT123), .Z(new_n848));
  NAND3_X1  g647(.A1(new_n819), .A2(new_n587), .A3(new_n821), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(KEYINPUT124), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT124), .ZN(new_n851));
  NAND4_X1  g650(.A1(new_n819), .A2(new_n851), .A3(new_n587), .A4(new_n821), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n808), .A2(new_n562), .A3(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT125), .ZN(new_n855));
  AND2_X1   g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(new_n846), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n857), .B1(new_n854), .B2(new_n855), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n848), .B1(new_n856), .B2(new_n858), .ZN(G1352gat));
  INV_X1    g658(.A(G204gat), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n845), .A2(new_n860), .A3(new_n346), .ZN(new_n861));
  XOR2_X1   g660(.A(new_n861), .B(KEYINPUT62), .Z(new_n862));
  NAND2_X1  g661(.A1(new_n808), .A2(new_n853), .ZN(new_n863));
  OAI21_X1  g662(.A(G204gat), .B1(new_n863), .B2(new_n347), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n862), .A2(new_n864), .ZN(G1353gat));
  INV_X1    g664(.A(G211gat), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n845), .A2(new_n866), .A3(new_n665), .ZN(new_n867));
  OAI211_X1 g666(.A(new_n665), .B(new_n853), .C1(new_n805), .C2(new_n807), .ZN(new_n868));
  AND3_X1   g667(.A1(new_n868), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n869));
  AOI21_X1  g668(.A(KEYINPUT63), .B1(new_n868), .B2(G211gat), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n867), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(KEYINPUT126), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT126), .ZN(new_n873));
  OAI211_X1 g672(.A(new_n873), .B(new_n867), .C1(new_n869), .C2(new_n870), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n872), .A2(new_n874), .ZN(G1354gat));
  AOI21_X1  g674(.A(G218gat), .B1(new_n845), .B2(new_n303), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT127), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n808), .A2(new_n877), .A3(new_n853), .ZN(new_n878));
  AND3_X1   g677(.A1(new_n878), .A2(new_n407), .A3(new_n303), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n863), .A2(KEYINPUT127), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n876), .B1(new_n879), .B2(new_n880), .ZN(G1355gat));
endmodule


