//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 0 1 1 1 0 0 1 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 1 0 1 1 0 0 0 1 0 0 0 1 1 1 0 0 1 0 0 0 0 1 0 0 0 1 1 0 1 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n737, new_n738, new_n739, new_n741, new_n742, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n774, new_n775,
    new_n776, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n840, new_n841,
    new_n843, new_n844, new_n845, new_n846, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n892, new_n893, new_n894, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n914, new_n915, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n958, new_n959, new_n960,
    new_n961, new_n962;
  INV_X1    g000(.A(KEYINPUT86), .ZN(new_n202));
  XNOR2_X1  g001(.A(G78gat), .B(G106gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(G22gat), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(G197gat), .B(G204gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT22), .ZN(new_n207));
  INV_X1    g006(.A(G211gat), .ZN(new_n208));
  INV_X1    g007(.A(G218gat), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n207), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n206), .A2(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(G211gat), .B(G218gat), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n212), .A2(new_n206), .A3(new_n210), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT29), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  XNOR2_X1  g017(.A(KEYINPUT78), .B(KEYINPUT3), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT75), .ZN(new_n221));
  INV_X1    g020(.A(G141gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(G148gat), .ZN(new_n223));
  INV_X1    g022(.A(G148gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(G141gat), .ZN(new_n225));
  AOI21_X1  g024(.A(KEYINPUT2), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  OR2_X1    g025(.A1(G155gat), .A2(G162gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(G155gat), .A2(G162gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n221), .B1(new_n226), .B2(new_n229), .ZN(new_n230));
  AND2_X1   g029(.A1(G155gat), .A2(G162gat), .ZN(new_n231));
  NOR2_X1   g030(.A1(G155gat), .A2(G162gat), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  XNOR2_X1  g032(.A(G141gat), .B(G148gat), .ZN(new_n234));
  OAI211_X1 g033(.A(new_n233), .B(KEYINPUT75), .C1(new_n234), .C2(KEYINPUT2), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT76), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n236), .B1(new_n222), .B2(G148gat), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n224), .A2(KEYINPUT76), .A3(G141gat), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n237), .A2(new_n223), .A3(new_n238), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n228), .B1(new_n227), .B2(KEYINPUT2), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n230), .A2(new_n235), .A3(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n220), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT72), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n216), .A2(new_n244), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n214), .A2(KEYINPUT72), .A3(new_n215), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND4_X1  g046(.A1(new_n230), .A2(new_n235), .A3(new_n241), .A4(new_n219), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(new_n217), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n243), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(G228gat), .ZN(new_n252));
  INV_X1    g051(.A(G233gat), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n251), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n250), .A2(KEYINPUT81), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n242), .A2(new_n217), .A3(new_n216), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n242), .A2(KEYINPUT3), .ZN(new_n257));
  AND4_X1   g056(.A1(G228gat), .A2(new_n256), .A3(G233gat), .A4(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT81), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n247), .A2(new_n259), .A3(new_n249), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n255), .A2(new_n258), .A3(new_n260), .ZN(new_n261));
  XOR2_X1   g060(.A(KEYINPUT31), .B(G50gat), .Z(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n254), .A2(new_n261), .A3(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n263), .B1(new_n254), .B2(new_n261), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n205), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n254), .A2(new_n261), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(new_n262), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n269), .A2(new_n264), .A3(new_n204), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n267), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n247), .ZN(new_n272));
  NAND2_X1  g071(.A1(G183gat), .A2(G190gat), .ZN(new_n273));
  NOR3_X1   g072(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n274));
  AOI21_X1  g073(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n275));
  NOR2_X1   g074(.A1(G169gat), .A2(G176gat), .ZN(new_n276));
  OAI22_X1  g075(.A1(new_n274), .A2(KEYINPUT68), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(G169gat), .ZN(new_n278));
  INV_X1    g077(.A(G176gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT68), .ZN(new_n281));
  NOR3_X1   g080(.A1(new_n280), .A2(new_n281), .A3(KEYINPUT26), .ZN(new_n282));
  OAI211_X1 g081(.A(KEYINPUT69), .B(new_n273), .C1(new_n277), .C2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(G190gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(KEYINPUT67), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT67), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(G190gat), .ZN(new_n287));
  AND2_X1   g086(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(KEYINPUT27), .B(G183gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(KEYINPUT28), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT28), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n288), .A2(new_n289), .A3(new_n292), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n283), .A2(new_n291), .A3(new_n293), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n281), .B1(new_n280), .B2(KEYINPUT26), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n274), .A2(KEYINPUT68), .ZN(new_n296));
  OAI211_X1 g095(.A(new_n295), .B(new_n296), .C1(new_n276), .C2(new_n275), .ZN(new_n297));
  AOI21_X1  g096(.A(KEYINPUT69), .B1(new_n297), .B2(new_n273), .ZN(new_n298));
  OAI21_X1  g097(.A(KEYINPUT66), .B1(G169gat), .B2(G176gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(KEYINPUT23), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT23), .ZN(new_n301));
  OAI211_X1 g100(.A(new_n301), .B(KEYINPUT66), .C1(G169gat), .C2(G176gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(G169gat), .A2(G176gat), .ZN(new_n303));
  AND3_X1   g102(.A1(new_n300), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(G183gat), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n285), .A2(new_n287), .A3(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT24), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n273), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g107(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n306), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  AND3_X1   g109(.A1(new_n304), .A2(new_n310), .A3(KEYINPUT25), .ZN(new_n311));
  XNOR2_X1  g110(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT65), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n308), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n273), .A2(KEYINPUT65), .A3(new_n307), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n305), .A2(new_n284), .ZN(new_n316));
  NAND4_X1  g115(.A1(new_n314), .A2(new_n315), .A3(new_n316), .A4(new_n309), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n312), .B1(new_n317), .B2(new_n304), .ZN(new_n318));
  OAI22_X1  g117(.A1(new_n294), .A2(new_n298), .B1(new_n311), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(G226gat), .A2(G233gat), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n217), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n273), .B1(new_n277), .B2(new_n282), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT69), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND4_X1  g124(.A1(new_n325), .A2(new_n283), .A3(new_n291), .A4(new_n293), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n304), .A2(new_n310), .A3(KEYINPUT25), .ZN(new_n327));
  AND2_X1   g126(.A1(new_n317), .A2(new_n304), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n327), .B1(new_n328), .B2(new_n312), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n322), .B1(new_n326), .B2(new_n329), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n272), .B1(new_n321), .B2(new_n330), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n319), .A2(new_n217), .A3(new_n320), .ZN(new_n332));
  NAND4_X1  g131(.A1(new_n326), .A2(new_n329), .A3(G226gat), .A4(G233gat), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n332), .A2(new_n247), .A3(new_n333), .ZN(new_n334));
  XNOR2_X1  g133(.A(G8gat), .B(G36gat), .ZN(new_n335));
  XNOR2_X1  g134(.A(G64gat), .B(G92gat), .ZN(new_n336));
  XOR2_X1   g135(.A(new_n335), .B(new_n336), .Z(new_n337));
  NAND3_X1  g136(.A1(new_n331), .A2(new_n334), .A3(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(KEYINPUT74), .B(KEYINPUT30), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(new_n337), .ZN(new_n341));
  NOR3_X1   g140(.A1(new_n321), .A2(new_n330), .A3(new_n272), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n247), .B1(new_n332), .B2(new_n333), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n341), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND4_X1  g143(.A1(new_n331), .A2(new_n334), .A3(KEYINPUT30), .A4(new_n337), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n340), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n271), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(G127gat), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n348), .A2(G134gat), .ZN(new_n349));
  INV_X1    g148(.A(G134gat), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n350), .A2(G127gat), .ZN(new_n351));
  OAI21_X1  g150(.A(KEYINPUT70), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n350), .A2(G127gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n348), .A2(G134gat), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT70), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(G113gat), .ZN(new_n357));
  INV_X1    g156(.A(G120gat), .ZN(new_n358));
  AOI21_X1  g157(.A(KEYINPUT1), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(G113gat), .A2(G120gat), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n352), .A2(new_n356), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n353), .A2(new_n354), .ZN(new_n363));
  NAND4_X1  g162(.A1(new_n363), .A2(KEYINPUT70), .A3(new_n360), .A4(new_n359), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n319), .A2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(G227gat), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n367), .A2(new_n253), .ZN(new_n368));
  AND2_X1   g167(.A1(new_n362), .A2(new_n364), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n326), .A2(new_n329), .A3(new_n369), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n366), .A2(new_n368), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(KEYINPUT32), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT33), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  XOR2_X1   g173(.A(G15gat), .B(G43gat), .Z(new_n375));
  XNOR2_X1  g174(.A(G71gat), .B(G99gat), .ZN(new_n376));
  XNOR2_X1  g175(.A(new_n375), .B(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n372), .A2(new_n374), .A3(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n377), .ZN(new_n379));
  OAI211_X1 g178(.A(new_n371), .B(KEYINPUT32), .C1(new_n373), .C2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(new_n368), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n319), .A2(new_n365), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n369), .B1(new_n326), .B2(new_n329), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n382), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(KEYINPUT34), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT34), .ZN(new_n387));
  OAI211_X1 g186(.A(new_n387), .B(new_n382), .C1(new_n383), .C2(new_n384), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n381), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n389), .A2(new_n378), .A3(new_n380), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT5), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n242), .A2(new_n364), .A3(new_n362), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n233), .B1(new_n234), .B2(KEYINPUT2), .ZN(new_n396));
  AOI22_X1  g195(.A1(new_n396), .A2(new_n221), .B1(new_n240), .B2(new_n239), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n365), .A2(new_n397), .A3(new_n235), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n395), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(G225gat), .A2(G233gat), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n394), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  AND3_X1   g201(.A1(new_n242), .A2(KEYINPUT77), .A3(KEYINPUT3), .ZN(new_n403));
  AOI21_X1  g202(.A(KEYINPUT77), .B1(new_n242), .B2(KEYINPUT3), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n369), .A2(new_n248), .ZN(new_n405));
  NOR3_X1   g204(.A1(new_n403), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  NAND4_X1  g205(.A1(new_n365), .A2(new_n397), .A3(KEYINPUT4), .A4(new_n235), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n369), .A2(new_n242), .ZN(new_n408));
  XNOR2_X1  g207(.A(KEYINPUT79), .B(KEYINPUT4), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  OAI211_X1 g209(.A(new_n400), .B(new_n407), .C1(new_n408), .C2(new_n410), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n402), .B1(new_n406), .B2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT77), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n257), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n242), .A2(KEYINPUT77), .A3(KEYINPUT3), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n414), .A2(new_n415), .A3(new_n369), .A4(new_n248), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n408), .A2(new_n410), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT4), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n398), .A2(new_n418), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n401), .A2(KEYINPUT5), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n416), .A2(new_n417), .A3(new_n419), .A4(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n412), .A2(new_n421), .ZN(new_n422));
  XNOR2_X1  g221(.A(G1gat), .B(G29gat), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n423), .B(KEYINPUT0), .ZN(new_n424));
  XNOR2_X1  g223(.A(G57gat), .B(G85gat), .ZN(new_n425));
  XOR2_X1   g224(.A(new_n424), .B(new_n425), .Z(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n422), .A2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT6), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n412), .A2(new_n421), .A3(new_n426), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  AOI211_X1 g230(.A(new_n429), .B(new_n426), .C1(new_n412), .C2(new_n421), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(KEYINPUT35), .B1(new_n431), .B2(new_n433), .ZN(new_n434));
  AND3_X1   g233(.A1(new_n347), .A2(new_n393), .A3(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT80), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n430), .A2(new_n429), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n426), .B1(new_n412), .B2(new_n421), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n340), .B1(new_n439), .B2(new_n432), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT73), .ZN(new_n441));
  AND3_X1   g240(.A1(new_n344), .A2(new_n345), .A3(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n441), .B1(new_n344), .B2(new_n345), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n436), .B1(new_n440), .B2(new_n444), .ZN(new_n445));
  AOI22_X1  g244(.A1(new_n431), .A2(new_n433), .B1(new_n338), .B2(new_n339), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n344), .A2(new_n345), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(KEYINPUT73), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n344), .A2(new_n441), .A3(new_n345), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n446), .A2(KEYINPUT80), .A3(new_n450), .ZN(new_n451));
  AOI22_X1  g250(.A1(KEYINPUT71), .A2(new_n389), .B1(new_n378), .B2(new_n380), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n389), .A2(new_n378), .A3(KEYINPUT71), .A4(new_n380), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n271), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n445), .A2(new_n451), .A3(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n435), .B1(new_n456), .B2(KEYINPUT35), .ZN(new_n457));
  AND2_X1   g256(.A1(new_n267), .A2(new_n270), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n458), .B1(new_n445), .B2(new_n451), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n419), .B1(new_n398), .B2(new_n409), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n401), .B1(new_n406), .B2(new_n460), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n399), .A2(new_n401), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT39), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  OAI211_X1 g264(.A(new_n463), .B(new_n401), .C1(new_n406), .C2(new_n460), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n465), .A2(new_n426), .A3(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT82), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n468), .A2(KEYINPUT40), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(new_n469), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n465), .A2(new_n426), .A3(new_n471), .A4(new_n466), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n346), .A2(new_n470), .A3(new_n428), .A4(new_n472), .ZN(new_n473));
  OAI21_X1  g272(.A(KEYINPUT37), .B1(new_n342), .B2(new_n343), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT37), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n331), .A2(new_n334), .A3(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n474), .A2(new_n341), .A3(new_n476), .ZN(new_n477));
  XOR2_X1   g276(.A(KEYINPUT83), .B(KEYINPUT38), .Z(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n474), .A2(new_n341), .A3(new_n478), .A4(new_n476), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n431), .A2(new_n433), .A3(new_n338), .ZN(new_n483));
  OAI211_X1 g282(.A(new_n473), .B(new_n458), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  AND4_X1   g283(.A1(KEYINPUT71), .A2(new_n389), .A3(new_n378), .A4(new_n380), .ZN(new_n485));
  OAI21_X1  g284(.A(KEYINPUT36), .B1(new_n485), .B2(new_n452), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT36), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n391), .A2(new_n487), .A3(new_n392), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n484), .A2(new_n489), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n459), .A2(new_n490), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n457), .A2(new_n491), .ZN(new_n492));
  XNOR2_X1  g291(.A(G43gat), .B(G50gat), .ZN(new_n493));
  OR2_X1    g292(.A1(new_n493), .A2(KEYINPUT15), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(KEYINPUT15), .ZN(new_n495));
  NAND2_X1  g294(.A1(G29gat), .A2(G36gat), .ZN(new_n496));
  NOR2_X1   g295(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n497));
  INV_X1    g296(.A(G36gat), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g298(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND4_X1  g300(.A1(new_n494), .A2(new_n495), .A3(new_n496), .A4(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(new_n500), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n503), .B1(KEYINPUT84), .B2(new_n499), .ZN(new_n504));
  OR2_X1    g303(.A1(new_n499), .A2(KEYINPUT84), .ZN(new_n505));
  AOI22_X1  g304(.A1(new_n504), .A2(new_n505), .B1(G29gat), .B2(G36gat), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n502), .B1(new_n506), .B2(new_n495), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT17), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  XNOR2_X1  g308(.A(G15gat), .B(G22gat), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT16), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n510), .B1(new_n511), .B2(G1gat), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n512), .B1(G1gat), .B2(new_n510), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT85), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n514), .B1(new_n510), .B2(G1gat), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n513), .A2(G8gat), .A3(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(G8gat), .ZN(new_n517));
  OAI221_X1 g316(.A(new_n512), .B1(new_n514), .B2(new_n517), .C1(G1gat), .C2(new_n510), .ZN(new_n518));
  AND2_X1   g317(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  OAI211_X1 g318(.A(new_n502), .B(KEYINPUT17), .C1(new_n506), .C2(new_n495), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n509), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(G229gat), .A2(G233gat), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n516), .A2(new_n518), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(new_n507), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n521), .A2(new_n522), .A3(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT18), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n521), .A2(KEYINPUT18), .A3(new_n522), .A4(new_n524), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n523), .B(new_n507), .ZN(new_n529));
  XOR2_X1   g328(.A(new_n522), .B(KEYINPUT13), .Z(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n527), .A2(new_n528), .A3(new_n531), .ZN(new_n532));
  XNOR2_X1  g331(.A(G113gat), .B(G141gat), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n533), .B(G197gat), .ZN(new_n534));
  XOR2_X1   g333(.A(KEYINPUT11), .B(G169gat), .Z(new_n535));
  XNOR2_X1  g334(.A(new_n534), .B(new_n535), .ZN(new_n536));
  XOR2_X1   g335(.A(new_n536), .B(KEYINPUT12), .Z(new_n537));
  NAND2_X1  g336(.A1(new_n532), .A2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n537), .ZN(new_n539));
  NAND4_X1  g338(.A1(new_n527), .A2(new_n539), .A3(new_n528), .A4(new_n531), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n202), .B1(new_n492), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n456), .A2(KEYINPUT35), .ZN(new_n544));
  INV_X1    g343(.A(new_n435), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AND2_X1   g345(.A1(new_n484), .A2(new_n489), .ZN(new_n547));
  NOR3_X1   g346(.A1(new_n440), .A2(new_n444), .A3(new_n436), .ZN(new_n548));
  AOI21_X1  g347(.A(KEYINPUT80), .B1(new_n446), .B2(new_n450), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n271), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n547), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n546), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n552), .A2(KEYINPUT86), .A3(new_n541), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n543), .A2(new_n553), .ZN(new_n554));
  XOR2_X1   g353(.A(G134gat), .B(G162gat), .Z(new_n555));
  XNOR2_X1  g354(.A(new_n555), .B(KEYINPUT90), .ZN(new_n556));
  AND2_X1   g355(.A1(G232gat), .A2(G233gat), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n557), .A2(KEYINPUT41), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n558), .B(KEYINPUT89), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n556), .B(new_n559), .ZN(new_n560));
  XOR2_X1   g359(.A(G99gat), .B(G106gat), .Z(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(G85gat), .ZN(new_n563));
  INV_X1    g362(.A(G92gat), .ZN(new_n564));
  OAI21_X1  g363(.A(KEYINPUT91), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT91), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n566), .A2(G85gat), .A3(G92gat), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n565), .A2(new_n567), .A3(KEYINPUT7), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT7), .ZN(new_n569));
  OAI211_X1 g368(.A(KEYINPUT91), .B(new_n569), .C1(new_n563), .C2(new_n564), .ZN(new_n570));
  NAND2_X1  g369(.A1(G99gat), .A2(G106gat), .ZN(new_n571));
  AOI22_X1  g370(.A1(KEYINPUT8), .A2(new_n571), .B1(new_n563), .B2(new_n564), .ZN(new_n572));
  NAND4_X1  g371(.A1(new_n562), .A2(new_n568), .A3(new_n570), .A4(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n568), .A2(new_n570), .A3(new_n572), .ZN(new_n575));
  AND2_X1   g374(.A1(new_n575), .A2(new_n561), .ZN(new_n576));
  OAI211_X1 g375(.A(new_n509), .B(new_n520), .C1(new_n574), .C2(new_n576), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n576), .A2(new_n574), .ZN(new_n578));
  AOI22_X1  g377(.A1(new_n578), .A2(new_n507), .B1(KEYINPUT41), .B2(new_n557), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(G190gat), .B(G218gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(KEYINPUT92), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n560), .B1(new_n584), .B2(KEYINPUT93), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n580), .B(new_n583), .ZN(new_n586));
  OR2_X1    g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n585), .A2(new_n586), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  XOR2_X1   g389(.A(G71gat), .B(G78gat), .Z(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT9), .ZN(new_n593));
  INV_X1    g392(.A(G71gat), .ZN(new_n594));
  INV_X1    g393(.A(G78gat), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n593), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  XOR2_X1   g395(.A(G57gat), .B(G64gat), .Z(new_n597));
  NAND3_X1  g396(.A1(new_n592), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n596), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(new_n591), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT21), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(G127gat), .B(G155gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n519), .B1(new_n602), .B2(new_n601), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(G231gat), .A2(G233gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(KEYINPUT87), .ZN(new_n609));
  XOR2_X1   g408(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  XOR2_X1   g410(.A(G183gat), .B(G211gat), .Z(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(KEYINPUT88), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n611), .B(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n607), .B(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n590), .A2(new_n615), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n601), .B1(new_n576), .B2(new_n574), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n575), .A2(new_n561), .ZN(new_n618));
  NAND4_X1  g417(.A1(new_n618), .A2(new_n573), .A3(new_n600), .A4(new_n598), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(G230gat), .A2(G233gat), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(G120gat), .B(G148gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(KEYINPUT95), .ZN(new_n625));
  XNOR2_X1  g424(.A(G176gat), .B(G204gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n623), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT10), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n617), .A2(new_n629), .A3(new_n619), .ZN(new_n630));
  OR2_X1    g429(.A1(new_n619), .A2(new_n629), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT94), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n622), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n630), .A2(new_n631), .A3(KEYINPUT94), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n628), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n632), .A2(new_n621), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n627), .B1(new_n637), .B2(new_n623), .ZN(new_n638));
  OR2_X1    g437(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n616), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n554), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n431), .A2(new_n433), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(KEYINPUT96), .B(G1gat), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n643), .B(new_n644), .ZN(G1324gat));
  INV_X1    g444(.A(KEYINPUT42), .ZN(new_n646));
  INV_X1    g445(.A(new_n346), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n641), .A2(new_n647), .ZN(new_n648));
  XOR2_X1   g447(.A(KEYINPUT16), .B(G8gat), .Z(new_n649));
  AOI21_X1  g448(.A(new_n646), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  OAI21_X1  g449(.A(G8gat), .B1(new_n641), .B2(new_n647), .ZN(new_n651));
  NOR2_X1   g450(.A1(KEYINPUT97), .A2(KEYINPUT42), .ZN(new_n652));
  MUX2_X1   g451(.A(KEYINPUT97), .B(new_n652), .S(new_n649), .Z(new_n653));
  AOI22_X1  g452(.A1(new_n650), .A2(new_n651), .B1(new_n648), .B2(new_n653), .ZN(G1325gat));
  INV_X1    g453(.A(new_n393), .ZN(new_n655));
  OR3_X1    g454(.A1(new_n641), .A2(G15gat), .A3(new_n655), .ZN(new_n656));
  OAI21_X1  g455(.A(G15gat), .B1(new_n641), .B2(new_n489), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(G1326gat));
  NAND3_X1  g457(.A1(new_n554), .A2(new_n271), .A3(new_n640), .ZN(new_n659));
  OR2_X1    g458(.A1(new_n659), .A2(KEYINPUT98), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(KEYINPUT98), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(KEYINPUT43), .B(G22gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n662), .B(new_n663), .ZN(G1327gat));
  NOR2_X1   g463(.A1(new_n615), .A2(new_n639), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n590), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n554), .A2(new_n667), .ZN(new_n668));
  NOR3_X1   g467(.A1(new_n668), .A2(G29gat), .A3(new_n642), .ZN(new_n669));
  XOR2_X1   g468(.A(new_n669), .B(KEYINPUT45), .Z(new_n670));
  INV_X1    g469(.A(KEYINPUT100), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT99), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n547), .B1(new_n459), .B2(new_n672), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n550), .A2(KEYINPUT99), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n546), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n590), .A2(KEYINPUT44), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n589), .B1(new_n457), .B2(new_n491), .ZN(new_n677));
  AOI22_X1  g476(.A1(new_n675), .A2(new_n676), .B1(new_n677), .B2(KEYINPUT44), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n666), .A2(new_n542), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n671), .B1(new_n678), .B2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT44), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n682), .B1(new_n552), .B2(new_n589), .ZN(new_n683));
  INV_X1    g482(.A(new_n676), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n550), .A2(KEYINPUT99), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n459), .A2(new_n672), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n685), .A2(new_n547), .A3(new_n686), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n684), .B1(new_n687), .B2(new_n546), .ZN(new_n688));
  OAI211_X1 g487(.A(KEYINPUT100), .B(new_n679), .C1(new_n683), .C2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n681), .A2(new_n689), .ZN(new_n690));
  OAI21_X1  g489(.A(G29gat), .B1(new_n690), .B2(new_n642), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n670), .A2(new_n691), .ZN(G1328gat));
  INV_X1    g491(.A(new_n667), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n693), .B1(new_n543), .B2(new_n553), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n694), .A2(new_n498), .A3(new_n346), .ZN(new_n695));
  XOR2_X1   g494(.A(new_n695), .B(KEYINPUT46), .Z(new_n696));
  OAI21_X1  g495(.A(G36gat), .B1(new_n690), .B2(new_n647), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(G1329gat));
  NAND2_X1  g497(.A1(new_n675), .A2(new_n676), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n677), .A2(KEYINPUT44), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(new_n679), .ZN(new_n702));
  OAI21_X1  g501(.A(G43gat), .B1(new_n702), .B2(new_n489), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT102), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n655), .A2(G43gat), .ZN(new_n705));
  AND3_X1   g504(.A1(new_n694), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n704), .B1(new_n694), .B2(new_n705), .ZN(new_n707));
  OAI211_X1 g506(.A(new_n703), .B(KEYINPUT47), .C1(new_n706), .C2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(new_n489), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n681), .A2(new_n709), .A3(new_n689), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT101), .ZN(new_n711));
  AND3_X1   g510(.A1(new_n710), .A2(new_n711), .A3(G43gat), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n711), .B1(new_n710), .B2(G43gat), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n706), .A2(new_n707), .ZN(new_n714));
  NOR3_X1   g513(.A1(new_n712), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n708), .B1(new_n715), .B2(KEYINPUT47), .ZN(G1330gat));
  NOR3_X1   g515(.A1(new_n668), .A2(G50gat), .A3(new_n458), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT48), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(G50gat), .B1(new_n702), .B2(new_n458), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n681), .A2(new_n271), .A3(new_n689), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n717), .B1(G50gat), .B2(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n721), .B1(KEYINPUT48), .B2(new_n723), .ZN(G1331gat));
  INV_X1    g523(.A(new_n675), .ZN(new_n725));
  INV_X1    g524(.A(new_n639), .ZN(new_n726));
  NOR4_X1   g525(.A1(new_n725), .A2(new_n541), .A3(new_n616), .A4(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(new_n642), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(G57gat), .ZN(G1332gat));
  XOR2_X1   g529(.A(new_n346), .B(KEYINPUT103), .Z(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n727), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n733), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n734));
  XOR2_X1   g533(.A(KEYINPUT49), .B(G64gat), .Z(new_n735));
  OAI21_X1  g534(.A(new_n734), .B1(new_n733), .B2(new_n735), .ZN(G1333gat));
  AOI21_X1  g535(.A(new_n594), .B1(new_n727), .B2(new_n709), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n655), .A2(G71gat), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n737), .B1(new_n727), .B2(new_n738), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g539(.A1(new_n727), .A2(new_n271), .ZN(new_n741));
  XNOR2_X1  g540(.A(KEYINPUT104), .B(G78gat), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n741), .B(new_n742), .ZN(G1335gat));
  NOR2_X1   g542(.A1(new_n541), .A2(new_n615), .ZN(new_n744));
  OAI211_X1 g543(.A(new_n639), .B(new_n744), .C1(new_n683), .C2(new_n688), .ZN(new_n745));
  OAI21_X1  g544(.A(G85gat), .B1(new_n745), .B2(new_n642), .ZN(new_n746));
  INV_X1    g545(.A(new_n744), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n590), .A2(new_n747), .ZN(new_n748));
  AOI21_X1  g547(.A(KEYINPUT51), .B1(new_n675), .B2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(new_n749), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n675), .A2(KEYINPUT51), .A3(new_n748), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n728), .A2(new_n563), .A3(new_n639), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(KEYINPUT105), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n746), .A2(new_n755), .ZN(G1336gat));
  INV_X1    g555(.A(KEYINPUT52), .ZN(new_n757));
  NOR3_X1   g556(.A1(new_n731), .A2(G92gat), .A3(new_n726), .ZN(new_n758));
  INV_X1    g557(.A(new_n751), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n758), .B1(new_n759), .B2(new_n749), .ZN(new_n760));
  OAI21_X1  g559(.A(KEYINPUT108), .B1(new_n745), .B2(new_n731), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(G92gat), .ZN(new_n762));
  NOR3_X1   g561(.A1(new_n745), .A2(KEYINPUT108), .A3(new_n731), .ZN(new_n763));
  OAI211_X1 g562(.A(new_n757), .B(new_n760), .C1(new_n762), .C2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n760), .A2(KEYINPUT106), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT106), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n752), .A2(new_n766), .A3(new_n758), .ZN(new_n767));
  OAI21_X1  g566(.A(G92gat), .B1(new_n745), .B2(new_n647), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n765), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT107), .ZN(new_n770));
  AND3_X1   g569(.A1(new_n769), .A2(new_n770), .A3(KEYINPUT52), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n770), .B1(new_n769), .B2(KEYINPUT52), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n764), .B1(new_n771), .B2(new_n772), .ZN(G1337gat));
  OAI21_X1  g572(.A(G99gat), .B1(new_n745), .B2(new_n489), .ZN(new_n774));
  NOR3_X1   g573(.A1(new_n655), .A2(G99gat), .A3(new_n726), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n752), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n774), .A2(new_n776), .ZN(G1338gat));
  OAI21_X1  g576(.A(G106gat), .B1(new_n745), .B2(new_n458), .ZN(new_n778));
  NOR3_X1   g577(.A1(new_n458), .A2(new_n726), .A3(G106gat), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n752), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(KEYINPUT110), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT110), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n778), .A2(new_n780), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n780), .A2(KEYINPUT109), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(KEYINPUT53), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n782), .A2(KEYINPUT53), .A3(new_n786), .A4(new_n784), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(G1339gat));
  INV_X1    g589(.A(KEYINPUT112), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n632), .A2(new_n633), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n792), .A2(new_n621), .A3(new_n635), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n630), .A2(new_n631), .A3(new_n622), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(KEYINPUT54), .ZN(new_n795));
  INV_X1    g594(.A(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n793), .A2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT54), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n632), .A2(new_n798), .A3(new_n621), .ZN(new_n799));
  INV_X1    g598(.A(new_n627), .ZN(new_n800));
  AND3_X1   g599(.A1(new_n799), .A2(KEYINPUT55), .A3(new_n800), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n636), .B1(new_n797), .B2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT55), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n795), .B1(new_n634), .B2(new_n635), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n799), .A2(new_n800), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n803), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n541), .A2(new_n802), .A3(new_n806), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n529), .A2(new_n530), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n522), .B1(new_n521), .B2(new_n524), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n536), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n540), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(new_n639), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n807), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(KEYINPUT111), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT111), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n807), .A2(new_n815), .A3(new_n812), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n814), .A2(new_n590), .A3(new_n816), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n589), .A2(new_n811), .A3(new_n806), .A4(new_n802), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n615), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NOR3_X1   g618(.A1(new_n616), .A2(new_n541), .A3(new_n639), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n791), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n816), .A2(new_n590), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n815), .B1(new_n807), .B2(new_n812), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n818), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(new_n615), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(new_n820), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n826), .A2(KEYINPUT112), .A3(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n821), .A2(new_n828), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n829), .A2(new_n642), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(new_n455), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n831), .A2(new_n732), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n541), .A2(new_n357), .ZN(new_n833));
  XNOR2_X1  g632(.A(new_n833), .B(KEYINPUT113), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n829), .A2(new_n271), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n836), .A2(new_n728), .A3(new_n393), .A4(new_n731), .ZN(new_n837));
  OAI21_X1  g636(.A(G113gat), .B1(new_n837), .B2(new_n542), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n835), .A2(new_n838), .ZN(G1340gat));
  NOR3_X1   g638(.A1(new_n837), .A2(new_n358), .A3(new_n726), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n832), .A2(new_n639), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n840), .B1(new_n841), .B2(new_n358), .ZN(G1341gat));
  NOR3_X1   g641(.A1(new_n837), .A2(new_n348), .A3(new_n825), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT114), .ZN(new_n844));
  XNOR2_X1  g643(.A(new_n843), .B(new_n844), .ZN(new_n845));
  AOI21_X1  g644(.A(G127gat), .B1(new_n832), .B2(new_n615), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n845), .A2(new_n846), .ZN(G1342gat));
  NAND2_X1  g646(.A1(new_n589), .A2(new_n647), .ZN(new_n848));
  XOR2_X1   g647(.A(new_n848), .B(KEYINPUT115), .Z(new_n849));
  OR3_X1    g648(.A1(new_n831), .A2(G134gat), .A3(new_n849), .ZN(new_n850));
  OR2_X1    g649(.A1(new_n850), .A2(KEYINPUT56), .ZN(new_n851));
  OAI21_X1  g650(.A(G134gat), .B1(new_n837), .B2(new_n590), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n850), .A2(KEYINPUT56), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(G1343gat));
  NOR3_X1   g653(.A1(new_n709), .A2(new_n732), .A3(new_n642), .ZN(new_n855));
  INV_X1    g654(.A(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n813), .A2(new_n590), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(new_n818), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n820), .B1(new_n825), .B2(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT57), .ZN(new_n860));
  NOR3_X1   g659(.A1(new_n859), .A2(new_n860), .A3(new_n458), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n821), .A2(new_n271), .A3(new_n828), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(new_n860), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT116), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n861), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n862), .A2(KEYINPUT116), .A3(new_n860), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n856), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n222), .B1(new_n867), .B2(new_n541), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n830), .A2(new_n271), .A3(new_n489), .ZN(new_n869));
  NOR4_X1   g668(.A1(new_n869), .A2(G141gat), .A3(new_n542), .A4(new_n732), .ZN(new_n870));
  OAI21_X1  g669(.A(KEYINPUT58), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(new_n870), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT58), .ZN(new_n873));
  AOI211_X1 g672(.A(new_n542), .B(new_n856), .C1(new_n865), .C2(new_n866), .ZN(new_n874));
  OAI211_X1 g673(.A(new_n872), .B(new_n873), .C1(new_n874), .C2(new_n222), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n871), .A2(new_n875), .ZN(G1344gat));
  NAND2_X1  g675(.A1(new_n224), .A2(KEYINPUT59), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n869), .A2(new_n732), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n877), .B1(new_n878), .B2(new_n639), .ZN(new_n879));
  NAND4_X1  g678(.A1(new_n821), .A2(new_n828), .A3(KEYINPUT57), .A4(new_n271), .ZN(new_n880));
  OR2_X1    g679(.A1(new_n858), .A2(KEYINPUT118), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n615), .B1(new_n858), .B2(KEYINPUT118), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n820), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n860), .B1(new_n883), .B2(new_n458), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n880), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n639), .A2(KEYINPUT59), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n886), .B1(new_n856), .B2(KEYINPUT117), .ZN(new_n887));
  OAI211_X1 g686(.A(new_n885), .B(new_n887), .C1(KEYINPUT117), .C2(new_n856), .ZN(new_n888));
  AOI211_X1 g687(.A(new_n726), .B(new_n856), .C1(new_n865), .C2(new_n866), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n888), .B1(new_n889), .B2(KEYINPUT59), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n879), .B1(new_n890), .B2(G148gat), .ZN(G1345gat));
  INV_X1    g690(.A(G155gat), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n878), .A2(new_n892), .A3(new_n615), .ZN(new_n893));
  AND2_X1   g692(.A1(new_n867), .A2(new_n615), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n893), .B1(new_n894), .B2(new_n892), .ZN(G1346gat));
  NAND2_X1  g694(.A1(new_n865), .A2(new_n866), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n896), .A2(new_n589), .A3(new_n855), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT119), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n867), .A2(KEYINPUT119), .A3(new_n589), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n899), .A2(G162gat), .A3(new_n900), .ZN(new_n901));
  OR3_X1    g700(.A1(new_n869), .A2(G162gat), .A3(new_n849), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(G1347gat));
  NAND2_X1  g702(.A1(new_n642), .A2(new_n346), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n655), .A2(new_n904), .ZN(new_n905));
  NAND4_X1  g704(.A1(new_n821), .A2(new_n828), .A3(new_n458), .A4(new_n905), .ZN(new_n906));
  NOR3_X1   g705(.A1(new_n906), .A2(new_n278), .A3(new_n542), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n829), .A2(new_n728), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n732), .A2(new_n455), .ZN(new_n909));
  XNOR2_X1  g708(.A(new_n909), .B(KEYINPUT120), .ZN(new_n910));
  AND2_X1   g709(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n911), .A2(new_n541), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n907), .B1(new_n912), .B2(new_n278), .ZN(G1348gat));
  NAND3_X1  g712(.A1(new_n911), .A2(new_n279), .A3(new_n639), .ZN(new_n914));
  OAI21_X1  g713(.A(G176gat), .B1(new_n906), .B2(new_n726), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(G1349gat));
  NOR2_X1   g715(.A1(KEYINPUT122), .A2(KEYINPUT60), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n911), .A2(new_n289), .A3(new_n615), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT121), .ZN(new_n919));
  OR3_X1    g718(.A1(new_n906), .A2(new_n919), .A3(new_n825), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n919), .B1(new_n906), .B2(new_n825), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n920), .A2(G183gat), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n917), .B1(new_n918), .B2(new_n922), .ZN(new_n923));
  AND2_X1   g722(.A1(KEYINPUT122), .A2(KEYINPUT60), .ZN(new_n924));
  XNOR2_X1  g723(.A(new_n923), .B(new_n924), .ZN(G1350gat));
  OAI21_X1  g724(.A(G190gat), .B1(new_n906), .B2(new_n590), .ZN(new_n926));
  XNOR2_X1  g725(.A(new_n926), .B(KEYINPUT61), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n911), .A2(new_n288), .A3(new_n589), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT123), .ZN(new_n929));
  AND2_X1   g728(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n928), .A2(new_n929), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n927), .B1(new_n930), .B2(new_n931), .ZN(G1351gat));
  NOR2_X1   g731(.A1(new_n709), .A2(new_n904), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n885), .A2(new_n933), .ZN(new_n934));
  INV_X1    g733(.A(new_n934), .ZN(new_n935));
  AND3_X1   g734(.A1(new_n935), .A2(G197gat), .A3(new_n541), .ZN(new_n936));
  NOR3_X1   g735(.A1(new_n709), .A2(new_n458), .A3(new_n731), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n908), .A2(new_n937), .ZN(new_n938));
  INV_X1    g737(.A(new_n938), .ZN(new_n939));
  AOI21_X1  g738(.A(G197gat), .B1(new_n939), .B2(new_n541), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n936), .A2(new_n940), .ZN(G1352gat));
  NOR3_X1   g740(.A1(new_n938), .A2(G204gat), .A3(new_n726), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT62), .ZN(new_n943));
  OR2_X1    g742(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  OAI21_X1  g743(.A(G204gat), .B1(new_n934), .B2(new_n726), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n942), .A2(new_n943), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(G1353gat));
  NAND3_X1  g746(.A1(new_n935), .A2(KEYINPUT125), .A3(new_n615), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT125), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n949), .B1(new_n934), .B2(new_n825), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n948), .A2(G211gat), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n951), .A2(KEYINPUT63), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT63), .ZN(new_n953));
  NAND4_X1  g752(.A1(new_n948), .A2(new_n953), .A3(new_n950), .A4(G211gat), .ZN(new_n954));
  NOR3_X1   g753(.A1(new_n938), .A2(G211gat), .A3(new_n825), .ZN(new_n955));
  XNOR2_X1  g754(.A(new_n955), .B(KEYINPUT124), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n952), .A2(new_n954), .A3(new_n956), .ZN(G1354gat));
  NOR2_X1   g756(.A1(new_n935), .A2(KEYINPUT126), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT126), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n589), .B1(new_n934), .B2(new_n959), .ZN(new_n960));
  OAI21_X1  g759(.A(G218gat), .B1(new_n958), .B2(new_n960), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n939), .A2(new_n209), .A3(new_n589), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n961), .A2(new_n962), .ZN(G1355gat));
endmodule


