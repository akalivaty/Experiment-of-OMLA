//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 1 0 1 0 0 1 0 0 0 0 0 0 0 0 1 1 0 1 1 1 0 0 1 1 0 1 0 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 0 0 0 0 0 0 0 1 0 0 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:04 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1287, new_n1288,
    new_n1289, new_n1290, new_n1291, new_n1292, new_n1293, new_n1294,
    new_n1295, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1308, new_n1309, new_n1310, new_n1311, new_n1312, new_n1313,
    new_n1314, new_n1315, new_n1316, new_n1317, new_n1319, new_n1320,
    new_n1321, new_n1322, new_n1323, new_n1324, new_n1325, new_n1326,
    new_n1327, new_n1329, new_n1330, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1379, new_n1380, new_n1381, new_n1382, new_n1383,
    new_n1384;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G13), .ZN(new_n204));
  OAI211_X1 g0004(.A(new_n204), .B(G250), .C1(G257), .C2(G264), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT0), .ZN(new_n206));
  OAI21_X1  g0006(.A(G50), .B1(G58), .B2(G68), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G1), .A2(G13), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n208), .A2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n213));
  INV_X1    g0013(.A(G77), .ZN(new_n214));
  INV_X1    g0014(.A(G244), .ZN(new_n215));
  INV_X1    g0015(.A(G87), .ZN(new_n216));
  INV_X1    g0016(.A(G250), .ZN(new_n217));
  OAI221_X1 g0017(.A(new_n213), .B1(new_n214), .B2(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n203), .B1(new_n218), .B2(new_n221), .ZN(new_n222));
  OAI211_X1 g0022(.A(new_n206), .B(new_n212), .C1(KEYINPUT1), .C2(new_n222), .ZN(new_n223));
  AOI21_X1  g0023(.A(new_n223), .B1(KEYINPUT1), .B2(new_n222), .ZN(G361));
  XOR2_X1   g0024(.A(G226), .B(G232), .Z(new_n225));
  XNOR2_X1  g0025(.A(G238), .B(G244), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n225), .B(new_n226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(KEYINPUT64), .B(KEYINPUT2), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XOR2_X1   g0029(.A(G264), .B(G270), .Z(new_n230));
  XNOR2_X1  g0030(.A(G250), .B(G257), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n229), .B(new_n232), .ZN(G358));
  XOR2_X1   g0033(.A(G87), .B(G97), .Z(new_n234));
  XOR2_X1   g0034(.A(G107), .B(G116), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G68), .B(G77), .Z(new_n237));
  XNOR2_X1  g0037(.A(G50), .B(G58), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n236), .B(new_n239), .Z(G351));
  INV_X1    g0040(.A(KEYINPUT8), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n241), .A2(G58), .ZN(new_n242));
  NOR2_X1   g0042(.A1(new_n242), .A2(KEYINPUT66), .ZN(new_n243));
  INV_X1    g0043(.A(G58), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n244), .A2(KEYINPUT8), .ZN(new_n245));
  AND2_X1   g0045(.A1(new_n242), .A2(new_n245), .ZN(new_n246));
  AOI21_X1  g0046(.A(new_n243), .B1(new_n246), .B2(KEYINPUT66), .ZN(new_n247));
  INV_X1    g0047(.A(G1), .ZN(new_n248));
  NAND3_X1  g0048(.A1(new_n248), .A2(G13), .A3(G20), .ZN(new_n249));
  INV_X1    g0049(.A(KEYINPUT68), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND4_X1  g0051(.A1(new_n248), .A2(KEYINPUT68), .A3(G13), .A4(G20), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n247), .A2(new_n253), .ZN(new_n254));
  AND2_X1   g0054(.A1(new_n251), .A2(new_n252), .ZN(new_n255));
  NAND3_X1  g0055(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(new_n209), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n210), .A2(G1), .ZN(new_n258));
  NOR3_X1   g0058(.A1(new_n255), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n254), .B1(new_n259), .B2(new_n247), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT16), .ZN(new_n261));
  INV_X1    g0061(.A(G68), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n244), .A2(new_n262), .ZN(new_n263));
  NOR2_X1   g0063(.A1(G58), .A2(G68), .ZN(new_n264));
  OAI21_X1  g0064(.A(G20), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NOR2_X1   g0065(.A1(G20), .A2(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G159), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  AND2_X1   g0068(.A1(KEYINPUT3), .A2(G33), .ZN(new_n269));
  NOR2_X1   g0069(.A1(KEYINPUT3), .A2(G33), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  AOI21_X1  g0071(.A(KEYINPUT7), .B1(new_n271), .B2(new_n210), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n262), .B1(new_n272), .B2(KEYINPUT80), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT3), .ZN(new_n274));
  INV_X1    g0074(.A(G33), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(KEYINPUT3), .A2(G33), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n276), .A2(new_n210), .A3(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT7), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT80), .ZN(new_n281));
  NAND4_X1  g0081(.A1(new_n276), .A2(KEYINPUT7), .A3(new_n210), .A4(new_n277), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n280), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  AOI211_X1 g0083(.A(new_n261), .B(new_n268), .C1(new_n273), .C2(new_n283), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n262), .B1(new_n280), .B2(new_n282), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n261), .B1(new_n285), .B2(new_n268), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(new_n257), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n260), .B1(new_n284), .B2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G169), .ZN(new_n289));
  NAND2_X1  g0089(.A1(G33), .A2(G41), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n290), .A2(G1), .A3(G13), .ZN(new_n291));
  INV_X1    g0091(.A(G223), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n292), .A2(G1698), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n293), .B1(new_n269), .B2(new_n270), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT81), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n276), .A2(new_n277), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n297), .A2(KEYINPUT81), .A3(new_n293), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  OAI211_X1 g0099(.A(G226), .B(G1698), .C1(new_n269), .C2(new_n270), .ZN(new_n300));
  NAND2_X1  g0100(.A1(G33), .A2(G87), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n291), .B1(new_n299), .B2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT65), .ZN(new_n305));
  AND2_X1   g0105(.A1(G33), .A2(G41), .ZN(new_n306));
  OAI21_X1  g0106(.A(G274), .B1(new_n306), .B2(new_n209), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n248), .B1(G41), .B2(G45), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n305), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n308), .ZN(new_n310));
  NAND4_X1  g0110(.A1(new_n310), .A2(new_n291), .A3(KEYINPUT65), .A4(G274), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n291), .A2(new_n308), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(G232), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n312), .A2(new_n315), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n289), .B1(new_n304), .B2(new_n316), .ZN(new_n317));
  AOI22_X1  g0117(.A1(new_n309), .A2(new_n311), .B1(new_n314), .B2(G232), .ZN(new_n318));
  INV_X1    g0118(.A(G179), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n302), .B1(new_n296), .B2(new_n298), .ZN(new_n320));
  OAI211_X1 g0120(.A(new_n318), .B(new_n319), .C1(new_n320), .C2(new_n291), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT82), .ZN(new_n322));
  AND3_X1   g0122(.A1(new_n317), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n322), .B1(new_n317), .B2(new_n321), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n288), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(KEYINPUT18), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n317), .A2(new_n321), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(KEYINPUT82), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n317), .A2(new_n321), .A3(new_n322), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT18), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n330), .A2(new_n331), .A3(new_n288), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT17), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n268), .B1(new_n273), .B2(new_n283), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(KEYINPUT16), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n335), .A2(new_n257), .A3(new_n286), .ZN(new_n336));
  OAI21_X1  g0136(.A(G200), .B1(new_n304), .B2(new_n316), .ZN(new_n337));
  OAI211_X1 g0137(.A(new_n318), .B(G190), .C1(new_n320), .C2(new_n291), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n336), .A2(new_n260), .A3(new_n337), .A4(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT83), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n333), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n337), .A2(new_n338), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n288), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n343), .A2(KEYINPUT83), .A3(KEYINPUT17), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n326), .A2(new_n332), .A3(new_n341), .A4(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(G238), .A2(G1698), .ZN(new_n346));
  INV_X1    g0146(.A(G232), .ZN(new_n347));
  OAI211_X1 g0147(.A(new_n297), .B(new_n346), .C1(new_n347), .C2(G1698), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n306), .A2(new_n209), .ZN(new_n349));
  OAI211_X1 g0149(.A(new_n348), .B(new_n349), .C1(G107), .C2(new_n297), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n350), .B1(new_n215), .B2(new_n313), .ZN(new_n351));
  INV_X1    g0151(.A(new_n312), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n353), .A2(G169), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT70), .ZN(new_n355));
  NOR3_X1   g0155(.A1(new_n351), .A2(G179), .A3(new_n352), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n354), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  OR2_X1    g0157(.A1(new_n356), .A2(new_n355), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n259), .A2(G77), .ZN(new_n359));
  INV_X1    g0159(.A(new_n257), .ZN(new_n360));
  XNOR2_X1  g0160(.A(KEYINPUT15), .B(G87), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n210), .A2(G33), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  AND3_X1   g0164(.A1(new_n362), .A2(KEYINPUT69), .A3(new_n364), .ZN(new_n365));
  AOI21_X1  g0165(.A(KEYINPUT69), .B1(new_n362), .B2(new_n364), .ZN(new_n366));
  INV_X1    g0166(.A(new_n266), .ZN(new_n367));
  OAI22_X1  g0167(.A1(new_n246), .A2(new_n367), .B1(new_n210), .B2(new_n214), .ZN(new_n368));
  NOR3_X1   g0168(.A1(new_n365), .A2(new_n366), .A3(new_n368), .ZN(new_n369));
  OAI221_X1 g0169(.A(new_n359), .B1(G77), .B2(new_n253), .C1(new_n360), .C2(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n357), .A2(new_n358), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n353), .A2(G190), .ZN(new_n372));
  INV_X1    g0172(.A(G200), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n372), .B1(new_n373), .B2(new_n353), .ZN(new_n374));
  OR2_X1    g0174(.A1(new_n374), .A2(new_n370), .ZN(new_n375));
  INV_X1    g0175(.A(G222), .ZN(new_n376));
  MUX2_X1   g0176(.A(new_n376), .B(new_n292), .S(G1698), .Z(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(new_n297), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n271), .A2(new_n214), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n378), .A2(new_n379), .A3(new_n349), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n314), .A2(G226), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n382), .A2(new_n352), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(new_n319), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n384), .B1(G169), .B2(new_n383), .ZN(new_n385));
  NOR2_X1   g0185(.A1(G50), .A2(G58), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n210), .B1(new_n386), .B2(new_n262), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n242), .A2(new_n245), .A3(KEYINPUT66), .ZN(new_n388));
  OAI211_X1 g0188(.A(new_n388), .B(new_n364), .C1(KEYINPUT66), .C2(new_n242), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n266), .A2(G150), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n387), .B1(new_n391), .B2(KEYINPUT67), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT67), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n389), .A2(new_n393), .A3(new_n390), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n360), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n253), .A2(G50), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n396), .B1(new_n259), .B2(G50), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n395), .A2(new_n398), .ZN(new_n399));
  OR2_X1    g0199(.A1(new_n385), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n371), .A2(new_n375), .A3(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT9), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n402), .B1(new_n395), .B2(new_n398), .ZN(new_n403));
  INV_X1    g0203(.A(new_n394), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n393), .B1(new_n389), .B2(new_n390), .ZN(new_n405));
  NOR3_X1   g0205(.A1(new_n404), .A2(new_n405), .A3(new_n387), .ZN(new_n406));
  OAI211_X1 g0206(.A(KEYINPUT9), .B(new_n397), .C1(new_n406), .C2(new_n360), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n312), .A2(new_n380), .A3(G190), .A4(new_n381), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(KEYINPUT72), .ZN(new_n409));
  OAI21_X1  g0209(.A(G200), .B1(new_n382), .B2(new_n352), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n291), .B1(new_n377), .B2(new_n297), .ZN(new_n411));
  AOI22_X1  g0211(.A1(new_n411), .A2(new_n379), .B1(G226), .B2(new_n314), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT72), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n412), .A2(new_n413), .A3(G190), .A4(new_n312), .ZN(new_n414));
  AND3_X1   g0214(.A1(new_n409), .A2(new_n410), .A3(new_n414), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n403), .A2(new_n407), .A3(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT71), .ZN(new_n417));
  AOI21_X1  g0217(.A(KEYINPUT10), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT10), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n409), .A2(new_n410), .A3(new_n414), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n420), .B1(new_n421), .B2(KEYINPUT71), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n422), .A2(new_n415), .A3(new_n407), .A4(new_n403), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n419), .A2(new_n423), .ZN(new_n424));
  NOR3_X1   g0224(.A1(new_n345), .A2(new_n401), .A3(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n309), .A2(KEYINPUT74), .A3(new_n311), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT75), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n313), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n291), .A2(KEYINPUT75), .A3(new_n308), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n428), .A2(G238), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n426), .A2(new_n430), .ZN(new_n431));
  AOI21_X1  g0231(.A(KEYINPUT74), .B1(new_n309), .B2(new_n311), .ZN(new_n432));
  OAI21_X1  g0232(.A(KEYINPUT76), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT74), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n312), .A2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT76), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n435), .A2(new_n436), .A3(new_n430), .A4(new_n426), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n433), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n347), .A2(G1698), .ZN(new_n439));
  OAI221_X1 g0239(.A(new_n439), .B1(G226), .B2(G1698), .C1(new_n269), .C2(new_n270), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT73), .ZN(new_n441));
  NAND2_X1  g0241(.A1(G33), .A2(G97), .ZN(new_n442));
  AND3_X1   g0242(.A1(new_n440), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n441), .B1(new_n440), .B2(new_n442), .ZN(new_n444));
  NOR3_X1   g0244(.A1(new_n443), .A2(new_n444), .A3(new_n291), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n438), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(KEYINPUT13), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT13), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n438), .A2(new_n449), .A3(new_n446), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n448), .A2(G190), .A3(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n449), .B1(new_n438), .B2(new_n446), .ZN(new_n452));
  AOI211_X1 g0252(.A(KEYINPUT13), .B(new_n445), .C1(new_n433), .C2(new_n437), .ZN(new_n453));
  OAI21_X1  g0253(.A(G200), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT12), .ZN(new_n455));
  OAI21_X1  g0255(.A(G68), .B1(new_n259), .B2(new_n455), .ZN(new_n456));
  AOI22_X1  g0256(.A1(new_n266), .A2(G50), .B1(G20), .B2(new_n262), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n457), .B1(new_n214), .B2(new_n363), .ZN(new_n458));
  AND2_X1   g0258(.A1(new_n458), .A2(new_n257), .ZN(new_n459));
  OR2_X1    g0259(.A1(new_n459), .A2(KEYINPUT11), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n255), .A2(KEYINPUT12), .A3(new_n262), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n458), .A2(KEYINPUT11), .A3(new_n257), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n253), .A2(new_n455), .ZN(new_n463));
  AND3_X1   g0263(.A1(new_n461), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n456), .A2(new_n460), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(KEYINPUT77), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT77), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n456), .A2(new_n460), .A3(new_n464), .A4(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n451), .A2(new_n454), .A3(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT78), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n451), .A2(new_n454), .A3(KEYINPUT78), .A4(new_n469), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT14), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n475), .B(G169), .C1(new_n452), .C2(new_n453), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n448), .A2(G179), .A3(new_n450), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT79), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n289), .B1(new_n448), .B2(new_n450), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n479), .B1(new_n480), .B2(new_n475), .ZN(new_n481));
  OAI21_X1  g0281(.A(G169), .B1(new_n452), .B2(new_n453), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n482), .A2(KEYINPUT79), .A3(KEYINPUT14), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n478), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  OAI211_X1 g0284(.A(new_n425), .B(new_n474), .C1(new_n469), .C2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(G41), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n248), .B(G45), .C1(new_n487), .C2(KEYINPUT5), .ZN(new_n488));
  AND2_X1   g0288(.A1(new_n487), .A2(KEYINPUT5), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n490), .A2(G274), .A3(new_n291), .ZN(new_n491));
  OAI211_X1 g0291(.A(G257), .B(new_n291), .C1(new_n488), .C2(new_n489), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n217), .B1(new_n276), .B2(new_n277), .ZN(new_n494));
  NOR2_X1   g0294(.A1(KEYINPUT85), .A2(KEYINPUT4), .ZN(new_n495));
  OAI21_X1  g0295(.A(G1698), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  OAI21_X1  g0296(.A(G244), .B1(new_n269), .B2(new_n270), .ZN(new_n497));
  AOI22_X1  g0297(.A1(new_n497), .A2(new_n495), .B1(G33), .B2(G283), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n215), .B1(new_n276), .B2(new_n277), .ZN(new_n499));
  INV_X1    g0299(.A(G1698), .ZN(new_n500));
  AOI21_X1  g0300(.A(KEYINPUT85), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT4), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n496), .B(new_n498), .C1(new_n501), .C2(new_n502), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n493), .B1(new_n503), .B2(new_n349), .ZN(new_n504));
  AND2_X1   g0304(.A1(new_n504), .A2(KEYINPUT86), .ZN(new_n505));
  OAI21_X1  g0305(.A(G200), .B1(new_n504), .B2(KEYINPUT86), .ZN(new_n506));
  OR2_X1    g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT6), .ZN(new_n508));
  AND2_X1   g0308(.A1(G97), .A2(G107), .ZN(new_n509));
  NOR2_X1   g0309(.A1(G97), .A2(G107), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(G107), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n512), .A2(KEYINPUT6), .A3(G97), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n210), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n367), .A2(new_n214), .ZN(new_n515));
  OAI21_X1  g0315(.A(KEYINPUT84), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT84), .ZN(new_n517));
  INV_X1    g0317(.A(new_n515), .ZN(new_n518));
  AND3_X1   g0318(.A1(new_n512), .A2(KEYINPUT6), .A3(G97), .ZN(new_n519));
  XNOR2_X1  g0319(.A(G97), .B(G107), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n519), .B1(new_n520), .B2(new_n508), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n517), .B(new_n518), .C1(new_n521), .C2(new_n210), .ZN(new_n522));
  INV_X1    g0322(.A(new_n282), .ZN(new_n523));
  OAI21_X1  g0323(.A(G107), .B1(new_n272), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n516), .A2(new_n522), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n257), .ZN(new_n526));
  AOI21_X1  g0326(.A(G97), .B1(new_n251), .B2(new_n252), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n248), .A2(G33), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n253), .A2(new_n360), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n527), .B1(new_n529), .B2(G97), .ZN(new_n530));
  INV_X1    g0330(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n526), .A2(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n532), .B1(G190), .B2(new_n504), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n496), .A2(new_n498), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n297), .A2(G244), .A3(new_n500), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT85), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n502), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n349), .B1(new_n534), .B2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(new_n493), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n538), .A2(new_n319), .A3(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT88), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n504), .A2(KEYINPUT88), .A3(new_n319), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n538), .A2(new_n539), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(new_n289), .ZN(new_n545));
  AND3_X1   g0345(.A1(new_n542), .A2(new_n543), .A3(new_n545), .ZN(new_n546));
  AOI21_X1  g0346(.A(KEYINPUT87), .B1(new_n526), .B2(new_n531), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT87), .ZN(new_n548));
  AOI211_X1 g0348(.A(new_n548), .B(new_n530), .C1(new_n525), .C2(new_n257), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  AOI22_X1  g0350(.A1(new_n507), .A2(new_n533), .B1(new_n546), .B2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT24), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n297), .A2(new_n210), .A3(G87), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(KEYINPUT22), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT22), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n297), .A2(new_n555), .A3(new_n210), .A4(G87), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT23), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n558), .B1(new_n210), .B2(G107), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n512), .A2(KEYINPUT23), .A3(G20), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(G116), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n275), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(new_n210), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(new_n565), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n552), .B1(new_n557), .B2(new_n566), .ZN(new_n567));
  AOI211_X1 g0367(.A(KEYINPUT24), .B(new_n565), .C1(new_n554), .C2(new_n556), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n257), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n529), .A2(new_n512), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT25), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n571), .B1(new_n255), .B2(new_n512), .ZN(new_n572));
  NOR3_X1   g0372(.A1(new_n253), .A2(KEYINPUT25), .A3(G107), .ZN(new_n573));
  NOR3_X1   g0373(.A1(new_n570), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  AND2_X1   g0374(.A1(new_n569), .A2(new_n574), .ZN(new_n575));
  OAI211_X1 g0375(.A(G257), .B(G1698), .C1(new_n269), .C2(new_n270), .ZN(new_n576));
  NAND2_X1  g0376(.A1(G33), .A2(G294), .ZN(new_n577));
  OAI21_X1  g0377(.A(G250), .B1(new_n269), .B2(new_n270), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n576), .B(new_n577), .C1(new_n578), .C2(G1698), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n349), .ZN(new_n580));
  OAI211_X1 g0380(.A(G264), .B(new_n291), .C1(new_n488), .C2(new_n489), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n580), .A2(new_n491), .A3(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(G190), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n584), .B1(G200), .B2(new_n582), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n575), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n569), .A2(new_n574), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n582), .A2(G169), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT91), .ZN(new_n589));
  INV_X1    g0389(.A(new_n581), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n590), .B1(new_n349), .B2(new_n579), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n591), .A2(G179), .A3(new_n491), .ZN(new_n592));
  AND3_X1   g0392(.A1(new_n588), .A2(new_n589), .A3(new_n592), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n589), .B1(new_n588), .B2(new_n592), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n587), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  AND2_X1   g0395(.A1(new_n586), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n255), .A2(new_n562), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n253), .A2(G116), .A3(new_n360), .A4(new_n528), .ZN(new_n598));
  AOI22_X1  g0398(.A1(new_n256), .A2(new_n209), .B1(G20), .B2(new_n562), .ZN(new_n599));
  AOI21_X1  g0399(.A(G20), .B1(G33), .B2(G283), .ZN(new_n600));
  INV_X1    g0400(.A(G97), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n600), .B1(G33), .B2(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(KEYINPUT20), .B1(new_n599), .B2(new_n602), .ZN(new_n603));
  AND3_X1   g0403(.A1(new_n599), .A2(new_n602), .A3(KEYINPUT20), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n597), .B(new_n598), .C1(new_n603), .C2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(G303), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n291), .B1(new_n271), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n500), .A2(G257), .ZN(new_n608));
  NAND2_X1  g0408(.A1(G264), .A2(G1698), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n297), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  OAI211_X1 g0411(.A(G270), .B(new_n291), .C1(new_n488), .C2(new_n489), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n611), .A2(new_n491), .A3(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n605), .A2(G169), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(KEYINPUT21), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT21), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n605), .A2(new_n616), .A3(G169), .A4(new_n613), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n613), .A2(new_n319), .ZN(new_n618));
  AOI22_X1  g0418(.A1(new_n615), .A2(new_n617), .B1(new_n605), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n215), .A2(G1698), .ZN(new_n620));
  OAI221_X1 g0420(.A(new_n620), .B1(G238), .B2(G1698), .C1(new_n269), .C2(new_n270), .ZN(new_n621));
  INV_X1    g0421(.A(new_n563), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n291), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(G45), .ZN(new_n624));
  OR3_X1    g0424(.A1(new_n624), .A2(G1), .A3(G274), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n217), .B1(new_n624), .B2(G1), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n625), .A2(new_n291), .A3(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  OAI21_X1  g0428(.A(G200), .B1(new_n623), .B2(new_n628), .ZN(new_n629));
  NOR2_X1   g0429(.A1(G238), .A2(G1698), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n630), .B1(new_n215), .B2(G1698), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n563), .B1(new_n631), .B2(new_n297), .ZN(new_n632));
  OAI211_X1 g0432(.A(G190), .B(new_n627), .C1(new_n632), .C2(new_n291), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n629), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n210), .A2(G33), .A3(G97), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT19), .ZN(new_n636));
  AND3_X1   g0436(.A1(new_n635), .A2(KEYINPUT89), .A3(new_n636), .ZN(new_n637));
  AOI21_X1  g0437(.A(KEYINPUT89), .B1(new_n635), .B2(new_n636), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n210), .B1(new_n442), .B2(new_n636), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n216), .A2(new_n601), .A3(new_n512), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  OAI211_X1 g0442(.A(new_n210), .B(G68), .C1(new_n269), .C2(new_n270), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n257), .B1(new_n639), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n255), .A2(new_n361), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n253), .A2(G87), .A3(new_n360), .A4(new_n528), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n645), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n634), .A2(new_n648), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n253), .A2(new_n360), .A3(new_n362), .A4(new_n528), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n645), .A2(new_n646), .A3(new_n650), .ZN(new_n651));
  OR2_X1    g0451(.A1(new_n651), .A2(KEYINPUT90), .ZN(new_n652));
  OAI21_X1  g0452(.A(G169), .B1(new_n623), .B2(new_n628), .ZN(new_n653));
  OAI211_X1 g0453(.A(G179), .B(new_n627), .C1(new_n632), .C2(new_n291), .ZN(new_n654));
  AOI22_X1  g0454(.A1(new_n651), .A2(KEYINPUT90), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n649), .B1(new_n652), .B2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n605), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n613), .A2(G200), .ZN(new_n658));
  OAI211_X1 g0458(.A(new_n657), .B(new_n658), .C1(new_n583), .C2(new_n613), .ZN(new_n659));
  AND3_X1   g0459(.A1(new_n619), .A2(new_n656), .A3(new_n659), .ZN(new_n660));
  AND4_X1   g0460(.A1(new_n486), .A2(new_n551), .A3(new_n596), .A4(new_n660), .ZN(G372));
  INV_X1    g0461(.A(new_n400), .ZN(new_n662));
  INV_X1    g0462(.A(new_n371), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n470), .A2(new_n663), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n664), .B1(new_n484), .B2(new_n469), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n341), .A2(new_n344), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  AND2_X1   g0467(.A1(new_n326), .A2(new_n332), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  AND3_X1   g0469(.A1(new_n419), .A2(new_n423), .A3(KEYINPUT94), .ZN(new_n670));
  AOI21_X1  g0470(.A(KEYINPUT94), .B1(new_n419), .B2(new_n423), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n662), .B1(new_n669), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n653), .A2(new_n654), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(new_n651), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n676), .B1(new_n648), .B2(new_n634), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n677), .B1(new_n575), .B2(new_n585), .ZN(new_n678));
  INV_X1    g0478(.A(new_n619), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n575), .B1(new_n588), .B2(new_n592), .ZN(new_n680));
  OAI211_X1 g0480(.A(new_n551), .B(new_n678), .C1(new_n679), .C2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT93), .ZN(new_n682));
  XOR2_X1   g0482(.A(KEYINPUT92), .B(KEYINPUT26), .Z(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n546), .A2(new_n550), .A3(new_n656), .A4(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT26), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n542), .A2(new_n532), .A3(new_n545), .A4(new_n543), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n686), .B1(new_n687), .B2(new_n677), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n682), .B1(new_n689), .B2(new_n676), .ZN(new_n690));
  INV_X1    g0490(.A(new_n676), .ZN(new_n691));
  AOI211_X1 g0491(.A(KEYINPUT93), .B(new_n691), .C1(new_n685), .C2(new_n688), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n681), .B1(new_n690), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n486), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n674), .A2(new_n694), .ZN(new_n695));
  XOR2_X1   g0495(.A(new_n695), .B(KEYINPUT95), .Z(G369));
  NAND3_X1  g0496(.A1(new_n248), .A2(new_n210), .A3(G13), .ZN(new_n697));
  OR2_X1    g0497(.A1(new_n697), .A2(KEYINPUT27), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(KEYINPUT27), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n698), .A2(G213), .A3(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(G343), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n679), .A2(new_n605), .A3(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n702), .ZN(new_n704));
  OAI211_X1 g0504(.A(new_n619), .B(new_n659), .C1(new_n657), .C2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(G330), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n596), .B1(new_n575), .B2(new_n704), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n710), .B1(new_n595), .B2(new_n704), .ZN(new_n711));
  AND2_X1   g0511(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n619), .A2(new_n702), .ZN(new_n714));
  AOI22_X1  g0514(.A1(new_n596), .A2(new_n714), .B1(new_n680), .B2(new_n704), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n713), .A2(new_n715), .ZN(G399));
  INV_X1    g0516(.A(new_n204), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n717), .A2(G41), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n641), .A2(G116), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n719), .A2(G1), .A3(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n721), .B1(new_n207), .B2(new_n719), .ZN(new_n722));
  XNOR2_X1  g0522(.A(new_n722), .B(KEYINPUT96), .ZN(new_n723));
  XNOR2_X1  g0523(.A(new_n723), .B(KEYINPUT28), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n551), .A2(new_n596), .A3(new_n660), .A4(new_n704), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT30), .ZN(new_n726));
  AND3_X1   g0526(.A1(new_n611), .A2(new_n491), .A3(new_n612), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n623), .A2(new_n628), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n727), .A2(G179), .A3(new_n591), .A4(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n726), .B1(new_n729), .B2(new_n544), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n613), .A2(new_n654), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n504), .A2(new_n731), .A3(KEYINPUT30), .A4(new_n591), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n728), .A2(G179), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n544), .A2(new_n582), .A3(new_n613), .A4(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n730), .A2(new_n732), .A3(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(KEYINPUT31), .B1(new_n735), .B2(new_n702), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n730), .A2(new_n734), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(KEYINPUT97), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT97), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n730), .A2(new_n739), .A3(new_n734), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n738), .A2(new_n732), .A3(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT31), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n704), .A2(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n736), .B1(new_n741), .B2(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n708), .B1(new_n725), .B2(new_n744), .ZN(new_n745));
  AOI21_X1  g0545(.A(KEYINPUT29), .B1(new_n693), .B2(new_n704), .ZN(new_n746));
  XNOR2_X1  g0546(.A(new_n746), .B(KEYINPUT98), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n649), .B1(new_n575), .B2(new_n585), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT100), .ZN(new_n749));
  AND3_X1   g0549(.A1(new_n595), .A2(new_n749), .A3(new_n619), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n749), .B1(new_n595), .B2(new_n619), .ZN(new_n751));
  OAI211_X1 g0551(.A(new_n551), .B(new_n748), .C1(new_n750), .C2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n547), .ZN(new_n753));
  AOI22_X1  g0553(.A1(new_n540), .A2(new_n541), .B1(new_n544), .B2(new_n289), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n530), .B1(new_n525), .B2(new_n257), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(KEYINPUT87), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n753), .A2(new_n754), .A3(new_n543), .A4(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n656), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n683), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(KEYINPUT99), .ZN(new_n760));
  INV_X1    g0560(.A(new_n634), .ZN(new_n761));
  INV_X1    g0561(.A(new_n648), .ZN(new_n762));
  AOI22_X1  g0562(.A1(new_n761), .A2(new_n762), .B1(new_n675), .B2(new_n651), .ZN(new_n763));
  NAND4_X1  g0563(.A1(new_n754), .A2(new_n763), .A3(new_n543), .A4(new_n532), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n760), .B1(new_n764), .B2(new_n686), .ZN(new_n765));
  INV_X1    g0565(.A(new_n687), .ZN(new_n766));
  NAND4_X1  g0566(.A1(new_n766), .A2(KEYINPUT99), .A3(KEYINPUT26), .A4(new_n763), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n759), .A2(new_n765), .A3(new_n767), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n752), .A2(new_n676), .A3(new_n768), .ZN(new_n769));
  AND2_X1   g0569(.A1(new_n769), .A2(new_n704), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(KEYINPUT29), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n745), .B1(new_n747), .B2(new_n771), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n724), .B1(new_n772), .B2(G1), .ZN(G364));
  AND2_X1   g0573(.A1(new_n210), .A2(G13), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G45), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n719), .A2(G1), .A3(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(G13), .A2(G33), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(G20), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n707), .A2(new_n779), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n209), .B1(G20), .B2(new_n289), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  XOR2_X1   g0582(.A(new_n782), .B(KEYINPUT102), .Z(new_n783));
  NOR2_X1   g0583(.A1(new_n239), .A2(new_n624), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n717), .A2(new_n297), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n785), .B1(G45), .B2(new_n207), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n784), .B1(KEYINPUT101), .B2(new_n786), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n787), .B1(KEYINPUT101), .B2(new_n786), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n717), .A2(new_n271), .ZN(new_n789));
  AOI22_X1  g0589(.A1(new_n789), .A2(G355), .B1(new_n562), .B2(new_n717), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n783), .B1(new_n788), .B2(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n210), .A2(G190), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n319), .A2(G200), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n373), .A2(G179), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n792), .A2(new_n795), .ZN(new_n796));
  OAI22_X1  g0596(.A1(new_n214), .A2(new_n794), .B1(new_n796), .B2(new_n512), .ZN(new_n797));
  NOR2_X1   g0597(.A1(G179), .A2(G200), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n210), .B1(new_n798), .B2(G190), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n210), .A2(new_n583), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(new_n793), .ZN(new_n801));
  OAI221_X1 g0601(.A(new_n297), .B1(new_n799), .B2(new_n601), .C1(new_n244), .C2(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n800), .A2(new_n795), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  AOI211_X1 g0604(.A(new_n797), .B(new_n802), .C1(G87), .C2(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n792), .A2(new_n798), .ZN(new_n806));
  INV_X1    g0606(.A(G159), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  XNOR2_X1  g0608(.A(new_n808), .B(KEYINPUT32), .ZN(new_n809));
  NAND3_X1  g0609(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n810));
  XNOR2_X1  g0610(.A(new_n810), .B(KEYINPUT103), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n811), .A2(new_n583), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n811), .A2(G190), .ZN(new_n813));
  AOI22_X1  g0613(.A1(G50), .A2(new_n812), .B1(new_n813), .B2(G68), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n805), .A2(new_n809), .A3(new_n814), .ZN(new_n815));
  OR2_X1    g0615(.A1(new_n815), .A2(KEYINPUT104), .ZN(new_n816));
  XNOR2_X1  g0616(.A(KEYINPUT33), .B(G317), .ZN(new_n817));
  AOI22_X1  g0617(.A1(G326), .A2(new_n812), .B1(new_n813), .B2(new_n817), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n806), .B(KEYINPUT105), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n819), .A2(G329), .ZN(new_n820));
  INV_X1    g0620(.A(G283), .ZN(new_n821));
  OAI22_X1  g0621(.A1(new_n803), .A2(new_n606), .B1(new_n796), .B2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n794), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n822), .B1(G311), .B2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(G322), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n271), .B1(new_n801), .B2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n799), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n826), .B1(G294), .B2(new_n827), .ZN(new_n828));
  NAND4_X1  g0628(.A1(new_n818), .A2(new_n820), .A3(new_n824), .A4(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n815), .A2(KEYINPUT104), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n816), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n791), .B1(new_n831), .B2(new_n781), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n776), .B1(new_n780), .B2(new_n832), .ZN(new_n833));
  XNOR2_X1  g0633(.A(new_n706), .B(G330), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n833), .B1(new_n834), .B2(new_n776), .ZN(new_n835));
  XNOR2_X1  g0635(.A(new_n835), .B(KEYINPUT106), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(G396));
  NAND2_X1  g0637(.A1(new_n693), .A2(new_n704), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n370), .A2(new_n702), .ZN(new_n839));
  OR2_X1    g0639(.A1(new_n371), .A2(new_n839), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n371), .A2(new_n375), .A3(new_n839), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n838), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n693), .A2(new_n704), .A3(new_n842), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n745), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n844), .A2(new_n745), .A3(new_n845), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n847), .A2(new_n776), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n846), .B1(new_n848), .B2(KEYINPUT109), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n849), .B1(KEYINPUT109), .B2(new_n848), .ZN(new_n850));
  INV_X1    g0650(.A(new_n781), .ZN(new_n851));
  INV_X1    g0651(.A(new_n801), .ZN(new_n852));
  AOI22_X1  g0652(.A1(G143), .A2(new_n852), .B1(new_n823), .B2(G159), .ZN(new_n853));
  INV_X1    g0653(.A(new_n813), .ZN(new_n854));
  INV_X1    g0654(.A(G150), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n853), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n856), .B1(G137), .B2(new_n812), .ZN(new_n857));
  XOR2_X1   g0657(.A(new_n857), .B(KEYINPUT34), .Z(new_n858));
  INV_X1    g0658(.A(G50), .ZN(new_n859));
  OAI221_X1 g0659(.A(new_n297), .B1(new_n796), .B2(new_n262), .C1(new_n859), .C2(new_n803), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n860), .B1(G58), .B2(new_n827), .ZN(new_n861));
  INV_X1    g0661(.A(G132), .ZN(new_n862));
  INV_X1    g0662(.A(new_n819), .ZN(new_n863));
  OAI211_X1 g0663(.A(new_n858), .B(new_n861), .C1(new_n862), .C2(new_n863), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n271), .B1(new_n803), .B2(new_n512), .ZN(new_n865));
  OAI22_X1  g0665(.A1(new_n216), .A2(new_n796), .B1(new_n794), .B2(new_n562), .ZN(new_n866));
  AOI211_X1 g0666(.A(new_n865), .B(new_n866), .C1(new_n819), .C2(G311), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n813), .A2(G283), .ZN(new_n868));
  INV_X1    g0668(.A(G294), .ZN(new_n869));
  OAI22_X1  g0669(.A1(new_n801), .A2(new_n869), .B1(new_n799), .B2(new_n601), .ZN(new_n870));
  OR2_X1    g0670(.A1(new_n870), .A2(KEYINPUT108), .ZN(new_n871));
  AOI22_X1  g0671(.A1(new_n812), .A2(G303), .B1(new_n870), .B2(KEYINPUT108), .ZN(new_n872));
  NAND4_X1  g0672(.A1(new_n867), .A2(new_n868), .A3(new_n871), .A4(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n851), .B1(new_n864), .B2(new_n873), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n781), .A2(new_n777), .ZN(new_n875));
  XOR2_X1   g0675(.A(new_n875), .B(KEYINPUT107), .Z(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(new_n877));
  AOI211_X1 g0677(.A(new_n776), .B(new_n874), .C1(new_n214), .C2(new_n877), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n878), .B1(new_n842), .B2(new_n778), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n850), .A2(new_n879), .ZN(G384));
  INV_X1    g0680(.A(new_n521), .ZN(new_n881));
  OR2_X1    g0681(.A1(new_n881), .A2(KEYINPUT35), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(KEYINPUT35), .ZN(new_n883));
  NAND4_X1  g0683(.A1(new_n882), .A2(new_n883), .A3(G116), .A4(new_n211), .ZN(new_n884));
  XOR2_X1   g0684(.A(new_n884), .B(KEYINPUT36), .Z(new_n885));
  OAI211_X1 g0685(.A(new_n208), .B(G77), .C1(new_n244), .C2(new_n262), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n859), .A2(G68), .ZN(new_n887));
  AOI211_X1 g0687(.A(new_n248), .B(G13), .C1(new_n886), .C2(new_n887), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n885), .A2(new_n888), .ZN(new_n889));
  AND3_X1   g0689(.A1(new_n735), .A2(KEYINPUT31), .A3(new_n702), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n890), .A2(new_n736), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n725), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(new_n842), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n466), .A2(new_n468), .A3(new_n702), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  AND2_X1   g0695(.A1(new_n472), .A2(new_n473), .ZN(new_n896));
  AND2_X1   g0696(.A1(new_n476), .A2(new_n477), .ZN(new_n897));
  AND3_X1   g0697(.A1(new_n482), .A2(KEYINPUT79), .A3(KEYINPUT14), .ZN(new_n898));
  AOI21_X1  g0698(.A(KEYINPUT79), .B1(new_n482), .B2(KEYINPUT14), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n897), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n895), .B1(new_n896), .B2(new_n900), .ZN(new_n901));
  XNOR2_X1  g0701(.A(new_n894), .B(KEYINPUT110), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n470), .B(new_n902), .C1(new_n484), .C2(new_n469), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n893), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT38), .ZN(new_n905));
  INV_X1    g0705(.A(new_n700), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n288), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n339), .A2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT113), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n325), .A2(new_n909), .ZN(new_n910));
  OAI211_X1 g0710(.A(KEYINPUT113), .B(new_n288), .C1(new_n323), .C2(new_n324), .ZN(new_n911));
  AOI211_X1 g0711(.A(KEYINPUT37), .B(new_n908), .C1(new_n910), .C2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT112), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT111), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n278), .A2(KEYINPUT80), .A3(new_n279), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n283), .A2(G68), .A3(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(new_n268), .ZN(new_n917));
  AOI21_X1  g0717(.A(KEYINPUT16), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n914), .B1(new_n918), .B2(new_n360), .ZN(new_n919));
  OAI211_X1 g0719(.A(KEYINPUT111), .B(new_n257), .C1(new_n334), .C2(KEYINPUT16), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n919), .A2(new_n335), .A3(new_n920), .ZN(new_n921));
  AOI22_X1  g0721(.A1(new_n921), .A2(new_n260), .B1(new_n328), .B2(new_n329), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n913), .B1(new_n922), .B2(new_n343), .ZN(new_n923));
  INV_X1    g0723(.A(new_n260), .ZN(new_n924));
  AND3_X1   g0724(.A1(new_n280), .A2(new_n281), .A3(new_n282), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n915), .A2(G68), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n917), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n360), .B1(new_n927), .B2(new_n261), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n284), .B1(new_n928), .B2(KEYINPUT111), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n924), .B1(new_n929), .B2(new_n919), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n323), .A2(new_n324), .ZN(new_n931));
  OAI211_X1 g0731(.A(KEYINPUT112), .B(new_n339), .C1(new_n930), .C2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n920), .A2(new_n335), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n927), .A2(new_n261), .ZN(new_n934));
  AOI21_X1  g0734(.A(KEYINPUT111), .B1(new_n934), .B2(new_n257), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n260), .B1(new_n933), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(new_n906), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n923), .A2(new_n932), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n912), .B1(new_n938), .B2(KEYINPUT37), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n937), .B1(new_n668), .B2(new_n666), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n905), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n930), .A2(new_n700), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n345), .A2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT37), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n339), .B1(new_n930), .B2(new_n931), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n942), .B1(new_n945), .B2(new_n913), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n944), .B1(new_n946), .B2(new_n932), .ZN(new_n947));
  OAI211_X1 g0747(.A(KEYINPUT38), .B(new_n943), .C1(new_n947), .C2(new_n912), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n941), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n904), .A2(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT40), .ZN(new_n951));
  AND2_X1   g0751(.A1(new_n892), .A2(new_n842), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n894), .B1(new_n474), .B2(new_n484), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n902), .A2(new_n470), .ZN(new_n954));
  INV_X1    g0754(.A(new_n469), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n954), .B1(new_n900), .B2(new_n955), .ZN(new_n956));
  OAI211_X1 g0756(.A(new_n952), .B(KEYINPUT40), .C1(new_n953), .C2(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n910), .A2(new_n911), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n908), .A2(KEYINPUT37), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n325), .A2(new_n339), .A3(new_n907), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(KEYINPUT37), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n345), .A2(new_n288), .A3(new_n906), .ZN(new_n965));
  AOI21_X1  g0765(.A(KEYINPUT38), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n948), .A2(new_n967), .ZN(new_n968));
  AOI22_X1  g0768(.A1(new_n950), .A2(new_n951), .B1(new_n958), .B2(new_n968), .ZN(new_n969));
  AND3_X1   g0769(.A1(new_n969), .A2(new_n486), .A3(new_n892), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n969), .B1(new_n486), .B2(new_n892), .ZN(new_n971));
  OR3_X1    g0771(.A1(new_n970), .A2(new_n971), .A3(new_n708), .ZN(new_n972));
  NOR3_X1   g0772(.A1(new_n484), .A2(new_n469), .A3(new_n702), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n949), .A2(KEYINPUT39), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n343), .B1(new_n936), .B2(new_n330), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n937), .B1(new_n976), .B2(KEYINPUT112), .ZN(new_n977));
  INV_X1    g0777(.A(new_n932), .ZN(new_n978));
  OAI21_X1  g0778(.A(KEYINPUT37), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n940), .B1(new_n979), .B2(new_n961), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n966), .B1(new_n980), .B2(KEYINPUT38), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT39), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n974), .B1(new_n975), .B2(new_n983), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n371), .A2(new_n702), .ZN(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n845), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n901), .A2(new_n903), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n987), .A2(new_n949), .A3(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(new_n668), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(new_n700), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n984), .A2(new_n992), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n990), .B1(new_n665), .B2(new_n666), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n400), .B1(new_n994), .B2(new_n672), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n485), .B1(KEYINPUT29), .B2(new_n770), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n995), .B1(new_n747), .B2(new_n996), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n993), .B(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n972), .A2(new_n998), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n999), .B1(new_n248), .B2(new_n774), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n972), .A2(new_n998), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n889), .B1(new_n1000), .B2(new_n1001), .ZN(G367));
  INV_X1    g0802(.A(new_n776), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n783), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1004), .B1(new_n204), .B2(new_n361), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n785), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n232), .A2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1003), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1008));
  OAI22_X1  g0808(.A1(new_n801), .A2(new_n855), .B1(new_n794), .B2(new_n859), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(KEYINPUT117), .B(G137), .ZN(new_n1010));
  OAI22_X1  g0810(.A1(new_n803), .A2(new_n244), .B1(new_n806), .B2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n297), .B1(new_n796), .B2(new_n214), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n799), .A2(new_n262), .ZN(new_n1013));
  NOR4_X1   g0813(.A1(new_n1009), .A2(new_n1011), .A3(new_n1012), .A4(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n812), .A2(G143), .ZN(new_n1015));
  OAI211_X1 g0815(.A(new_n1014), .B(new_n1015), .C1(new_n807), .C2(new_n854), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n804), .A2(G116), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1017), .B(KEYINPUT46), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n794), .A2(new_n821), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n796), .A2(new_n601), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n806), .ZN(new_n1021));
  AOI211_X1 g0821(.A(new_n1019), .B(new_n1020), .C1(G317), .C2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n271), .B1(new_n801), .B2(new_n606), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1023), .B1(G107), .B2(new_n827), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1018), .A2(new_n1022), .A3(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n812), .ZN(new_n1026));
  INV_X1    g0826(.A(G311), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n869), .A2(new_n854), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1016), .B1(new_n1025), .B2(new_n1028), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT47), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1008), .B1(new_n1030), .B2(new_n781), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n762), .A2(new_n704), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1032), .A2(new_n691), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n677), .B2(new_n1032), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n779), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1031), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n551), .B1(new_n755), .B2(new_n704), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n766), .A2(new_n702), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n596), .A2(new_n714), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT42), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n757), .B1(new_n1040), .B2(new_n595), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1044), .A2(new_n704), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT114), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1034), .A2(KEYINPUT43), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1046), .A2(new_n1047), .A3(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1047), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n1050), .A2(new_n1051), .B1(KEYINPUT43), .B2(new_n1034), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n1051), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n1034), .A2(KEYINPUT43), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1053), .A2(new_n1054), .A3(new_n1049), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1052), .A2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1056), .B1(new_n713), .B2(new_n1040), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n713), .A2(new_n1040), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1052), .A2(new_n1055), .A3(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1059), .A2(KEYINPUT115), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT115), .ZN(new_n1061));
  NAND4_X1  g0861(.A1(new_n1052), .A2(new_n1055), .A3(new_n1061), .A4(new_n1058), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1057), .A2(new_n1060), .A3(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n775), .A2(G1), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1039), .A2(new_n715), .ZN(new_n1065));
  XOR2_X1   g0865(.A(new_n1065), .B(KEYINPUT45), .Z(new_n1066));
  NOR2_X1   g0866(.A1(new_n1039), .A2(new_n715), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1067), .B(KEYINPUT44), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n712), .A2(KEYINPUT116), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1066), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n712), .A2(KEYINPUT116), .ZN(new_n1071));
  XOR2_X1   g0871(.A(new_n1070), .B(new_n1071), .Z(new_n1072));
  OAI21_X1  g0872(.A(new_n1041), .B1(new_n711), .B2(new_n714), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n709), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n1073), .B(new_n1074), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n772), .B1(new_n1072), .B2(new_n1075), .ZN(new_n1076));
  XOR2_X1   g0876(.A(new_n718), .B(KEYINPUT41), .Z(new_n1077));
  INV_X1    g0877(.A(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1064), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1036), .B1(new_n1063), .B2(new_n1079), .ZN(G387));
  INV_X1    g0880(.A(new_n1075), .ZN(new_n1081));
  OR2_X1    g0881(.A1(new_n711), .A2(new_n1035), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n720), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n789), .A2(new_n1083), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1084), .B1(G107), .B2(new_n204), .ZN(new_n1085));
  OR2_X1    g0885(.A1(new_n229), .A2(new_n624), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n246), .A2(G50), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(new_n1087), .B(KEYINPUT50), .ZN(new_n1088));
  AOI211_X1 g0888(.A(G45), .B(new_n1083), .C1(G68), .C2(G77), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1006), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1085), .B1(new_n1086), .B2(new_n1090), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1003), .B1(new_n1091), .B2(new_n783), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n803), .A2(new_n214), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(KEYINPUT118), .B(G150), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1093), .B1(new_n1021), .B2(new_n1094), .ZN(new_n1095));
  OAI221_X1 g0895(.A(new_n1095), .B1(new_n859), .B2(new_n801), .C1(new_n262), .C2(new_n794), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n799), .A2(new_n361), .ZN(new_n1097));
  NOR4_X1   g0897(.A1(new_n1096), .A2(new_n271), .A3(new_n1020), .A4(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n812), .A2(G159), .ZN(new_n1099));
  XOR2_X1   g0899(.A(new_n1099), .B(KEYINPUT119), .Z(new_n1100));
  NAND2_X1  g0900(.A1(new_n813), .A2(new_n247), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1098), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n803), .A2(new_n869), .B1(new_n799), .B2(new_n821), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(G317), .A2(new_n852), .B1(new_n823), .B2(G303), .ZN(new_n1104));
  OAI221_X1 g0904(.A(new_n1104), .B1(new_n854), .B2(new_n1027), .C1(new_n825), .C2(new_n1026), .ZN(new_n1105));
  INV_X1    g0905(.A(KEYINPUT48), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1103), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1107), .B1(new_n1106), .B2(new_n1105), .ZN(new_n1108));
  XOR2_X1   g0908(.A(new_n1108), .B(KEYINPUT49), .Z(new_n1109));
  AOI21_X1  g0909(.A(new_n297), .B1(new_n1021), .B2(G326), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1110), .B1(new_n562), .B2(new_n796), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1102), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1092), .B1(new_n1112), .B2(new_n781), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n1081), .A2(new_n1064), .B1(new_n1082), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n772), .A2(new_n1081), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1115), .A2(new_n718), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n772), .A2(new_n1081), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1114), .B1(new_n1116), .B2(new_n1117), .ZN(G393));
  INV_X1    g0918(.A(new_n1064), .ZN(new_n1119));
  OR2_X1    g0919(.A1(new_n1072), .A2(new_n1119), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n1039), .A2(new_n1035), .ZN(new_n1121));
  XNOR2_X1  g0921(.A(new_n1121), .B(KEYINPUT120), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n783), .B1(G97), .B2(new_n717), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n236), .A2(new_n785), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n776), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n812), .A2(G317), .B1(G311), .B2(new_n852), .ZN(new_n1126));
  XOR2_X1   g0926(.A(new_n1126), .B(KEYINPUT52), .Z(new_n1127));
  OAI221_X1 g0927(.A(new_n271), .B1(new_n799), .B2(new_n562), .C1(new_n512), .C2(new_n796), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(G283), .A2(new_n804), .B1(new_n1021), .B2(G322), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1129), .B1(new_n869), .B2(new_n794), .ZN(new_n1130));
  AOI211_X1 g0930(.A(new_n1128), .B(new_n1130), .C1(G303), .C2(new_n813), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n812), .A2(G150), .B1(G159), .B2(new_n852), .ZN(new_n1132));
  XOR2_X1   g0932(.A(new_n1132), .B(KEYINPUT51), .Z(new_n1133));
  OAI221_X1 g0933(.A(new_n297), .B1(new_n799), .B2(new_n214), .C1(new_n216), .C2(new_n796), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(G68), .A2(new_n804), .B1(new_n1021), .B2(G143), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1135), .B1(new_n246), .B2(new_n794), .ZN(new_n1136));
  AOI211_X1 g0936(.A(new_n1134), .B(new_n1136), .C1(G50), .C2(new_n813), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(new_n1127), .A2(new_n1131), .B1(new_n1133), .B2(new_n1137), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n1122), .B(new_n1125), .C1(new_n851), .C2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1120), .A2(new_n1139), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n1072), .A2(new_n1115), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n1141), .A2(new_n719), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1072), .A2(new_n1115), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1140), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(G390));
  INV_X1    g0945(.A(KEYINPUT122), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n708), .B1(new_n725), .B2(new_n891), .ZN(new_n1147));
  INV_X1    g0947(.A(KEYINPUT121), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n842), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  AOI211_X1 g0949(.A(KEYINPUT121), .B(new_n708), .C1(new_n725), .C2(new_n891), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  OR2_X1    g0951(.A1(new_n1151), .A2(new_n988), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n769), .A2(new_n704), .A3(new_n842), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(new_n986), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n745), .A2(new_n842), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1154), .B1(new_n988), .B2(new_n1156), .ZN(new_n1157));
  OAI211_X1 g0957(.A(new_n952), .B(G330), .C1(new_n953), .C2(new_n956), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n901), .A2(new_n903), .A3(new_n1155), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n1152), .A2(new_n1157), .B1(new_n987), .B2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(KEYINPUT29), .ZN(new_n1162));
  AOI21_X1  g0962(.A(KEYINPUT98), .B1(new_n838), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(KEYINPUT98), .ZN(new_n1164));
  AOI211_X1 g0964(.A(new_n1164), .B(KEYINPUT29), .C1(new_n693), .C2(new_n704), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n996), .B1(new_n1163), .B2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n486), .A2(new_n1147), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1166), .A2(new_n674), .A3(new_n1167), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1146), .B1(new_n1161), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1160), .A2(new_n987), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1156), .B1(new_n953), .B2(new_n956), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1154), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n1171), .B(new_n1172), .C1(new_n1151), .C2(new_n988), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1170), .A2(new_n1173), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n997), .A2(new_n1174), .A3(KEYINPUT122), .A4(new_n1167), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1169), .A2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n988), .A2(new_n1154), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1177), .A2(new_n974), .A3(new_n968), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n975), .A2(new_n983), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n973), .B1(new_n987), .B2(new_n988), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1171), .B(new_n1178), .C1(new_n1179), .C2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(new_n845), .A2(new_n986), .B1(new_n901), .B2(new_n903), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n975), .B(new_n983), .C1(new_n1183), .C2(new_n973), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1158), .B1(new_n1184), .B2(new_n1178), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n1182), .A2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1176), .A2(new_n1186), .ZN(new_n1187));
  NOR3_X1   g0987(.A1(new_n939), .A2(new_n905), .A3(new_n940), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n974), .B1(new_n1188), .B2(new_n966), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(new_n901), .A2(new_n903), .B1(new_n1153), .B2(new_n986), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  AND3_X1   g0991(.A1(new_n948), .A2(new_n967), .A3(new_n982), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n982), .B1(new_n941), .B2(new_n948), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n987), .A2(new_n988), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1195), .A2(new_n974), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1191), .B1(new_n1194), .B2(new_n1196), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1181), .B1(new_n1197), .B2(new_n1158), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1198), .A2(new_n1169), .A3(new_n1175), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1187), .A2(new_n718), .A3(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1194), .A2(new_n777), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1003), .B1(new_n876), .B2(new_n247), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(G107), .A2(new_n813), .B1(new_n812), .B2(G283), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n819), .A2(G294), .ZN(new_n1204));
  OAI22_X1  g1004(.A1(new_n801), .A2(new_n562), .B1(new_n796), .B2(new_n262), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1205), .B1(G97), .B2(new_n823), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n271), .B1(new_n803), .B2(new_n216), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1207), .B1(G77), .B2(new_n827), .ZN(new_n1208));
  NAND4_X1  g1008(.A1(new_n1203), .A2(new_n1204), .A3(new_n1206), .A4(new_n1208), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n801), .A2(new_n862), .B1(new_n796), .B2(new_n859), .ZN(new_n1210));
  XOR2_X1   g1010(.A(KEYINPUT54), .B(G143), .Z(new_n1211));
  AOI211_X1 g1011(.A(new_n271), .B(new_n1210), .C1(new_n823), .C2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n804), .A2(new_n1094), .ZN(new_n1213));
  OR2_X1    g1013(.A1(new_n1213), .A2(KEYINPUT53), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n1213), .A2(KEYINPUT53), .B1(G159), .B2(new_n827), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n819), .A2(G125), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1212), .A2(new_n1214), .A3(new_n1215), .A4(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n812), .A2(G128), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1218), .B1(new_n854), .B2(new_n1010), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1209), .B1(new_n1217), .B2(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1202), .B1(new_n1220), .B2(new_n781), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n1186), .A2(new_n1064), .B1(new_n1201), .B2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1200), .A2(new_n1222), .ZN(G378));
  INV_X1    g1023(.A(KEYINPUT57), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1168), .B1(new_n1176), .B2(new_n1186), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n400), .B1(new_n670), .B2(new_n671), .ZN(new_n1226));
  XNOR2_X1  g1026(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n399), .A2(new_n700), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1227), .ZN(new_n1230));
  OAI211_X1 g1030(.A(new_n400), .B(new_n1230), .C1(new_n670), .C2(new_n671), .ZN(new_n1231));
  AND3_X1   g1031(.A1(new_n1228), .A2(new_n1229), .A3(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1229), .B1(new_n1228), .B2(new_n1231), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1235), .B1(new_n969), .B2(G330), .ZN(new_n1236));
  AOI21_X1  g1036(.A(KEYINPUT40), .B1(new_n904), .B2(new_n949), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n957), .A2(new_n981), .ZN(new_n1238));
  NOR4_X1   g1038(.A1(new_n1237), .A2(new_n1238), .A3(new_n708), .A4(new_n1234), .ZN(new_n1239));
  OAI211_X1 g1039(.A(new_n989), .B(new_n991), .C1(new_n1194), .C2(new_n974), .ZN(new_n1240));
  NOR3_X1   g1040(.A1(new_n1236), .A2(new_n1239), .A3(new_n1240), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n904), .A2(KEYINPUT40), .A3(new_n968), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n952), .B1(new_n953), .B2(new_n956), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1243), .B1(new_n948), .B2(new_n941), .ZN(new_n1244));
  OAI211_X1 g1044(.A(G330), .B(new_n1242), .C1(new_n1244), .C2(KEYINPUT40), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1245), .A2(new_n1234), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n969), .A2(G330), .A3(new_n1235), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n993), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1241), .A2(new_n1248), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1224), .B1(new_n1225), .B2(new_n1249), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1240), .B1(new_n1236), .B2(new_n1239), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1246), .A2(new_n1247), .A3(new_n993), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1198), .B1(new_n1169), .B2(new_n1175), .ZN(new_n1254));
  OAI211_X1 g1054(.A(KEYINPUT57), .B(new_n1253), .C1(new_n1254), .C2(new_n1168), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1250), .A2(new_n718), .A3(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1119), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1234), .A2(new_n777), .ZN(new_n1258));
  NOR3_X1   g1058(.A1(new_n781), .A2(G50), .A3(new_n777), .ZN(new_n1259));
  OAI211_X1 g1059(.A(new_n275), .B(new_n487), .C1(new_n796), .C2(new_n807), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n813), .A2(G132), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n823), .A2(G137), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n804), .A2(new_n1211), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n852), .A2(G128), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1261), .A2(new_n1262), .A3(new_n1263), .A4(new_n1264), .ZN(new_n1265));
  AOI22_X1  g1065(.A1(new_n812), .A2(G125), .B1(G150), .B2(new_n827), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1266), .A2(KEYINPUT123), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1266), .A2(KEYINPUT123), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1265), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  AND2_X1   g1071(.A1(new_n1271), .A2(KEYINPUT59), .ZN(new_n1272));
  AOI211_X1 g1072(.A(new_n1260), .B(new_n1272), .C1(G124), .C2(new_n1021), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1273), .B1(KEYINPUT59), .B2(new_n1271), .ZN(new_n1274));
  AOI21_X1  g1074(.A(G50), .B1(new_n277), .B2(new_n487), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n796), .ZN(new_n1276));
  AOI22_X1  g1076(.A1(G107), .A2(new_n852), .B1(new_n1276), .B2(G58), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1277), .B1(new_n361), .B2(new_n794), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n271), .A2(new_n487), .ZN(new_n1279));
  NOR4_X1   g1079(.A1(new_n1278), .A2(new_n1013), .A3(new_n1093), .A4(new_n1279), .ZN(new_n1280));
  AOI22_X1  g1080(.A1(G97), .A2(new_n813), .B1(new_n812), .B2(G116), .ZN(new_n1281));
  OAI211_X1 g1081(.A(new_n1280), .B(new_n1281), .C1(new_n821), .C2(new_n863), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT58), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1275), .B1(new_n1282), .B2(new_n1283), .ZN(new_n1284));
  OAI211_X1 g1084(.A(new_n1274), .B(new_n1284), .C1(new_n1283), .C2(new_n1282), .ZN(new_n1285));
  AOI211_X1 g1085(.A(new_n776), .B(new_n1259), .C1(new_n1285), .C2(new_n781), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1258), .A2(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1287), .ZN(new_n1288));
  OAI21_X1  g1088(.A(KEYINPUT124), .B1(new_n1257), .B2(new_n1288), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1064), .B1(new_n1241), .B2(new_n1248), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT124), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1290), .A2(new_n1291), .A3(new_n1287), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1289), .A2(new_n1292), .ZN(new_n1293));
  AND3_X1   g1093(.A1(new_n1256), .A2(KEYINPUT125), .A3(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(KEYINPUT125), .B1(new_n1256), .B2(new_n1293), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1294), .A2(new_n1295), .ZN(G375));
  NAND3_X1  g1096(.A1(new_n901), .A2(new_n777), .A3(new_n903), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(new_n876), .A2(G68), .ZN(new_n1298));
  AOI22_X1  g1098(.A1(G116), .A2(new_n813), .B1(new_n812), .B2(G294), .ZN(new_n1299));
  AOI211_X1 g1099(.A(new_n297), .B(new_n1097), .C1(G77), .C2(new_n1276), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n819), .A2(G303), .ZN(new_n1301));
  OAI22_X1  g1101(.A1(new_n803), .A2(new_n601), .B1(new_n794), .B2(new_n512), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1302), .B1(G283), .B2(new_n852), .ZN(new_n1303));
  NAND4_X1  g1103(.A1(new_n1299), .A2(new_n1300), .A3(new_n1301), .A4(new_n1303), .ZN(new_n1304));
  OAI22_X1  g1104(.A1(new_n1026), .A2(new_n862), .B1(new_n801), .B2(new_n1010), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1305), .B1(new_n813), .B2(new_n1211), .ZN(new_n1306));
  XNOR2_X1  g1106(.A(new_n1306), .B(KEYINPUT126), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n819), .A2(G128), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n827), .A2(G50), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n271), .B1(new_n1276), .B2(G58), .ZN(new_n1310));
  AOI22_X1  g1110(.A1(G159), .A2(new_n804), .B1(new_n823), .B2(G150), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1308), .A2(new_n1309), .A3(new_n1310), .A4(new_n1311), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1304), .B1(new_n1307), .B2(new_n1312), .ZN(new_n1313));
  AOI211_X1 g1113(.A(new_n776), .B(new_n1298), .C1(new_n1313), .C2(new_n781), .ZN(new_n1314));
  AOI22_X1  g1114(.A1(new_n1174), .A2(new_n1064), .B1(new_n1297), .B2(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1161), .A2(new_n1168), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1316), .A2(new_n1078), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1315), .B1(new_n1176), .B2(new_n1317), .ZN(G381));
  INV_X1    g1118(.A(new_n1295), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1256), .A2(KEYINPUT125), .A3(new_n1293), .ZN(new_n1320));
  AOI21_X1  g1120(.A(G378), .B1(new_n1319), .B2(new_n1320), .ZN(new_n1321));
  OAI211_X1 g1121(.A(new_n1144), .B(new_n1036), .C1(new_n1063), .C2(new_n1079), .ZN(new_n1322));
  INV_X1    g1122(.A(new_n1322), .ZN(new_n1323));
  NOR3_X1   g1123(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1324), .A2(KEYINPUT127), .ZN(new_n1325));
  NOR2_X1   g1125(.A1(new_n1324), .A2(KEYINPUT127), .ZN(new_n1326));
  NOR2_X1   g1126(.A1(new_n1326), .A2(G381), .ZN(new_n1327));
  NAND4_X1  g1127(.A1(new_n1321), .A2(new_n1323), .A3(new_n1325), .A4(new_n1327), .ZN(G407));
  INV_X1    g1128(.A(G378), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1329), .B1(new_n1294), .B2(new_n1295), .ZN(new_n1330));
  OAI211_X1 g1130(.A(G407), .B(G213), .C1(G343), .C2(new_n1330), .ZN(G409));
  NAND2_X1  g1131(.A1(G387), .A2(G390), .ZN(new_n1332));
  XNOR2_X1  g1132(.A(G393), .B(new_n836), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1332), .A2(new_n1322), .A3(new_n1333), .ZN(new_n1334));
  INV_X1    g1134(.A(new_n1334), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n1333), .B1(new_n1332), .B2(new_n1322), .ZN(new_n1336));
  NOR2_X1   g1136(.A1(new_n1335), .A2(new_n1336), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT60), .ZN(new_n1338));
  OAI21_X1  g1138(.A(new_n718), .B1(new_n1316), .B2(new_n1338), .ZN(new_n1339));
  NAND3_X1  g1139(.A1(new_n1169), .A2(new_n1175), .A3(KEYINPUT60), .ZN(new_n1340));
  AOI21_X1  g1140(.A(new_n1339), .B1(new_n1340), .B2(new_n1316), .ZN(new_n1341));
  INV_X1    g1141(.A(new_n1341), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1342), .A2(G384), .A3(new_n1315), .ZN(new_n1343));
  INV_X1    g1143(.A(new_n1315), .ZN(new_n1344));
  OAI211_X1 g1144(.A(new_n850), .B(new_n879), .C1(new_n1341), .C2(new_n1344), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1343), .A2(new_n1345), .ZN(new_n1346));
  INV_X1    g1146(.A(G213), .ZN(new_n1347));
  NOR2_X1   g1147(.A1(new_n1347), .A2(G343), .ZN(new_n1348));
  NAND3_X1  g1148(.A1(new_n1346), .A2(G2897), .A3(new_n1348), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1348), .A2(G2897), .ZN(new_n1350));
  NAND3_X1  g1150(.A1(new_n1343), .A2(new_n1345), .A3(new_n1350), .ZN(new_n1351));
  AOI21_X1  g1151(.A(new_n1329), .B1(new_n1256), .B2(new_n1293), .ZN(new_n1352));
  NAND4_X1  g1152(.A1(new_n1200), .A2(new_n1222), .A3(new_n1290), .A4(new_n1287), .ZN(new_n1353));
  NOR3_X1   g1153(.A1(new_n1225), .A2(new_n1249), .A3(new_n1077), .ZN(new_n1354));
  OAI22_X1  g1154(.A1(new_n1353), .A2(new_n1354), .B1(new_n1347), .B2(G343), .ZN(new_n1355));
  OAI211_X1 g1155(.A(new_n1349), .B(new_n1351), .C1(new_n1352), .C2(new_n1355), .ZN(new_n1356));
  INV_X1    g1156(.A(KEYINPUT61), .ZN(new_n1357));
  NOR3_X1   g1157(.A1(new_n1352), .A2(new_n1355), .A3(new_n1346), .ZN(new_n1358));
  INV_X1    g1158(.A(KEYINPUT62), .ZN(new_n1359));
  OAI211_X1 g1159(.A(new_n1356), .B(new_n1357), .C1(new_n1358), .C2(new_n1359), .ZN(new_n1360));
  INV_X1    g1160(.A(new_n1352), .ZN(new_n1361));
  INV_X1    g1161(.A(new_n1355), .ZN(new_n1362));
  INV_X1    g1162(.A(new_n1346), .ZN(new_n1363));
  NAND3_X1  g1163(.A1(new_n1361), .A2(new_n1362), .A3(new_n1363), .ZN(new_n1364));
  NOR2_X1   g1164(.A1(new_n1364), .A2(KEYINPUT62), .ZN(new_n1365));
  OAI21_X1  g1165(.A(new_n1337), .B1(new_n1360), .B2(new_n1365), .ZN(new_n1366));
  AND2_X1   g1166(.A1(new_n1349), .A2(new_n1351), .ZN(new_n1367));
  NAND2_X1  g1167(.A1(new_n1361), .A2(new_n1362), .ZN(new_n1368));
  AOI21_X1  g1168(.A(KEYINPUT61), .B1(new_n1367), .B2(new_n1368), .ZN(new_n1369));
  NAND2_X1  g1169(.A1(new_n1332), .A2(new_n1322), .ZN(new_n1370));
  INV_X1    g1170(.A(new_n1333), .ZN(new_n1371));
  NAND2_X1  g1171(.A1(new_n1370), .A2(new_n1371), .ZN(new_n1372));
  NAND2_X1  g1172(.A1(new_n1372), .A2(new_n1334), .ZN(new_n1373));
  INV_X1    g1173(.A(KEYINPUT63), .ZN(new_n1374));
  NAND2_X1  g1174(.A1(new_n1364), .A2(new_n1374), .ZN(new_n1375));
  NAND2_X1  g1175(.A1(new_n1358), .A2(KEYINPUT63), .ZN(new_n1376));
  NAND4_X1  g1176(.A1(new_n1369), .A2(new_n1373), .A3(new_n1375), .A4(new_n1376), .ZN(new_n1377));
  NAND2_X1  g1177(.A1(new_n1366), .A2(new_n1377), .ZN(G405));
  AND3_X1   g1178(.A1(new_n1330), .A2(new_n1346), .A3(new_n1361), .ZN(new_n1379));
  AOI21_X1  g1179(.A(new_n1346), .B1(new_n1330), .B2(new_n1361), .ZN(new_n1380));
  OAI21_X1  g1180(.A(new_n1373), .B1(new_n1379), .B2(new_n1380), .ZN(new_n1381));
  OAI21_X1  g1181(.A(new_n1363), .B1(new_n1321), .B2(new_n1352), .ZN(new_n1382));
  NAND3_X1  g1182(.A1(new_n1330), .A2(new_n1346), .A3(new_n1361), .ZN(new_n1383));
  NAND3_X1  g1183(.A1(new_n1382), .A2(new_n1337), .A3(new_n1383), .ZN(new_n1384));
  NAND2_X1  g1184(.A1(new_n1381), .A2(new_n1384), .ZN(G402));
endmodule


