

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583;

  XOR2_X1 U324 ( .A(KEYINPUT45), .B(KEYINPUT113), .Z(n292) );
  XNOR2_X1 U325 ( .A(n404), .B(n292), .ZN(n405) );
  INV_X1 U326 ( .A(KEYINPUT114), .ZN(n407) );
  XNOR2_X1 U327 ( .A(n430), .B(KEYINPUT55), .ZN(n449) );
  INV_X1 U328 ( .A(G169GAT), .ZN(n451) );
  XNOR2_X1 U329 ( .A(n365), .B(n364), .ZN(n549) );
  XOR2_X1 U330 ( .A(n462), .B(KEYINPUT28), .Z(n520) );
  XNOR2_X1 U331 ( .A(n451), .B(KEYINPUT118), .ZN(n452) );
  XNOR2_X1 U332 ( .A(n453), .B(n452), .ZN(G1348GAT) );
  XOR2_X1 U333 ( .A(KEYINPUT66), .B(KEYINPUT29), .Z(n294) );
  XNOR2_X1 U334 ( .A(KEYINPUT69), .B(KEYINPUT68), .ZN(n293) );
  XNOR2_X1 U335 ( .A(n294), .B(n293), .ZN(n304) );
  XOR2_X1 U336 ( .A(G197GAT), .B(G113GAT), .Z(n296) );
  XOR2_X1 U337 ( .A(G169GAT), .B(G8GAT), .Z(n332) );
  XOR2_X1 U338 ( .A(G15GAT), .B(G1GAT), .Z(n396) );
  XNOR2_X1 U339 ( .A(n332), .B(n396), .ZN(n295) );
  XNOR2_X1 U340 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U341 ( .A(G141GAT), .B(G22GAT), .Z(n416) );
  XOR2_X1 U342 ( .A(n297), .B(n416), .Z(n302) );
  XOR2_X1 U343 ( .A(KEYINPUT30), .B(KEYINPUT70), .Z(n299) );
  NAND2_X1 U344 ( .A1(G229GAT), .A2(G233GAT), .ZN(n298) );
  XNOR2_X1 U345 ( .A(n299), .B(n298), .ZN(n300) );
  XNOR2_X1 U346 ( .A(KEYINPUT67), .B(n300), .ZN(n301) );
  XNOR2_X1 U347 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U348 ( .A(n304), .B(n303), .ZN(n309) );
  XOR2_X1 U349 ( .A(G29GAT), .B(KEYINPUT8), .Z(n306) );
  XNOR2_X1 U350 ( .A(G43GAT), .B(G36GAT), .ZN(n305) );
  XNOR2_X1 U351 ( .A(n306), .B(n305), .ZN(n308) );
  XOR2_X1 U352 ( .A(G50GAT), .B(KEYINPUT7), .Z(n307) );
  XOR2_X1 U353 ( .A(n308), .B(n307), .Z(n360) );
  XOR2_X1 U354 ( .A(n309), .B(n360), .Z(n381) );
  INV_X1 U355 ( .A(n381), .ZN(n566) );
  XOR2_X1 U356 ( .A(KEYINPUT71), .B(n566), .Z(n450) );
  XOR2_X1 U357 ( .A(KEYINPUT6), .B(KEYINPUT92), .Z(n311) );
  XNOR2_X1 U358 ( .A(G141GAT), .B(G148GAT), .ZN(n310) );
  XNOR2_X1 U359 ( .A(n311), .B(n310), .ZN(n315) );
  XOR2_X1 U360 ( .A(KEYINPUT4), .B(KEYINPUT91), .Z(n313) );
  XNOR2_X1 U361 ( .A(KEYINPUT1), .B(KEYINPUT5), .ZN(n312) );
  XNOR2_X1 U362 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U363 ( .A(n315), .B(n314), .Z(n320) );
  XOR2_X1 U364 ( .A(G57GAT), .B(KEYINPUT93), .Z(n317) );
  NAND2_X1 U365 ( .A1(G225GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U366 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U367 ( .A(G1GAT), .B(n318), .ZN(n319) );
  XNOR2_X1 U368 ( .A(n320), .B(n319), .ZN(n326) );
  XOR2_X1 U369 ( .A(G155GAT), .B(KEYINPUT3), .Z(n322) );
  XNOR2_X1 U370 ( .A(G162GAT), .B(KEYINPUT2), .ZN(n321) );
  XNOR2_X1 U371 ( .A(n322), .B(n321), .ZN(n419) );
  XOR2_X1 U372 ( .A(G85GAT), .B(n419), .Z(n324) );
  XNOR2_X1 U373 ( .A(G134GAT), .B(G120GAT), .ZN(n323) );
  XNOR2_X1 U374 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U375 ( .A(n326), .B(n325), .Z(n331) );
  XOR2_X1 U376 ( .A(KEYINPUT81), .B(KEYINPUT0), .Z(n328) );
  XNOR2_X1 U377 ( .A(KEYINPUT82), .B(G127GAT), .ZN(n327) );
  XNOR2_X1 U378 ( .A(n328), .B(n327), .ZN(n329) );
  XOR2_X1 U379 ( .A(G113GAT), .B(n329), .Z(n436) );
  XNOR2_X1 U380 ( .A(G29GAT), .B(n436), .ZN(n330) );
  XOR2_X1 U381 ( .A(n331), .B(n330), .Z(n466) );
  XOR2_X1 U382 ( .A(G190GAT), .B(n332), .Z(n334) );
  NAND2_X1 U383 ( .A1(G226GAT), .A2(G233GAT), .ZN(n333) );
  XNOR2_X1 U384 ( .A(n334), .B(n333), .ZN(n338) );
  XOR2_X1 U385 ( .A(G92GAT), .B(G64GAT), .Z(n336) );
  XNOR2_X1 U386 ( .A(G176GAT), .B(KEYINPUT73), .ZN(n335) );
  XNOR2_X1 U387 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U388 ( .A(G204GAT), .B(n337), .Z(n377) );
  XOR2_X1 U389 ( .A(n338), .B(n377), .Z(n343) );
  XOR2_X1 U390 ( .A(KEYINPUT89), .B(G218GAT), .Z(n340) );
  XNOR2_X1 U391 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n339) );
  XNOR2_X1 U392 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U393 ( .A(G197GAT), .B(n341), .Z(n427) );
  XNOR2_X1 U394 ( .A(G36GAT), .B(n427), .ZN(n342) );
  XNOR2_X1 U395 ( .A(n343), .B(n342), .ZN(n348) );
  XOR2_X1 U396 ( .A(KEYINPUT85), .B(KEYINPUT17), .Z(n345) );
  XNOR2_X1 U397 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n344) );
  XNOR2_X1 U398 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U399 ( .A(KEYINPUT19), .B(n346), .ZN(n446) );
  INV_X1 U400 ( .A(n446), .ZN(n347) );
  XOR2_X1 U401 ( .A(n348), .B(n347), .Z(n455) );
  XNOR2_X1 U402 ( .A(KEYINPUT115), .B(KEYINPUT48), .ZN(n412) );
  XOR2_X1 U403 ( .A(KEYINPUT9), .B(KEYINPUT11), .Z(n350) );
  XNOR2_X1 U404 ( .A(G92GAT), .B(KEYINPUT77), .ZN(n349) );
  XOR2_X1 U405 ( .A(n350), .B(n349), .Z(n365) );
  XOR2_X1 U406 ( .A(KEYINPUT78), .B(KEYINPUT79), .Z(n352) );
  XNOR2_X1 U407 ( .A(G162GAT), .B(G106GAT), .ZN(n351) );
  XNOR2_X1 U408 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U409 ( .A(n353), .B(KEYINPUT10), .Z(n355) );
  XOR2_X1 U410 ( .A(G99GAT), .B(G85GAT), .Z(n372) );
  XNOR2_X1 U411 ( .A(G218GAT), .B(n372), .ZN(n354) );
  XNOR2_X1 U412 ( .A(n355), .B(n354), .ZN(n359) );
  XOR2_X1 U413 ( .A(KEYINPUT65), .B(KEYINPUT76), .Z(n357) );
  NAND2_X1 U414 ( .A1(G232GAT), .A2(G233GAT), .ZN(n356) );
  XNOR2_X1 U415 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U416 ( .A(n359), .B(n358), .Z(n363) );
  INV_X1 U417 ( .A(n360), .ZN(n361) );
  XOR2_X1 U418 ( .A(G190GAT), .B(G134GAT), .Z(n431) );
  XOR2_X1 U419 ( .A(n361), .B(n431), .Z(n362) );
  XNOR2_X1 U420 ( .A(n363), .B(n362), .ZN(n364) );
  XOR2_X1 U421 ( .A(KEYINPUT33), .B(KEYINPUT32), .Z(n371) );
  XNOR2_X1 U422 ( .A(G106GAT), .B(G78GAT), .ZN(n366) );
  XNOR2_X1 U423 ( .A(n366), .B(G148GAT), .ZN(n415) );
  XOR2_X1 U424 ( .A(KEYINPUT72), .B(KEYINPUT74), .Z(n368) );
  XNOR2_X1 U425 ( .A(KEYINPUT75), .B(KEYINPUT31), .ZN(n367) );
  XNOR2_X1 U426 ( .A(n368), .B(n367), .ZN(n369) );
  XNOR2_X1 U427 ( .A(n415), .B(n369), .ZN(n370) );
  XNOR2_X1 U428 ( .A(n371), .B(n370), .ZN(n376) );
  XOR2_X1 U429 ( .A(G57GAT), .B(KEYINPUT13), .Z(n386) );
  XOR2_X1 U430 ( .A(n386), .B(n372), .Z(n374) );
  NAND2_X1 U431 ( .A1(G230GAT), .A2(G233GAT), .ZN(n373) );
  XNOR2_X1 U432 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U433 ( .A(n376), .B(n375), .Z(n379) );
  XOR2_X1 U434 ( .A(G120GAT), .B(G71GAT), .Z(n432) );
  XNOR2_X1 U435 ( .A(n432), .B(n377), .ZN(n378) );
  XNOR2_X1 U436 ( .A(n379), .B(n378), .ZN(n571) );
  XNOR2_X1 U437 ( .A(KEYINPUT41), .B(KEYINPUT64), .ZN(n380) );
  XOR2_X1 U438 ( .A(n571), .B(n380), .Z(n552) );
  INV_X1 U439 ( .A(n552), .ZN(n530) );
  NAND2_X1 U440 ( .A1(n381), .A2(n530), .ZN(n382) );
  XNOR2_X1 U441 ( .A(n382), .B(KEYINPUT112), .ZN(n383) );
  XNOR2_X1 U442 ( .A(KEYINPUT46), .B(n383), .ZN(n401) );
  XOR2_X1 U443 ( .A(G155GAT), .B(G71GAT), .Z(n385) );
  XNOR2_X1 U444 ( .A(G183GAT), .B(G127GAT), .ZN(n384) );
  XNOR2_X1 U445 ( .A(n385), .B(n384), .ZN(n400) );
  XOR2_X1 U446 ( .A(n386), .B(KEYINPUT14), .Z(n388) );
  NAND2_X1 U447 ( .A1(G231GAT), .A2(G233GAT), .ZN(n387) );
  XNOR2_X1 U448 ( .A(n388), .B(n387), .ZN(n392) );
  XOR2_X1 U449 ( .A(KEYINPUT12), .B(KEYINPUT15), .Z(n390) );
  XNOR2_X1 U450 ( .A(G8GAT), .B(KEYINPUT80), .ZN(n389) );
  XNOR2_X1 U451 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U452 ( .A(n392), .B(n391), .Z(n398) );
  XOR2_X1 U453 ( .A(G64GAT), .B(G78GAT), .Z(n394) );
  XNOR2_X1 U454 ( .A(G22GAT), .B(G211GAT), .ZN(n393) );
  XNOR2_X1 U455 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U456 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U457 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U458 ( .A(n400), .B(n399), .ZN(n533) );
  INV_X1 U459 ( .A(n533), .ZN(n576) );
  NAND2_X1 U460 ( .A1(n401), .A2(n576), .ZN(n402) );
  NOR2_X1 U461 ( .A1(n549), .A2(n402), .ZN(n403) );
  XNOR2_X1 U462 ( .A(KEYINPUT47), .B(n403), .ZN(n410) );
  INV_X1 U463 ( .A(n450), .ZN(n528) );
  XOR2_X1 U464 ( .A(KEYINPUT36), .B(n549), .Z(n580) );
  NOR2_X1 U465 ( .A1(n576), .A2(n580), .ZN(n404) );
  NAND2_X1 U466 ( .A1(n405), .A2(n571), .ZN(n406) );
  NOR2_X1 U467 ( .A1(n528), .A2(n406), .ZN(n408) );
  XNOR2_X1 U468 ( .A(n408), .B(n407), .ZN(n409) );
  NAND2_X1 U469 ( .A1(n410), .A2(n409), .ZN(n411) );
  XNOR2_X1 U470 ( .A(n412), .B(n411), .ZN(n540) );
  NOR2_X1 U471 ( .A1(n455), .A2(n540), .ZN(n413) );
  XNOR2_X1 U472 ( .A(n413), .B(KEYINPUT54), .ZN(n414) );
  AND2_X1 U473 ( .A1(n466), .A2(n414), .ZN(n565) );
  XOR2_X1 U474 ( .A(n415), .B(KEYINPUT88), .Z(n418) );
  XNOR2_X1 U475 ( .A(G50GAT), .B(n416), .ZN(n417) );
  XNOR2_X1 U476 ( .A(n418), .B(n417), .ZN(n423) );
  XOR2_X1 U477 ( .A(n419), .B(KEYINPUT24), .Z(n421) );
  NAND2_X1 U478 ( .A1(G228GAT), .A2(G233GAT), .ZN(n420) );
  XNOR2_X1 U479 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U480 ( .A(n423), .B(n422), .Z(n429) );
  XOR2_X1 U481 ( .A(KEYINPUT22), .B(G204GAT), .Z(n425) );
  XNOR2_X1 U482 ( .A(KEYINPUT23), .B(KEYINPUT90), .ZN(n424) );
  XNOR2_X1 U483 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U484 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U485 ( .A(n429), .B(n428), .ZN(n462) );
  NAND2_X1 U486 ( .A1(n565), .A2(n462), .ZN(n430) );
  XOR2_X1 U487 ( .A(n432), .B(n431), .Z(n434) );
  NAND2_X1 U488 ( .A1(G227GAT), .A2(G233GAT), .ZN(n433) );
  XNOR2_X1 U489 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U490 ( .A(n435), .B(G99GAT), .Z(n438) );
  XNOR2_X1 U491 ( .A(G43GAT), .B(n436), .ZN(n437) );
  XNOR2_X1 U492 ( .A(n438), .B(n437), .ZN(n442) );
  XOR2_X1 U493 ( .A(G176GAT), .B(KEYINPUT84), .Z(n440) );
  XNOR2_X1 U494 ( .A(G169GAT), .B(KEYINPUT20), .ZN(n439) );
  XNOR2_X1 U495 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U496 ( .A(n442), .B(n441), .Z(n448) );
  XOR2_X1 U497 ( .A(KEYINPUT87), .B(KEYINPUT86), .Z(n444) );
  XNOR2_X1 U498 ( .A(G15GAT), .B(KEYINPUT83), .ZN(n443) );
  XNOR2_X1 U499 ( .A(n444), .B(n443), .ZN(n445) );
  XOR2_X1 U500 ( .A(n446), .B(n445), .Z(n447) );
  XOR2_X1 U501 ( .A(n448), .B(n447), .Z(n458) );
  INV_X1 U502 ( .A(n458), .ZN(n526) );
  NAND2_X1 U503 ( .A1(n449), .A2(n526), .ZN(n560) );
  NOR2_X1 U504 ( .A1(n450), .A2(n560), .ZN(n453) );
  XOR2_X1 U505 ( .A(KEYINPUT34), .B(KEYINPUT96), .Z(n472) );
  NAND2_X1 U506 ( .A1(n571), .A2(n528), .ZN(n486) );
  NOR2_X1 U507 ( .A1(n549), .A2(n576), .ZN(n454) );
  XNOR2_X1 U508 ( .A(n454), .B(KEYINPUT16), .ZN(n470) );
  INV_X1 U509 ( .A(n455), .ZN(n516) );
  XNOR2_X1 U510 ( .A(n516), .B(KEYINPUT94), .ZN(n456) );
  XNOR2_X1 U511 ( .A(KEYINPUT27), .B(n456), .ZN(n460) );
  INV_X1 U512 ( .A(n466), .ZN(n514) );
  NAND2_X1 U513 ( .A1(n460), .A2(n514), .ZN(n457) );
  XOR2_X1 U514 ( .A(KEYINPUT95), .B(n457), .Z(n539) );
  NOR2_X1 U515 ( .A1(n520), .A2(n539), .ZN(n525) );
  NAND2_X1 U516 ( .A1(n525), .A2(n458), .ZN(n469) );
  NOR2_X1 U517 ( .A1(n462), .A2(n526), .ZN(n459) );
  XNOR2_X1 U518 ( .A(n459), .B(KEYINPUT26), .ZN(n564) );
  NAND2_X1 U519 ( .A1(n460), .A2(n564), .ZN(n465) );
  NAND2_X1 U520 ( .A1(n526), .A2(n516), .ZN(n461) );
  NAND2_X1 U521 ( .A1(n462), .A2(n461), .ZN(n463) );
  XOR2_X1 U522 ( .A(KEYINPUT25), .B(n463), .Z(n464) );
  NAND2_X1 U523 ( .A1(n465), .A2(n464), .ZN(n467) );
  NAND2_X1 U524 ( .A1(n467), .A2(n466), .ZN(n468) );
  NAND2_X1 U525 ( .A1(n469), .A2(n468), .ZN(n482) );
  NAND2_X1 U526 ( .A1(n470), .A2(n482), .ZN(n502) );
  NOR2_X1 U527 ( .A1(n486), .A2(n502), .ZN(n480) );
  NAND2_X1 U528 ( .A1(n480), .A2(n514), .ZN(n471) );
  XNOR2_X1 U529 ( .A(n472), .B(n471), .ZN(n473) );
  XOR2_X1 U530 ( .A(G1GAT), .B(n473), .Z(G1324GAT) );
  NAND2_X1 U531 ( .A1(n516), .A2(n480), .ZN(n474) );
  XNOR2_X1 U532 ( .A(n474), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U533 ( .A(KEYINPUT98), .B(KEYINPUT99), .Z(n476) );
  XNOR2_X1 U534 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n475) );
  XNOR2_X1 U535 ( .A(n476), .B(n475), .ZN(n479) );
  NAND2_X1 U536 ( .A1(n480), .A2(n526), .ZN(n477) );
  XNOR2_X1 U537 ( .A(n477), .B(KEYINPUT97), .ZN(n478) );
  XNOR2_X1 U538 ( .A(n479), .B(n478), .ZN(G1326GAT) );
  NAND2_X1 U539 ( .A1(n480), .A2(n520), .ZN(n481) );
  XNOR2_X1 U540 ( .A(n481), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U541 ( .A1(n576), .A2(n482), .ZN(n483) );
  NOR2_X1 U542 ( .A1(n580), .A2(n483), .ZN(n484) );
  XOR2_X1 U543 ( .A(n484), .B(KEYINPUT101), .Z(n485) );
  XNOR2_X1 U544 ( .A(KEYINPUT37), .B(n485), .ZN(n512) );
  NOR2_X1 U545 ( .A1(n512), .A2(n486), .ZN(n488) );
  XNOR2_X1 U546 ( .A(KEYINPUT102), .B(KEYINPUT38), .ZN(n487) );
  XNOR2_X1 U547 ( .A(n488), .B(n487), .ZN(n499) );
  NAND2_X1 U548 ( .A1(n514), .A2(n499), .ZN(n490) );
  XOR2_X1 U549 ( .A(KEYINPUT100), .B(KEYINPUT39), .Z(n489) );
  XNOR2_X1 U550 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U551 ( .A(G29GAT), .B(n491), .ZN(G1328GAT) );
  XOR2_X1 U552 ( .A(KEYINPUT103), .B(KEYINPUT104), .Z(n493) );
  NAND2_X1 U553 ( .A1(n499), .A2(n516), .ZN(n492) );
  XNOR2_X1 U554 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U555 ( .A(G36GAT), .B(n494), .ZN(G1329GAT) );
  XNOR2_X1 U556 ( .A(G43GAT), .B(KEYINPUT106), .ZN(n498) );
  XOR2_X1 U557 ( .A(KEYINPUT40), .B(KEYINPUT105), .Z(n496) );
  NAND2_X1 U558 ( .A1(n499), .A2(n526), .ZN(n495) );
  XNOR2_X1 U559 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U560 ( .A(n498), .B(n497), .ZN(G1330GAT) );
  XOR2_X1 U561 ( .A(G50GAT), .B(KEYINPUT107), .Z(n501) );
  NAND2_X1 U562 ( .A1(n499), .A2(n520), .ZN(n500) );
  XNOR2_X1 U563 ( .A(n501), .B(n500), .ZN(G1331GAT) );
  XOR2_X1 U564 ( .A(KEYINPUT108), .B(KEYINPUT42), .Z(n504) );
  NAND2_X1 U565 ( .A1(n566), .A2(n530), .ZN(n511) );
  NOR2_X1 U566 ( .A1(n511), .A2(n502), .ZN(n508) );
  NAND2_X1 U567 ( .A1(n508), .A2(n514), .ZN(n503) );
  XNOR2_X1 U568 ( .A(n504), .B(n503), .ZN(n505) );
  XOR2_X1 U569 ( .A(G57GAT), .B(n505), .Z(G1332GAT) );
  NAND2_X1 U570 ( .A1(n516), .A2(n508), .ZN(n506) );
  XNOR2_X1 U571 ( .A(n506), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U572 ( .A1(n508), .A2(n526), .ZN(n507) );
  XNOR2_X1 U573 ( .A(n507), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U574 ( .A(G78GAT), .B(KEYINPUT43), .Z(n510) );
  NAND2_X1 U575 ( .A1(n508), .A2(n520), .ZN(n509) );
  XNOR2_X1 U576 ( .A(n510), .B(n509), .ZN(G1335GAT) );
  NOR2_X1 U577 ( .A1(n512), .A2(n511), .ZN(n513) );
  XOR2_X1 U578 ( .A(KEYINPUT109), .B(n513), .Z(n521) );
  NAND2_X1 U579 ( .A1(n514), .A2(n521), .ZN(n515) );
  XNOR2_X1 U580 ( .A(G85GAT), .B(n515), .ZN(G1336GAT) );
  NAND2_X1 U581 ( .A1(n516), .A2(n521), .ZN(n517) );
  XNOR2_X1 U582 ( .A(n517), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U583 ( .A1(n521), .A2(n526), .ZN(n518) );
  XNOR2_X1 U584 ( .A(n518), .B(KEYINPUT110), .ZN(n519) );
  XNOR2_X1 U585 ( .A(G99GAT), .B(n519), .ZN(G1338GAT) );
  XOR2_X1 U586 ( .A(KEYINPUT111), .B(KEYINPUT44), .Z(n523) );
  NAND2_X1 U587 ( .A1(n521), .A2(n520), .ZN(n522) );
  XNOR2_X1 U588 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U589 ( .A(G106GAT), .B(n524), .ZN(G1339GAT) );
  NAND2_X1 U590 ( .A1(n526), .A2(n525), .ZN(n527) );
  NOR2_X1 U591 ( .A1(n540), .A2(n527), .ZN(n536) );
  NAND2_X1 U592 ( .A1(n528), .A2(n536), .ZN(n529) );
  XNOR2_X1 U593 ( .A(n529), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U594 ( .A(G120GAT), .B(KEYINPUT49), .Z(n532) );
  NAND2_X1 U595 ( .A1(n536), .A2(n530), .ZN(n531) );
  XNOR2_X1 U596 ( .A(n532), .B(n531), .ZN(G1341GAT) );
  NAND2_X1 U597 ( .A1(n533), .A2(n536), .ZN(n534) );
  XNOR2_X1 U598 ( .A(n534), .B(KEYINPUT50), .ZN(n535) );
  XNOR2_X1 U599 ( .A(G127GAT), .B(n535), .ZN(G1342GAT) );
  XOR2_X1 U600 ( .A(G134GAT), .B(KEYINPUT51), .Z(n538) );
  NAND2_X1 U601 ( .A1(n536), .A2(n549), .ZN(n537) );
  XNOR2_X1 U602 ( .A(n538), .B(n537), .ZN(G1343GAT) );
  NOR2_X1 U603 ( .A1(n540), .A2(n539), .ZN(n541) );
  NAND2_X1 U604 ( .A1(n541), .A2(n564), .ZN(n550) );
  NOR2_X1 U605 ( .A1(n566), .A2(n550), .ZN(n542) );
  XOR2_X1 U606 ( .A(KEYINPUT116), .B(n542), .Z(n543) );
  XNOR2_X1 U607 ( .A(G141GAT), .B(n543), .ZN(G1344GAT) );
  NOR2_X1 U608 ( .A1(n550), .A2(n552), .ZN(n547) );
  XOR2_X1 U609 ( .A(KEYINPUT52), .B(KEYINPUT117), .Z(n545) );
  XNOR2_X1 U610 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n544) );
  XNOR2_X1 U611 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U612 ( .A(n547), .B(n546), .ZN(G1345GAT) );
  NOR2_X1 U613 ( .A1(n576), .A2(n550), .ZN(n548) );
  XOR2_X1 U614 ( .A(G155GAT), .B(n548), .Z(G1346GAT) );
  INV_X1 U615 ( .A(n549), .ZN(n561) );
  NOR2_X1 U616 ( .A1(n561), .A2(n550), .ZN(n551) );
  XOR2_X1 U617 ( .A(G162GAT), .B(n551), .Z(G1347GAT) );
  NOR2_X1 U618 ( .A1(n560), .A2(n552), .ZN(n556) );
  XOR2_X1 U619 ( .A(KEYINPUT119), .B(KEYINPUT56), .Z(n554) );
  XNOR2_X1 U620 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n553) );
  XNOR2_X1 U621 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n556), .B(n555), .ZN(G1349GAT) );
  NOR2_X1 U623 ( .A1(n576), .A2(n560), .ZN(n557) );
  XOR2_X1 U624 ( .A(G183GAT), .B(n557), .Z(G1350GAT) );
  XOR2_X1 U625 ( .A(KEYINPUT120), .B(KEYINPUT58), .Z(n559) );
  XNOR2_X1 U626 ( .A(G190GAT), .B(KEYINPUT121), .ZN(n558) );
  XNOR2_X1 U627 ( .A(n559), .B(n558), .ZN(n563) );
  NOR2_X1 U628 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U629 ( .A(n563), .B(n562), .Z(G1351GAT) );
  NAND2_X1 U630 ( .A1(n565), .A2(n564), .ZN(n579) );
  OR2_X1 U631 ( .A1(n566), .A2(n579), .ZN(n570) );
  XOR2_X1 U632 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n568) );
  XNOR2_X1 U633 ( .A(G197GAT), .B(KEYINPUT122), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(G1352GAT) );
  NOR2_X1 U636 ( .A1(n579), .A2(n571), .ZN(n575) );
  XOR2_X1 U637 ( .A(KEYINPUT123), .B(KEYINPUT61), .Z(n573) );
  XNOR2_X1 U638 ( .A(G204GAT), .B(KEYINPUT124), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n573), .B(n572), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(G1353GAT) );
  NOR2_X1 U641 ( .A1(n576), .A2(n579), .ZN(n578) );
  XNOR2_X1 U642 ( .A(G211GAT), .B(KEYINPUT125), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(G1354GAT) );
  NOR2_X1 U644 ( .A1(n580), .A2(n579), .ZN(n582) );
  XNOR2_X1 U645 ( .A(KEYINPUT62), .B(KEYINPUT126), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n582), .B(n581), .ZN(n583) );
  XOR2_X1 U647 ( .A(G218GAT), .B(n583), .Z(G1355GAT) );
endmodule

