//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 1 1 1 0 1 0 0 1 0 0 0 1 0 1 1 0 0 0 1 1 1 1 0 0 0 0 0 0 0 0 1 0 1 1 1 1 1 1 1 1 1 1 1 1 1 0 0 0 1 0 0 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:14 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n689,
    new_n690, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n707, new_n708, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n727, new_n728, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n894, new_n895, new_n896, new_n897, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n926, new_n927, new_n928, new_n929,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961;
  INV_X1    g000(.A(G237), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n187), .A2(new_n188), .A3(G214), .ZN(new_n189));
  OR2_X1    g003(.A1(KEYINPUT95), .A2(G143), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n189), .B(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT18), .ZN(new_n192));
  INV_X1    g006(.A(G131), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n191), .B1(new_n192), .B2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT96), .ZN(new_n195));
  XNOR2_X1  g009(.A(new_n194), .B(new_n195), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n191), .A2(new_n193), .ZN(new_n197));
  XNOR2_X1  g011(.A(G125), .B(G140), .ZN(new_n198));
  INV_X1    g012(.A(G146), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  XOR2_X1   g014(.A(G125), .B(G140), .Z(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G146), .ZN(new_n202));
  AOI22_X1  g016(.A1(new_n197), .A2(KEYINPUT18), .B1(new_n200), .B2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n196), .A2(new_n203), .ZN(new_n204));
  XNOR2_X1  g018(.A(G113), .B(G122), .ZN(new_n205));
  INV_X1    g019(.A(G104), .ZN(new_n206));
  XNOR2_X1  g020(.A(new_n205), .B(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G125), .ZN(new_n208));
  OR3_X1    g022(.A1(new_n208), .A2(KEYINPUT16), .A3(G140), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT16), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n209), .B1(new_n201), .B2(new_n210), .ZN(new_n211));
  XNOR2_X1  g025(.A(new_n211), .B(G146), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n197), .A2(KEYINPUT17), .ZN(new_n213));
  XNOR2_X1  g027(.A(new_n191), .B(new_n193), .ZN(new_n214));
  OAI211_X1 g028(.A(new_n212), .B(new_n213), .C1(new_n214), .C2(KEYINPUT17), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n204), .A2(new_n207), .A3(new_n215), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n211), .A2(new_n199), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n201), .A2(KEYINPUT97), .ZN(new_n218));
  XNOR2_X1  g032(.A(new_n218), .B(KEYINPUT19), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n217), .B1(new_n219), .B2(new_n199), .ZN(new_n220));
  AOI22_X1  g034(.A1(new_n203), .A2(new_n196), .B1(new_n220), .B2(new_n214), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n216), .B1(new_n221), .B2(new_n207), .ZN(new_n222));
  NOR2_X1   g036(.A1(G475), .A2(G902), .ZN(new_n223));
  XOR2_X1   g037(.A(new_n223), .B(KEYINPUT98), .Z(new_n224));
  NAND3_X1  g038(.A1(new_n222), .A2(KEYINPUT20), .A3(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  AOI21_X1  g040(.A(KEYINPUT20), .B1(new_n222), .B2(new_n224), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(G122), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(G116), .ZN(new_n230));
  XNOR2_X1  g044(.A(KEYINPUT69), .B(G116), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n230), .B1(new_n231), .B2(new_n229), .ZN(new_n232));
  XNOR2_X1  g046(.A(new_n232), .B(G107), .ZN(new_n233));
  OR2_X1    g047(.A1(KEYINPUT64), .A2(G134), .ZN(new_n234));
  NAND2_X1  g048(.A1(KEYINPUT64), .A2(G134), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(G143), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(G128), .ZN(new_n239));
  XNOR2_X1  g053(.A(KEYINPUT66), .B(G128), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n239), .B1(new_n240), .B2(new_n238), .ZN(new_n241));
  INV_X1    g055(.A(G134), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT13), .ZN(new_n243));
  OAI22_X1  g057(.A1(new_n240), .A2(new_n238), .B1(new_n243), .B2(new_n239), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n244), .B1(new_n243), .B2(new_n239), .ZN(new_n245));
  OAI221_X1 g059(.A(new_n233), .B1(new_n237), .B2(new_n241), .C1(new_n242), .C2(new_n245), .ZN(new_n246));
  XNOR2_X1  g060(.A(new_n241), .B(new_n237), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n231), .A2(new_n229), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(KEYINPUT14), .ZN(new_n249));
  OAI211_X1 g063(.A(new_n249), .B(G107), .C1(KEYINPUT14), .C2(new_n232), .ZN(new_n250));
  OAI211_X1 g064(.A(new_n247), .B(new_n250), .C1(G107), .C2(new_n232), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n246), .A2(new_n251), .ZN(new_n252));
  XOR2_X1   g066(.A(KEYINPUT9), .B(G234), .Z(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(G217), .ZN(new_n255));
  NOR3_X1   g069(.A1(new_n254), .A2(new_n255), .A3(G953), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n252), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n246), .A2(new_n251), .A3(new_n256), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n258), .A2(KEYINPUT99), .A3(new_n259), .ZN(new_n260));
  OR3_X1    g074(.A1(new_n252), .A2(KEYINPUT99), .A3(new_n257), .ZN(new_n261));
  INV_X1    g075(.A(G902), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n260), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(G478), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n264), .A2(KEYINPUT15), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(new_n265), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n260), .A2(new_n261), .A3(new_n262), .A4(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n216), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n207), .B1(new_n204), .B2(new_n215), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n262), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(G475), .ZN(new_n272));
  NAND4_X1  g086(.A1(new_n228), .A2(new_n266), .A3(new_n268), .A4(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(G234), .A2(G237), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n274), .A2(G952), .A3(new_n188), .ZN(new_n275));
  XOR2_X1   g089(.A(KEYINPUT21), .B(G898), .Z(new_n276));
  NAND3_X1  g090(.A1(new_n274), .A2(G902), .A3(G953), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n275), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  NOR3_X1   g093(.A1(new_n273), .A2(KEYINPUT100), .A3(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT100), .ZN(new_n281));
  INV_X1    g095(.A(new_n227), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n282), .A2(new_n272), .A3(new_n225), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n266), .A2(new_n268), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n281), .B1(new_n285), .B2(new_n278), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n280), .A2(new_n286), .ZN(new_n287));
  OAI21_X1  g101(.A(G210), .B1(G237), .B2(G902), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n199), .A2(G143), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n238), .A2(G146), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  AND2_X1   g106(.A1(KEYINPUT0), .A2(G128), .ZN(new_n293));
  NOR2_X1   g107(.A1(KEYINPUT0), .A2(G128), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n292), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n295), .B1(new_n292), .B2(new_n293), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(G125), .ZN(new_n297));
  AND2_X1   g111(.A1(new_n290), .A2(new_n291), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT1), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n298), .A2(new_n299), .A3(G128), .ZN(new_n300));
  INV_X1    g114(.A(G128), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(KEYINPUT66), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT66), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(G128), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n299), .B1(G143), .B2(new_n199), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n292), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n300), .A2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n297), .B1(new_n309), .B2(G125), .ZN(new_n310));
  XNOR2_X1  g124(.A(new_n310), .B(KEYINPUT92), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n188), .A2(G224), .ZN(new_n312));
  XNOR2_X1  g126(.A(new_n311), .B(new_n312), .ZN(new_n313));
  XOR2_X1   g127(.A(G110), .B(G122), .Z(new_n314));
  OAI21_X1  g128(.A(KEYINPUT3), .B1(new_n206), .B2(G107), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT3), .ZN(new_n316));
  INV_X1    g130(.A(G107), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n316), .A2(new_n317), .A3(G104), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n206), .A2(G107), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n315), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT80), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND4_X1  g136(.A1(new_n315), .A2(new_n318), .A3(KEYINPUT80), .A4(new_n319), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n322), .A2(G101), .A3(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(G101), .ZN(new_n325));
  NAND4_X1  g139(.A1(new_n315), .A2(new_n318), .A3(new_n325), .A4(new_n319), .ZN(new_n326));
  AND2_X1   g140(.A1(new_n326), .A2(KEYINPUT4), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n324), .A2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT81), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n324), .A2(KEYINPUT81), .A3(new_n327), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(G119), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(G116), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n334), .B1(new_n231), .B2(new_n333), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT68), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT2), .ZN(new_n337));
  INV_X1    g151(.A(G113), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n337), .A2(new_n338), .A3(KEYINPUT67), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT67), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n340), .B1(KEYINPUT2), .B2(G113), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  AND2_X1   g156(.A1(KEYINPUT2), .A2(G113), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n336), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  AOI211_X1 g159(.A(KEYINPUT68), .B(new_n343), .C1(new_n339), .C2(new_n341), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n335), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT70), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n342), .A2(new_n344), .ZN(new_n350));
  OR2_X1    g164(.A1(new_n335), .A2(new_n350), .ZN(new_n351));
  OAI211_X1 g165(.A(KEYINPUT70), .B(new_n335), .C1(new_n345), .C2(new_n346), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n349), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  AND2_X1   g167(.A1(new_n322), .A2(new_n323), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT82), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT4), .ZN(new_n356));
  NAND4_X1  g170(.A1(new_n354), .A2(new_n355), .A3(new_n356), .A4(G101), .ZN(new_n357));
  OAI21_X1  g171(.A(KEYINPUT82), .B1(new_n324), .B2(KEYINPUT4), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n332), .A2(new_n353), .A3(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT5), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n361), .A2(new_n333), .A3(G116), .ZN(new_n362));
  OAI211_X1 g176(.A(G113), .B(new_n362), .C1(new_n335), .C2(new_n361), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n351), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT83), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n365), .A2(new_n317), .A3(G104), .ZN(new_n366));
  OAI21_X1  g180(.A(KEYINPUT83), .B1(new_n317), .B2(G104), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n206), .A2(G107), .ZN(new_n368));
  OAI211_X1 g182(.A(G101), .B(new_n366), .C1(new_n367), .C2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(new_n326), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT86), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n369), .A2(new_n326), .A3(KEYINPUT86), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  OAI21_X1  g188(.A(KEYINPUT90), .B1(new_n364), .B2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n373), .ZN(new_n376));
  AOI21_X1  g190(.A(KEYINPUT86), .B1(new_n369), .B2(new_n326), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT90), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n378), .A2(new_n379), .A3(new_n351), .A4(new_n363), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n375), .A2(new_n380), .ZN(new_n381));
  AND3_X1   g195(.A1(new_n360), .A2(new_n381), .A3(KEYINPUT91), .ZN(new_n382));
  AOI21_X1  g196(.A(KEYINPUT91), .B1(new_n360), .B2(new_n381), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n314), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(new_n314), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n360), .A2(new_n381), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(KEYINPUT6), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n384), .A2(new_n387), .ZN(new_n388));
  OAI211_X1 g202(.A(KEYINPUT6), .B(new_n314), .C1(new_n382), .C2(new_n383), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n313), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n312), .A2(KEYINPUT7), .ZN(new_n391));
  XNOR2_X1  g205(.A(new_n310), .B(new_n391), .ZN(new_n392));
  XOR2_X1   g206(.A(new_n314), .B(KEYINPUT8), .Z(new_n393));
  AND2_X1   g207(.A1(new_n364), .A2(new_n370), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n364), .A2(new_n374), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n393), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n386), .A2(new_n392), .A3(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT93), .ZN(new_n398));
  AND3_X1   g212(.A1(new_n397), .A2(new_n398), .A3(new_n262), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n398), .B1(new_n397), .B2(new_n262), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n289), .B1(new_n390), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n360), .A2(new_n381), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT91), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n360), .A2(new_n381), .A3(KEYINPUT91), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n385), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(new_n387), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n389), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(new_n313), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(new_n400), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n397), .A2(new_n398), .A3(new_n262), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n411), .A2(new_n288), .A3(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT94), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n402), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n288), .B1(new_n411), .B2(new_n414), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(KEYINPUT94), .ZN(new_n419));
  OAI21_X1  g233(.A(G214), .B1(G237), .B2(G902), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n417), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n287), .A2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(G472), .ZN(new_n423));
  XNOR2_X1  g237(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n424));
  XNOR2_X1  g238(.A(new_n424), .B(G101), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n187), .A2(new_n188), .A3(G210), .ZN(new_n426));
  XNOR2_X1  g240(.A(new_n425), .B(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT28), .ZN(new_n429));
  INV_X1    g243(.A(new_n235), .ZN(new_n430));
  NOR2_X1   g244(.A1(KEYINPUT64), .A2(G134), .ZN(new_n431));
  INV_X1    g245(.A(G137), .ZN(new_n432));
  NOR3_X1   g246(.A1(new_n430), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  NOR2_X1   g247(.A1(G134), .A2(G137), .ZN(new_n434));
  OAI21_X1  g248(.A(KEYINPUT11), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NOR4_X1   g249(.A1(new_n430), .A2(new_n431), .A3(KEYINPUT11), .A4(G137), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  AOI21_X1  g251(.A(G131), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT11), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n234), .A2(G137), .A3(new_n235), .ZN(new_n440));
  INV_X1    g254(.A(new_n434), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n439), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NOR3_X1   g256(.A1(new_n442), .A2(new_n193), .A3(new_n436), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n296), .B1(new_n438), .B2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT65), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n435), .A2(new_n437), .A3(G131), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n193), .B1(new_n442), .B2(new_n436), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n449), .A2(KEYINPUT65), .A3(new_n296), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n236), .A2(G137), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n432), .A2(G134), .ZN(new_n452));
  OAI21_X1  g266(.A(G131), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n448), .A2(new_n308), .A3(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n446), .A2(new_n450), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(new_n353), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n444), .A2(new_n454), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n457), .A2(new_n353), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n429), .B1(new_n456), .B2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT71), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n461), .B1(new_n458), .B2(KEYINPUT28), .ZN(new_n462));
  OAI211_X1 g276(.A(KEYINPUT71), .B(new_n429), .C1(new_n457), .C2(new_n353), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n428), .B1(new_n460), .B2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT30), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n455), .A2(new_n466), .ZN(new_n467));
  OAI211_X1 g281(.A(new_n467), .B(new_n353), .C1(new_n466), .C2(new_n457), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT31), .ZN(new_n469));
  NAND4_X1  g283(.A1(new_n468), .A2(new_n469), .A3(new_n459), .A4(new_n427), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n465), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n457), .A2(new_n466), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n472), .B1(new_n455), .B2(new_n466), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n458), .B1(new_n473), .B2(new_n353), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n469), .B1(new_n474), .B2(new_n427), .ZN(new_n475));
  OAI211_X1 g289(.A(new_n423), .B(new_n262), .C1(new_n471), .C2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(KEYINPUT32), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n468), .A2(new_n459), .ZN(new_n478));
  OAI21_X1  g292(.A(KEYINPUT31), .B1(new_n478), .B2(new_n428), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n479), .A2(new_n470), .A3(new_n465), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT32), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n480), .A2(new_n481), .A3(new_n423), .A4(new_n262), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n477), .A2(new_n482), .ZN(new_n483));
  OR2_X1    g297(.A1(new_n460), .A2(new_n464), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n427), .B1(new_n484), .B2(KEYINPUT29), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n474), .A2(new_n428), .ZN(new_n486));
  AOI21_X1  g300(.A(KEYINPUT29), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n457), .A2(new_n353), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n429), .B1(new_n459), .B2(new_n488), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n464), .A2(new_n489), .ZN(new_n490));
  OAI211_X1 g304(.A(new_n427), .B(new_n490), .C1(new_n484), .C2(KEYINPUT29), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(new_n262), .ZN(new_n492));
  OAI21_X1  g306(.A(G472), .B1(new_n487), .B2(new_n492), .ZN(new_n493));
  AND2_X1   g307(.A1(KEYINPUT76), .A2(KEYINPUT25), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n301), .A2(G119), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n496), .B1(new_n240), .B2(new_n333), .ZN(new_n497));
  XNOR2_X1  g311(.A(KEYINPUT24), .B(G110), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n497), .A2(KEYINPUT73), .A3(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  AOI21_X1  g314(.A(KEYINPUT73), .B1(new_n497), .B2(new_n498), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g316(.A(KEYINPUT23), .B1(new_n301), .B2(G119), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n495), .B1(new_n305), .B2(G119), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT23), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  OAI21_X1  g321(.A(KEYINPUT72), .B1(new_n507), .B2(G110), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n503), .B1(new_n497), .B2(KEYINPUT23), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT72), .ZN(new_n510));
  INV_X1    g324(.A(G110), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n509), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n502), .A2(new_n508), .A3(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(new_n217), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n513), .A2(new_n514), .A3(new_n200), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n497), .A2(new_n498), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n212), .A2(new_n516), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n517), .B1(new_n511), .B2(new_n509), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n519), .B(KEYINPUT22), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n520), .B(G137), .ZN(new_n521));
  AND4_X1   g335(.A1(KEYINPUT75), .A2(new_n515), .A3(new_n518), .A4(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n515), .A2(new_n518), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT74), .ZN(new_n524));
  XNOR2_X1  g338(.A(new_n521), .B(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(KEYINPUT75), .B1(new_n523), .B2(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n515), .A2(new_n518), .A3(new_n521), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n522), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n494), .B1(new_n529), .B2(G902), .ZN(new_n530));
  NOR2_X1   g344(.A1(KEYINPUT76), .A2(KEYINPUT25), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n494), .A2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(new_n528), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n525), .B1(new_n515), .B2(new_n518), .ZN(new_n534));
  NOR3_X1   g348(.A1(new_n533), .A2(new_n534), .A3(KEYINPUT75), .ZN(new_n535));
  OAI211_X1 g349(.A(new_n262), .B(new_n532), .C1(new_n535), .C2(new_n522), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n255), .B1(G234), .B2(new_n262), .ZN(new_n537));
  AND3_X1   g351(.A1(new_n530), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n529), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT77), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n537), .A2(G902), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n541), .ZN(new_n543));
  OAI21_X1  g357(.A(KEYINPUT77), .B1(new_n529), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  OAI21_X1  g359(.A(KEYINPUT78), .B1(new_n538), .B2(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n530), .A2(new_n536), .A3(new_n537), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT78), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n547), .A2(new_n548), .A3(new_n544), .A4(new_n542), .ZN(new_n549));
  AOI22_X1  g363(.A1(new_n483), .A2(new_n493), .B1(new_n546), .B2(new_n549), .ZN(new_n550));
  XNOR2_X1  g364(.A(G110), .B(G140), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n188), .A2(G227), .ZN(new_n552));
  XNOR2_X1  g366(.A(new_n551), .B(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n332), .A2(new_n359), .A3(new_n296), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT85), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT84), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n301), .B1(new_n306), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n290), .A2(KEYINPUT1), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(KEYINPUT84), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(new_n292), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n370), .B1(new_n561), .B2(new_n300), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n555), .B1(new_n562), .B2(KEYINPUT10), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n298), .B1(new_n557), .B2(new_n559), .ZN(new_n564));
  INV_X1    g378(.A(new_n300), .ZN(new_n565));
  OAI211_X1 g379(.A(new_n326), .B(new_n369), .C1(new_n564), .C2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT10), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n566), .A2(KEYINPUT85), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n563), .A2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n449), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n378), .A2(KEYINPUT10), .A3(new_n308), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n554), .A2(new_n569), .A3(new_n570), .A4(new_n571), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n309), .B1(new_n376), .B2(new_n377), .ZN(new_n573));
  AOI22_X1  g387(.A1(new_n573), .A2(new_n566), .B1(new_n447), .B2(new_n448), .ZN(new_n574));
  OAI21_X1  g388(.A(KEYINPUT88), .B1(new_n574), .B2(KEYINPUT12), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n308), .B1(new_n372), .B2(new_n373), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n449), .B1(new_n576), .B2(new_n562), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT88), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT12), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  OAI211_X1 g394(.A(new_n449), .B(KEYINPUT12), .C1(new_n576), .C2(new_n562), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(KEYINPUT87), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n573), .A2(new_n566), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT87), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n583), .A2(new_n584), .A3(KEYINPUT12), .A4(new_n449), .ZN(new_n585));
  AOI22_X1  g399(.A1(new_n575), .A2(new_n580), .B1(new_n582), .B2(new_n585), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n572), .B1(new_n586), .B2(KEYINPUT89), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n575), .A2(new_n580), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n582), .A2(new_n585), .ZN(new_n589));
  AND3_X1   g403(.A1(new_n588), .A2(new_n589), .A3(KEYINPUT89), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n553), .B1(new_n587), .B2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(G469), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n554), .A2(new_n569), .A3(new_n571), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(new_n449), .ZN(new_n594));
  INV_X1    g408(.A(new_n553), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n594), .A2(new_n595), .A3(new_n572), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n591), .A2(new_n592), .A3(new_n262), .A4(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(G469), .A2(G902), .ZN(new_n598));
  INV_X1    g412(.A(new_n572), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n595), .B1(new_n586), .B2(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n594), .A2(new_n553), .A3(new_n572), .ZN(new_n601));
  AND2_X1   g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(G469), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n597), .A2(new_n598), .A3(new_n603), .ZN(new_n604));
  OAI21_X1  g418(.A(G221), .B1(new_n254), .B2(G902), .ZN(new_n605));
  XOR2_X1   g419(.A(new_n605), .B(KEYINPUT79), .Z(new_n606));
  AND2_X1   g420(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n422), .A2(new_n550), .A3(new_n607), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n608), .B(G101), .ZN(G3));
  NOR3_X1   g423(.A1(new_n390), .A2(new_n401), .A3(new_n289), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n420), .B1(new_n610), .B2(new_n418), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(KEYINPUT102), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n402), .A2(new_n415), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT102), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n613), .A2(new_n614), .A3(new_n420), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT33), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n260), .A2(new_n261), .A3(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n258), .A2(KEYINPUT33), .A3(new_n259), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n264), .A2(G902), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n617), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n263), .A2(new_n264), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  AND3_X1   g437(.A1(new_n282), .A2(new_n272), .A3(new_n225), .ZN(new_n624));
  NOR3_X1   g438(.A1(new_n623), .A2(new_n279), .A3(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n612), .A2(new_n615), .A3(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT103), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n612), .A2(KEYINPUT103), .A3(new_n615), .A4(new_n625), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n546), .A2(new_n549), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n262), .B1(new_n471), .B2(new_n475), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(G472), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n633), .A2(KEYINPUT101), .A3(new_n476), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT101), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n632), .A2(new_n635), .A3(G472), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n630), .A2(new_n631), .A3(new_n607), .A4(new_n637), .ZN(new_n638));
  XOR2_X1   g452(.A(KEYINPUT34), .B(G104), .Z(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G6));
  AOI21_X1  g454(.A(new_n614), .B1(new_n613), .B2(new_n420), .ZN(new_n641));
  INV_X1    g455(.A(new_n420), .ZN(new_n642));
  AOI211_X1 g456(.A(KEYINPUT102), .B(new_n642), .C1(new_n402), .C2(new_n415), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  XOR2_X1   g459(.A(new_n278), .B(KEYINPUT104), .Z(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n637), .A2(new_n631), .A3(new_n607), .A4(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n624), .A2(new_n284), .ZN(new_n649));
  NOR3_X1   g463(.A1(new_n645), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(KEYINPUT35), .B(G107), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G9));
  NOR2_X1   g466(.A1(new_n526), .A2(KEYINPUT36), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(new_n523), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(new_n541), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n547), .A2(new_n655), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n422), .A2(new_n607), .A3(new_n637), .A4(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(KEYINPUT37), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(new_n511), .ZN(G12));
  NAND2_X1  g473(.A1(new_n604), .A2(new_n606), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n660), .B1(new_n483), .B2(new_n493), .ZN(new_n661));
  OR2_X1    g475(.A1(new_n277), .A2(G900), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n283), .B1(new_n275), .B2(new_n662), .ZN(new_n663));
  AND2_X1   g477(.A1(new_n663), .A2(new_n284), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n644), .A2(new_n656), .A3(new_n661), .A4(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(G128), .ZN(G30));
  NAND2_X1  g480(.A1(new_n417), .A2(new_n419), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(KEYINPUT38), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n283), .A2(new_n284), .ZN(new_n669));
  OR2_X1    g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n662), .A2(new_n275), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(KEYINPUT39), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n607), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(KEYINPUT40), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT105), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n478), .A2(new_n427), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n459), .A2(new_n428), .A3(new_n488), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(new_n262), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n423), .B1(new_n676), .B2(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n675), .B1(new_n483), .B2(new_n681), .ZN(new_n682));
  AOI211_X1 g496(.A(KEYINPUT105), .B(new_n680), .C1(new_n477), .C2(new_n482), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(new_n656), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(new_n420), .ZN(new_n686));
  NOR4_X1   g500(.A1(new_n670), .A2(new_n674), .A3(new_n684), .A4(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(new_n238), .ZN(G45));
  AND3_X1   g502(.A1(new_n622), .A2(new_n283), .A3(new_n671), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n644), .A2(new_n656), .A3(new_n661), .A4(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G146), .ZN(G48));
  NAND3_X1  g505(.A1(new_n591), .A2(new_n262), .A3(new_n596), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(G469), .ZN(new_n693));
  AND3_X1   g507(.A1(new_n693), .A2(new_n605), .A3(new_n597), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n550), .A2(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  AOI21_X1  g510(.A(KEYINPUT103), .B1(new_n644), .B2(new_n625), .ZN(new_n697));
  INV_X1    g511(.A(new_n629), .ZN(new_n698));
  OAI21_X1  g512(.A(new_n696), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(KEYINPUT106), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT106), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n630), .A2(new_n701), .A3(new_n696), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(KEYINPUT41), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G113), .ZN(G15));
  NOR2_X1   g519(.A1(new_n645), .A2(new_n649), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n695), .A2(new_n646), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G116), .ZN(G18));
  NAND2_X1  g523(.A1(new_n483), .A2(new_n493), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(new_n694), .ZN(new_n712));
  NOR3_X1   g526(.A1(new_n711), .A2(new_n712), .A3(new_n287), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n612), .A2(new_n615), .A3(new_n656), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G119), .ZN(G21));
  NOR2_X1   g531(.A1(new_n645), .A2(new_n712), .ZN(new_n718));
  INV_X1    g532(.A(new_n669), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n470), .B1(new_n490), .B2(new_n427), .ZN(new_n720));
  OAI211_X1 g534(.A(new_n423), .B(new_n262), .C1(new_n720), .C2(new_n475), .ZN(new_n721));
  AND2_X1   g535(.A1(new_n633), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n538), .A2(new_n545), .ZN(new_n723));
  AND3_X1   g537(.A1(new_n722), .A2(new_n723), .A3(new_n647), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n718), .A2(new_n719), .A3(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G122), .ZN(G24));
  AND4_X1   g540(.A1(new_n633), .A2(new_n656), .A3(new_n689), .A4(new_n721), .ZN(new_n727));
  AND4_X1   g541(.A1(new_n615), .A2(new_n612), .A3(new_n727), .A4(new_n694), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(new_n208), .ZN(G27));
  AOI21_X1  g543(.A(new_n642), .B1(new_n417), .B2(new_n419), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n598), .B(KEYINPUT107), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT108), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n600), .A2(new_n732), .ZN(new_n733));
  OAI211_X1 g547(.A(KEYINPUT108), .B(new_n595), .C1(new_n586), .C2(new_n599), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n733), .A2(G469), .A3(new_n601), .A4(new_n734), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n597), .A2(new_n731), .A3(new_n735), .ZN(new_n736));
  AND2_X1   g550(.A1(new_n736), .A2(new_n605), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n550), .A2(new_n689), .A3(new_n730), .A4(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT42), .ZN(new_n739));
  AND3_X1   g553(.A1(new_n736), .A2(KEYINPUT42), .A3(new_n605), .ZN(new_n740));
  AND3_X1   g554(.A1(new_n730), .A2(new_n740), .A3(new_n689), .ZN(new_n741));
  AND2_X1   g555(.A1(new_n710), .A2(new_n723), .ZN(new_n742));
  AOI22_X1  g556(.A1(new_n738), .A2(new_n739), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(new_n193), .ZN(G33));
  AND4_X1   g558(.A1(new_n550), .A2(new_n664), .A3(new_n730), .A4(new_n737), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(new_n242), .ZN(G36));
  INV_X1    g560(.A(KEYINPUT109), .ZN(new_n747));
  AOI21_X1  g561(.A(KEYINPUT43), .B1(new_n624), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n624), .A2(new_n622), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n748), .B(new_n749), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n750), .A2(new_n636), .A3(new_n634), .A4(new_n656), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT44), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n730), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  XOR2_X1   g567(.A(new_n753), .B(KEYINPUT110), .Z(new_n754));
  NAND4_X1  g568(.A1(new_n733), .A2(KEYINPUT45), .A3(new_n601), .A4(new_n734), .ZN(new_n755));
  OAI211_X1 g569(.A(new_n755), .B(G469), .C1(KEYINPUT45), .C2(new_n602), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(new_n731), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT46), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n756), .A2(KEYINPUT46), .A3(new_n731), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n759), .A2(new_n597), .A3(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n761), .A2(new_n605), .A3(new_n672), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n762), .B1(new_n752), .B2(new_n751), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n754), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G137), .ZN(G39));
  NAND2_X1  g579(.A1(new_n761), .A2(new_n605), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT47), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n761), .A2(KEYINPUT47), .A3(new_n605), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(new_n730), .ZN(new_n771));
  INV_X1    g585(.A(new_n689), .ZN(new_n772));
  NOR3_X1   g586(.A1(new_n771), .A2(new_n631), .A3(new_n772), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n770), .A2(new_n711), .A3(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G140), .ZN(G42));
  NAND2_X1  g589(.A1(new_n693), .A2(new_n597), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(KEYINPUT111), .ZN(new_n777));
  XOR2_X1   g591(.A(new_n777), .B(KEYINPUT49), .Z(new_n778));
  AND4_X1   g592(.A1(new_n606), .A2(new_n778), .A3(new_n668), .A4(new_n684), .ZN(new_n779));
  INV_X1    g593(.A(new_n749), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n779), .A2(new_n723), .A3(new_n420), .A4(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n188), .A2(G952), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n771), .A2(new_n712), .ZN(new_n783));
  INV_X1    g597(.A(new_n275), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n783), .A2(new_n784), .A3(new_n750), .ZN(new_n785));
  INV_X1    g599(.A(new_n742), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  XOR2_X1   g601(.A(new_n787), .B(KEYINPUT119), .Z(new_n788));
  AOI21_X1  g602(.A(new_n782), .B1(new_n788), .B2(KEYINPUT48), .ZN(new_n789));
  AND4_X1   g603(.A1(new_n723), .A2(new_n750), .A3(new_n784), .A4(new_n722), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n790), .A2(new_n668), .A3(new_n642), .A4(new_n694), .ZN(new_n791));
  NOR2_X1   g605(.A1(KEYINPUT116), .A2(KEYINPUT50), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n791), .B(new_n792), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n777), .A2(new_n606), .ZN(new_n794));
  OAI211_X1 g608(.A(new_n730), .B(new_n790), .C1(new_n770), .C2(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n722), .A2(new_n656), .ZN(new_n796));
  OAI211_X1 g610(.A(new_n793), .B(new_n795), .C1(new_n796), .C2(new_n785), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n680), .B1(new_n477), .B2(new_n482), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(new_n675), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n799), .A2(new_n275), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT117), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n800), .A2(new_n801), .A3(new_n631), .A4(new_n783), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n684), .A2(new_n784), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n783), .A2(new_n631), .ZN(new_n804));
  OAI21_X1  g618(.A(KEYINPUT117), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n802), .A2(new_n805), .A3(new_n624), .A4(new_n623), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT118), .ZN(new_n807));
  OR2_X1    g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n806), .A2(new_n807), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n797), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n789), .B1(new_n810), .B2(KEYINPUT51), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT51), .ZN(new_n812));
  AOI211_X1 g626(.A(new_n812), .B(new_n797), .C1(new_n809), .C2(new_n808), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n685), .A2(new_n284), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n661), .A2(new_n663), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n727), .A2(new_n737), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n771), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NOR3_X1   g632(.A1(new_n743), .A2(new_n818), .A3(new_n745), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n710), .A2(new_n607), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n714), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n728), .B1(new_n821), .B2(new_n664), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT52), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n671), .B(KEYINPUT113), .ZN(new_n824));
  AOI21_X1  g638(.A(KEYINPUT114), .B1(new_n685), .B2(new_n824), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n547), .A2(KEYINPUT114), .A3(new_n655), .A4(new_n824), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n826), .A2(new_n736), .A3(new_n605), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n799), .A2(new_n644), .A3(new_n719), .A4(new_n828), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n822), .A2(new_n823), .A3(new_n829), .A4(new_n690), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n644), .A2(new_n694), .A3(new_n727), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n665), .A2(new_n690), .A3(new_n831), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n828), .B1(new_n682), .B2(new_n683), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n644), .A2(new_n719), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  OAI21_X1  g649(.A(KEYINPUT52), .B1(new_n832), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n657), .A2(new_n608), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n623), .A2(new_n624), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n838), .B1(new_n284), .B2(new_n624), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n648), .A2(new_n421), .A3(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT53), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n837), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n819), .A2(new_n830), .A3(new_n836), .A4(new_n842), .ZN(new_n843));
  AOI22_X1  g657(.A1(new_n706), .A2(new_n707), .B1(new_n715), .B2(new_n713), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n701), .B1(new_n630), .B2(new_n696), .ZN(new_n845));
  AOI211_X1 g659(.A(KEYINPUT106), .B(new_n695), .C1(new_n628), .C2(new_n629), .ZN(new_n846));
  OAI211_X1 g660(.A(new_n725), .B(new_n844), .C1(new_n845), .C2(new_n846), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n843), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n847), .A2(KEYINPUT112), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT112), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n703), .A2(new_n850), .A3(new_n725), .A4(new_n844), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n819), .A2(new_n830), .A3(new_n836), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n837), .A2(new_n840), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n849), .A2(new_n851), .A3(new_n852), .A4(new_n853), .ZN(new_n854));
  AOI211_X1 g668(.A(KEYINPUT54), .B(new_n848), .C1(new_n854), .C2(new_n841), .ZN(new_n855));
  INV_X1    g669(.A(new_n855), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n849), .A2(new_n851), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n857), .A2(KEYINPUT115), .A3(new_n852), .A4(new_n842), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT115), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n849), .A2(new_n851), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n859), .B1(new_n860), .B2(new_n843), .ZN(new_n861));
  AOI22_X1  g675(.A1(new_n858), .A2(new_n861), .B1(new_n841), .B2(new_n854), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT54), .ZN(new_n863));
  OAI211_X1 g677(.A(new_n814), .B(new_n856), .C1(new_n862), .C2(new_n863), .ZN(new_n864));
  OR3_X1    g678(.A1(new_n787), .A2(KEYINPUT119), .A3(KEYINPUT48), .ZN(new_n865));
  INV_X1    g679(.A(new_n865), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n802), .A2(new_n838), .A3(new_n805), .ZN(new_n867));
  AND2_X1   g681(.A1(new_n718), .A2(new_n790), .ZN(new_n868));
  NOR4_X1   g682(.A1(new_n864), .A2(new_n866), .A3(new_n867), .A4(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(G952), .A2(G953), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n781), .B1(new_n869), .B2(new_n870), .ZN(G75));
  AOI21_X1  g685(.A(new_n848), .B1(new_n854), .B2(new_n841), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n872), .A2(new_n262), .ZN(new_n873));
  AOI21_X1  g687(.A(KEYINPUT56), .B1(new_n873), .B2(G210), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n409), .B(new_n410), .ZN(new_n875));
  XOR2_X1   g689(.A(KEYINPUT120), .B(KEYINPUT55), .Z(new_n876));
  XNOR2_X1  g690(.A(new_n875), .B(new_n876), .ZN(new_n877));
  AND2_X1   g691(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n874), .A2(new_n877), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n188), .A2(G952), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(G51));
  XOR2_X1   g695(.A(new_n731), .B(KEYINPUT57), .Z(new_n882));
  NAND2_X1  g696(.A1(new_n854), .A2(new_n841), .ZN(new_n883));
  INV_X1    g697(.A(new_n848), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n863), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n882), .B1(new_n885), .B2(new_n855), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT121), .ZN(new_n887));
  AND2_X1   g701(.A1(new_n591), .A2(new_n596), .ZN(new_n888));
  AND3_X1   g702(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n887), .B1(new_n886), .B2(new_n888), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  OR3_X1    g705(.A1(new_n872), .A2(new_n262), .A3(new_n756), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n880), .B1(new_n891), .B2(new_n892), .ZN(G54));
  NAND3_X1  g707(.A1(new_n873), .A2(KEYINPUT58), .A3(G475), .ZN(new_n894));
  INV_X1    g708(.A(new_n222), .ZN(new_n895));
  AND2_X1   g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n894), .A2(new_n895), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n896), .A2(new_n897), .A3(new_n880), .ZN(G60));
  AND2_X1   g712(.A1(new_n617), .A2(new_n618), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n856), .B1(new_n862), .B2(new_n863), .ZN(new_n900));
  XNOR2_X1  g714(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n264), .A2(new_n262), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n901), .B(new_n902), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n899), .B1(new_n900), .B2(new_n903), .ZN(new_n904));
  OAI211_X1 g718(.A(new_n899), .B(new_n903), .C1(new_n885), .C2(new_n855), .ZN(new_n905));
  INV_X1    g719(.A(new_n905), .ZN(new_n906));
  NOR3_X1   g720(.A1(new_n904), .A2(new_n880), .A3(new_n906), .ZN(G63));
  INV_X1    g721(.A(KEYINPUT61), .ZN(new_n908));
  NAND2_X1  g722(.A1(G217), .A2(G902), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n909), .B(KEYINPUT60), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n872), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(new_n654), .ZN(new_n912));
  INV_X1    g726(.A(new_n880), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n529), .B1(new_n872), .B2(new_n910), .ZN(new_n915));
  INV_X1    g729(.A(new_n915), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n908), .B1(new_n914), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(KEYINPUT123), .ZN(new_n918));
  INV_X1    g732(.A(new_n914), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT124), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n908), .B1(new_n915), .B2(new_n920), .ZN(new_n921));
  OAI211_X1 g735(.A(new_n919), .B(new_n921), .C1(new_n920), .C2(new_n915), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT123), .ZN(new_n923));
  OAI211_X1 g737(.A(new_n923), .B(new_n908), .C1(new_n914), .C2(new_n916), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n918), .A2(new_n922), .A3(new_n924), .ZN(G66));
  AOI21_X1  g739(.A(new_n188), .B1(new_n276), .B2(G224), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n857), .A2(new_n853), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n926), .B1(new_n927), .B2(new_n188), .ZN(new_n928));
  OAI211_X1 g742(.A(new_n388), .B(new_n389), .C1(G898), .C2(new_n188), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n928), .B(new_n929), .Z(G69));
  XOR2_X1   g744(.A(new_n473), .B(new_n219), .Z(new_n931));
  NAND3_X1  g745(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n687), .A2(new_n832), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(KEYINPUT62), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n550), .A2(new_n730), .ZN(new_n935));
  NOR3_X1   g749(.A1(new_n935), .A2(new_n673), .A3(new_n839), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(KEYINPUT125), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n934), .A2(new_n764), .A3(new_n774), .A4(new_n937), .ZN(new_n938));
  OAI211_X1 g752(.A(new_n931), .B(new_n932), .C1(new_n938), .C2(G953), .ZN(new_n939));
  INV_X1    g753(.A(G900), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n940), .A2(new_n188), .A3(G227), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n931), .A2(new_n941), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n764), .A2(new_n690), .A3(new_n774), .A4(new_n822), .ZN(new_n943));
  NOR3_X1   g757(.A1(new_n762), .A2(new_n786), .A3(new_n834), .ZN(new_n944));
  NOR4_X1   g758(.A1(new_n943), .A2(new_n743), .A3(new_n745), .A4(new_n944), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n942), .B1(new_n945), .B2(G953), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n939), .A2(new_n946), .ZN(G72));
  NAND2_X1  g761(.A1(G472), .A2(G902), .ZN(new_n948));
  XOR2_X1   g762(.A(new_n948), .B(KEYINPUT63), .Z(new_n949));
  OAI21_X1  g763(.A(new_n949), .B1(new_n938), .B2(new_n927), .ZN(new_n950));
  INV_X1    g764(.A(new_n676), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT126), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n950), .A2(KEYINPUT126), .A3(new_n951), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n945), .A2(new_n853), .A3(new_n857), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n486), .B1(new_n957), .B2(new_n949), .ZN(new_n958));
  INV_X1    g772(.A(new_n486), .ZN(new_n959));
  INV_X1    g773(.A(new_n949), .ZN(new_n960));
  NOR4_X1   g774(.A1(new_n862), .A2(new_n959), .A3(new_n951), .A4(new_n960), .ZN(new_n961));
  NOR4_X1   g775(.A1(new_n956), .A2(new_n880), .A3(new_n958), .A4(new_n961), .ZN(G57));
endmodule


