

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581;

  XNOR2_X1 U323 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n373) );
  XNOR2_X1 U324 ( .A(n438), .B(n310), .ZN(n311) );
  XNOR2_X1 U325 ( .A(n312), .B(n311), .ZN(n320) );
  XNOR2_X1 U326 ( .A(KEYINPUT120), .B(KEYINPUT55), .ZN(n435) );
  XNOR2_X1 U327 ( .A(n374), .B(n373), .ZN(n537) );
  XNOR2_X1 U328 ( .A(KEYINPUT104), .B(KEYINPUT36), .ZN(n329) );
  XNOR2_X1 U329 ( .A(n436), .B(n435), .ZN(n451) );
  XNOR2_X1 U330 ( .A(n559), .B(n329), .ZN(n579) );
  XOR2_X1 U331 ( .A(n450), .B(n449), .Z(n517) );
  XNOR2_X1 U332 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U333 ( .A(n455), .B(n454), .ZN(G1349GAT) );
  XOR2_X1 U334 ( .A(G85GAT), .B(G92GAT), .Z(n309) );
  XOR2_X1 U335 ( .A(KEYINPUT32), .B(KEYINPUT33), .Z(n292) );
  XNOR2_X1 U336 ( .A(KEYINPUT72), .B(KEYINPUT31), .ZN(n291) );
  XNOR2_X1 U337 ( .A(n292), .B(n291), .ZN(n295) );
  XOR2_X1 U338 ( .A(G64GAT), .B(KEYINPUT71), .Z(n294) );
  XNOR2_X1 U339 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n293) );
  XNOR2_X1 U340 ( .A(n294), .B(n293), .ZN(n342) );
  XOR2_X1 U341 ( .A(n295), .B(n342), .Z(n301) );
  XOR2_X1 U342 ( .A(G71GAT), .B(G120GAT), .Z(n297) );
  XNOR2_X1 U343 ( .A(G99GAT), .B(G176GAT), .ZN(n296) );
  XNOR2_X1 U344 ( .A(n297), .B(n296), .ZN(n437) );
  XOR2_X1 U345 ( .A(G78GAT), .B(G148GAT), .Z(n299) );
  XNOR2_X1 U346 ( .A(G106GAT), .B(G204GAT), .ZN(n298) );
  XNOR2_X1 U347 ( .A(n299), .B(n298), .ZN(n427) );
  XNOR2_X1 U348 ( .A(n437), .B(n427), .ZN(n300) );
  XNOR2_X1 U349 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U350 ( .A(n309), .B(n302), .ZN(n304) );
  AND2_X1 U351 ( .A1(G230GAT), .A2(G233GAT), .ZN(n303) );
  XNOR2_X1 U352 ( .A(n304), .B(n303), .ZN(n569) );
  INV_X1 U353 ( .A(G162GAT), .ZN(n305) );
  NAND2_X1 U354 ( .A1(G50GAT), .A2(n305), .ZN(n308) );
  INV_X1 U355 ( .A(G50GAT), .ZN(n306) );
  NAND2_X1 U356 ( .A1(n306), .A2(G162GAT), .ZN(n307) );
  NAND2_X1 U357 ( .A1(n308), .A2(n307), .ZN(n422) );
  XNOR2_X1 U358 ( .A(n309), .B(n422), .ZN(n312) );
  XOR2_X1 U359 ( .A(G43GAT), .B(G134GAT), .Z(n438) );
  AND2_X1 U360 ( .A1(G232GAT), .A2(G233GAT), .ZN(n310) );
  XOR2_X1 U361 ( .A(KEYINPUT9), .B(KEYINPUT66), .Z(n314) );
  XNOR2_X1 U362 ( .A(KEYINPUT73), .B(KEYINPUT74), .ZN(n313) );
  XNOR2_X1 U363 ( .A(n314), .B(n313), .ZN(n318) );
  XOR2_X1 U364 ( .A(KEYINPUT75), .B(G106GAT), .Z(n316) );
  XNOR2_X1 U365 ( .A(G190GAT), .B(G99GAT), .ZN(n315) );
  XNOR2_X1 U366 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U367 ( .A(n318), .B(n317), .Z(n319) );
  XNOR2_X1 U368 ( .A(n320), .B(n319), .ZN(n324) );
  XOR2_X1 U369 ( .A(KEYINPUT77), .B(KEYINPUT11), .Z(n322) );
  XNOR2_X1 U370 ( .A(KEYINPUT10), .B(KEYINPUT67), .ZN(n321) );
  XNOR2_X1 U371 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U372 ( .A(n324), .B(n323), .ZN(n328) );
  XNOR2_X1 U373 ( .A(G29GAT), .B(KEYINPUT8), .ZN(n325) );
  XNOR2_X1 U374 ( .A(n325), .B(KEYINPUT7), .ZN(n351) );
  XNOR2_X1 U375 ( .A(G36GAT), .B(G218GAT), .ZN(n326) );
  XNOR2_X1 U376 ( .A(n326), .B(KEYINPUT76), .ZN(n378) );
  XOR2_X1 U377 ( .A(n351), .B(n378), .Z(n327) );
  XNOR2_X1 U378 ( .A(n328), .B(n327), .ZN(n559) );
  XOR2_X1 U379 ( .A(G15GAT), .B(G127GAT), .Z(n446) );
  XOR2_X1 U380 ( .A(G78GAT), .B(G211GAT), .Z(n331) );
  XNOR2_X1 U381 ( .A(G183GAT), .B(G155GAT), .ZN(n330) );
  XNOR2_X1 U382 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U383 ( .A(n446), .B(n332), .Z(n334) );
  NAND2_X1 U384 ( .A1(G231GAT), .A2(G233GAT), .ZN(n333) );
  XNOR2_X1 U385 ( .A(n334), .B(n333), .ZN(n346) );
  XOR2_X1 U386 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n336) );
  XNOR2_X1 U387 ( .A(KEYINPUT81), .B(KEYINPUT15), .ZN(n335) );
  XNOR2_X1 U388 ( .A(n336), .B(n335), .ZN(n340) );
  XOR2_X1 U389 ( .A(KEYINPUT79), .B(KEYINPUT80), .Z(n338) );
  XNOR2_X1 U390 ( .A(G71GAT), .B(KEYINPUT78), .ZN(n337) );
  XNOR2_X1 U391 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U392 ( .A(n340), .B(n339), .Z(n344) );
  XNOR2_X1 U393 ( .A(G22GAT), .B(G1GAT), .ZN(n341) );
  XNOR2_X1 U394 ( .A(n341), .B(G8GAT), .ZN(n355) );
  XNOR2_X1 U395 ( .A(n355), .B(n342), .ZN(n343) );
  XNOR2_X1 U396 ( .A(n344), .B(n343), .ZN(n345) );
  XNOR2_X1 U397 ( .A(n346), .B(n345), .ZN(n554) );
  NOR2_X1 U398 ( .A1(n579), .A2(n554), .ZN(n348) );
  XNOR2_X1 U399 ( .A(KEYINPUT45), .B(KEYINPUT114), .ZN(n347) );
  XNOR2_X1 U400 ( .A(n348), .B(n347), .ZN(n365) );
  XOR2_X1 U401 ( .A(KEYINPUT29), .B(KEYINPUT69), .Z(n354) );
  XOR2_X1 U402 ( .A(KEYINPUT70), .B(KEYINPUT30), .Z(n350) );
  XNOR2_X1 U403 ( .A(G15GAT), .B(G113GAT), .ZN(n349) );
  XNOR2_X1 U404 ( .A(n350), .B(n349), .ZN(n352) );
  XNOR2_X1 U405 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U406 ( .A(n354), .B(n353), .ZN(n359) );
  XOR2_X1 U407 ( .A(G43GAT), .B(n355), .Z(n357) );
  NAND2_X1 U408 ( .A1(G229GAT), .A2(G233GAT), .ZN(n356) );
  XNOR2_X1 U409 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U410 ( .A(n359), .B(n358), .Z(n364) );
  XOR2_X1 U411 ( .A(G141GAT), .B(G197GAT), .Z(n361) );
  XNOR2_X1 U412 ( .A(G169GAT), .B(G36GAT), .ZN(n360) );
  XNOR2_X1 U413 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U414 ( .A(n362), .B(G50GAT), .ZN(n363) );
  XOR2_X1 U415 ( .A(n364), .B(n363), .Z(n495) );
  INV_X1 U416 ( .A(n495), .ZN(n565) );
  NAND2_X1 U417 ( .A1(n365), .A2(n565), .ZN(n366) );
  NOR2_X1 U418 ( .A1(n569), .A2(n366), .ZN(n372) );
  INV_X1 U419 ( .A(n554), .ZN(n573) );
  XNOR2_X1 U420 ( .A(n569), .B(KEYINPUT41), .ZN(n542) );
  NOR2_X1 U421 ( .A1(n565), .A2(n542), .ZN(n367) );
  XNOR2_X1 U422 ( .A(n367), .B(KEYINPUT46), .ZN(n368) );
  NOR2_X1 U423 ( .A1(n573), .A2(n368), .ZN(n369) );
  NAND2_X1 U424 ( .A1(n559), .A2(n369), .ZN(n370) );
  XNOR2_X1 U425 ( .A(KEYINPUT47), .B(n370), .ZN(n371) );
  NOR2_X1 U426 ( .A1(n372), .A2(n371), .ZN(n374) );
  XOR2_X1 U427 ( .A(KEYINPUT98), .B(KEYINPUT97), .Z(n380) );
  XOR2_X1 U428 ( .A(KEYINPUT99), .B(G64GAT), .Z(n376) );
  XNOR2_X1 U429 ( .A(G8GAT), .B(G176GAT), .ZN(n375) );
  XNOR2_X1 U430 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U431 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U432 ( .A(n380), .B(n379), .ZN(n384) );
  XOR2_X1 U433 ( .A(G92GAT), .B(G204GAT), .Z(n382) );
  NAND2_X1 U434 ( .A1(G226GAT), .A2(G233GAT), .ZN(n381) );
  XNOR2_X1 U435 ( .A(n382), .B(n381), .ZN(n383) );
  XOR2_X1 U436 ( .A(n384), .B(n383), .Z(n392) );
  XNOR2_X1 U437 ( .A(G183GAT), .B(KEYINPUT18), .ZN(n385) );
  XNOR2_X1 U438 ( .A(n385), .B(KEYINPUT19), .ZN(n386) );
  XOR2_X1 U439 ( .A(n386), .B(KEYINPUT17), .Z(n388) );
  XNOR2_X1 U440 ( .A(G169GAT), .B(G190GAT), .ZN(n387) );
  XNOR2_X1 U441 ( .A(n388), .B(n387), .ZN(n450) );
  XOR2_X1 U442 ( .A(G211GAT), .B(KEYINPUT89), .Z(n390) );
  XNOR2_X1 U443 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n389) );
  XNOR2_X1 U444 ( .A(n390), .B(n389), .ZN(n429) );
  XNOR2_X1 U445 ( .A(n450), .B(n429), .ZN(n391) );
  XNOR2_X1 U446 ( .A(n392), .B(n391), .ZN(n514) );
  NOR2_X1 U447 ( .A1(n537), .A2(n514), .ZN(n393) );
  XNOR2_X1 U448 ( .A(n393), .B(KEYINPUT54), .ZN(n417) );
  XOR2_X1 U449 ( .A(KEYINPUT1), .B(KEYINPUT6), .Z(n395) );
  XNOR2_X1 U450 ( .A(G1GAT), .B(G57GAT), .ZN(n394) );
  XNOR2_X1 U451 ( .A(n395), .B(n394), .ZN(n399) );
  XOR2_X1 U452 ( .A(KEYINPUT96), .B(KEYINPUT4), .Z(n397) );
  XNOR2_X1 U453 ( .A(KEYINPUT93), .B(KEYINPUT5), .ZN(n396) );
  XNOR2_X1 U454 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U455 ( .A(n399), .B(n398), .Z(n404) );
  XOR2_X1 U456 ( .A(G113GAT), .B(KEYINPUT0), .Z(n445) );
  XOR2_X1 U457 ( .A(KEYINPUT95), .B(KEYINPUT94), .Z(n401) );
  NAND2_X1 U458 ( .A1(G225GAT), .A2(G233GAT), .ZN(n400) );
  XNOR2_X1 U459 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U460 ( .A(n445), .B(n402), .ZN(n403) );
  XNOR2_X1 U461 ( .A(n404), .B(n403), .ZN(n408) );
  XOR2_X1 U462 ( .A(KEYINPUT75), .B(G162GAT), .Z(n406) );
  XNOR2_X1 U463 ( .A(G29GAT), .B(G134GAT), .ZN(n405) );
  XNOR2_X1 U464 ( .A(n406), .B(n405), .ZN(n407) );
  XOR2_X1 U465 ( .A(n408), .B(n407), .Z(n416) );
  XOR2_X1 U466 ( .A(KEYINPUT2), .B(KEYINPUT90), .Z(n410) );
  XNOR2_X1 U467 ( .A(KEYINPUT3), .B(G155GAT), .ZN(n409) );
  XNOR2_X1 U468 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U469 ( .A(G141GAT), .B(n411), .Z(n430) );
  XOR2_X1 U470 ( .A(G85GAT), .B(G148GAT), .Z(n413) );
  XNOR2_X1 U471 ( .A(G127GAT), .B(G120GAT), .ZN(n412) );
  XNOR2_X1 U472 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U473 ( .A(n430), .B(n414), .ZN(n415) );
  XNOR2_X1 U474 ( .A(n416), .B(n415), .ZN(n511) );
  NAND2_X1 U475 ( .A1(n417), .A2(n511), .ZN(n418) );
  XNOR2_X1 U476 ( .A(n418), .B(KEYINPUT65), .ZN(n562) );
  XOR2_X1 U477 ( .A(KEYINPUT22), .B(KEYINPUT24), .Z(n420) );
  XNOR2_X1 U478 ( .A(G218GAT), .B(KEYINPUT88), .ZN(n419) );
  XNOR2_X1 U479 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U480 ( .A(n422), .B(n421), .Z(n424) );
  NAND2_X1 U481 ( .A1(G228GAT), .A2(G233GAT), .ZN(n423) );
  XNOR2_X1 U482 ( .A(n424), .B(n423), .ZN(n434) );
  XOR2_X1 U483 ( .A(KEYINPUT23), .B(KEYINPUT92), .Z(n426) );
  XNOR2_X1 U484 ( .A(G22GAT), .B(KEYINPUT91), .ZN(n425) );
  XNOR2_X1 U485 ( .A(n426), .B(n425), .ZN(n428) );
  XOR2_X1 U486 ( .A(n428), .B(n427), .Z(n432) );
  XNOR2_X1 U487 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U488 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U489 ( .A(n434), .B(n433), .ZN(n465) );
  NAND2_X1 U490 ( .A1(n562), .A2(n465), .ZN(n436) );
  XOR2_X1 U491 ( .A(n438), .B(n437), .Z(n440) );
  NAND2_X1 U492 ( .A1(G227GAT), .A2(G233GAT), .ZN(n439) );
  XNOR2_X1 U493 ( .A(n440), .B(n439), .ZN(n444) );
  XOR2_X1 U494 ( .A(KEYINPUT86), .B(KEYINPUT84), .Z(n442) );
  XNOR2_X1 U495 ( .A(KEYINPUT85), .B(KEYINPUT20), .ZN(n441) );
  XNOR2_X1 U496 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U497 ( .A(n444), .B(n443), .Z(n448) );
  XNOR2_X1 U498 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U499 ( .A(n448), .B(n447), .ZN(n449) );
  INV_X1 U500 ( .A(n517), .ZN(n525) );
  NAND2_X1 U501 ( .A1(n451), .A2(n525), .ZN(n558) );
  XOR2_X1 U502 ( .A(KEYINPUT105), .B(n542), .Z(n528) );
  NOR2_X1 U503 ( .A1(n558), .A2(n528), .ZN(n455) );
  XNOR2_X1 U504 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n453) );
  XNOR2_X1 U505 ( .A(G176GAT), .B(KEYINPUT122), .ZN(n452) );
  NOR2_X1 U506 ( .A1(n565), .A2(n569), .ZN(n486) );
  NAND2_X1 U507 ( .A1(n559), .A2(n573), .ZN(n458) );
  XNOR2_X1 U508 ( .A(KEYINPUT82), .B(KEYINPUT16), .ZN(n456) );
  XNOR2_X1 U509 ( .A(n456), .B(KEYINPUT83), .ZN(n457) );
  XNOR2_X1 U510 ( .A(n458), .B(n457), .ZN(n473) );
  XNOR2_X1 U511 ( .A(n514), .B(KEYINPUT27), .ZN(n467) );
  NOR2_X1 U512 ( .A1(n511), .A2(n467), .ZN(n539) );
  XNOR2_X1 U513 ( .A(KEYINPUT28), .B(KEYINPUT68), .ZN(n459) );
  XNOR2_X1 U514 ( .A(n459), .B(n465), .ZN(n520) );
  NAND2_X1 U515 ( .A1(n539), .A2(n520), .ZN(n524) );
  XNOR2_X1 U516 ( .A(KEYINPUT87), .B(n517), .ZN(n460) );
  NOR2_X1 U517 ( .A1(n524), .A2(n460), .ZN(n461) );
  XOR2_X1 U518 ( .A(KEYINPUT100), .B(n461), .Z(n472) );
  OR2_X1 U519 ( .A1(n517), .A2(n514), .ZN(n462) );
  NAND2_X1 U520 ( .A1(n462), .A2(n465), .ZN(n463) );
  XNOR2_X1 U521 ( .A(n463), .B(KEYINPUT101), .ZN(n464) );
  XNOR2_X1 U522 ( .A(n464), .B(KEYINPUT25), .ZN(n469) );
  NOR2_X1 U523 ( .A1(n465), .A2(n525), .ZN(n466) );
  XOR2_X1 U524 ( .A(n466), .B(KEYINPUT26), .Z(n563) );
  OR2_X1 U525 ( .A1(n467), .A2(n563), .ZN(n468) );
  NAND2_X1 U526 ( .A1(n469), .A2(n468), .ZN(n470) );
  NAND2_X1 U527 ( .A1(n511), .A2(n470), .ZN(n471) );
  NAND2_X1 U528 ( .A1(n472), .A2(n471), .ZN(n484) );
  AND2_X1 U529 ( .A1(n473), .A2(n484), .ZN(n496) );
  NAND2_X1 U530 ( .A1(n486), .A2(n496), .ZN(n480) );
  NOR2_X1 U531 ( .A1(n511), .A2(n480), .ZN(n474) );
  XOR2_X1 U532 ( .A(n474), .B(KEYINPUT34), .Z(n475) );
  XNOR2_X1 U533 ( .A(G1GAT), .B(n475), .ZN(G1324GAT) );
  NOR2_X1 U534 ( .A1(n514), .A2(n480), .ZN(n476) );
  XOR2_X1 U535 ( .A(G8GAT), .B(n476), .Z(G1325GAT) );
  NOR2_X1 U536 ( .A1(n517), .A2(n480), .ZN(n478) );
  XNOR2_X1 U537 ( .A(KEYINPUT35), .B(KEYINPUT102), .ZN(n477) );
  XNOR2_X1 U538 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U539 ( .A(G15GAT), .B(n479), .ZN(G1326GAT) );
  NOR2_X1 U540 ( .A1(n520), .A2(n480), .ZN(n482) );
  XNOR2_X1 U541 ( .A(G22GAT), .B(KEYINPUT103), .ZN(n481) );
  XNOR2_X1 U542 ( .A(n482), .B(n481), .ZN(G1327GAT) );
  NOR2_X1 U543 ( .A1(n579), .A2(n573), .ZN(n483) );
  NAND2_X1 U544 ( .A1(n484), .A2(n483), .ZN(n485) );
  XNOR2_X1 U545 ( .A(KEYINPUT37), .B(n485), .ZN(n510) );
  NAND2_X1 U546 ( .A1(n510), .A2(n486), .ZN(n487) );
  XNOR2_X1 U547 ( .A(KEYINPUT38), .B(n487), .ZN(n493) );
  NOR2_X1 U548 ( .A1(n511), .A2(n493), .ZN(n488) );
  XNOR2_X1 U549 ( .A(n488), .B(KEYINPUT39), .ZN(n489) );
  XNOR2_X1 U550 ( .A(G29GAT), .B(n489), .ZN(G1328GAT) );
  NOR2_X1 U551 ( .A1(n514), .A2(n493), .ZN(n490) );
  XOR2_X1 U552 ( .A(G36GAT), .B(n490), .Z(G1329GAT) );
  NOR2_X1 U553 ( .A1(n517), .A2(n493), .ZN(n491) );
  XOR2_X1 U554 ( .A(n491), .B(KEYINPUT40), .Z(n492) );
  XNOR2_X1 U555 ( .A(G43GAT), .B(n492), .ZN(G1330GAT) );
  NOR2_X1 U556 ( .A1(n493), .A2(n520), .ZN(n494) );
  XOR2_X1 U557 ( .A(G50GAT), .B(n494), .Z(G1331GAT) );
  NOR2_X1 U558 ( .A1(n495), .A2(n528), .ZN(n509) );
  AND2_X1 U559 ( .A1(n509), .A2(n496), .ZN(n497) );
  XOR2_X1 U560 ( .A(KEYINPUT106), .B(n497), .Z(n505) );
  NOR2_X1 U561 ( .A1(n511), .A2(n505), .ZN(n498) );
  XOR2_X1 U562 ( .A(KEYINPUT42), .B(n498), .Z(n499) );
  XNOR2_X1 U563 ( .A(G57GAT), .B(n499), .ZN(G1332GAT) );
  XNOR2_X1 U564 ( .A(G64GAT), .B(KEYINPUT107), .ZN(n501) );
  NOR2_X1 U565 ( .A1(n514), .A2(n505), .ZN(n500) );
  XNOR2_X1 U566 ( .A(n501), .B(n500), .ZN(G1333GAT) );
  XNOR2_X1 U567 ( .A(KEYINPUT108), .B(KEYINPUT109), .ZN(n503) );
  NOR2_X1 U568 ( .A1(n517), .A2(n505), .ZN(n502) );
  XNOR2_X1 U569 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U570 ( .A(G71GAT), .B(n504), .ZN(G1334GAT) );
  NOR2_X1 U571 ( .A1(n505), .A2(n520), .ZN(n507) );
  XNOR2_X1 U572 ( .A(KEYINPUT43), .B(KEYINPUT110), .ZN(n506) );
  XNOR2_X1 U573 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U574 ( .A(G78GAT), .B(n508), .ZN(G1335GAT) );
  NAND2_X1 U575 ( .A1(n510), .A2(n509), .ZN(n519) );
  NOR2_X1 U576 ( .A1(n511), .A2(n519), .ZN(n513) );
  XNOR2_X1 U577 ( .A(G85GAT), .B(KEYINPUT111), .ZN(n512) );
  XNOR2_X1 U578 ( .A(n513), .B(n512), .ZN(G1336GAT) );
  NOR2_X1 U579 ( .A1(n514), .A2(n519), .ZN(n515) );
  XOR2_X1 U580 ( .A(KEYINPUT112), .B(n515), .Z(n516) );
  XNOR2_X1 U581 ( .A(G92GAT), .B(n516), .ZN(G1337GAT) );
  NOR2_X1 U582 ( .A1(n517), .A2(n519), .ZN(n518) );
  XOR2_X1 U583 ( .A(G99GAT), .B(n518), .Z(G1338GAT) );
  NOR2_X1 U584 ( .A1(n520), .A2(n519), .ZN(n522) );
  XNOR2_X1 U585 ( .A(KEYINPUT44), .B(KEYINPUT113), .ZN(n521) );
  XNOR2_X1 U586 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U587 ( .A(G106GAT), .B(n523), .ZN(G1339GAT) );
  NOR2_X1 U588 ( .A1(n537), .A2(n524), .ZN(n526) );
  NAND2_X1 U589 ( .A1(n526), .A2(n525), .ZN(n533) );
  NOR2_X1 U590 ( .A1(n565), .A2(n533), .ZN(n527) );
  XOR2_X1 U591 ( .A(G113GAT), .B(n527), .Z(G1340GAT) );
  NOR2_X1 U592 ( .A1(n528), .A2(n533), .ZN(n530) );
  XNOR2_X1 U593 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n529) );
  XNOR2_X1 U594 ( .A(n530), .B(n529), .ZN(G1341GAT) );
  NOR2_X1 U595 ( .A1(n554), .A2(n533), .ZN(n531) );
  XOR2_X1 U596 ( .A(KEYINPUT50), .B(n531), .Z(n532) );
  XNOR2_X1 U597 ( .A(G127GAT), .B(n532), .ZN(G1342GAT) );
  NOR2_X1 U598 ( .A1(n559), .A2(n533), .ZN(n535) );
  XNOR2_X1 U599 ( .A(KEYINPUT51), .B(KEYINPUT115), .ZN(n534) );
  XNOR2_X1 U600 ( .A(n535), .B(n534), .ZN(n536) );
  XOR2_X1 U601 ( .A(G134GAT), .B(n536), .Z(G1343GAT) );
  NOR2_X1 U602 ( .A1(n537), .A2(n563), .ZN(n538) );
  NAND2_X1 U603 ( .A1(n539), .A2(n538), .ZN(n549) );
  NOR2_X1 U604 ( .A1(n565), .A2(n549), .ZN(n540) );
  XOR2_X1 U605 ( .A(G141GAT), .B(n540), .Z(n541) );
  XNOR2_X1 U606 ( .A(KEYINPUT116), .B(n541), .ZN(G1344GAT) );
  NOR2_X1 U607 ( .A1(n542), .A2(n549), .ZN(n544) );
  XNOR2_X1 U608 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n543) );
  XNOR2_X1 U609 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U610 ( .A(G148GAT), .B(n545), .ZN(G1345GAT) );
  NOR2_X1 U611 ( .A1(n554), .A2(n549), .ZN(n547) );
  XNOR2_X1 U612 ( .A(KEYINPUT117), .B(KEYINPUT118), .ZN(n546) );
  XNOR2_X1 U613 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U614 ( .A(G155GAT), .B(n548), .ZN(G1346GAT) );
  NOR2_X1 U615 ( .A1(n559), .A2(n549), .ZN(n551) );
  XNOR2_X1 U616 ( .A(G162GAT), .B(KEYINPUT119), .ZN(n550) );
  XNOR2_X1 U617 ( .A(n551), .B(n550), .ZN(G1347GAT) );
  NOR2_X1 U618 ( .A1(n565), .A2(n558), .ZN(n553) );
  XNOR2_X1 U619 ( .A(G169GAT), .B(KEYINPUT121), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n553), .B(n552), .ZN(G1348GAT) );
  NOR2_X1 U621 ( .A1(n554), .A2(n558), .ZN(n555) );
  XOR2_X1 U622 ( .A(G183GAT), .B(n555), .Z(G1350GAT) );
  XOR2_X1 U623 ( .A(KEYINPUT123), .B(KEYINPUT58), .Z(n557) );
  XNOR2_X1 U624 ( .A(G190GAT), .B(KEYINPUT124), .ZN(n556) );
  XNOR2_X1 U625 ( .A(n557), .B(n556), .ZN(n561) );
  NOR2_X1 U626 ( .A1(n559), .A2(n558), .ZN(n560) );
  XOR2_X1 U627 ( .A(n561), .B(n560), .Z(G1351GAT) );
  INV_X1 U628 ( .A(n563), .ZN(n564) );
  NAND2_X1 U629 ( .A1(n562), .A2(n564), .ZN(n578) );
  NOR2_X1 U630 ( .A1(n565), .A2(n578), .ZN(n567) );
  XNOR2_X1 U631 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U633 ( .A(G197GAT), .B(n568), .ZN(G1352GAT) );
  XOR2_X1 U634 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n571) );
  INV_X1 U635 ( .A(n578), .ZN(n574) );
  NAND2_X1 U636 ( .A1(n574), .A2(n569), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(n572) );
  XOR2_X1 U638 ( .A(G204GAT), .B(n572), .Z(G1353GAT) );
  NAND2_X1 U639 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n575), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U641 ( .A(KEYINPUT62), .B(KEYINPUT126), .Z(n577) );
  XNOR2_X1 U642 ( .A(G218GAT), .B(KEYINPUT127), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(n581) );
  NOR2_X1 U644 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U645 ( .A(n581), .B(n580), .Z(G1355GAT) );
endmodule

