

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763;

  NOR2_X1 U368 ( .A1(G953), .A2(G237), .ZN(n485) );
  XNOR2_X1 U369 ( .A(n415), .B(n395), .ZN(n470) );
  INV_X1 U370 ( .A(G953), .ZN(n751) );
  INV_X1 U371 ( .A(n660), .ZN(n663) );
  XNOR2_X1 U372 ( .A(n597), .B(n596), .ZN(n761) );
  OR2_X1 U373 ( .A1(n728), .A2(G902), .ZN(n346) );
  INV_X2 U374 ( .A(n716), .ZN(n727) );
  NOR2_X2 U375 ( .A1(n601), .A2(n368), .ZN(n591) );
  NOR2_X1 U376 ( .A1(n584), .A2(n434), .ZN(n435) );
  INV_X4 U377 ( .A(G116), .ZN(n488) );
  XNOR2_X1 U378 ( .A(n371), .B(n513), .ZN(n762) );
  NOR2_X1 U379 ( .A1(n512), .A2(n355), .ZN(n379) );
  XNOR2_X1 U380 ( .A(n435), .B(n357), .ZN(n520) );
  XNOR2_X1 U381 ( .A(n741), .B(n401), .ZN(n637) );
  XNOR2_X1 U382 ( .A(n373), .B(n420), .ZN(n481) );
  XNOR2_X1 U383 ( .A(G128), .B(KEYINPUT78), .ZN(n415) );
  XNOR2_X1 U384 ( .A(KEYINPUT74), .B(KEYINPUT16), .ZN(n419) );
  AND2_X1 U385 ( .A1(n556), .A2(n548), .ZN(n347) );
  NOR2_X1 U386 ( .A1(n360), .A2(n348), .ZN(n405) );
  NOR2_X1 U387 ( .A1(n762), .A2(KEYINPUT44), .ZN(n370) );
  INV_X1 U388 ( .A(n679), .ZN(n543) );
  NOR2_X1 U389 ( .A1(n688), .A2(n689), .ZN(n685) );
  NAND2_X1 U390 ( .A1(n351), .A2(n370), .ZN(n554) );
  NAND2_X1 U391 ( .A1(n546), .A2(n380), .ZN(n547) );
  XNOR2_X1 U392 ( .A(n450), .B(n390), .ZN(n748) );
  INV_X1 U393 ( .A(KEYINPUT10), .ZN(n390) );
  XNOR2_X1 U394 ( .A(G125), .B(G140), .ZN(n450) );
  XNOR2_X1 U395 ( .A(n374), .B(G110), .ZN(n373) );
  XNOR2_X1 U396 ( .A(G107), .B(G104), .ZN(n374) );
  INV_X1 U397 ( .A(G143), .ZN(n395) );
  XNOR2_X1 U398 ( .A(G125), .B(KEYINPUT18), .ZN(n412) );
  XNOR2_X1 U399 ( .A(n394), .B(G146), .ZN(n476) );
  INV_X1 U400 ( .A(KEYINPUT4), .ZN(n394) );
  NAND2_X1 U401 ( .A1(n677), .A2(n356), .ZN(n366) );
  XNOR2_X1 U402 ( .A(n426), .B(n425), .ZN(n673) );
  XNOR2_X1 U403 ( .A(n386), .B(n354), .ZN(n689) );
  OR2_X1 U404 ( .A1(n733), .A2(G902), .ZN(n386) );
  XNOR2_X1 U405 ( .A(n749), .B(n495), .ZN(n626) );
  XNOR2_X1 U406 ( .A(n499), .B(n500), .ZN(n389) );
  XOR2_X1 U407 ( .A(KEYINPUT70), .B(KEYINPUT24), .Z(n499) );
  XNOR2_X1 U408 ( .A(n498), .B(KEYINPUT23), .ZN(n388) );
  XNOR2_X1 U409 ( .A(G119), .B(G110), .ZN(n498) );
  XNOR2_X1 U410 ( .A(n748), .B(G146), .ZN(n501) );
  XNOR2_X1 U411 ( .A(n379), .B(n378), .ZN(n360) );
  INV_X1 U412 ( .A(KEYINPUT66), .ZN(n378) );
  INV_X1 U413 ( .A(n689), .ZN(n568) );
  XNOR2_X1 U414 ( .A(G113), .B(G104), .ZN(n440) );
  INV_X1 U415 ( .A(KEYINPUT77), .ZN(n409) );
  XNOR2_X1 U416 ( .A(KEYINPUT15), .B(G902), .ZN(n611) );
  XNOR2_X1 U417 ( .A(n473), .B(KEYINPUT67), .ZN(n474) );
  XOR2_X1 U418 ( .A(KEYINPUT93), .B(KEYINPUT5), .Z(n487) );
  XNOR2_X1 U419 ( .A(G101), .B(KEYINPUT92), .ZN(n489) );
  INV_X1 U420 ( .A(KEYINPUT48), .ZN(n603) );
  AND2_X1 U421 ( .A1(n384), .A2(n383), .ZN(n382) );
  XNOR2_X1 U422 ( .A(n376), .B(G113), .ZN(n492) );
  XNOR2_X1 U423 ( .A(KEYINPUT3), .B(G119), .ZN(n376) );
  XOR2_X1 U424 ( .A(KEYINPUT76), .B(G140), .Z(n479) );
  XNOR2_X1 U425 ( .A(n476), .B(n392), .ZN(n391) );
  XNOR2_X1 U426 ( .A(n393), .B(G131), .ZN(n392) );
  INV_X1 U427 ( .A(G137), .ZN(n393) );
  INV_X1 U428 ( .A(KEYINPUT38), .ZN(n369) );
  AND2_X1 U429 ( .A1(n689), .A2(n385), .ZN(n578) );
  INV_X1 U430 ( .A(n688), .ZN(n385) );
  XNOR2_X1 U431 ( .A(G107), .B(KEYINPUT7), .ZN(n460) );
  NAND2_X1 U432 ( .A1(G234), .A2(G237), .ZN(n430) );
  XNOR2_X1 U433 ( .A(n519), .B(n518), .ZN(n683) );
  NAND2_X2 U434 ( .A1(n365), .A2(n363), .ZN(n700) );
  NAND2_X1 U435 ( .A1(n364), .A2(n349), .ZN(n363) );
  AND2_X1 U436 ( .A1(n367), .A2(n366), .ZN(n365) );
  NOR2_X1 U437 ( .A1(n588), .A2(n580), .ZN(n399) );
  XNOR2_X1 U438 ( .A(n398), .B(n397), .ZN(n396) );
  INV_X1 U439 ( .A(KEYINPUT30), .ZN(n397) );
  XNOR2_X1 U440 ( .A(n428), .B(n427), .ZN(n584) );
  XNOR2_X1 U441 ( .A(n501), .B(n387), .ZN(n504) );
  XNOR2_X1 U442 ( .A(n389), .B(n388), .ZN(n387) );
  BUF_X1 U443 ( .A(n727), .Z(n731) );
  XNOR2_X1 U444 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U445 ( .A(KEYINPUT36), .B(KEYINPUT113), .ZN(n575) );
  NAND2_X1 U446 ( .A1(n372), .A2(n352), .ZN(n371) );
  XNOR2_X1 U447 ( .A(n536), .B(KEYINPUT31), .ZN(n666) );
  NAND2_X1 U448 ( .A1(n535), .A2(n534), .ZN(n536) );
  INV_X1 U449 ( .A(n540), .ZN(n534) );
  NAND2_X1 U450 ( .A1(n404), .A2(n403), .ZN(n634) );
  NOR2_X1 U451 ( .A1(n405), .A2(n350), .ZN(n404) );
  NAND2_X1 U452 ( .A1(n381), .A2(n568), .ZN(n380) );
  XNOR2_X1 U453 ( .A(n545), .B(n544), .ZN(n381) );
  NOR2_X1 U454 ( .A1(n630), .A2(n735), .ZN(n632) );
  OR2_X1 U455 ( .A1(n568), .A2(KEYINPUT106), .ZN(n348) );
  NOR2_X1 U456 ( .A1(n677), .A2(n356), .ZN(n349) );
  AND2_X1 U457 ( .A1(n568), .A2(KEYINPUT106), .ZN(n350) );
  XOR2_X1 U458 ( .A(n551), .B(n550), .Z(n351) );
  AND2_X1 U459 ( .A1(n511), .A2(n567), .ZN(n352) );
  XNOR2_X1 U460 ( .A(n594), .B(KEYINPUT110), .ZN(n678) );
  OR2_X1 U461 ( .A1(n666), .A2(n653), .ZN(n353) );
  XOR2_X1 U462 ( .A(n508), .B(n507), .Z(n354) );
  NAND2_X1 U463 ( .A1(n497), .A2(n606), .ZN(n355) );
  XOR2_X1 U464 ( .A(KEYINPUT111), .B(KEYINPUT41), .Z(n356) );
  XNOR2_X1 U465 ( .A(n593), .B(n592), .ZN(n763) );
  XOR2_X1 U466 ( .A(KEYINPUT85), .B(KEYINPUT0), .Z(n357) );
  NAND2_X1 U467 ( .A1(n615), .A2(KEYINPUT2), .ZN(n358) );
  XNOR2_X1 U468 ( .A(n475), .B(n474), .ZN(n359) );
  XNOR2_X1 U469 ( .A(n475), .B(n474), .ZN(n512) );
  INV_X1 U470 ( .A(G116), .ZN(n402) );
  NAND2_X1 U471 ( .A1(n360), .A2(KEYINPUT106), .ZN(n403) );
  NAND2_X1 U472 ( .A1(n637), .A2(n611), .ZN(n400) );
  AND2_X2 U473 ( .A1(n382), .A2(n361), .ZN(n604) );
  XNOR2_X1 U474 ( .A(n362), .B(KEYINPUT46), .ZN(n361) );
  NOR2_X1 U475 ( .A1(n761), .A2(n763), .ZN(n362) );
  NAND2_X1 U476 ( .A1(n595), .A2(n700), .ZN(n597) );
  INV_X1 U477 ( .A(n678), .ZN(n364) );
  NAND2_X1 U478 ( .A1(n678), .A2(n356), .ZN(n367) );
  INV_X1 U479 ( .A(n674), .ZN(n368) );
  XNOR2_X2 U480 ( .A(n599), .B(n369), .ZN(n674) );
  INV_X1 U481 ( .A(n359), .ZN(n372) );
  XNOR2_X2 U482 ( .A(n375), .B(n481), .ZN(n741) );
  XNOR2_X2 U483 ( .A(n377), .B(n492), .ZN(n375) );
  XNOR2_X2 U484 ( .A(n461), .B(n419), .ZN(n377) );
  XNOR2_X2 U485 ( .A(n488), .B(G122), .ZN(n461) );
  INV_X1 U486 ( .A(n380), .ZN(n651) );
  XNOR2_X1 U487 ( .A(n586), .B(KEYINPUT47), .ZN(n383) );
  NOR2_X1 U488 ( .A1(n668), .A2(n760), .ZN(n384) );
  XNOR2_X2 U489 ( .A(n477), .B(n391), .ZN(n749) );
  XNOR2_X2 U490 ( .A(n470), .B(G134), .ZN(n477) );
  NAND2_X1 U491 ( .A1(n399), .A2(n396), .ZN(n601) );
  NAND2_X1 U492 ( .A1(n587), .A2(n673), .ZN(n398) );
  XNOR2_X2 U493 ( .A(n400), .B(n423), .ZN(n574) );
  XNOR2_X1 U494 ( .A(n417), .B(n418), .ZN(n401) );
  NAND2_X1 U495 ( .A1(n406), .A2(n528), .ZN(n527) );
  NAND2_X1 U496 ( .A1(n634), .A2(n514), .ZN(n406) );
  NOR2_X1 U497 ( .A1(n359), .A2(n484), .ZN(n407) );
  NAND2_X1 U498 ( .A1(n407), .A2(n567), .ZN(n545) );
  BUF_X1 U499 ( .A(n621), .Z(n736) );
  XNOR2_X1 U500 ( .A(n558), .B(n557), .ZN(n621) );
  XNOR2_X1 U501 ( .A(KEYINPUT35), .B(KEYINPUT69), .ZN(n550) );
  INV_X1 U502 ( .A(KEYINPUT11), .ZN(n442) );
  XNOR2_X1 U503 ( .A(n489), .B(n402), .ZN(n490) );
  XNOR2_X1 U504 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U505 ( .A(n491), .B(n490), .ZN(n494) );
  XNOR2_X1 U506 ( .A(n445), .B(n444), .ZN(n449) );
  XNOR2_X1 U507 ( .A(n517), .B(KEYINPUT33), .ZN(n518) );
  XNOR2_X1 U508 ( .A(n461), .B(n460), .ZN(n465) );
  NOR2_X1 U509 ( .A1(n716), .A2(n624), .ZN(n628) );
  INV_X1 U510 ( .A(KEYINPUT63), .ZN(n631) );
  INV_X1 U511 ( .A(KEYINPUT17), .ZN(n408) );
  NAND2_X1 U512 ( .A1(KEYINPUT77), .A2(n408), .ZN(n411) );
  NAND2_X1 U513 ( .A1(n409), .A2(KEYINPUT17), .ZN(n410) );
  NAND2_X1 U514 ( .A1(n411), .A2(n410), .ZN(n413) );
  XNOR2_X1 U515 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U516 ( .A(n414), .B(n476), .ZN(n418) );
  AND2_X1 U517 ( .A1(G224), .A2(n751), .ZN(n416) );
  XNOR2_X1 U518 ( .A(n470), .B(n416), .ZN(n417) );
  XNOR2_X1 U519 ( .A(G101), .B(KEYINPUT87), .ZN(n420) );
  OR2_X1 U520 ( .A1(G237), .A2(G902), .ZN(n424) );
  NAND2_X1 U521 ( .A1(n424), .A2(G210), .ZN(n422) );
  XNOR2_X1 U522 ( .A(KEYINPUT79), .B(KEYINPUT88), .ZN(n421) );
  XNOR2_X1 U523 ( .A(n422), .B(n421), .ZN(n423) );
  NAND2_X1 U524 ( .A1(n424), .A2(G214), .ZN(n426) );
  INV_X1 U525 ( .A(KEYINPUT89), .ZN(n425) );
  NAND2_X1 U526 ( .A1(n574), .A2(n673), .ZN(n428) );
  INV_X1 U527 ( .A(KEYINPUT19), .ZN(n427) );
  INV_X1 U528 ( .A(KEYINPUT14), .ZN(n429) );
  XNOR2_X1 U529 ( .A(n430), .B(n429), .ZN(n706) );
  INV_X1 U530 ( .A(n706), .ZN(n561) );
  NAND2_X1 U531 ( .A1(G953), .A2(G902), .ZN(n559) );
  NOR2_X1 U532 ( .A1(G898), .A2(n559), .ZN(n432) );
  NAND2_X1 U533 ( .A1(G952), .A2(n751), .ZN(n563) );
  INV_X1 U534 ( .A(n563), .ZN(n431) );
  OR2_X1 U535 ( .A1(n432), .A2(n431), .ZN(n433) );
  NAND2_X1 U536 ( .A1(n561), .A2(n433), .ZN(n434) );
  NAND2_X1 U537 ( .A1(n611), .A2(G234), .ZN(n437) );
  XNOR2_X1 U538 ( .A(KEYINPUT90), .B(KEYINPUT20), .ZN(n436) );
  XNOR2_X1 U539 ( .A(n437), .B(n436), .ZN(n505) );
  AND2_X1 U540 ( .A1(n505), .A2(G221), .ZN(n439) );
  INV_X1 U541 ( .A(KEYINPUT21), .ZN(n438) );
  XNOR2_X1 U542 ( .A(n439), .B(n438), .ZN(n688) );
  XNOR2_X1 U543 ( .A(KEYINPUT13), .B(G475), .ZN(n459) );
  INV_X1 U544 ( .A(G902), .ZN(n457) );
  XOR2_X1 U545 ( .A(KEYINPUT12), .B(G122), .Z(n441) );
  XNOR2_X1 U546 ( .A(n441), .B(n440), .ZN(n445) );
  XNOR2_X1 U547 ( .A(G131), .B(G143), .ZN(n443) );
  XOR2_X1 U548 ( .A(KEYINPUT96), .B(KEYINPUT95), .Z(n447) );
  NAND2_X1 U549 ( .A1(G214), .A2(n485), .ZN(n446) );
  XNOR2_X1 U550 ( .A(n447), .B(n446), .ZN(n448) );
  XOR2_X1 U551 ( .A(n449), .B(n448), .Z(n455) );
  XOR2_X1 U552 ( .A(KEYINPUT100), .B(KEYINPUT97), .Z(n452) );
  XNOR2_X1 U553 ( .A(KEYINPUT99), .B(KEYINPUT98), .ZN(n451) );
  XNOR2_X1 U554 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U555 ( .A(n501), .B(n453), .ZN(n454) );
  XNOR2_X1 U556 ( .A(n455), .B(n454), .ZN(n645) );
  INV_X1 U557 ( .A(n645), .ZN(n456) );
  NAND2_X1 U558 ( .A1(n457), .A2(n456), .ZN(n458) );
  XNOR2_X1 U559 ( .A(n459), .B(n458), .ZN(n542) );
  XOR2_X1 U560 ( .A(KEYINPUT102), .B(KEYINPUT9), .Z(n463) );
  XNOR2_X1 U561 ( .A(KEYINPUT101), .B(KEYINPUT103), .ZN(n462) );
  XNOR2_X1 U562 ( .A(n463), .B(n462), .ZN(n464) );
  XOR2_X1 U563 ( .A(n465), .B(n464), .Z(n469) );
  XOR2_X1 U564 ( .A(KEYINPUT82), .B(KEYINPUT8), .Z(n467) );
  NAND2_X1 U565 ( .A1(G234), .A2(n751), .ZN(n466) );
  XNOR2_X1 U566 ( .A(n467), .B(n466), .ZN(n502) );
  NAND2_X1 U567 ( .A1(G217), .A2(n502), .ZN(n468) );
  XNOR2_X1 U568 ( .A(n469), .B(n468), .ZN(n471) );
  XNOR2_X1 U569 ( .A(n471), .B(n477), .ZN(n728) );
  XNOR2_X1 U570 ( .A(G478), .B(n346), .ZN(n541) );
  INV_X1 U571 ( .A(n541), .ZN(n515) );
  NAND2_X1 U572 ( .A1(n542), .A2(n515), .ZN(n677) );
  NOR2_X1 U573 ( .A1(n688), .A2(n677), .ZN(n472) );
  NAND2_X1 U574 ( .A1(n520), .A2(n472), .ZN(n475) );
  XNOR2_X1 U575 ( .A(KEYINPUT73), .B(KEYINPUT22), .ZN(n473) );
  NAND2_X1 U576 ( .A1(G227), .A2(n751), .ZN(n478) );
  XNOR2_X1 U577 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U578 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U579 ( .A(n749), .B(n482), .ZN(n721) );
  OR2_X1 U580 ( .A1(n721), .A2(G902), .ZN(n483) );
  INV_X1 U581 ( .A(G469), .ZN(n717) );
  XNOR2_X2 U582 ( .A(n483), .B(n717), .ZN(n582) );
  XNOR2_X2 U583 ( .A(n582), .B(KEYINPUT1), .ZN(n606) );
  INV_X1 U584 ( .A(n606), .ZN(n484) );
  NAND2_X1 U585 ( .A1(n485), .A2(G210), .ZN(n486) );
  XNOR2_X1 U586 ( .A(n487), .B(n486), .ZN(n491) );
  INV_X1 U587 ( .A(n492), .ZN(n493) );
  XNOR2_X1 U588 ( .A(n494), .B(n493), .ZN(n495) );
  NAND2_X1 U589 ( .A1(n626), .A2(n457), .ZN(n496) );
  INV_X1 U590 ( .A(G472), .ZN(n624) );
  XNOR2_X1 U591 ( .A(n496), .B(n624), .ZN(n509) );
  XNOR2_X1 U592 ( .A(n509), .B(KEYINPUT105), .ZN(n587) );
  INV_X1 U593 ( .A(n587), .ZN(n497) );
  XNOR2_X1 U594 ( .A(G128), .B(G137), .ZN(n500) );
  NAND2_X1 U595 ( .A1(G221), .A2(n502), .ZN(n503) );
  XNOR2_X1 U596 ( .A(n504), .B(n503), .ZN(n733) );
  NAND2_X1 U597 ( .A1(G217), .A2(n505), .ZN(n508) );
  XOR2_X1 U598 ( .A(KEYINPUT25), .B(KEYINPUT75), .Z(n506) );
  XNOR2_X1 U599 ( .A(n506), .B(KEYINPUT91), .ZN(n507) );
  NOR2_X1 U600 ( .A1(n606), .A2(n568), .ZN(n511) );
  BUF_X1 U601 ( .A(n509), .Z(n695) );
  INV_X1 U602 ( .A(KEYINPUT6), .ZN(n510) );
  XNOR2_X1 U603 ( .A(n695), .B(n510), .ZN(n567) );
  INV_X1 U604 ( .A(KEYINPUT32), .ZN(n513) );
  NOR2_X1 U605 ( .A1(n762), .A2(KEYINPUT69), .ZN(n514) );
  INV_X1 U606 ( .A(KEYINPUT65), .ZN(n528) );
  INV_X1 U607 ( .A(KEYINPUT35), .ZN(n525) );
  NOR2_X1 U608 ( .A1(n542), .A2(n515), .ZN(n598) );
  INV_X1 U609 ( .A(n598), .ZN(n524) );
  INV_X1 U610 ( .A(n606), .ZN(n516) );
  NAND2_X1 U611 ( .A1(n516), .A2(n685), .ZN(n532) );
  NOR2_X1 U612 ( .A1(n532), .A2(n567), .ZN(n519) );
  XNOR2_X1 U613 ( .A(KEYINPUT71), .B(KEYINPUT107), .ZN(n517) );
  INV_X1 U614 ( .A(n520), .ZN(n540) );
  NOR2_X1 U615 ( .A1(n683), .A2(n540), .ZN(n522) );
  XOR2_X1 U616 ( .A(KEYINPUT72), .B(KEYINPUT34), .Z(n521) );
  XNOR2_X1 U617 ( .A(n522), .B(n521), .ZN(n523) );
  NOR2_X2 U618 ( .A1(n524), .A2(n523), .ZN(n551) );
  XNOR2_X1 U619 ( .A(n525), .B(n551), .ZN(n759) );
  INV_X1 U620 ( .A(KEYINPUT44), .ZN(n529) );
  NOR2_X1 U621 ( .A1(n759), .A2(n529), .ZN(n526) );
  NAND2_X1 U622 ( .A1(n527), .A2(n526), .ZN(n531) );
  NAND2_X1 U623 ( .A1(n529), .A2(n528), .ZN(n530) );
  NAND2_X1 U624 ( .A1(n531), .A2(n530), .ZN(n549) );
  OR2_X1 U625 ( .A1(n532), .A2(n695), .ZN(n533) );
  XNOR2_X1 U626 ( .A(n533), .B(KEYINPUT94), .ZN(n698) );
  INV_X1 U627 ( .A(n698), .ZN(n535) );
  INV_X1 U628 ( .A(n582), .ZN(n537) );
  NAND2_X1 U629 ( .A1(n537), .A2(n685), .ZN(n588) );
  INV_X1 U630 ( .A(n588), .ZN(n538) );
  NAND2_X1 U631 ( .A1(n538), .A2(n695), .ZN(n539) );
  NOR2_X1 U632 ( .A1(n540), .A2(n539), .ZN(n653) );
  OR2_X1 U633 ( .A1(n542), .A2(n541), .ZN(n660) );
  AND2_X1 U634 ( .A1(n542), .A2(n541), .ZN(n665) );
  NOR2_X1 U635 ( .A1(n663), .A2(n665), .ZN(n679) );
  NAND2_X1 U636 ( .A1(n353), .A2(n543), .ZN(n546) );
  INV_X1 U637 ( .A(KEYINPUT84), .ZN(n544) );
  XOR2_X1 U638 ( .A(n547), .B(KEYINPUT104), .Z(n548) );
  INV_X1 U639 ( .A(n762), .ZN(n552) );
  NAND2_X1 U640 ( .A1(n552), .A2(KEYINPUT65), .ZN(n553) );
  NAND2_X1 U641 ( .A1(n554), .A2(n553), .ZN(n555) );
  NAND2_X1 U642 ( .A1(n555), .A2(n634), .ZN(n556) );
  NAND2_X1 U643 ( .A1(n347), .A2(n549), .ZN(n558) );
  INV_X1 U644 ( .A(KEYINPUT45), .ZN(n557) );
  NOR2_X1 U645 ( .A1(G900), .A2(n559), .ZN(n560) );
  NAND2_X1 U646 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U647 ( .A(KEYINPUT108), .B(n562), .Z(n565) );
  NOR2_X1 U648 ( .A1(n706), .A2(n563), .ZN(n564) );
  NOR2_X1 U649 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U650 ( .A(KEYINPUT80), .B(n566), .ZN(n580) );
  INV_X1 U651 ( .A(n580), .ZN(n589) );
  INV_X1 U652 ( .A(n673), .ZN(n572) );
  INV_X1 U653 ( .A(n567), .ZN(n570) );
  AND2_X1 U654 ( .A1(n663), .A2(n578), .ZN(n569) );
  NAND2_X1 U655 ( .A1(n570), .A2(n569), .ZN(n571) );
  NOR2_X1 U656 ( .A1(n572), .A2(n571), .ZN(n573) );
  NAND2_X1 U657 ( .A1(n589), .A2(n573), .ZN(n607) );
  BUF_X2 U658 ( .A(n574), .Z(n599) );
  INV_X1 U659 ( .A(n599), .ZN(n609) );
  NOR2_X1 U660 ( .A1(n607), .A2(n609), .ZN(n576) );
  NOR2_X1 U661 ( .A1(n577), .A2(n606), .ZN(n668) );
  NAND2_X1 U662 ( .A1(n578), .A2(n587), .ZN(n579) );
  NOR2_X1 U663 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U664 ( .A(KEYINPUT28), .B(n581), .Z(n583) );
  NOR2_X1 U665 ( .A1(n583), .A2(n582), .ZN(n595) );
  INV_X1 U666 ( .A(n584), .ZN(n585) );
  NAND2_X1 U667 ( .A1(n595), .A2(n585), .ZN(n661) );
  NOR2_X1 U668 ( .A1(n661), .A2(n679), .ZN(n586) );
  INV_X1 U669 ( .A(KEYINPUT39), .ZN(n590) );
  XNOR2_X1 U670 ( .A(n591), .B(n590), .ZN(n605) );
  NAND2_X1 U671 ( .A1(n605), .A2(n663), .ZN(n593) );
  INV_X1 U672 ( .A(KEYINPUT40), .ZN(n592) );
  NAND2_X1 U673 ( .A1(n674), .A2(n673), .ZN(n594) );
  XOR2_X1 U674 ( .A(KEYINPUT112), .B(KEYINPUT42), .Z(n596) );
  NAND2_X1 U675 ( .A1(n599), .A2(n598), .ZN(n600) );
  OR2_X1 U676 ( .A1(n601), .A2(n600), .ZN(n602) );
  XNOR2_X1 U677 ( .A(KEYINPUT109), .B(n602), .ZN(n760) );
  XNOR2_X1 U678 ( .A(n604), .B(n603), .ZN(n618) );
  NAND2_X1 U679 ( .A1(n605), .A2(n665), .ZN(n671) );
  NOR2_X1 U680 ( .A1(n484), .A2(n607), .ZN(n608) );
  XOR2_X1 U681 ( .A(n608), .B(KEYINPUT43), .Z(n610) );
  NAND2_X1 U682 ( .A1(n610), .A2(n609), .ZN(n633) );
  AND2_X1 U683 ( .A1(n671), .A2(n633), .ZN(n619) );
  INV_X1 U684 ( .A(n611), .ZN(n615) );
  NAND2_X1 U685 ( .A1(n619), .A2(n615), .ZN(n612) );
  OR2_X2 U686 ( .A1(n618), .A2(n612), .ZN(n613) );
  NOR2_X1 U687 ( .A1(n621), .A2(n613), .ZN(n614) );
  INV_X1 U688 ( .A(n614), .ZN(n616) );
  NAND2_X1 U689 ( .A1(n616), .A2(n358), .ZN(n617) );
  XNOR2_X1 U690 ( .A(n617), .B(KEYINPUT64), .ZN(n623) );
  INV_X1 U691 ( .A(n618), .ZN(n620) );
  NAND2_X1 U692 ( .A1(n620), .A2(n619), .ZN(n750) );
  NOR2_X1 U693 ( .A1(n750), .A2(n736), .ZN(n710) );
  NAND2_X1 U694 ( .A1(n710), .A2(KEYINPUT2), .ZN(n622) );
  NAND2_X1 U695 ( .A1(n623), .A2(n622), .ZN(n716) );
  XNOR2_X1 U696 ( .A(KEYINPUT114), .B(KEYINPUT62), .ZN(n625) );
  XNOR2_X1 U697 ( .A(n626), .B(n625), .ZN(n627) );
  XNOR2_X1 U698 ( .A(n628), .B(n627), .ZN(n630) );
  INV_X1 U699 ( .A(G952), .ZN(n629) );
  AND2_X1 U700 ( .A1(n629), .A2(G953), .ZN(n735) );
  XNOR2_X1 U701 ( .A(n632), .B(n631), .ZN(G57) );
  XNOR2_X1 U702 ( .A(n633), .B(G140), .ZN(G42) );
  XNOR2_X1 U703 ( .A(G110), .B(KEYINPUT115), .ZN(n635) );
  XOR2_X1 U704 ( .A(n635), .B(n634), .Z(G12) );
  NAND2_X1 U705 ( .A1(n727), .A2(G210), .ZN(n639) );
  XNOR2_X1 U706 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n636) );
  XNOR2_X1 U707 ( .A(n637), .B(n636), .ZN(n638) );
  XNOR2_X1 U708 ( .A(n639), .B(n638), .ZN(n640) );
  NOR2_X2 U709 ( .A1(n640), .A2(n735), .ZN(n642) );
  XOR2_X1 U710 ( .A(KEYINPUT83), .B(KEYINPUT56), .Z(n641) );
  XNOR2_X1 U711 ( .A(n642), .B(n641), .ZN(G51) );
  NAND2_X1 U712 ( .A1(n727), .A2(G475), .ZN(n647) );
  XNOR2_X1 U713 ( .A(KEYINPUT86), .B(KEYINPUT125), .ZN(n643) );
  XNOR2_X1 U714 ( .A(n643), .B(KEYINPUT59), .ZN(n644) );
  XNOR2_X1 U715 ( .A(n645), .B(n644), .ZN(n646) );
  XNOR2_X1 U716 ( .A(n647), .B(n646), .ZN(n648) );
  NOR2_X2 U717 ( .A1(n648), .A2(n735), .ZN(n650) );
  XNOR2_X1 U718 ( .A(KEYINPUT68), .B(KEYINPUT60), .ZN(n649) );
  XNOR2_X1 U719 ( .A(n650), .B(n649), .ZN(G60) );
  XOR2_X1 U720 ( .A(G101), .B(n651), .Z(G3) );
  NAND2_X1 U721 ( .A1(n653), .A2(n663), .ZN(n652) );
  XNOR2_X1 U722 ( .A(n652), .B(G104), .ZN(G6) );
  XOR2_X1 U723 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n655) );
  NAND2_X1 U724 ( .A1(n653), .A2(n665), .ZN(n654) );
  XNOR2_X1 U725 ( .A(n655), .B(n654), .ZN(n656) );
  XNOR2_X1 U726 ( .A(G107), .B(n656), .ZN(G9) );
  INV_X1 U727 ( .A(n665), .ZN(n657) );
  NOR2_X1 U728 ( .A1(n661), .A2(n657), .ZN(n659) );
  XNOR2_X1 U729 ( .A(G128), .B(KEYINPUT29), .ZN(n658) );
  XNOR2_X1 U730 ( .A(n659), .B(n658), .ZN(G30) );
  NOR2_X1 U731 ( .A1(n661), .A2(n660), .ZN(n662) );
  XOR2_X1 U732 ( .A(G146), .B(n662), .Z(G48) );
  NAND2_X1 U733 ( .A1(n666), .A2(n663), .ZN(n664) );
  XNOR2_X1 U734 ( .A(n664), .B(G113), .ZN(G15) );
  NAND2_X1 U735 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U736 ( .A(n667), .B(G116), .ZN(G18) );
  XNOR2_X1 U737 ( .A(n668), .B(KEYINPUT116), .ZN(n669) );
  XNOR2_X1 U738 ( .A(n669), .B(KEYINPUT37), .ZN(n670) );
  XNOR2_X1 U739 ( .A(G125), .B(n670), .ZN(G27) );
  XNOR2_X1 U740 ( .A(G134), .B(n671), .ZN(G36) );
  INV_X1 U741 ( .A(n683), .ZN(n672) );
  NAND2_X1 U742 ( .A1(n672), .A2(n700), .ZN(n709) );
  NOR2_X1 U743 ( .A1(n674), .A2(n673), .ZN(n675) );
  XNOR2_X1 U744 ( .A(n675), .B(KEYINPUT120), .ZN(n676) );
  NOR2_X1 U745 ( .A1(n677), .A2(n676), .ZN(n681) );
  NOR2_X1 U746 ( .A1(n679), .A2(n678), .ZN(n680) );
  NOR2_X1 U747 ( .A1(n681), .A2(n680), .ZN(n682) );
  NOR2_X1 U748 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X1 U749 ( .A(n684), .B(KEYINPUT121), .ZN(n703) );
  NOR2_X1 U750 ( .A1(n685), .A2(n484), .ZN(n686) );
  XOR2_X1 U751 ( .A(KEYINPUT50), .B(n686), .Z(n687) );
  XNOR2_X1 U752 ( .A(KEYINPUT119), .B(n687), .ZN(n694) );
  XOR2_X1 U753 ( .A(KEYINPUT118), .B(KEYINPUT117), .Z(n691) );
  NAND2_X1 U754 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U755 ( .A(n691), .B(n690), .ZN(n692) );
  XNOR2_X1 U756 ( .A(KEYINPUT49), .B(n692), .ZN(n693) );
  NOR2_X1 U757 ( .A1(n694), .A2(n693), .ZN(n696) );
  NAND2_X1 U758 ( .A1(n696), .A2(n695), .ZN(n697) );
  NAND2_X1 U759 ( .A1(n698), .A2(n697), .ZN(n699) );
  XOR2_X1 U760 ( .A(KEYINPUT51), .B(n699), .Z(n701) );
  NAND2_X1 U761 ( .A1(n701), .A2(n700), .ZN(n702) );
  NAND2_X1 U762 ( .A1(n703), .A2(n702), .ZN(n704) );
  XOR2_X1 U763 ( .A(KEYINPUT52), .B(n704), .Z(n705) );
  NOR2_X1 U764 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U765 ( .A1(n707), .A2(G952), .ZN(n708) );
  NAND2_X1 U766 ( .A1(n709), .A2(n708), .ZN(n713) );
  NOR2_X1 U767 ( .A1(n710), .A2(KEYINPUT81), .ZN(n711) );
  XNOR2_X1 U768 ( .A(n711), .B(KEYINPUT2), .ZN(n712) );
  NOR2_X1 U769 ( .A1(n713), .A2(n712), .ZN(n714) );
  NAND2_X1 U770 ( .A1(n751), .A2(n714), .ZN(n715) );
  XOR2_X1 U771 ( .A(KEYINPUT53), .B(n715), .Z(G75) );
  BUF_X1 U772 ( .A(n716), .Z(n718) );
  NOR2_X1 U773 ( .A1(n718), .A2(n717), .ZN(n725) );
  XNOR2_X1 U774 ( .A(KEYINPUT123), .B(KEYINPUT124), .ZN(n719) );
  XNOR2_X1 U775 ( .A(n719), .B(KEYINPUT122), .ZN(n720) );
  XOR2_X1 U776 ( .A(n720), .B(KEYINPUT57), .Z(n723) );
  XNOR2_X1 U777 ( .A(n721), .B(KEYINPUT58), .ZN(n722) );
  XNOR2_X1 U778 ( .A(n723), .B(n722), .ZN(n724) );
  XNOR2_X1 U779 ( .A(n725), .B(n724), .ZN(n726) );
  NOR2_X1 U780 ( .A1(n735), .A2(n726), .ZN(G54) );
  NAND2_X1 U781 ( .A1(n731), .A2(G478), .ZN(n729) );
  XNOR2_X1 U782 ( .A(n729), .B(n728), .ZN(n730) );
  NOR2_X1 U783 ( .A1(n735), .A2(n730), .ZN(G63) );
  NAND2_X1 U784 ( .A1(n731), .A2(G217), .ZN(n732) );
  XNOR2_X1 U785 ( .A(n733), .B(n732), .ZN(n734) );
  NOR2_X1 U786 ( .A1(n735), .A2(n734), .ZN(G66) );
  NOR2_X1 U787 ( .A1(n736), .A2(G953), .ZN(n740) );
  INV_X1 U788 ( .A(G898), .ZN(n742) );
  NAND2_X1 U789 ( .A1(G953), .A2(G224), .ZN(n737) );
  XOR2_X1 U790 ( .A(KEYINPUT61), .B(n737), .Z(n738) );
  NOR2_X1 U791 ( .A1(n742), .A2(n738), .ZN(n739) );
  NOR2_X1 U792 ( .A1(n740), .A2(n739), .ZN(n747) );
  INV_X1 U793 ( .A(n741), .ZN(n744) );
  NAND2_X1 U794 ( .A1(n742), .A2(G953), .ZN(n743) );
  NAND2_X1 U795 ( .A1(n744), .A2(n743), .ZN(n745) );
  XNOR2_X1 U796 ( .A(n745), .B(KEYINPUT126), .ZN(n746) );
  XNOR2_X1 U797 ( .A(n747), .B(n746), .ZN(G69) );
  XOR2_X1 U798 ( .A(n749), .B(n748), .Z(n753) );
  XNOR2_X1 U799 ( .A(n750), .B(n753), .ZN(n752) );
  NAND2_X1 U800 ( .A1(n752), .A2(n751), .ZN(n758) );
  XNOR2_X1 U801 ( .A(G227), .B(n753), .ZN(n754) );
  NAND2_X1 U802 ( .A1(n754), .A2(G900), .ZN(n755) );
  NAND2_X1 U803 ( .A1(G953), .A2(n755), .ZN(n756) );
  XOR2_X1 U804 ( .A(KEYINPUT127), .B(n756), .Z(n757) );
  NAND2_X1 U805 ( .A1(n758), .A2(n757), .ZN(G72) );
  XOR2_X1 U806 ( .A(G122), .B(n759), .Z(G24) );
  XOR2_X1 U807 ( .A(G143), .B(n760), .Z(G45) );
  XOR2_X1 U808 ( .A(n761), .B(G137), .Z(G39) );
  XOR2_X1 U809 ( .A(G119), .B(n762), .Z(G21) );
  XOR2_X1 U810 ( .A(G131), .B(n763), .Z(G33) );
endmodule

