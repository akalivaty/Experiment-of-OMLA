

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n792, n793, n794, n795,
         n796, n797, n798;

  AND2_X1 U375 ( .A1(n661), .A2(n660), .ZN(n372) );
  XNOR2_X1 U376 ( .A(n721), .B(KEYINPUT77), .ZN(n659) );
  NOR2_X1 U377 ( .A1(n362), .A2(n363), .ZN(n382) );
  XNOR2_X1 U378 ( .A(n644), .B(n643), .ZN(n797) );
  INV_X1 U379 ( .A(KEYINPUT85), .ZN(n357) );
  XNOR2_X1 U380 ( .A(n365), .B(KEYINPUT75), .ZN(n631) );
  BUF_X1 U381 ( .A(n727), .Z(n355) );
  XNOR2_X1 U382 ( .A(n364), .B(n354), .ZN(n624) );
  XNOR2_X1 U383 ( .A(n557), .B(KEYINPUT1), .ZN(n727) );
  INV_X1 U384 ( .A(KEYINPUT108), .ZN(n354) );
  XNOR2_X1 U385 ( .A(n352), .B(n499), .ZN(n726) );
  NAND2_X1 U386 ( .A1(n609), .A2(n571), .ZN(n352) );
  XNOR2_X1 U387 ( .A(n469), .B(G134), .ZN(n502) );
  BUF_X2 U388 ( .A(G128), .Z(n361) );
  NOR2_X1 U389 ( .A1(G953), .A2(G237), .ZN(n511) );
  XNOR2_X2 U390 ( .A(n495), .B(n494), .ZN(n581) );
  OR2_X2 U391 ( .A1(n600), .A2(n599), .ZN(n737) );
  NAND2_X1 U392 ( .A1(n353), .A2(n649), .ZN(n652) );
  NAND2_X1 U393 ( .A1(n418), .A2(n419), .ZN(n353) );
  AND2_X1 U394 ( .A1(n624), .A2(n623), .ZN(n707) );
  XNOR2_X2 U395 ( .A(n524), .B(n523), .ZN(n599) );
  NAND2_X1 U396 ( .A1(n373), .A2(n356), .ZN(n435) );
  NAND2_X1 U397 ( .A1(n358), .A2(n357), .ZN(n356) );
  INV_X1 U398 ( .A(n796), .ZN(n358) );
  AND2_X1 U399 ( .A1(n797), .A2(n645), .ZN(n648) );
  XNOR2_X1 U400 ( .A(G131), .B(G143), .ZN(n462) );
  AND2_X1 U401 ( .A1(n428), .A2(n638), .ZN(n359) );
  NAND2_X2 U402 ( .A1(n417), .A2(n415), .ZN(n414) );
  NOR2_X1 U403 ( .A1(n742), .A2(n605), .ZN(n589) );
  OR2_X1 U404 ( .A1(n577), .A2(n576), .ZN(n578) );
  NAND2_X1 U405 ( .A1(n394), .A2(n390), .ZN(n623) );
  AND2_X1 U406 ( .A1(n398), .A2(n395), .ZN(n394) );
  XNOR2_X1 U407 ( .A(n447), .B(n446), .ZN(n771) );
  XNOR2_X1 U408 ( .A(n518), .B(n471), .ZN(n447) );
  XNOR2_X1 U409 ( .A(n441), .B(G146), .ZN(n459) );
  INV_X1 U410 ( .A(G125), .ZN(n441) );
  NAND2_X1 U411 ( .A1(n416), .A2(KEYINPUT83), .ZN(n415) );
  INV_X1 U412 ( .A(n725), .ZN(n413) );
  NOR2_X1 U413 ( .A1(n666), .A2(n720), .ZN(n725) );
  NAND2_X1 U414 ( .A1(n617), .A2(n619), .ZN(n620) );
  AND2_X1 U415 ( .A1(n618), .A2(KEYINPUT65), .ZN(n619) );
  XNOR2_X1 U416 ( .A(n589), .B(KEYINPUT34), .ZN(n592) );
  NOR2_X1 U417 ( .A1(n737), .A2(n602), .ZN(n604) );
  AND2_X1 U418 ( .A1(n629), .A2(n377), .ZN(n630) );
  XNOR2_X1 U419 ( .A(n459), .B(n440), .ZN(n490) );
  XNOR2_X1 U420 ( .A(KEYINPUT16), .B(G110), .ZN(n445) );
  AND2_X1 U421 ( .A1(n414), .A2(n413), .ZN(n360) );
  AND2_X2 U422 ( .A1(n414), .A2(n413), .ZN(n686) );
  AND2_X1 U423 ( .A1(n796), .A2(KEYINPUT85), .ZN(n362) );
  NAND2_X1 U424 ( .A1(n616), .A2(n620), .ZN(n363) );
  NAND2_X1 U425 ( .A1(n543), .A2(n542), .ZN(n364) );
  NAND2_X1 U426 ( .A1(n707), .A2(n630), .ZN(n365) );
  NOR2_X1 U427 ( .A1(n695), .A2(G902), .ZN(n510) );
  XNOR2_X1 U428 ( .A(n783), .B(G146), .ZN(n366) );
  XNOR2_X1 U429 ( .A(n521), .B(n508), .ZN(n695) );
  XNOR2_X1 U430 ( .A(n783), .B(G146), .ZN(n521) );
  INV_X1 U431 ( .A(n582), .ZN(n367) );
  XNOR2_X1 U432 ( .A(n491), .B(n784), .ZN(n368) );
  XNOR2_X1 U433 ( .A(n491), .B(n784), .ZN(n687) );
  XNOR2_X2 U434 ( .A(n502), .B(n501), .ZN(n783) );
  XNOR2_X2 U435 ( .A(n489), .B(n488), .ZN(n491) );
  NAND2_X1 U436 ( .A1(n621), .A2(n382), .ZN(n622) );
  AND2_X1 U437 ( .A1(n716), .A2(n427), .ZN(n424) );
  NAND2_X1 U438 ( .A1(n384), .A2(KEYINPUT74), .ZN(n427) );
  AND2_X1 U439 ( .A1(n641), .A2(n653), .ZN(n746) );
  INV_X1 U440 ( .A(G902), .ZN(n522) );
  XNOR2_X1 U441 ( .A(G902), .B(KEYINPUT88), .ZN(n455) );
  INV_X1 U442 ( .A(KEYINPUT82), .ZN(n430) );
  AND2_X1 U443 ( .A1(n422), .A2(n420), .ZN(n419) );
  INV_X1 U444 ( .A(KEYINPUT76), .ZN(n438) );
  NOR2_X1 U445 ( .A1(n726), .A2(n727), .ZN(n439) );
  NAND2_X1 U446 ( .A1(n402), .A2(n400), .ZN(n399) );
  NOR2_X1 U447 ( .A1(n401), .A2(n747), .ZN(n400) );
  XNOR2_X1 U448 ( .A(G113), .B(G137), .ZN(n515) );
  XOR2_X1 U449 ( .A(KEYINPUT5), .B(KEYINPUT94), .Z(n513) );
  XNOR2_X1 U450 ( .A(G131), .B(KEYINPUT4), .ZN(n501) );
  XNOR2_X1 U451 ( .A(G113), .B(G104), .ZN(n461) );
  NAND2_X1 U452 ( .A1(n383), .A2(n655), .ZN(n721) );
  XNOR2_X1 U453 ( .A(n468), .B(n467), .ZN(n552) );
  NOR2_X1 U454 ( .A1(n405), .A2(n397), .ZN(n396) );
  INV_X1 U455 ( .A(KEYINPUT19), .ZN(n397) );
  INV_X1 U456 ( .A(n399), .ZN(n393) );
  NOR2_X1 U457 ( .A1(n599), .A2(n555), .ZN(n541) );
  NAND2_X1 U458 ( .A1(n426), .A2(n425), .ZN(n423) );
  NAND2_X1 U459 ( .A1(n421), .A2(KEYINPUT71), .ZN(n420) );
  NAND2_X1 U460 ( .A1(G234), .A2(G237), .ZN(n528) );
  INV_X1 U461 ( .A(G237), .ZN(n456) );
  INV_X1 U462 ( .A(KEYINPUT8), .ZN(n476) );
  NAND2_X1 U463 ( .A1(n475), .A2(G234), .ZN(n477) );
  XNOR2_X1 U464 ( .A(KEYINPUT96), .B(KEYINPUT11), .ZN(n408) );
  XNOR2_X1 U465 ( .A(G140), .B(KEYINPUT12), .ZN(n409) );
  XNOR2_X1 U466 ( .A(G122), .B(KEYINPUT99), .ZN(n411) );
  NAND2_X1 U467 ( .A1(n381), .A2(n380), .ZN(n615) );
  INV_X1 U468 ( .A(n700), .ZN(n380) );
  XNOR2_X1 U469 ( .A(n652), .B(n651), .ZN(n383) );
  NAND2_X1 U470 ( .A1(n406), .A2(n657), .ZN(n404) );
  OR2_X1 U471 ( .A1(n681), .A2(n403), .ZN(n402) );
  NAND2_X1 U472 ( .A1(n442), .A2(n656), .ZN(n403) );
  XNOR2_X1 U473 ( .A(n493), .B(n443), .ZN(n494) );
  XNOR2_X1 U474 ( .A(G469), .B(KEYINPUT72), .ZN(n509) );
  XNOR2_X1 U475 ( .A(n366), .B(n520), .ZN(n674) );
  XOR2_X1 U476 ( .A(KEYINPUT23), .B(KEYINPUT92), .Z(n485) );
  XNOR2_X1 U477 ( .A(G119), .B(n361), .ZN(n486) );
  INV_X1 U478 ( .A(G116), .ZN(n470) );
  XNOR2_X1 U479 ( .A(KEYINPUT101), .B(KEYINPUT7), .ZN(n473) );
  XOR2_X1 U480 ( .A(KEYINPUT102), .B(KEYINPUT9), .Z(n474) );
  XNOR2_X1 U481 ( .A(G122), .B(G107), .ZN(n471) );
  XNOR2_X1 U482 ( .A(n410), .B(n407), .ZN(n464) );
  XNOR2_X1 U483 ( .A(n412), .B(n411), .ZN(n410) );
  XNOR2_X1 U484 ( .A(n409), .B(n408), .ZN(n407) );
  XNOR2_X1 U485 ( .A(KEYINPUT97), .B(KEYINPUT98), .ZN(n412) );
  INV_X1 U486 ( .A(KEYINPUT10), .ZN(n440) );
  AND2_X1 U487 ( .A1(n661), .A2(n657), .ZN(n658) );
  XNOR2_X1 U488 ( .A(G101), .B(G110), .ZN(n503) );
  XOR2_X1 U489 ( .A(G104), .B(G107), .Z(n504) );
  XNOR2_X1 U490 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n448) );
  XNOR2_X1 U491 ( .A(KEYINPUT79), .B(KEYINPUT4), .ZN(n451) );
  NAND2_X1 U492 ( .A1(n393), .A2(n391), .ZN(n390) );
  NOR2_X1 U493 ( .A1(n392), .A2(KEYINPUT19), .ZN(n391) );
  NAND2_X1 U494 ( .A1(n431), .A2(n553), .ZN(n641) );
  INV_X1 U495 ( .A(n599), .ZN(n732) );
  INV_X1 U496 ( .A(n581), .ZN(n609) );
  XOR2_X1 U497 ( .A(KEYINPUT87), .B(n671), .Z(n698) );
  OR2_X1 U498 ( .A1(n711), .A2(n703), .ZN(n369) );
  AND2_X1 U499 ( .A1(n627), .A2(n429), .ZN(n370) );
  XNOR2_X1 U500 ( .A(G137), .B(G140), .ZN(n371) );
  AND2_X1 U501 ( .A1(n437), .A2(KEYINPUT44), .ZN(n373) );
  AND2_X1 U502 ( .A1(n359), .A2(n424), .ZN(n374) );
  AND2_X1 U503 ( .A1(n425), .A2(KEYINPUT71), .ZN(n375) );
  AND2_X1 U504 ( .A1(n402), .A2(n404), .ZN(n376) );
  XNOR2_X1 U505 ( .A(n746), .B(n430), .ZN(n629) );
  XOR2_X1 U506 ( .A(KEYINPUT70), .B(KEYINPUT47), .Z(n377) );
  INV_X1 U507 ( .A(KEYINPUT74), .ZN(n429) );
  AND2_X1 U508 ( .A1(n596), .A2(n595), .ZN(n378) );
  XNOR2_X1 U509 ( .A(n455), .B(KEYINPUT15), .ZN(n656) );
  XNOR2_X2 U510 ( .A(n379), .B(n485), .ZN(n489) );
  NAND2_X2 U511 ( .A1(n484), .A2(G221), .ZN(n379) );
  XNOR2_X1 U512 ( .A(n439), .B(n438), .ZN(n600) );
  NAND2_X1 U513 ( .A1(n369), .A2(n629), .ZN(n381) );
  NOR2_X2 U514 ( .A1(n677), .A2(n698), .ZN(n679) );
  NOR2_X2 U515 ( .A1(n672), .A2(n698), .ZN(n673) );
  NOR2_X2 U516 ( .A1(n684), .A2(n698), .ZN(n685) );
  AND2_X1 U517 ( .A1(n383), .A2(n662), .ZN(n665) );
  NAND2_X1 U518 ( .A1(n628), .A2(n627), .ZN(n384) );
  AND2_X1 U519 ( .A1(n628), .A2(n370), .ZN(n425) );
  NAND2_X1 U520 ( .A1(n385), .A2(n657), .ZN(n417) );
  NAND2_X1 U521 ( .A1(n386), .A2(n389), .ZN(n385) );
  NAND2_X1 U522 ( .A1(n372), .A2(n659), .ZN(n386) );
  XNOR2_X2 U523 ( .A(n388), .B(n387), .ZN(n518) );
  XNOR2_X2 U524 ( .A(KEYINPUT3), .B(G119), .ZN(n387) );
  XNOR2_X2 U525 ( .A(G101), .B(G116), .ZN(n388) );
  INV_X1 U526 ( .A(KEYINPUT2), .ZN(n389) );
  NAND2_X1 U527 ( .A1(n393), .A2(n405), .ZN(n632) );
  INV_X1 U528 ( .A(n405), .ZN(n392) );
  INV_X1 U529 ( .A(n396), .ZN(n395) );
  NAND2_X1 U530 ( .A1(n399), .A2(KEYINPUT19), .ZN(n398) );
  NAND2_X1 U531 ( .A1(n405), .A2(n376), .ZN(n562) );
  INV_X1 U532 ( .A(n404), .ZN(n401) );
  NAND2_X1 U533 ( .A1(n681), .A2(n406), .ZN(n405) );
  INV_X1 U534 ( .A(n442), .ZN(n406) );
  NAND2_X1 U535 ( .A1(n623), .A2(n567), .ZN(n570) );
  NAND2_X1 U536 ( .A1(n658), .A2(n659), .ZN(n416) );
  NAND2_X1 U537 ( .A1(n375), .A2(n426), .ZN(n422) );
  NAND2_X1 U538 ( .A1(n374), .A2(n423), .ZN(n418) );
  NAND2_X1 U539 ( .A1(n424), .A2(n428), .ZN(n421) );
  INV_X1 U540 ( .A(n631), .ZN(n426) );
  NAND2_X1 U541 ( .A1(n631), .A2(KEYINPUT74), .ZN(n428) );
  INV_X1 U542 ( .A(n653), .ZN(n702) );
  NAND2_X1 U543 ( .A1(n598), .A2(n597), .ZN(n653) );
  INV_X1 U544 ( .A(n598), .ZN(n431) );
  NAND2_X1 U545 ( .A1(n435), .A2(n432), .ZN(n621) );
  NAND2_X1 U546 ( .A1(n433), .A2(n378), .ZN(n432) );
  NAND2_X1 U547 ( .A1(n796), .A2(n434), .ZN(n433) );
  AND2_X1 U548 ( .A1(n617), .A2(n618), .ZN(n434) );
  XNOR2_X2 U549 ( .A(n594), .B(n593), .ZN(n796) );
  NAND2_X1 U550 ( .A1(n587), .A2(n586), .ZN(n437) );
  NOR2_X1 U551 ( .A1(n600), .A2(n611), .ZN(n588) );
  XOR2_X1 U552 ( .A(n458), .B(n457), .Z(n442) );
  AND2_X1 U553 ( .A1(n496), .A2(G217), .ZN(n443) );
  AND2_X1 U554 ( .A1(n355), .A2(n599), .ZN(n444) );
  INV_X1 U555 ( .A(n656), .ZN(n657) );
  INV_X1 U556 ( .A(KEYINPUT93), .ZN(n514) );
  XNOR2_X1 U557 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U558 ( .A(n517), .B(n516), .ZN(n519) );
  INV_X1 U559 ( .A(KEYINPUT69), .ZN(n499) );
  BUF_X1 U560 ( .A(n721), .Z(n785) );
  XNOR2_X1 U561 ( .A(n461), .B(n445), .ZN(n446) );
  INV_X4 U562 ( .A(G953), .ZN(n475) );
  NAND2_X1 U563 ( .A1(n475), .A2(G224), .ZN(n449) );
  XNOR2_X1 U564 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U565 ( .A(n450), .B(n459), .ZN(n453) );
  XNOR2_X2 U566 ( .A(G143), .B(G128), .ZN(n469) );
  XNOR2_X1 U567 ( .A(n469), .B(n451), .ZN(n452) );
  XNOR2_X1 U568 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U569 ( .A(n771), .B(n454), .ZN(n681) );
  NAND2_X1 U570 ( .A1(n522), .A2(n456), .ZN(n525) );
  NAND2_X1 U571 ( .A1(n525), .A2(G210), .ZN(n458) );
  INV_X1 U572 ( .A(KEYINPUT89), .ZN(n457) );
  INV_X1 U573 ( .A(n562), .ZN(n537) );
  NAND2_X1 U574 ( .A1(G214), .A2(n511), .ZN(n460) );
  XNOR2_X1 U575 ( .A(n460), .B(n490), .ZN(n466) );
  XNOR2_X1 U576 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U577 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U578 ( .A(n466), .B(n465), .ZN(n667) );
  NAND2_X1 U579 ( .A1(n667), .A2(n522), .ZN(n468) );
  XNOR2_X1 U580 ( .A(KEYINPUT13), .B(G475), .ZN(n467) );
  XNOR2_X1 U581 ( .A(n471), .B(n470), .ZN(n472) );
  XNOR2_X1 U582 ( .A(n502), .B(n472), .ZN(n481) );
  XNOR2_X1 U583 ( .A(n474), .B(n473), .ZN(n479) );
  XNOR2_X2 U584 ( .A(n477), .B(n476), .ZN(n484) );
  NAND2_X1 U585 ( .A1(G217), .A2(n484), .ZN(n478) );
  XNOR2_X1 U586 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U587 ( .A(n481), .B(n480), .ZN(n692) );
  NAND2_X1 U588 ( .A1(n692), .A2(n522), .ZN(n483) );
  XNOR2_X1 U589 ( .A(KEYINPUT103), .B(G478), .ZN(n482) );
  XNOR2_X1 U590 ( .A(n483), .B(n482), .ZN(n553) );
  OR2_X1 U591 ( .A1(n552), .A2(n553), .ZN(n590) );
  XOR2_X1 U592 ( .A(KEYINPUT24), .B(G110), .Z(n487) );
  XOR2_X1 U593 ( .A(n487), .B(n486), .Z(n488) );
  XNOR2_X1 U594 ( .A(n490), .B(n371), .ZN(n784) );
  NAND2_X1 U595 ( .A1(n687), .A2(n522), .ZN(n495) );
  XOR2_X1 U596 ( .A(KEYINPUT25), .B(KEYINPUT78), .Z(n493) );
  NAND2_X1 U597 ( .A1(G234), .A2(n656), .ZN(n492) );
  XNOR2_X1 U598 ( .A(n492), .B(KEYINPUT20), .ZN(n496) );
  AND2_X1 U599 ( .A1(n496), .A2(G221), .ZN(n498) );
  INV_X1 U600 ( .A(KEYINPUT21), .ZN(n497) );
  XNOR2_X1 U601 ( .A(n498), .B(n497), .ZN(n729) );
  INV_X1 U602 ( .A(n729), .ZN(n571) );
  XNOR2_X1 U603 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U604 ( .A(n371), .B(n505), .ZN(n507) );
  NAND2_X1 U605 ( .A1(G227), .A2(n475), .ZN(n506) );
  XNOR2_X1 U606 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X2 U607 ( .A(n510), .B(n509), .ZN(n557) );
  NOR2_X1 U608 ( .A1(n726), .A2(n557), .ZN(n606) );
  XOR2_X1 U609 ( .A(KEYINPUT30), .B(KEYINPUT107), .Z(n527) );
  NAND2_X1 U610 ( .A1(n511), .A2(G210), .ZN(n512) );
  XNOR2_X1 U611 ( .A(n513), .B(n512), .ZN(n517) );
  XNOR2_X1 U612 ( .A(n519), .B(n518), .ZN(n520) );
  NAND2_X1 U613 ( .A1(n674), .A2(n522), .ZN(n524) );
  XNOR2_X1 U614 ( .A(G472), .B(KEYINPUT73), .ZN(n523) );
  NAND2_X1 U615 ( .A1(n525), .A2(G214), .ZN(n743) );
  NAND2_X1 U616 ( .A1(n732), .A2(n743), .ZN(n526) );
  XNOR2_X1 U617 ( .A(n527), .B(n526), .ZN(n534) );
  XNOR2_X1 U618 ( .A(n528), .B(KEYINPUT90), .ZN(n529) );
  XNOR2_X1 U619 ( .A(KEYINPUT14), .B(n529), .ZN(n530) );
  NAND2_X1 U620 ( .A1(G952), .A2(n530), .ZN(n759) );
  NOR2_X1 U621 ( .A1(n759), .A2(G953), .ZN(n563) );
  AND2_X1 U622 ( .A1(n530), .A2(G953), .ZN(n531) );
  NAND2_X1 U623 ( .A1(G902), .A2(n531), .ZN(n564) );
  NOR2_X1 U624 ( .A1(G900), .A2(n564), .ZN(n532) );
  XNOR2_X1 U625 ( .A(n532), .B(KEYINPUT106), .ZN(n533) );
  NOR2_X1 U626 ( .A1(n563), .A2(n533), .ZN(n539) );
  NOR2_X1 U627 ( .A1(n534), .A2(n539), .ZN(n535) );
  NAND2_X1 U628 ( .A1(n606), .A2(n535), .ZN(n639) );
  NOR2_X1 U629 ( .A1(n590), .A2(n639), .ZN(n536) );
  NAND2_X1 U630 ( .A1(n537), .A2(n536), .ZN(n627) );
  XNOR2_X1 U631 ( .A(G143), .B(KEYINPUT114), .ZN(n538) );
  XNOR2_X1 U632 ( .A(n627), .B(n538), .ZN(G45) );
  NOR2_X1 U633 ( .A1(n729), .A2(n539), .ZN(n540) );
  NAND2_X1 U634 ( .A1(n540), .A2(n581), .ZN(n555) );
  XNOR2_X1 U635 ( .A(n541), .B(KEYINPUT28), .ZN(n543) );
  INV_X1 U636 ( .A(n557), .ZN(n542) );
  AND2_X1 U637 ( .A1(n552), .A2(n553), .ZN(n749) );
  NAND2_X1 U638 ( .A1(n749), .A2(n743), .ZN(n545) );
  INV_X1 U639 ( .A(KEYINPUT38), .ZN(n544) );
  XNOR2_X1 U640 ( .A(n562), .B(n544), .ZN(n748) );
  OR2_X1 U641 ( .A1(n545), .A2(n748), .ZN(n549) );
  XNOR2_X1 U642 ( .A(KEYINPUT111), .B(KEYINPUT41), .ZN(n547) );
  INV_X1 U643 ( .A(KEYINPUT110), .ZN(n546) );
  XNOR2_X1 U644 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U645 ( .A(n549), .B(n548), .ZN(n740) );
  NAND2_X1 U646 ( .A1(n624), .A2(n740), .ZN(n551) );
  XNOR2_X1 U647 ( .A(KEYINPUT112), .B(KEYINPUT42), .ZN(n550) );
  XNOR2_X1 U648 ( .A(n551), .B(n550), .ZN(n645) );
  XNOR2_X1 U649 ( .A(n645), .B(G137), .ZN(G39) );
  XNOR2_X1 U650 ( .A(n552), .B(KEYINPUT100), .ZN(n598) );
  INV_X1 U651 ( .A(n553), .ZN(n597) );
  INV_X1 U652 ( .A(n641), .ZN(n712) );
  INV_X1 U653 ( .A(KEYINPUT6), .ZN(n554) );
  XNOR2_X1 U654 ( .A(n599), .B(n554), .ZN(n611) );
  NOR2_X1 U655 ( .A1(n611), .A2(n555), .ZN(n556) );
  NAND2_X1 U656 ( .A1(n712), .A2(n556), .ZN(n633) );
  INV_X1 U657 ( .A(n355), .ZN(n636) );
  NAND2_X1 U658 ( .A1(n743), .A2(n355), .ZN(n558) );
  NOR2_X1 U659 ( .A1(n633), .A2(n558), .ZN(n560) );
  INV_X1 U660 ( .A(KEYINPUT43), .ZN(n559) );
  XNOR2_X1 U661 ( .A(n560), .B(n559), .ZN(n561) );
  NAND2_X1 U662 ( .A1(n561), .A2(n562), .ZN(n662) );
  XNOR2_X1 U663 ( .A(n662), .B(G140), .ZN(G42) );
  INV_X1 U664 ( .A(n743), .ZN(n747) );
  INV_X1 U665 ( .A(n563), .ZN(n566) );
  OR2_X1 U666 ( .A1(n564), .A2(G898), .ZN(n565) );
  NAND2_X1 U667 ( .A1(n566), .A2(n565), .ZN(n567) );
  INV_X1 U668 ( .A(KEYINPUT68), .ZN(n568) );
  XNOR2_X1 U669 ( .A(n568), .B(KEYINPUT0), .ZN(n569) );
  XNOR2_X2 U670 ( .A(n570), .B(n569), .ZN(n601) );
  AND2_X1 U671 ( .A1(n749), .A2(n571), .ZN(n572) );
  NAND2_X1 U672 ( .A1(n601), .A2(n572), .ZN(n574) );
  INV_X1 U673 ( .A(KEYINPUT22), .ZN(n573) );
  XNOR2_X2 U674 ( .A(n574), .B(n573), .ZN(n613) );
  INV_X1 U675 ( .A(n613), .ZN(n577) );
  NOR2_X1 U676 ( .A1(n355), .A2(n367), .ZN(n575) );
  NAND2_X1 U677 ( .A1(n575), .A2(n611), .ZN(n576) );
  XNOR2_X2 U678 ( .A(n578), .B(KEYINPUT32), .ZN(n618) );
  XNOR2_X1 U679 ( .A(n618), .B(G119), .ZN(G21) );
  NAND2_X1 U680 ( .A1(n613), .A2(n444), .ZN(n580) );
  INV_X1 U681 ( .A(KEYINPUT66), .ZN(n579) );
  XNOR2_X1 U682 ( .A(n580), .B(n579), .ZN(n583) );
  BUF_X1 U683 ( .A(n581), .Z(n582) );
  NAND2_X1 U684 ( .A1(n583), .A2(n582), .ZN(n585) );
  INV_X1 U685 ( .A(KEYINPUT105), .ZN(n584) );
  XNOR2_X2 U686 ( .A(n585), .B(n584), .ZN(n617) );
  NAND2_X1 U687 ( .A1(n617), .A2(n618), .ZN(n587) );
  INV_X1 U688 ( .A(KEYINPUT65), .ZN(n586) );
  XNOR2_X1 U689 ( .A(n588), .B(KEYINPUT33), .ZN(n742) );
  XNOR2_X1 U690 ( .A(n601), .B(KEYINPUT91), .ZN(n605) );
  INV_X1 U691 ( .A(n590), .ZN(n591) );
  NAND2_X1 U692 ( .A1(n592), .A2(n591), .ZN(n594) );
  INV_X1 U693 ( .A(KEYINPUT35), .ZN(n593) );
  NOR2_X1 U694 ( .A1(KEYINPUT85), .A2(KEYINPUT65), .ZN(n596) );
  INV_X1 U695 ( .A(KEYINPUT44), .ZN(n595) );
  INV_X1 U696 ( .A(n601), .ZN(n602) );
  XNOR2_X1 U697 ( .A(KEYINPUT31), .B(KEYINPUT95), .ZN(n603) );
  XNOR2_X1 U698 ( .A(n604), .B(n603), .ZN(n711) );
  INV_X1 U699 ( .A(n605), .ZN(n607) );
  NAND2_X1 U700 ( .A1(n607), .A2(n606), .ZN(n608) );
  NOR2_X1 U701 ( .A1(n732), .A2(n608), .ZN(n703) );
  AND2_X1 U702 ( .A1(n355), .A2(n367), .ZN(n610) );
  AND2_X1 U703 ( .A1(n611), .A2(n610), .ZN(n612) );
  AND2_X1 U704 ( .A1(n613), .A2(n612), .ZN(n700) );
  INV_X1 U705 ( .A(KEYINPUT104), .ZN(n614) );
  XNOR2_X1 U706 ( .A(n615), .B(n614), .ZN(n616) );
  XNOR2_X2 U707 ( .A(n622), .B(KEYINPUT45), .ZN(n661) );
  INV_X1 U708 ( .A(n746), .ZN(n625) );
  NAND2_X1 U709 ( .A1(n707), .A2(n625), .ZN(n626) );
  NAND2_X1 U710 ( .A1(n626), .A2(KEYINPUT47), .ZN(n628) );
  OR2_X1 U711 ( .A1(n633), .A2(n632), .ZN(n635) );
  XNOR2_X1 U712 ( .A(KEYINPUT113), .B(KEYINPUT36), .ZN(n634) );
  XNOR2_X1 U713 ( .A(n635), .B(n634), .ZN(n637) );
  NAND2_X1 U714 ( .A1(n637), .A2(n636), .ZN(n716) );
  INV_X1 U715 ( .A(KEYINPUT71), .ZN(n638) );
  NOR2_X1 U716 ( .A1(n639), .A2(n748), .ZN(n640) );
  XNOR2_X1 U717 ( .A(n640), .B(KEYINPUT39), .ZN(n654) );
  OR2_X1 U718 ( .A1(n654), .A2(n641), .ZN(n644) );
  INV_X1 U719 ( .A(KEYINPUT109), .ZN(n642) );
  XNOR2_X1 U720 ( .A(n642), .B(KEYINPUT40), .ZN(n643) );
  XNOR2_X1 U721 ( .A(KEYINPUT84), .B(KEYINPUT46), .ZN(n646) );
  XNOR2_X1 U722 ( .A(n646), .B(KEYINPUT64), .ZN(n647) );
  XNOR2_X1 U723 ( .A(n648), .B(n647), .ZN(n649) );
  INV_X1 U724 ( .A(KEYINPUT48), .ZN(n651) );
  OR2_X1 U725 ( .A1(n654), .A2(n653), .ZN(n719) );
  AND2_X1 U726 ( .A1(n662), .A2(n719), .ZN(n655) );
  INV_X1 U727 ( .A(KEYINPUT83), .ZN(n660) );
  INV_X1 U728 ( .A(n661), .ZN(n666) );
  NAND2_X1 U729 ( .A1(n719), .A2(KEYINPUT2), .ZN(n663) );
  XOR2_X1 U730 ( .A(n663), .B(KEYINPUT80), .Z(n664) );
  NAND2_X1 U731 ( .A1(n665), .A2(n664), .ZN(n720) );
  NAND2_X1 U732 ( .A1(n686), .A2(G475), .ZN(n670) );
  XOR2_X1 U733 ( .A(KEYINPUT67), .B(KEYINPUT59), .Z(n668) );
  XNOR2_X1 U734 ( .A(n667), .B(n668), .ZN(n669) );
  XNOR2_X1 U735 ( .A(n670), .B(n669), .ZN(n672) );
  NOR2_X1 U736 ( .A1(n475), .A2(G952), .ZN(n671) );
  XNOR2_X1 U737 ( .A(n673), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U738 ( .A1(n686), .A2(G472), .ZN(n676) );
  XOR2_X1 U739 ( .A(KEYINPUT62), .B(n674), .Z(n675) );
  XNOR2_X1 U740 ( .A(n676), .B(n675), .ZN(n677) );
  XOR2_X1 U741 ( .A(KEYINPUT86), .B(KEYINPUT63), .Z(n678) );
  XNOR2_X1 U742 ( .A(n679), .B(n678), .ZN(G57) );
  NAND2_X1 U743 ( .A1(n686), .A2(G210), .ZN(n683) );
  XOR2_X1 U744 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n680) );
  XNOR2_X1 U745 ( .A(n681), .B(n680), .ZN(n682) );
  XNOR2_X1 U746 ( .A(n683), .B(n682), .ZN(n684) );
  XNOR2_X1 U747 ( .A(n685), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U748 ( .A(n617), .B(G110), .ZN(G12) );
  NAND2_X1 U749 ( .A1(n360), .A2(G217), .ZN(n689) );
  XOR2_X1 U750 ( .A(n368), .B(KEYINPUT120), .Z(n688) );
  XNOR2_X1 U751 ( .A(n689), .B(n688), .ZN(n690) );
  NOR2_X1 U752 ( .A1(n690), .A2(n698), .ZN(G66) );
  NAND2_X1 U753 ( .A1(n360), .A2(G478), .ZN(n691) );
  XOR2_X1 U754 ( .A(n692), .B(n691), .Z(n693) );
  NOR2_X1 U755 ( .A1(n693), .A2(n698), .ZN(G63) );
  NAND2_X1 U756 ( .A1(n360), .A2(G469), .ZN(n697) );
  XOR2_X1 U757 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n694) );
  XNOR2_X1 U758 ( .A(n695), .B(n694), .ZN(n696) );
  XNOR2_X1 U759 ( .A(n697), .B(n696), .ZN(n699) );
  NOR2_X1 U760 ( .A1(n699), .A2(n698), .ZN(G54) );
  XOR2_X1 U761 ( .A(G101), .B(n700), .Z(G3) );
  NAND2_X1 U762 ( .A1(n703), .A2(n712), .ZN(n701) );
  XNOR2_X1 U763 ( .A(n701), .B(G104), .ZN(G6) );
  XOR2_X1 U764 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n705) );
  NAND2_X1 U765 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U766 ( .A(n705), .B(n704), .ZN(n706) );
  XNOR2_X1 U767 ( .A(G107), .B(n706), .ZN(G9) );
  XOR2_X1 U768 ( .A(n361), .B(KEYINPUT29), .Z(n709) );
  NAND2_X1 U769 ( .A1(n707), .A2(n702), .ZN(n708) );
  XNOR2_X1 U770 ( .A(n709), .B(n708), .ZN(G30) );
  NAND2_X1 U771 ( .A1(n707), .A2(n712), .ZN(n710) );
  XNOR2_X1 U772 ( .A(n710), .B(G146), .ZN(G48) );
  BUF_X1 U773 ( .A(n711), .Z(n714) );
  NAND2_X1 U774 ( .A1(n714), .A2(n712), .ZN(n713) );
  XNOR2_X1 U775 ( .A(n713), .B(G113), .ZN(G15) );
  NAND2_X1 U776 ( .A1(n714), .A2(n702), .ZN(n715) );
  XNOR2_X1 U777 ( .A(n715), .B(G116), .ZN(G18) );
  INV_X1 U778 ( .A(n716), .ZN(n717) );
  XNOR2_X1 U779 ( .A(G125), .B(n717), .ZN(n718) );
  XNOR2_X1 U780 ( .A(n718), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U781 ( .A(G134), .B(n719), .ZN(G36) );
  INV_X1 U782 ( .A(n720), .ZN(n722) );
  NOR2_X1 U783 ( .A1(n722), .A2(n785), .ZN(n723) );
  NAND2_X1 U784 ( .A1(n661), .A2(n723), .ZN(n768) );
  XNOR2_X1 U785 ( .A(KEYINPUT81), .B(KEYINPUT2), .ZN(n724) );
  NOR2_X1 U786 ( .A1(n725), .A2(n724), .ZN(n766) );
  NAND2_X1 U787 ( .A1(n355), .A2(n726), .ZN(n728) );
  XNOR2_X1 U788 ( .A(KEYINPUT50), .B(n728), .ZN(n735) );
  XOR2_X1 U789 ( .A(KEYINPUT115), .B(KEYINPUT49), .Z(n731) );
  NAND2_X1 U790 ( .A1(n729), .A2(n582), .ZN(n730) );
  XNOR2_X1 U791 ( .A(n731), .B(n730), .ZN(n733) );
  NOR2_X1 U792 ( .A1(n733), .A2(n732), .ZN(n734) );
  NAND2_X1 U793 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U794 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U795 ( .A(n738), .B(KEYINPUT51), .ZN(n739) );
  XNOR2_X1 U796 ( .A(KEYINPUT116), .B(n739), .ZN(n741) );
  INV_X1 U797 ( .A(n740), .ZN(n761) );
  NOR2_X1 U798 ( .A1(n741), .A2(n761), .ZN(n755) );
  INV_X1 U799 ( .A(n748), .ZN(n744) );
  NAND2_X1 U800 ( .A1(n744), .A2(n743), .ZN(n745) );
  NOR2_X1 U801 ( .A1(n746), .A2(n745), .ZN(n752) );
  NAND2_X1 U802 ( .A1(n748), .A2(n747), .ZN(n750) );
  AND2_X1 U803 ( .A1(n750), .A2(n749), .ZN(n751) );
  NOR2_X1 U804 ( .A1(n752), .A2(n751), .ZN(n753) );
  NOR2_X1 U805 ( .A1(n742), .A2(n753), .ZN(n754) );
  NOR2_X1 U806 ( .A1(n755), .A2(n754), .ZN(n756) );
  XOR2_X1 U807 ( .A(n756), .B(KEYINPUT52), .Z(n757) );
  XNOR2_X1 U808 ( .A(KEYINPUT117), .B(n757), .ZN(n758) );
  NOR2_X1 U809 ( .A1(n759), .A2(n758), .ZN(n760) );
  XOR2_X1 U810 ( .A(KEYINPUT118), .B(n760), .Z(n764) );
  NOR2_X1 U811 ( .A1(n742), .A2(n761), .ZN(n762) );
  NOR2_X1 U812 ( .A1(n762), .A2(G953), .ZN(n763) );
  NAND2_X1 U813 ( .A1(n764), .A2(n763), .ZN(n765) );
  NOR2_X1 U814 ( .A1(n766), .A2(n765), .ZN(n767) );
  NAND2_X1 U815 ( .A1(n768), .A2(n767), .ZN(n769) );
  XNOR2_X1 U816 ( .A(n769), .B(KEYINPUT119), .ZN(n770) );
  XNOR2_X1 U817 ( .A(KEYINPUT53), .B(n770), .ZN(G75) );
  XNOR2_X1 U818 ( .A(n771), .B(KEYINPUT122), .ZN(n773) );
  NOR2_X1 U819 ( .A1(G898), .A2(n475), .ZN(n772) );
  NOR2_X1 U820 ( .A1(n773), .A2(n772), .ZN(n774) );
  XOR2_X1 U821 ( .A(KEYINPUT124), .B(n774), .Z(n775) );
  XNOR2_X1 U822 ( .A(KEYINPUT123), .B(n775), .ZN(n782) );
  NAND2_X1 U823 ( .A1(n661), .A2(n475), .ZN(n780) );
  XOR2_X1 U824 ( .A(KEYINPUT121), .B(KEYINPUT61), .Z(n777) );
  NAND2_X1 U825 ( .A1(G224), .A2(G953), .ZN(n776) );
  XNOR2_X1 U826 ( .A(n777), .B(n776), .ZN(n778) );
  NAND2_X1 U827 ( .A1(n778), .A2(G898), .ZN(n779) );
  NAND2_X1 U828 ( .A1(n780), .A2(n779), .ZN(n781) );
  XNOR2_X1 U829 ( .A(n782), .B(n781), .ZN(G69) );
  XOR2_X1 U830 ( .A(n783), .B(n784), .Z(n788) );
  INV_X1 U831 ( .A(n788), .ZN(n786) );
  XOR2_X1 U832 ( .A(n786), .B(n785), .Z(n787) );
  NAND2_X1 U833 ( .A1(n787), .A2(n475), .ZN(n794) );
  XOR2_X1 U834 ( .A(n788), .B(G227), .Z(n789) );
  XNOR2_X1 U835 ( .A(n789), .B(KEYINPUT125), .ZN(n790) );
  NAND2_X1 U836 ( .A1(n790), .A2(G900), .ZN(n792) );
  NAND2_X1 U837 ( .A1(n792), .A2(G953), .ZN(n793) );
  NAND2_X1 U838 ( .A1(n794), .A2(n793), .ZN(n795) );
  XNOR2_X1 U839 ( .A(KEYINPUT126), .B(n795), .ZN(G72) );
  XNOR2_X1 U840 ( .A(n796), .B(G122), .ZN(G24) );
  XOR2_X1 U841 ( .A(G131), .B(n797), .Z(n798) );
  XNOR2_X1 U842 ( .A(KEYINPUT127), .B(n798), .ZN(G33) );
endmodule

