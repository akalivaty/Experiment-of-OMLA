//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 0 1 1 0 1 0 1 1 1 1 0 1 0 0 1 1 1 1 1 1 0 1 0 1 1 0 0 0 1 0 1 1 0 0 1 0 1 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:32 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n696, new_n698, new_n699,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n717, new_n718, new_n719, new_n720, new_n721, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n736, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995;
  INV_X1    g000(.A(KEYINPUT97), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  INV_X1    g002(.A(G146), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT16), .ZN(new_n190));
  INV_X1    g004(.A(G125), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G140), .ZN(new_n192));
  INV_X1    g006(.A(G140), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G125), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n192), .A2(new_n194), .A3(KEYINPUT73), .ZN(new_n195));
  OR3_X1    g009(.A1(new_n193), .A2(KEYINPUT73), .A3(G125), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n190), .B1(new_n195), .B2(new_n196), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n194), .A2(KEYINPUT16), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n189), .B1(new_n197), .B2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(new_n198), .ZN(new_n200));
  NOR3_X1   g014(.A1(new_n193), .A2(KEYINPUT73), .A3(G125), .ZN(new_n201));
  XNOR2_X1  g015(.A(G125), .B(G140), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n201), .B1(new_n202), .B2(KEYINPUT73), .ZN(new_n203));
  OAI211_X1 g017(.A(G146), .B(new_n200), .C1(new_n203), .C2(new_n190), .ZN(new_n204));
  INV_X1    g018(.A(G237), .ZN(new_n205));
  INV_X1    g019(.A(G953), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n205), .A2(new_n206), .A3(G214), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT85), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G143), .ZN(new_n209));
  INV_X1    g023(.A(G143), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(KEYINPUT85), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n207), .A2(new_n209), .A3(new_n211), .ZN(new_n212));
  NOR2_X1   g026(.A1(G237), .A2(G953), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n213), .A2(KEYINPUT85), .A3(new_n210), .A4(G214), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n212), .A2(KEYINPUT17), .A3(G131), .A4(new_n214), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n199), .A2(new_n204), .A3(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT89), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT17), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n212), .A2(G131), .A3(new_n214), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(KEYINPUT88), .ZN(new_n221));
  AOI21_X1  g035(.A(G131), .B1(new_n212), .B2(new_n214), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  AOI211_X1 g037(.A(KEYINPUT88), .B(G131), .C1(new_n212), .C2(new_n214), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n219), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n199), .A2(new_n204), .A3(KEYINPUT89), .A4(new_n215), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n218), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  XNOR2_X1  g041(.A(G113), .B(G122), .ZN(new_n228));
  INV_X1    g042(.A(G104), .ZN(new_n229));
  XNOR2_X1  g043(.A(new_n228), .B(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n195), .A2(new_n196), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT86), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  AOI21_X1  g047(.A(KEYINPUT86), .B1(new_n195), .B2(new_n196), .ZN(new_n234));
  OAI21_X1  g048(.A(G146), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n202), .A2(new_n189), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n235), .A2(KEYINPUT87), .A3(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT87), .ZN(new_n238));
  OAI211_X1 g052(.A(new_n238), .B(G146), .C1(new_n233), .C2(new_n234), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n212), .A2(new_n214), .ZN(new_n240));
  NAND2_X1  g054(.A1(KEYINPUT18), .A2(G131), .ZN(new_n241));
  XOR2_X1   g055(.A(new_n240), .B(new_n241), .Z(new_n242));
  NAND3_X1  g056(.A1(new_n237), .A2(new_n239), .A3(new_n242), .ZN(new_n243));
  AND3_X1   g057(.A1(new_n227), .A2(new_n230), .A3(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n230), .B1(new_n227), .B2(new_n243), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n188), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G475), .ZN(new_n247));
  NOR2_X1   g061(.A1(G475), .A2(G902), .ZN(new_n248));
  OAI21_X1  g062(.A(KEYINPUT19), .B1(new_n233), .B2(new_n234), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT19), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n202), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n249), .A2(new_n189), .A3(new_n251), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n223), .A2(new_n224), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n252), .A2(new_n253), .A3(new_n204), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n230), .B1(new_n254), .B2(new_n243), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n248), .B1(new_n244), .B2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT20), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n227), .A2(new_n230), .A3(new_n243), .ZN(new_n259));
  AND2_X1   g073(.A1(new_n254), .A2(new_n243), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n259), .B1(new_n260), .B2(new_n230), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n261), .A2(KEYINPUT20), .A3(new_n248), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n247), .A2(new_n258), .A3(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT90), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n247), .A2(new_n258), .A3(new_n262), .A4(KEYINPUT90), .ZN(new_n266));
  AND2_X1   g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(G128), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(G143), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n268), .A2(G143), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n269), .B1(new_n270), .B2(KEYINPUT13), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT92), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n210), .A2(G128), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT13), .ZN(new_n275));
  OAI21_X1  g089(.A(KEYINPUT92), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  OAI211_X1 g090(.A(new_n273), .B(G134), .C1(new_n271), .C2(new_n276), .ZN(new_n277));
  AND2_X1   g091(.A1(new_n269), .A2(new_n274), .ZN(new_n278));
  INV_X1    g092(.A(G134), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT91), .ZN(new_n281));
  INV_X1    g095(.A(G122), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n281), .B1(new_n282), .B2(G116), .ZN(new_n283));
  INV_X1    g097(.A(G116), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n284), .A2(KEYINPUT91), .A3(G122), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(G107), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n282), .A2(G116), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n286), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n287), .B1(new_n286), .B2(new_n288), .ZN(new_n291));
  OAI211_X1 g105(.A(new_n277), .B(new_n280), .C1(new_n290), .C2(new_n291), .ZN(new_n292));
  AND3_X1   g106(.A1(new_n284), .A2(KEYINPUT91), .A3(G122), .ZN(new_n293));
  AOI21_X1  g107(.A(KEYINPUT91), .B1(new_n284), .B2(G122), .ZN(new_n294));
  OAI21_X1  g108(.A(KEYINPUT14), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT14), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n283), .A2(new_n296), .A3(new_n285), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n295), .A2(new_n288), .A3(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n298), .A2(KEYINPUT93), .A3(G107), .ZN(new_n299));
  XNOR2_X1  g113(.A(new_n278), .B(new_n279), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  AOI22_X1  g115(.A1(new_n298), .A2(G107), .B1(new_n289), .B2(KEYINPUT93), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n292), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  XOR2_X1   g117(.A(KEYINPUT9), .B(G234), .Z(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(G217), .ZN(new_n306));
  NOR3_X1   g120(.A1(new_n305), .A2(new_n306), .A3(G953), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n303), .A2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT94), .ZN(new_n310));
  OAI211_X1 g124(.A(new_n292), .B(new_n307), .C1(new_n301), .C2(new_n302), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n309), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n303), .A2(KEYINPUT94), .A3(new_n308), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n312), .A2(new_n188), .A3(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(G478), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n315), .A2(KEYINPUT15), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(new_n316), .ZN(new_n318));
  NAND4_X1  g132(.A1(new_n312), .A2(new_n188), .A3(new_n313), .A4(new_n318), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n317), .A2(KEYINPUT95), .A3(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(KEYINPUT95), .B1(new_n317), .B2(new_n319), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(G952), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n324), .A2(G953), .ZN(new_n325));
  NAND2_X1  g139(.A1(G234), .A2(G237), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n326), .A2(G902), .A3(G953), .ZN(new_n329));
  XNOR2_X1  g143(.A(new_n329), .B(KEYINPUT96), .ZN(new_n330));
  XNOR2_X1  g144(.A(KEYINPUT21), .B(G898), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n328), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n323), .A2(new_n333), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n187), .B1(new_n267), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n265), .A2(new_n266), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n336), .A2(KEYINPUT97), .A3(new_n323), .A4(new_n333), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(G469), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n279), .A2(G137), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT11), .ZN(new_n341));
  INV_X1    g155(.A(G137), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n341), .B1(G134), .B2(new_n342), .ZN(new_n343));
  NOR3_X1   g157(.A1(new_n279), .A2(KEYINPUT11), .A3(G137), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n340), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(G131), .ZN(new_n346));
  INV_X1    g160(.A(G131), .ZN(new_n347));
  OAI211_X1 g161(.A(new_n347), .B(new_n340), .C1(new_n343), .C2(new_n344), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n346), .A2(KEYINPUT66), .A3(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT66), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n345), .A2(new_n350), .A3(G131), .ZN(new_n351));
  AND2_X1   g165(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT81), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n189), .A2(G143), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n268), .B1(new_n354), .B2(KEYINPUT1), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  OAI21_X1  g170(.A(KEYINPUT64), .B1(new_n189), .B2(G143), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT64), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n358), .A2(new_n210), .A3(G146), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(new_n354), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n210), .A2(G146), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n354), .A2(new_n362), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n363), .A2(new_n268), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT1), .ZN(new_n365));
  AOI22_X1  g179(.A1(new_n356), .A2(new_n361), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT79), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n367), .A2(new_n287), .A3(G104), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(KEYINPUT3), .ZN(new_n369));
  INV_X1    g183(.A(G101), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n229), .A2(G107), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT3), .ZN(new_n372));
  NAND4_X1  g186(.A1(new_n367), .A2(new_n372), .A3(new_n287), .A4(G104), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n369), .A2(new_n370), .A3(new_n371), .A4(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n287), .A2(G104), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n371), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(G101), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n374), .A2(KEYINPUT80), .A3(new_n377), .ZN(new_n378));
  OR2_X1    g192(.A1(new_n377), .A2(KEYINPUT80), .ZN(new_n379));
  AND3_X1   g193(.A1(new_n366), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n356), .A2(new_n363), .ZN(new_n381));
  AND2_X1   g195(.A1(new_n354), .A2(new_n362), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n382), .A2(new_n365), .A3(G128), .ZN(new_n383));
  AOI22_X1  g197(.A1(new_n378), .A2(new_n379), .B1(new_n381), .B2(new_n383), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n352), .B(new_n353), .C1(new_n380), .C2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(KEYINPUT12), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n378), .A2(new_n379), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n381), .A2(new_n383), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT10), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(new_n352), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n369), .A2(new_n371), .A3(new_n373), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(G101), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n394), .A2(KEYINPUT4), .A3(new_n374), .ZN(new_n395));
  NAND4_X1  g209(.A1(new_n354), .A2(new_n362), .A3(KEYINPUT0), .A4(G128), .ZN(new_n396));
  AOI22_X1  g210(.A1(new_n357), .A2(new_n359), .B1(G143), .B2(new_n189), .ZN(new_n397));
  XNOR2_X1  g211(.A(KEYINPUT0), .B(G128), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n396), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT4), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n393), .A2(new_n401), .A3(G101), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n395), .A2(new_n400), .A3(new_n402), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n383), .B1(new_n397), .B2(new_n355), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n387), .A2(KEYINPUT10), .A3(new_n404), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n391), .A2(new_n392), .A3(new_n403), .A4(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n366), .A2(new_n378), .A3(new_n379), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n389), .A2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT12), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n408), .A2(new_n353), .A3(new_n409), .A4(new_n352), .ZN(new_n410));
  XNOR2_X1  g224(.A(G110), .B(G140), .ZN(new_n411));
  AND2_X1   g225(.A1(new_n206), .A2(G227), .ZN(new_n412));
  XOR2_X1   g226(.A(new_n411), .B(new_n412), .Z(new_n413));
  NAND4_X1  g227(.A1(new_n386), .A2(new_n406), .A3(new_n410), .A4(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n391), .A2(new_n403), .A3(new_n405), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(new_n352), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n413), .B1(new_n417), .B2(new_n406), .ZN(new_n418));
  OAI211_X1 g232(.A(new_n339), .B(new_n188), .C1(new_n415), .C2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(G469), .A2(G902), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n386), .A2(new_n406), .A3(new_n410), .ZN(new_n421));
  INV_X1    g235(.A(new_n413), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n417), .A2(new_n406), .A3(new_n413), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n423), .A2(new_n424), .A3(G469), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n419), .A2(new_n420), .A3(new_n425), .ZN(new_n426));
  OAI21_X1  g240(.A(G221), .B1(new_n305), .B2(G902), .ZN(new_n427));
  AND2_X1   g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(G214), .B1(G237), .B2(G902), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(G224), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n431), .A2(G953), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n399), .A2(G125), .ZN(new_n433));
  XNOR2_X1  g247(.A(new_n433), .B(KEYINPUT82), .ZN(new_n434));
  OAI211_X1 g248(.A(new_n383), .B(new_n191), .C1(new_n355), .C2(new_n397), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT83), .ZN(new_n436));
  XNOR2_X1  g250(.A(new_n435), .B(new_n436), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n432), .B1(new_n434), .B2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT82), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n433), .B(new_n439), .ZN(new_n440));
  XNOR2_X1  g254(.A(new_n435), .B(KEYINPUT83), .ZN(new_n441));
  INV_X1    g255(.A(new_n432), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n440), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n438), .A2(new_n443), .ZN(new_n444));
  XOR2_X1   g258(.A(KEYINPUT2), .B(G113), .Z(new_n445));
  XNOR2_X1  g259(.A(G116), .B(G119), .ZN(new_n446));
  XNOR2_X1  g260(.A(new_n445), .B(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n395), .A2(new_n402), .A3(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(G119), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(G116), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n450), .A2(KEYINPUT5), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n451), .B1(KEYINPUT5), .B2(new_n446), .ZN(new_n452));
  AOI22_X1  g266(.A1(new_n452), .A2(G113), .B1(new_n446), .B2(new_n445), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n387), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n448), .A2(new_n454), .ZN(new_n455));
  XOR2_X1   g269(.A(G110), .B(G122), .Z(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(new_n456), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n448), .A2(new_n454), .A3(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n457), .A2(KEYINPUT6), .A3(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT6), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n455), .A2(new_n461), .A3(new_n456), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n444), .A2(new_n460), .A3(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT7), .ZN(new_n464));
  OAI22_X1  g278(.A1(new_n434), .A2(new_n437), .B1(new_n464), .B2(new_n432), .ZN(new_n465));
  NAND4_X1  g279(.A1(new_n440), .A2(new_n441), .A3(KEYINPUT7), .A4(new_n442), .ZN(new_n466));
  XOR2_X1   g280(.A(KEYINPUT84), .B(KEYINPUT8), .Z(new_n467));
  XNOR2_X1  g281(.A(new_n456), .B(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(new_n454), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n387), .A2(new_n453), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND4_X1  g285(.A1(new_n465), .A2(new_n466), .A3(new_n459), .A4(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n463), .A2(new_n188), .A3(new_n472), .ZN(new_n473));
  OAI21_X1  g287(.A(G210), .B1(G237), .B2(G902), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n463), .A2(new_n188), .A3(new_n474), .A4(new_n472), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n430), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  XOR2_X1   g292(.A(KEYINPUT69), .B(KEYINPUT27), .Z(new_n479));
  NAND2_X1  g293(.A1(new_n213), .A2(G210), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n479), .B(new_n480), .ZN(new_n481));
  XNOR2_X1  g295(.A(KEYINPUT26), .B(G101), .ZN(new_n482));
  XNOR2_X1  g296(.A(new_n481), .B(new_n482), .ZN(new_n483));
  XNOR2_X1  g297(.A(KEYINPUT70), .B(KEYINPUT28), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n279), .A2(KEYINPUT67), .A3(G137), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n342), .A2(G134), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(KEYINPUT67), .B1(new_n279), .B2(G137), .ZN(new_n488));
  OAI21_X1  g302(.A(G131), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(new_n348), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT68), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n489), .A2(new_n348), .A3(KEYINPUT68), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n492), .A2(new_n404), .A3(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n349), .A2(new_n400), .A3(new_n351), .ZN(new_n495));
  INV_X1    g309(.A(new_n447), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n398), .B1(new_n360), .B2(new_n354), .ZN(new_n499));
  INV_X1    g313(.A(new_n396), .ZN(new_n500));
  OAI21_X1  g314(.A(KEYINPUT65), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT65), .ZN(new_n502));
  OAI211_X1 g316(.A(new_n396), .B(new_n502), .C1(new_n397), .C2(new_n398), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n349), .A2(new_n501), .A3(new_n351), .A4(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n404), .A2(new_n348), .A3(new_n489), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n496), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n484), .B1(new_n498), .B2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT28), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n497), .A2(new_n508), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n483), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  AND3_X1   g325(.A1(new_n494), .A2(new_n495), .A3(KEYINPUT30), .ZN(new_n512));
  AOI21_X1  g326(.A(KEYINPUT30), .B1(new_n504), .B2(new_n505), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n498), .B1(new_n514), .B2(new_n447), .ZN(new_n515));
  AOI21_X1  g329(.A(KEYINPUT31), .B1(new_n515), .B2(new_n483), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n504), .A2(new_n505), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT30), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n494), .A2(new_n495), .A3(KEYINPUT30), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n519), .A2(new_n447), .A3(new_n520), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n521), .A2(KEYINPUT31), .A3(new_n483), .A4(new_n497), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n511), .B1(new_n516), .B2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT32), .ZN(new_n525));
  NOR2_X1   g339(.A1(G472), .A2(G902), .ZN(new_n526));
  XOR2_X1   g340(.A(new_n526), .B(KEYINPUT71), .Z(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n524), .A2(new_n525), .A3(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n521), .A2(new_n483), .A3(new_n497), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT31), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n510), .B1(new_n532), .B2(new_n522), .ZN(new_n533));
  OAI21_X1  g347(.A(KEYINPUT32), .B1(new_n533), .B2(new_n527), .ZN(new_n534));
  INV_X1    g348(.A(new_n509), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n496), .B1(new_n494), .B2(new_n495), .ZN(new_n536));
  OR2_X1    g350(.A1(new_n498), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n535), .B1(new_n537), .B2(KEYINPUT28), .ZN(new_n538));
  INV_X1    g352(.A(new_n483), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT29), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(G902), .B1(new_n538), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n521), .A2(new_n497), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(new_n539), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n507), .A2(new_n483), .A3(new_n509), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n544), .A2(new_n540), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n542), .A2(new_n546), .ZN(new_n547));
  AOI22_X1  g361(.A1(new_n529), .A2(new_n534), .B1(G472), .B2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT25), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(KEYINPUT77), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT23), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n551), .B1(new_n449), .B2(G128), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n449), .A2(G128), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n268), .A2(KEYINPUT23), .A3(G119), .ZN(new_n554));
  AND3_X1   g368(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(G110), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT72), .ZN(new_n558));
  NOR3_X1   g372(.A1(new_n558), .A2(new_n449), .A3(G128), .ZN(new_n559));
  AOI21_X1  g373(.A(KEYINPUT72), .B1(new_n268), .B2(G119), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n553), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  XNOR2_X1  g375(.A(KEYINPUT24), .B(G110), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  AOI211_X1 g377(.A(new_n557), .B(new_n563), .C1(new_n199), .C2(new_n204), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT74), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n555), .A2(new_n565), .A3(new_n556), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n561), .A2(new_n562), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n568));
  OAI21_X1  g382(.A(KEYINPUT74), .B1(new_n568), .B2(G110), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n566), .A2(new_n567), .A3(new_n569), .ZN(new_n570));
  AND3_X1   g384(.A1(new_n570), .A2(new_n236), .A3(new_n204), .ZN(new_n571));
  OAI21_X1  g385(.A(KEYINPUT75), .B1(new_n564), .B2(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n206), .A2(G221), .A3(G234), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n573), .B(KEYINPUT76), .ZN(new_n574));
  AND2_X1   g388(.A1(new_n574), .A2(KEYINPUT22), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n574), .A2(KEYINPUT22), .ZN(new_n576));
  OR3_X1    g390(.A1(new_n575), .A2(new_n576), .A3(new_n342), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n342), .B1(new_n575), .B2(new_n576), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n563), .B1(new_n199), .B2(new_n204), .ZN(new_n580));
  INV_X1    g394(.A(new_n557), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT75), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n570), .A2(new_n236), .A3(new_n204), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n572), .A2(new_n579), .A3(new_n585), .ZN(new_n586));
  OAI211_X1 g400(.A(new_n577), .B(new_n578), .C1(new_n564), .C2(new_n571), .ZN(new_n587));
  AND2_X1   g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n550), .B1(new_n588), .B2(G902), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n306), .B1(G234), .B2(new_n188), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n586), .A2(new_n587), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n591), .A2(KEYINPUT77), .A3(new_n549), .A4(new_n188), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n589), .A2(new_n590), .A3(new_n592), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n590), .A2(G902), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n594), .B(KEYINPUT78), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n593), .B1(new_n596), .B2(new_n588), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n548), .A2(new_n597), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n338), .A2(new_n428), .A3(new_n478), .A4(new_n598), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n599), .B(KEYINPUT98), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n600), .B(new_n370), .ZN(G3));
  NAND2_X1  g415(.A1(new_n478), .A2(new_n333), .ZN(new_n602));
  OAI21_X1  g416(.A(G472), .B1(new_n533), .B2(G902), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n524), .A2(new_n528), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n426), .A2(new_n427), .ZN(new_n606));
  NOR4_X1   g420(.A1(new_n602), .A2(new_n605), .A3(new_n597), .A4(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT33), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n312), .A2(new_n608), .A3(new_n313), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n309), .A2(KEYINPUT33), .A3(new_n311), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n609), .A2(G478), .A3(new_n188), .A4(new_n610), .ZN(new_n611));
  XOR2_X1   g425(.A(KEYINPUT99), .B(G478), .Z(new_n612));
  NAND2_X1  g426(.A1(new_n314), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n265), .A2(new_n266), .A3(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n607), .A2(new_n616), .ZN(new_n617));
  XNOR2_X1  g431(.A(KEYINPUT100), .B(KEYINPUT34), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(new_n229), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n617), .B(new_n619), .ZN(G6));
  NOR2_X1   g434(.A1(new_n323), .A2(new_n263), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n607), .A2(new_n621), .ZN(new_n622));
  XOR2_X1   g436(.A(KEYINPUT35), .B(G107), .Z(new_n623));
  XNOR2_X1  g437(.A(new_n622), .B(new_n623), .ZN(G9));
  INV_X1    g438(.A(new_n605), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT36), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n577), .A2(new_n626), .A3(new_n578), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT101), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n627), .B(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n572), .A2(new_n585), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n627), .B(KEYINPUT101), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(new_n630), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n596), .B1(new_n632), .B2(new_n634), .ZN(new_n635));
  AOI22_X1  g449(.A1(new_n591), .A2(new_n188), .B1(KEYINPUT77), .B2(new_n549), .ZN(new_n636));
  AOI211_X1 g450(.A(G902), .B(new_n550), .C1(new_n586), .C2(new_n587), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n635), .B1(new_n638), .B2(new_n590), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n606), .A2(new_n639), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n338), .A2(new_n478), .A3(new_n625), .A4(new_n640), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(KEYINPUT37), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(new_n556), .ZN(G12));
  XOR2_X1   g457(.A(new_n327), .B(KEYINPUT103), .Z(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(G900), .ZN(new_n646));
  AND3_X1   g460(.A1(new_n330), .A2(KEYINPUT102), .A3(new_n646), .ZN(new_n647));
  AOI21_X1  g461(.A(KEYINPUT102), .B1(new_n330), .B2(new_n646), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n645), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  NOR3_X1   g464(.A1(new_n323), .A2(new_n263), .A3(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n547), .A2(G472), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n525), .B1(new_n524), .B2(new_n528), .ZN(new_n653));
  NOR3_X1   g467(.A1(new_n533), .A2(KEYINPUT32), .A3(new_n527), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n652), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n651), .A2(new_n655), .A3(new_n640), .A4(new_n478), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(G128), .ZN(G30));
  XOR2_X1   g471(.A(new_n649), .B(KEYINPUT39), .Z(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n428), .A2(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT40), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n539), .B1(new_n498), .B2(new_n536), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n530), .A2(G472), .A3(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(G472), .A2(G902), .ZN(new_n665));
  AND3_X1   g479(.A1(new_n664), .A2(KEYINPUT104), .A3(new_n665), .ZN(new_n666));
  AOI21_X1  g480(.A(KEYINPUT104), .B1(new_n664), .B2(new_n665), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n668), .B1(new_n653), .B2(new_n654), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(KEYINPUT105), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT105), .ZN(new_n671));
  OAI211_X1 g485(.A(new_n671), .B(new_n668), .C1(new_n653), .C2(new_n654), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n322), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(new_n320), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n675), .A2(new_n639), .A3(new_n265), .A4(new_n266), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n662), .A2(new_n673), .A3(new_n677), .ZN(new_n678));
  AND3_X1   g492(.A1(new_n476), .A2(KEYINPUT38), .A3(new_n477), .ZN(new_n679));
  AOI21_X1  g493(.A(KEYINPUT38), .B1(new_n476), .B2(new_n477), .ZN(new_n680));
  OR2_X1    g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  OR2_X1    g495(.A1(new_n681), .A2(new_n430), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n678), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(new_n210), .ZN(G45));
  AND4_X1   g498(.A1(new_n265), .A2(new_n266), .A3(new_n614), .A4(new_n649), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n685), .A2(new_n655), .A3(new_n640), .A4(new_n478), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G146), .ZN(G48));
  NOR2_X1   g501(.A1(new_n415), .A2(new_n418), .ZN(new_n688));
  OAI21_X1  g502(.A(G469), .B1(new_n688), .B2(G902), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n689), .A2(new_n427), .A3(new_n419), .ZN(new_n690));
  NOR4_X1   g504(.A1(new_n548), .A2(new_n602), .A3(new_n597), .A4(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n616), .ZN(new_n692));
  XNOR2_X1  g506(.A(KEYINPUT41), .B(G113), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(KEYINPUT106), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n692), .B(new_n694), .ZN(G15));
  NAND2_X1  g509(.A1(new_n691), .A2(new_n621), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G116), .ZN(G18));
  INV_X1    g511(.A(new_n635), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n593), .A2(new_n698), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n548), .A2(new_n690), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n338), .A2(new_n478), .A3(new_n699), .A4(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G119), .ZN(G21));
  AOI22_X1  g516(.A1(new_n638), .A2(new_n590), .B1(new_n595), .B2(new_n591), .ZN(new_n703));
  OAI22_X1  g517(.A1(new_n516), .A2(new_n523), .B1(new_n483), .B2(new_n538), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(new_n528), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n703), .A2(new_n333), .A3(new_n603), .A4(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n675), .A2(new_n265), .A3(new_n266), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n417), .A2(new_n406), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(new_n422), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(new_n414), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n339), .B1(new_n710), .B2(new_n188), .ZN(new_n711));
  INV_X1    g525(.A(new_n419), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n713), .A2(new_n478), .A3(new_n427), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n706), .A2(new_n707), .A3(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(new_n282), .ZN(G24));
  AND3_X1   g530(.A1(new_n699), .A2(new_n603), .A3(new_n705), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n476), .A2(new_n477), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(new_n429), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n719), .A2(new_n690), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n717), .A2(new_n685), .A3(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G125), .ZN(G27));
  XNOR2_X1  g536(.A(new_n606), .B(KEYINPUT107), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT108), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n724), .B1(new_n718), .B2(new_n430), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n476), .A2(KEYINPUT108), .A3(new_n429), .A4(new_n477), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  INV_X1    g541(.A(new_n727), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n723), .A2(new_n598), .A3(new_n728), .A4(new_n685), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT42), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NOR3_X1   g545(.A1(new_n727), .A2(new_n548), .A3(new_n597), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n732), .A2(KEYINPUT42), .A3(new_n685), .A4(new_n723), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G131), .ZN(G33));
  AND3_X1   g549(.A1(new_n732), .A2(new_n651), .A3(new_n723), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(new_n279), .ZN(G36));
  INV_X1    g551(.A(KEYINPUT43), .ZN(new_n738));
  INV_X1    g552(.A(new_n614), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n738), .B1(new_n267), .B2(new_n739), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n336), .A2(KEYINPUT43), .A3(new_n614), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n742), .A2(new_n605), .A3(new_n699), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT44), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n742), .A2(KEYINPUT44), .A3(new_n605), .A4(new_n699), .ZN(new_n746));
  XOR2_X1   g560(.A(new_n727), .B(KEYINPUT109), .Z(new_n747));
  NAND3_X1  g561(.A1(new_n745), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(KEYINPUT110), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n423), .A2(new_n424), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(KEYINPUT45), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(G469), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n752), .A2(KEYINPUT46), .A3(new_n420), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT46), .ZN(new_n754));
  OAI211_X1 g568(.A(new_n754), .B(G469), .C1(new_n751), .C2(G902), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n753), .A2(new_n419), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(new_n427), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n757), .A2(new_n658), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT110), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n745), .A2(new_n746), .A3(new_n759), .A4(new_n747), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n749), .A2(new_n758), .A3(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G137), .ZN(G39));
  NAND4_X1  g576(.A1(new_n728), .A2(new_n597), .A3(new_n548), .A4(new_n685), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(KEYINPUT111), .ZN(new_n764));
  AOI21_X1  g578(.A(KEYINPUT47), .B1(new_n756), .B2(new_n427), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n756), .A2(KEYINPUT47), .A3(new_n427), .ZN(new_n766));
  INV_X1    g580(.A(new_n766), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n764), .B1(new_n765), .B2(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G140), .ZN(G42));
  OAI21_X1  g583(.A(new_n430), .B1(new_n679), .B2(new_n680), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT119), .ZN(new_n771));
  OR3_X1    g585(.A1(new_n770), .A2(new_n771), .A3(new_n690), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n771), .B1(new_n770), .B2(new_n690), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  AND3_X1   g588(.A1(new_n703), .A2(new_n603), .A3(new_n705), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n645), .B1(new_n740), .B2(new_n741), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n774), .A2(KEYINPUT50), .A3(new_n775), .A4(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT50), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n776), .A2(new_n775), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n772), .A2(new_n773), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n778), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n777), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n727), .A2(new_n690), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n776), .A2(new_n717), .A3(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(new_n672), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n529), .A2(new_n534), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n671), .B1(new_n786), .B2(new_n668), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n788), .A2(new_n328), .A3(new_n703), .A4(new_n783), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n789), .A2(new_n267), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n790), .A2(new_n739), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n782), .A2(KEYINPUT51), .A3(new_n784), .A4(new_n791), .ZN(new_n792));
  AND3_X1   g606(.A1(new_n747), .A2(new_n776), .A3(new_n775), .ZN(new_n793));
  INV_X1    g607(.A(new_n765), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n711), .A2(new_n712), .A3(new_n427), .ZN(new_n795));
  INV_X1    g609(.A(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n794), .A2(new_n766), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n793), .A2(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(new_n798), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n325), .B1(new_n792), .B2(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT51), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT118), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n803), .B1(new_n767), .B2(new_n765), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n794), .A2(KEYINPUT118), .A3(new_n766), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n804), .A2(new_n805), .A3(new_n796), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n806), .A2(new_n793), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  AOI22_X1  g622(.A1(new_n777), .A2(new_n781), .B1(new_n790), .B2(new_n739), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n809), .A2(new_n784), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n802), .B1(new_n808), .B2(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n776), .A2(new_n775), .A3(new_n720), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n789), .A2(new_n615), .ZN(new_n813));
  INV_X1    g627(.A(new_n813), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n801), .A2(new_n811), .A3(new_n812), .A4(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n776), .A2(new_n598), .A3(new_n783), .ZN(new_n816));
  XOR2_X1   g630(.A(new_n816), .B(KEYINPUT48), .Z(new_n817));
  OAI21_X1  g631(.A(KEYINPUT120), .B1(new_n815), .B2(new_n817), .ZN(new_n818));
  AND3_X1   g632(.A1(new_n782), .A2(new_n784), .A3(new_n791), .ZN(new_n819));
  AOI21_X1  g633(.A(KEYINPUT51), .B1(new_n819), .B2(new_n807), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n820), .A2(new_n800), .A3(new_n813), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT120), .ZN(new_n822));
  INV_X1    g636(.A(new_n817), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n821), .A2(new_n822), .A3(new_n823), .A4(new_n812), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT115), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT113), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n428), .A2(new_n478), .A3(new_n649), .ZN(new_n827));
  AOI211_X1 g641(.A(new_n676), .B(new_n827), .C1(new_n670), .C2(new_n672), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n686), .A2(new_n656), .A3(new_n721), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n826), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT52), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n719), .A2(new_n606), .A3(new_n650), .ZN(new_n832));
  OAI211_X1 g646(.A(new_n677), .B(new_n832), .C1(new_n785), .C2(new_n787), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n719), .B1(new_n786), .B2(new_n652), .ZN(new_n834));
  OAI211_X1 g648(.A(new_n834), .B(new_n640), .C1(new_n651), .C2(new_n685), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n833), .A2(KEYINPUT113), .A3(new_n721), .A4(new_n835), .ZN(new_n836));
  AND3_X1   g650(.A1(new_n830), .A2(new_n831), .A3(new_n836), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n831), .B1(new_n830), .B2(new_n836), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n825), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT112), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n317), .A2(new_n319), .ZN(new_n841));
  AOI22_X1  g655(.A1(new_n615), .A2(new_n840), .B1(new_n336), .B2(new_n841), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n842), .B1(new_n840), .B2(new_n615), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n843), .A2(new_n607), .ZN(new_n844));
  AND3_X1   g658(.A1(new_n599), .A2(new_n641), .A3(new_n844), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n715), .B1(new_n691), .B2(new_n616), .ZN(new_n846));
  AND3_X1   g660(.A1(new_n701), .A2(new_n846), .A3(new_n696), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n736), .B1(new_n733), .B2(new_n731), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n723), .A2(new_n685), .A3(new_n717), .ZN(new_n849));
  INV_X1    g663(.A(new_n263), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n655), .A2(new_n640), .A3(new_n850), .A4(new_n649), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n849), .B1(new_n841), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n852), .A2(new_n728), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n845), .A2(new_n847), .A3(new_n848), .A4(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(new_n854), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n686), .A2(new_n656), .A3(new_n721), .ZN(new_n856));
  AOI21_X1  g670(.A(KEYINPUT113), .B1(new_n856), .B2(new_n833), .ZN(new_n857));
  AND4_X1   g671(.A1(KEYINPUT113), .A2(new_n833), .A3(new_n721), .A4(new_n835), .ZN(new_n858));
  OAI21_X1  g672(.A(KEYINPUT52), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n830), .A2(new_n831), .A3(new_n836), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n859), .A2(KEYINPUT115), .A3(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n839), .A2(new_n855), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n862), .A2(KEYINPUT53), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT53), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT114), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n856), .A2(KEYINPUT52), .A3(new_n833), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n860), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n865), .B1(new_n860), .B2(new_n866), .ZN(new_n868));
  OAI211_X1 g682(.A(new_n855), .B(new_n864), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n863), .A2(KEYINPUT54), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n862), .A2(new_n864), .ZN(new_n871));
  XNOR2_X1  g685(.A(KEYINPUT117), .B(KEYINPUT54), .ZN(new_n872));
  INV_X1    g686(.A(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n599), .A2(new_n641), .A3(new_n844), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n701), .A2(new_n846), .A3(new_n696), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(KEYINPUT116), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT116), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n701), .A2(new_n846), .A3(new_n877), .A4(new_n696), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n874), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  AND3_X1   g693(.A1(new_n848), .A2(KEYINPUT53), .A3(new_n853), .ZN(new_n880));
  OAI211_X1 g694(.A(new_n879), .B(new_n880), .C1(new_n867), .C2(new_n868), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n871), .A2(new_n873), .A3(new_n881), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n818), .A2(new_n824), .A3(new_n870), .A4(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n324), .A2(new_n206), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n713), .B(KEYINPUT49), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n267), .A2(new_n739), .ZN(new_n887));
  AND2_X1   g701(.A1(new_n427), .A2(new_n429), .ZN(new_n888));
  AND3_X1   g702(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n889), .A2(new_n703), .A3(new_n681), .A4(new_n788), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n885), .A2(new_n890), .ZN(G75));
  NOR2_X1   g705(.A1(new_n206), .A2(G952), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n859), .A2(new_n860), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n854), .B1(new_n893), .B2(new_n825), .ZN(new_n894));
  AOI21_X1  g708(.A(KEYINPUT53), .B1(new_n894), .B2(new_n861), .ZN(new_n895));
  INV_X1    g709(.A(new_n881), .ZN(new_n896));
  OAI211_X1 g710(.A(G210), .B(G902), .C1(new_n895), .C2(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT56), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n460), .A2(new_n462), .ZN(new_n900));
  XOR2_X1   g714(.A(new_n900), .B(new_n444), .Z(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(KEYINPUT55), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n892), .B1(new_n899), .B2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT121), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n897), .A2(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(new_n902), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n871), .A2(new_n881), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n907), .A2(KEYINPUT121), .A3(G210), .A4(G902), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n905), .A2(new_n898), .A3(new_n906), .A4(new_n908), .ZN(new_n909));
  AND2_X1   g723(.A1(new_n903), .A2(new_n909), .ZN(G51));
  XOR2_X1   g724(.A(new_n420), .B(KEYINPUT57), .Z(new_n911));
  INV_X1    g725(.A(new_n882), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n873), .B1(new_n871), .B2(new_n881), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n911), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(new_n710), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n907), .A2(G469), .A3(G902), .A4(new_n751), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n892), .B1(new_n915), .B2(new_n916), .ZN(G54));
  INV_X1    g731(.A(new_n892), .ZN(new_n918));
  AND2_X1   g732(.A1(KEYINPUT58), .A2(G475), .ZN(new_n919));
  AND3_X1   g733(.A1(new_n907), .A2(G902), .A3(new_n919), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n918), .B1(new_n920), .B2(new_n261), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n907), .A2(G902), .A3(new_n261), .A4(new_n919), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT122), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n920), .A2(KEYINPUT122), .A3(new_n261), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n921), .B1(new_n924), .B2(new_n925), .ZN(G60));
  AND2_X1   g740(.A1(new_n609), .A2(new_n610), .ZN(new_n927));
  INV_X1    g741(.A(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(G478), .A2(G902), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n929), .B(KEYINPUT59), .Z(new_n930));
  INV_X1    g744(.A(new_n913), .ZN(new_n931));
  AOI211_X1 g745(.A(new_n928), .B(new_n930), .C1(new_n931), .C2(new_n882), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n930), .B1(new_n870), .B2(new_n882), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n918), .B1(new_n933), .B2(new_n927), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n932), .A2(new_n934), .ZN(G63));
  NAND2_X1  g749(.A1(G217), .A2(G902), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(KEYINPUT60), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n937), .B1(new_n871), .B2(new_n881), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n918), .B1(new_n938), .B2(new_n591), .ZN(new_n939));
  INV_X1    g753(.A(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(new_n632), .ZN(new_n941));
  INV_X1    g755(.A(new_n634), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n938), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n940), .A2(KEYINPUT61), .A3(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT61), .ZN(new_n945));
  INV_X1    g759(.A(new_n938), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n941), .A2(new_n942), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n945), .B1(new_n948), .B2(new_n939), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n944), .A2(new_n949), .ZN(G66));
  NAND2_X1  g764(.A1(new_n845), .A2(new_n847), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(new_n206), .ZN(new_n952));
  OAI21_X1  g766(.A(G953), .B1(new_n331), .B2(new_n431), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(KEYINPUT123), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n900), .B1(G898), .B2(new_n206), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n955), .B(new_n956), .ZN(G69));
  NAND2_X1  g771(.A1(new_n249), .A2(new_n251), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n514), .B(new_n958), .Z(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(new_n960));
  OAI22_X1  g774(.A1(new_n683), .A2(new_n829), .B1(KEYINPUT124), .B2(KEYINPUT62), .ZN(new_n961));
  XNOR2_X1  g775(.A(KEYINPUT124), .B(KEYINPUT62), .ZN(new_n962));
  OAI211_X1 g776(.A(new_n856), .B(new_n962), .C1(new_n678), .C2(new_n682), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n761), .A2(new_n768), .A3(new_n961), .A4(new_n963), .ZN(new_n964));
  AND4_X1   g778(.A1(new_n428), .A2(new_n843), .A3(new_n659), .A4(new_n732), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n960), .B1(new_n966), .B2(G953), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n967), .A2(KEYINPUT125), .ZN(new_n968));
  NAND2_X1  g782(.A1(G900), .A2(G953), .ZN(new_n969));
  INV_X1    g783(.A(new_n707), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n758), .A2(new_n478), .A3(new_n598), .A4(new_n970), .ZN(new_n971));
  AND2_X1   g785(.A1(new_n848), .A2(new_n856), .ZN(new_n972));
  NAND4_X1  g786(.A1(new_n761), .A2(new_n768), .A3(new_n971), .A4(new_n972), .ZN(new_n973));
  OAI211_X1 g787(.A(new_n959), .B(new_n969), .C1(new_n973), .C2(G953), .ZN(new_n974));
  AND2_X1   g788(.A1(new_n974), .A2(KEYINPUT126), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT125), .ZN(new_n976));
  OAI211_X1 g790(.A(new_n976), .B(new_n960), .C1(new_n966), .C2(G953), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n968), .A2(new_n975), .A3(new_n977), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n206), .B1(G227), .B2(G900), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  INV_X1    g794(.A(new_n979), .ZN(new_n981));
  NAND4_X1  g795(.A1(new_n968), .A2(new_n981), .A3(new_n975), .A4(new_n977), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n980), .A2(new_n982), .ZN(G72));
  XNOR2_X1  g797(.A(new_n665), .B(KEYINPUT63), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n984), .B1(new_n544), .B2(new_n530), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n863), .A2(new_n869), .A3(new_n985), .ZN(new_n986));
  AND2_X1   g800(.A1(new_n986), .A2(new_n918), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n973), .A2(new_n951), .ZN(new_n988));
  OAI211_X1 g802(.A(new_n539), .B(new_n515), .C1(new_n988), .C2(new_n984), .ZN(new_n989));
  NOR3_X1   g803(.A1(new_n964), .A2(new_n951), .A3(new_n965), .ZN(new_n990));
  OAI211_X1 g804(.A(new_n483), .B(new_n543), .C1(new_n990), .C2(new_n984), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n987), .A2(new_n989), .A3(new_n991), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n992), .A2(KEYINPUT127), .ZN(new_n993));
  INV_X1    g807(.A(KEYINPUT127), .ZN(new_n994));
  NAND4_X1  g808(.A1(new_n987), .A2(new_n994), .A3(new_n989), .A4(new_n991), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n993), .A2(new_n995), .ZN(G57));
endmodule


