

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579;

  XOR2_X1 U320 ( .A(KEYINPUT38), .B(n474), .Z(n504) );
  XOR2_X1 U321 ( .A(n428), .B(KEYINPUT54), .Z(n288) );
  INV_X1 U322 ( .A(KEYINPUT99), .ZN(n459) );
  NOR2_X1 U323 ( .A1(n521), .A2(n467), .ZN(n468) );
  XNOR2_X1 U324 ( .A(n327), .B(KEYINPUT70), .ZN(n328) );
  XNOR2_X1 U325 ( .A(n329), .B(n328), .ZN(n333) );
  XNOR2_X1 U326 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U327 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U328 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U329 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U330 ( .A(n455), .B(G204GAT), .ZN(n456) );
  XNOR2_X1 U331 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U332 ( .A(n457), .B(n456), .ZN(G1353GAT) );
  XNOR2_X1 U333 ( .A(n478), .B(n477), .ZN(G1330GAT) );
  XOR2_X1 U334 ( .A(KEYINPUT81), .B(KEYINPUT82), .Z(n290) );
  XNOR2_X1 U335 ( .A(G190GAT), .B(KEYINPUT83), .ZN(n289) );
  XNOR2_X1 U336 ( .A(n290), .B(n289), .ZN(n291) );
  XOR2_X1 U337 ( .A(n291), .B(G99GAT), .Z(n293) );
  XOR2_X1 U338 ( .A(G15GAT), .B(G127GAT), .Z(n372) );
  XNOR2_X1 U339 ( .A(G43GAT), .B(n372), .ZN(n292) );
  XNOR2_X1 U340 ( .A(n293), .B(n292), .ZN(n299) );
  XOR2_X1 U341 ( .A(G120GAT), .B(G71GAT), .Z(n337) );
  XOR2_X1 U342 ( .A(KEYINPUT80), .B(KEYINPUT0), .Z(n295) );
  XNOR2_X1 U343 ( .A(G113GAT), .B(G134GAT), .ZN(n294) );
  XNOR2_X1 U344 ( .A(n295), .B(n294), .ZN(n441) );
  XOR2_X1 U345 ( .A(n337), .B(n441), .Z(n297) );
  NAND2_X1 U346 ( .A1(G227GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U347 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U348 ( .A(n299), .B(n298), .Z(n307) );
  XOR2_X1 U349 ( .A(KEYINPUT17), .B(KEYINPUT84), .Z(n301) );
  XNOR2_X1 U350 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n300) );
  XNOR2_X1 U351 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U352 ( .A(G169GAT), .B(n302), .Z(n421) );
  XOR2_X1 U353 ( .A(G176GAT), .B(KEYINPUT85), .Z(n304) );
  XNOR2_X1 U354 ( .A(G183GAT), .B(KEYINPUT20), .ZN(n303) );
  XNOR2_X1 U355 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U356 ( .A(n421), .B(n305), .ZN(n306) );
  XNOR2_X1 U357 ( .A(n307), .B(n306), .ZN(n531) );
  XOR2_X1 U358 ( .A(KEYINPUT86), .B(G218GAT), .Z(n309) );
  XNOR2_X1 U359 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n308) );
  XNOR2_X1 U360 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U361 ( .A(G197GAT), .B(n310), .Z(n417) );
  XOR2_X1 U362 ( .A(KEYINPUT3), .B(KEYINPUT2), .Z(n312) );
  XNOR2_X1 U363 ( .A(KEYINPUT87), .B(G155GAT), .ZN(n311) );
  XNOR2_X1 U364 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U365 ( .A(KEYINPUT88), .B(n313), .Z(n445) );
  XNOR2_X1 U366 ( .A(n417), .B(n445), .ZN(n325) );
  XOR2_X1 U367 ( .A(KEYINPUT22), .B(KEYINPUT23), .Z(n315) );
  XNOR2_X1 U368 ( .A(G204GAT), .B(KEYINPUT24), .ZN(n314) );
  XNOR2_X1 U369 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U370 ( .A(G50GAT), .B(G162GAT), .Z(n385) );
  XOR2_X1 U371 ( .A(n316), .B(n385), .Z(n323) );
  XOR2_X1 U372 ( .A(G141GAT), .B(G22GAT), .Z(n348) );
  XOR2_X1 U373 ( .A(G78GAT), .B(G148GAT), .Z(n318) );
  XNOR2_X1 U374 ( .A(G106GAT), .B(KEYINPUT71), .ZN(n317) );
  XNOR2_X1 U375 ( .A(n318), .B(n317), .ZN(n329) );
  XOR2_X1 U376 ( .A(KEYINPUT89), .B(n329), .Z(n320) );
  NAND2_X1 U377 ( .A1(G228GAT), .A2(G233GAT), .ZN(n319) );
  XNOR2_X1 U378 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U379 ( .A(n348), .B(n321), .ZN(n322) );
  XNOR2_X1 U380 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U381 ( .A(n325), .B(n324), .ZN(n479) );
  NOR2_X1 U382 ( .A1(n531), .A2(n479), .ZN(n326) );
  XOR2_X1 U383 ( .A(KEYINPUT26), .B(n326), .Z(n548) );
  INV_X1 U384 ( .A(n548), .ZN(n463) );
  AND2_X1 U385 ( .A1(G230GAT), .A2(G233GAT), .ZN(n327) );
  XOR2_X1 U386 ( .A(KEYINPUT32), .B(KEYINPUT31), .Z(n331) );
  XNOR2_X1 U387 ( .A(KEYINPUT33), .B(KEYINPUT72), .ZN(n330) );
  XOR2_X1 U388 ( .A(n331), .B(n330), .Z(n332) );
  XNOR2_X1 U389 ( .A(n333), .B(n332), .ZN(n340) );
  XOR2_X1 U390 ( .A(G64GAT), .B(G92GAT), .Z(n335) );
  XNOR2_X1 U391 ( .A(G176GAT), .B(G204GAT), .ZN(n334) );
  XNOR2_X1 U392 ( .A(n335), .B(n334), .ZN(n412) );
  XNOR2_X1 U393 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n336) );
  XNOR2_X1 U394 ( .A(n336), .B(KEYINPUT69), .ZN(n369) );
  XNOR2_X1 U395 ( .A(n412), .B(n369), .ZN(n338) );
  XOR2_X1 U396 ( .A(G99GAT), .B(G85GAT), .Z(n386) );
  XOR2_X1 U397 ( .A(n341), .B(n386), .Z(n404) );
  XNOR2_X1 U398 ( .A(n404), .B(KEYINPUT41), .ZN(n568) );
  INV_X1 U399 ( .A(n568), .ZN(n507) );
  XOR2_X1 U400 ( .A(KEYINPUT67), .B(G8GAT), .Z(n343) );
  XNOR2_X1 U401 ( .A(G113GAT), .B(G15GAT), .ZN(n342) );
  XNOR2_X1 U402 ( .A(n343), .B(n342), .ZN(n347) );
  XOR2_X1 U403 ( .A(KEYINPUT66), .B(KEYINPUT64), .Z(n345) );
  XNOR2_X1 U404 ( .A(KEYINPUT29), .B(KEYINPUT30), .ZN(n344) );
  XNOR2_X1 U405 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U406 ( .A(n347), .B(n346), .ZN(n360) );
  XOR2_X1 U407 ( .A(G50GAT), .B(G36GAT), .Z(n350) );
  XOR2_X1 U408 ( .A(G1GAT), .B(KEYINPUT68), .Z(n373) );
  XNOR2_X1 U409 ( .A(n348), .B(n373), .ZN(n349) );
  XNOR2_X1 U410 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U411 ( .A(n351), .B(G197GAT), .Z(n358) );
  XOR2_X1 U412 ( .A(G29GAT), .B(G43GAT), .Z(n353) );
  XNOR2_X1 U413 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n352) );
  XNOR2_X1 U414 ( .A(n353), .B(n352), .ZN(n388) );
  XOR2_X1 U415 ( .A(n388), .B(KEYINPUT65), .Z(n355) );
  NAND2_X1 U416 ( .A1(G229GAT), .A2(G233GAT), .ZN(n354) );
  XNOR2_X1 U417 ( .A(n355), .B(n354), .ZN(n356) );
  XNOR2_X1 U418 ( .A(G169GAT), .B(n356), .ZN(n357) );
  XNOR2_X1 U419 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U420 ( .A(n360), .B(n359), .ZN(n564) );
  INV_X1 U421 ( .A(n564), .ZN(n552) );
  NAND2_X1 U422 ( .A1(n507), .A2(n552), .ZN(n362) );
  XNOR2_X1 U423 ( .A(KEYINPUT46), .B(KEYINPUT111), .ZN(n361) );
  XNOR2_X1 U424 ( .A(n362), .B(n361), .ZN(n382) );
  XOR2_X1 U425 ( .A(KEYINPUT15), .B(KEYINPUT78), .Z(n364) );
  XNOR2_X1 U426 ( .A(G71GAT), .B(G64GAT), .ZN(n363) );
  XNOR2_X1 U427 ( .A(n364), .B(n363), .ZN(n381) );
  XOR2_X1 U428 ( .A(KEYINPUT14), .B(KEYINPUT77), .Z(n366) );
  NAND2_X1 U429 ( .A1(G231GAT), .A2(G233GAT), .ZN(n365) );
  XNOR2_X1 U430 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U431 ( .A(n367), .B(KEYINPUT12), .Z(n371) );
  XNOR2_X1 U432 ( .A(G8GAT), .B(G183GAT), .ZN(n368) );
  XNOR2_X1 U433 ( .A(n368), .B(KEYINPUT76), .ZN(n413) );
  XNOR2_X1 U434 ( .A(n413), .B(n369), .ZN(n370) );
  XNOR2_X1 U435 ( .A(n371), .B(n370), .ZN(n377) );
  XOR2_X1 U436 ( .A(G78GAT), .B(G155GAT), .Z(n375) );
  XNOR2_X1 U437 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U438 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U439 ( .A(n377), .B(n376), .Z(n379) );
  XNOR2_X1 U440 ( .A(G22GAT), .B(G211GAT), .ZN(n378) );
  XNOR2_X1 U441 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U442 ( .A(n381), .B(n380), .ZN(n574) );
  NOR2_X1 U443 ( .A1(n382), .A2(n574), .ZN(n383) );
  XNOR2_X1 U444 ( .A(KEYINPUT112), .B(n383), .ZN(n401) );
  XNOR2_X1 U445 ( .A(G36GAT), .B(G190GAT), .ZN(n384) );
  XNOR2_X1 U446 ( .A(n384), .B(KEYINPUT75), .ZN(n419) );
  XNOR2_X1 U447 ( .A(n385), .B(n419), .ZN(n387) );
  XNOR2_X1 U448 ( .A(n387), .B(n386), .ZN(n392) );
  XOR2_X1 U449 ( .A(G92GAT), .B(n388), .Z(n390) );
  NAND2_X1 U450 ( .A1(G232GAT), .A2(G233GAT), .ZN(n389) );
  XNOR2_X1 U451 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U452 ( .A(n392), .B(n391), .Z(n400) );
  XOR2_X1 U453 ( .A(KEYINPUT11), .B(KEYINPUT74), .Z(n394) );
  XNOR2_X1 U454 ( .A(G218GAT), .B(KEYINPUT73), .ZN(n393) );
  XNOR2_X1 U455 ( .A(n394), .B(n393), .ZN(n398) );
  XOR2_X1 U456 ( .A(KEYINPUT10), .B(KEYINPUT9), .Z(n396) );
  XNOR2_X1 U457 ( .A(G134GAT), .B(G106GAT), .ZN(n395) );
  XNOR2_X1 U458 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U459 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U460 ( .A(n400), .B(n399), .ZN(n542) );
  NAND2_X1 U461 ( .A1(n401), .A2(n542), .ZN(n403) );
  XNOR2_X1 U462 ( .A(KEYINPUT113), .B(KEYINPUT47), .ZN(n402) );
  XNOR2_X1 U463 ( .A(n403), .B(n402), .ZN(n410) );
  XOR2_X1 U464 ( .A(n542), .B(KEYINPUT36), .Z(n576) );
  NAND2_X1 U465 ( .A1(n574), .A2(n576), .ZN(n405) );
  XNOR2_X1 U466 ( .A(n405), .B(KEYINPUT114), .ZN(n406) );
  XNOR2_X1 U467 ( .A(n406), .B(KEYINPUT45), .ZN(n407) );
  NOR2_X1 U468 ( .A1(n404), .A2(n407), .ZN(n408) );
  NAND2_X1 U469 ( .A1(n408), .A2(n564), .ZN(n409) );
  NAND2_X1 U470 ( .A1(n410), .A2(n409), .ZN(n411) );
  XNOR2_X1 U471 ( .A(n411), .B(KEYINPUT48), .ZN(n549) );
  XNOR2_X1 U472 ( .A(n413), .B(n412), .ZN(n425) );
  XOR2_X1 U473 ( .A(KEYINPUT94), .B(KEYINPUT96), .Z(n415) );
  NAND2_X1 U474 ( .A1(G226GAT), .A2(G233GAT), .ZN(n414) );
  XNOR2_X1 U475 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U476 ( .A(n417), .B(n416), .ZN(n423) );
  XOR2_X1 U477 ( .A(KEYINPUT95), .B(KEYINPUT97), .Z(n418) );
  XNOR2_X1 U478 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U479 ( .A(n425), .B(n424), .ZN(n523) );
  NAND2_X1 U480 ( .A1(n549), .A2(n523), .ZN(n427) );
  XOR2_X1 U481 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n426) );
  XNOR2_X1 U482 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U483 ( .A(KEYINPUT92), .B(G148GAT), .Z(n430) );
  XNOR2_X1 U484 ( .A(G120GAT), .B(G127GAT), .ZN(n429) );
  XNOR2_X1 U485 ( .A(n430), .B(n429), .ZN(n434) );
  XOR2_X1 U486 ( .A(G85GAT), .B(G162GAT), .Z(n432) );
  XNOR2_X1 U487 ( .A(G29GAT), .B(G141GAT), .ZN(n431) );
  XNOR2_X1 U488 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U489 ( .A(n434), .B(n433), .ZN(n449) );
  XOR2_X1 U490 ( .A(KEYINPUT90), .B(KEYINPUT93), .Z(n436) );
  XNOR2_X1 U491 ( .A(G57GAT), .B(KEYINPUT5), .ZN(n435) );
  XNOR2_X1 U492 ( .A(n436), .B(n435), .ZN(n440) );
  XOR2_X1 U493 ( .A(KEYINPUT6), .B(KEYINPUT91), .Z(n438) );
  XNOR2_X1 U494 ( .A(KEYINPUT4), .B(KEYINPUT1), .ZN(n437) );
  XNOR2_X1 U495 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U496 ( .A(n440), .B(n439), .Z(n447) );
  XOR2_X1 U497 ( .A(n441), .B(G1GAT), .Z(n443) );
  NAND2_X1 U498 ( .A1(G225GAT), .A2(G233GAT), .ZN(n442) );
  XNOR2_X1 U499 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U500 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U501 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U502 ( .A(n449), .B(n448), .ZN(n521) );
  INV_X1 U503 ( .A(n521), .ZN(n480) );
  AND2_X1 U504 ( .A1(n288), .A2(n480), .ZN(n450) );
  NAND2_X1 U505 ( .A1(n463), .A2(n450), .ZN(n451) );
  XNOR2_X1 U506 ( .A(n451), .B(KEYINPUT125), .ZN(n577) );
  NAND2_X1 U507 ( .A1(n577), .A2(n552), .ZN(n454) );
  XOR2_X1 U508 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n452) );
  XNOR2_X1 U509 ( .A(n452), .B(G197GAT), .ZN(n453) );
  XNOR2_X1 U510 ( .A(n454), .B(n453), .ZN(G1352GAT) );
  NAND2_X1 U511 ( .A1(n577), .A2(n404), .ZN(n457) );
  XOR2_X1 U512 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n455) );
  XOR2_X1 U513 ( .A(n479), .B(KEYINPUT28), .Z(n526) );
  XNOR2_X1 U514 ( .A(n523), .B(KEYINPUT27), .ZN(n464) );
  NAND2_X1 U515 ( .A1(n521), .A2(n464), .ZN(n547) );
  NOR2_X1 U516 ( .A1(n526), .A2(n547), .ZN(n532) );
  XOR2_X1 U517 ( .A(n532), .B(KEYINPUT98), .Z(n458) );
  NOR2_X1 U518 ( .A1(n531), .A2(n458), .ZN(n470) );
  NAND2_X1 U519 ( .A1(n523), .A2(n531), .ZN(n460) );
  XNOR2_X1 U520 ( .A(n460), .B(n459), .ZN(n461) );
  NAND2_X1 U521 ( .A1(n479), .A2(n461), .ZN(n462) );
  XNOR2_X1 U522 ( .A(n462), .B(KEYINPUT25), .ZN(n466) );
  AND2_X1 U523 ( .A1(n464), .A2(n463), .ZN(n465) );
  NOR2_X1 U524 ( .A1(n466), .A2(n465), .ZN(n467) );
  XNOR2_X1 U525 ( .A(n468), .B(KEYINPUT100), .ZN(n469) );
  NOR2_X1 U526 ( .A1(n470), .A2(n469), .ZN(n471) );
  XOR2_X1 U527 ( .A(KEYINPUT101), .B(n471), .Z(n490) );
  NOR2_X1 U528 ( .A1(n574), .A2(n490), .ZN(n472) );
  NAND2_X1 U529 ( .A1(n576), .A2(n472), .ZN(n473) );
  XOR2_X1 U530 ( .A(KEYINPUT37), .B(n473), .Z(n520) );
  OR2_X1 U531 ( .A1(n564), .A2(n404), .ZN(n492) );
  OR2_X1 U532 ( .A1(n520), .A2(n492), .ZN(n474) );
  NAND2_X1 U533 ( .A1(n531), .A2(n504), .ZN(n478) );
  XOR2_X1 U534 ( .A(KEYINPUT40), .B(KEYINPUT104), .Z(n476) );
  XNOR2_X1 U535 ( .A(G43GAT), .B(KEYINPUT105), .ZN(n475) );
  AND2_X1 U536 ( .A1(n480), .A2(n479), .ZN(n481) );
  NAND2_X1 U537 ( .A1(n288), .A2(n481), .ZN(n482) );
  XNOR2_X1 U538 ( .A(n482), .B(KEYINPUT55), .ZN(n483) );
  NAND2_X1 U539 ( .A1(n483), .A2(n531), .ZN(n571) );
  NOR2_X1 U540 ( .A1(n542), .A2(n571), .ZN(n484) );
  XNOR2_X1 U541 ( .A(KEYINPUT58), .B(n484), .ZN(n486) );
  INV_X1 U542 ( .A(G190GAT), .ZN(n485) );
  XNOR2_X1 U543 ( .A(n486), .B(n485), .ZN(G1351GAT) );
  XNOR2_X1 U544 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n494) );
  XOR2_X1 U545 ( .A(KEYINPUT79), .B(KEYINPUT16), .Z(n488) );
  NAND2_X1 U546 ( .A1(n542), .A2(n574), .ZN(n487) );
  XNOR2_X1 U547 ( .A(n488), .B(n487), .ZN(n489) );
  NOR2_X1 U548 ( .A1(n490), .A2(n489), .ZN(n491) );
  XOR2_X1 U549 ( .A(KEYINPUT102), .B(n491), .Z(n508) );
  NOR2_X1 U550 ( .A1(n508), .A2(n492), .ZN(n499) );
  NAND2_X1 U551 ( .A1(n521), .A2(n499), .ZN(n493) );
  XNOR2_X1 U552 ( .A(n494), .B(n493), .ZN(G1324GAT) );
  NAND2_X1 U553 ( .A1(n499), .A2(n523), .ZN(n495) );
  XNOR2_X1 U554 ( .A(n495), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U555 ( .A(KEYINPUT103), .B(KEYINPUT35), .Z(n497) );
  NAND2_X1 U556 ( .A1(n499), .A2(n531), .ZN(n496) );
  XNOR2_X1 U557 ( .A(n497), .B(n496), .ZN(n498) );
  XOR2_X1 U558 ( .A(G15GAT), .B(n498), .Z(G1326GAT) );
  NAND2_X1 U559 ( .A1(n499), .A2(n526), .ZN(n500) );
  XNOR2_X1 U560 ( .A(n500), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U561 ( .A1(n521), .A2(n504), .ZN(n502) );
  XOR2_X1 U562 ( .A(G29GAT), .B(KEYINPUT39), .Z(n501) );
  XNOR2_X1 U563 ( .A(n502), .B(n501), .ZN(G1328GAT) );
  NAND2_X1 U564 ( .A1(n504), .A2(n523), .ZN(n503) );
  XNOR2_X1 U565 ( .A(n503), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U566 ( .A1(n504), .A2(n526), .ZN(n505) );
  XNOR2_X1 U567 ( .A(n505), .B(KEYINPUT106), .ZN(n506) );
  XNOR2_X1 U568 ( .A(G50GAT), .B(n506), .ZN(G1331GAT) );
  XNOR2_X1 U569 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n510) );
  NAND2_X1 U570 ( .A1(n564), .A2(n507), .ZN(n519) );
  NOR2_X1 U571 ( .A1(n508), .A2(n519), .ZN(n515) );
  NAND2_X1 U572 ( .A1(n521), .A2(n515), .ZN(n509) );
  XNOR2_X1 U573 ( .A(n510), .B(n509), .ZN(G1332GAT) );
  XOR2_X1 U574 ( .A(G64GAT), .B(KEYINPUT107), .Z(n512) );
  NAND2_X1 U575 ( .A1(n515), .A2(n523), .ZN(n511) );
  XNOR2_X1 U576 ( .A(n512), .B(n511), .ZN(G1333GAT) );
  NAND2_X1 U577 ( .A1(n515), .A2(n531), .ZN(n513) );
  XNOR2_X1 U578 ( .A(n513), .B(KEYINPUT108), .ZN(n514) );
  XNOR2_X1 U579 ( .A(G71GAT), .B(n514), .ZN(G1334GAT) );
  XOR2_X1 U580 ( .A(KEYINPUT109), .B(KEYINPUT43), .Z(n517) );
  NAND2_X1 U581 ( .A1(n515), .A2(n526), .ZN(n516) );
  XNOR2_X1 U582 ( .A(n517), .B(n516), .ZN(n518) );
  XOR2_X1 U583 ( .A(G78GAT), .B(n518), .Z(G1335GAT) );
  NOR2_X1 U584 ( .A1(n520), .A2(n519), .ZN(n527) );
  NAND2_X1 U585 ( .A1(n521), .A2(n527), .ZN(n522) );
  XNOR2_X1 U586 ( .A(G85GAT), .B(n522), .ZN(G1336GAT) );
  NAND2_X1 U587 ( .A1(n527), .A2(n523), .ZN(n524) );
  XNOR2_X1 U588 ( .A(n524), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U589 ( .A1(n527), .A2(n531), .ZN(n525) );
  XNOR2_X1 U590 ( .A(n525), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U591 ( .A(KEYINPUT44), .B(KEYINPUT110), .Z(n529) );
  NAND2_X1 U592 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U593 ( .A(n529), .B(n528), .ZN(n530) );
  XOR2_X1 U594 ( .A(G106GAT), .B(n530), .Z(G1339GAT) );
  INV_X1 U595 ( .A(n531), .ZN(n534) );
  NAND2_X1 U596 ( .A1(n549), .A2(n532), .ZN(n533) );
  NOR2_X1 U597 ( .A1(n534), .A2(n533), .ZN(n543) );
  NAND2_X1 U598 ( .A1(n543), .A2(n552), .ZN(n535) );
  XNOR2_X1 U599 ( .A(G113GAT), .B(n535), .ZN(G1340GAT) );
  XOR2_X1 U600 ( .A(G120GAT), .B(KEYINPUT49), .Z(n537) );
  NAND2_X1 U601 ( .A1(n543), .A2(n507), .ZN(n536) );
  XNOR2_X1 U602 ( .A(n537), .B(n536), .ZN(G1341GAT) );
  XNOR2_X1 U603 ( .A(G127GAT), .B(KEYINPUT115), .ZN(n541) );
  XOR2_X1 U604 ( .A(KEYINPUT116), .B(KEYINPUT50), .Z(n539) );
  NAND2_X1 U605 ( .A1(n543), .A2(n574), .ZN(n538) );
  XNOR2_X1 U606 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U607 ( .A(n541), .B(n540), .ZN(G1342GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT51), .B(KEYINPUT117), .Z(n545) );
  INV_X1 U609 ( .A(n542), .ZN(n562) );
  NAND2_X1 U610 ( .A1(n543), .A2(n562), .ZN(n544) );
  XNOR2_X1 U611 ( .A(n545), .B(n544), .ZN(n546) );
  XOR2_X1 U612 ( .A(G134GAT), .B(n546), .Z(G1343GAT) );
  XOR2_X1 U613 ( .A(G141GAT), .B(KEYINPUT119), .Z(n554) );
  NOR2_X1 U614 ( .A1(n548), .A2(n547), .ZN(n550) );
  NAND2_X1 U615 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U616 ( .A(KEYINPUT118), .B(n551), .Z(n561) );
  NAND2_X1 U617 ( .A1(n561), .A2(n552), .ZN(n553) );
  XNOR2_X1 U618 ( .A(n554), .B(n553), .ZN(G1344GAT) );
  XOR2_X1 U619 ( .A(KEYINPUT53), .B(KEYINPUT121), .Z(n556) );
  XNOR2_X1 U620 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n555) );
  XNOR2_X1 U621 ( .A(n556), .B(n555), .ZN(n557) );
  XOR2_X1 U622 ( .A(KEYINPUT120), .B(n557), .Z(n559) );
  NAND2_X1 U623 ( .A1(n561), .A2(n507), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n559), .B(n558), .ZN(G1345GAT) );
  NAND2_X1 U625 ( .A1(n561), .A2(n574), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n560), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U627 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U628 ( .A(G162GAT), .B(n563), .ZN(G1347GAT) );
  NOR2_X1 U629 ( .A1(n564), .A2(n571), .ZN(n565) );
  XOR2_X1 U630 ( .A(G169GAT), .B(n565), .Z(G1348GAT) );
  XOR2_X1 U631 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n567) );
  XNOR2_X1 U632 ( .A(G176GAT), .B(KEYINPUT124), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n567), .B(n566), .ZN(n570) );
  NOR2_X1 U634 ( .A1(n568), .A2(n571), .ZN(n569) );
  XOR2_X1 U635 ( .A(n570), .B(n569), .Z(G1349GAT) );
  INV_X1 U636 ( .A(n574), .ZN(n572) );
  NOR2_X1 U637 ( .A1(n572), .A2(n571), .ZN(n573) );
  XOR2_X1 U638 ( .A(G183GAT), .B(n573), .Z(G1350GAT) );
  NAND2_X1 U639 ( .A1(n574), .A2(n577), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n575), .B(G211GAT), .ZN(G1354GAT) );
  NAND2_X1 U641 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U642 ( .A(n578), .B(KEYINPUT62), .ZN(n579) );
  XNOR2_X1 U643 ( .A(G218GAT), .B(n579), .ZN(G1355GAT) );
endmodule

