

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U546 ( .A1(n639), .A2(n553), .ZN(n652) );
  OR2_X1 U547 ( .A1(KEYINPUT26), .A2(G1996), .ZN(n513) );
  XOR2_X1 U548 ( .A(n745), .B(KEYINPUT32), .Z(n514) );
  NAND2_X1 U549 ( .A1(n692), .A2(n691), .ZN(n712) );
  INV_X1 U550 ( .A(n736), .ZN(n720) );
  XNOR2_X1 U551 ( .A(n717), .B(KEYINPUT99), .ZN(n718) );
  NOR2_X1 U552 ( .A1(G164), .A2(G1384), .ZN(n777) );
  NOR2_X1 U553 ( .A1(n799), .A2(n754), .ZN(n755) );
  NOR2_X1 U554 ( .A1(G651), .A2(n639), .ZN(n647) );
  INV_X1 U555 ( .A(G2105), .ZN(n518) );
  AND2_X2 U556 ( .A1(n518), .A2(G2104), .ZN(n886) );
  NAND2_X1 U557 ( .A1(G102), .A2(n886), .ZN(n517) );
  NOR2_X1 U558 ( .A1(G2104), .A2(G2105), .ZN(n515) );
  XOR2_X2 U559 ( .A(n515), .B(KEYINPUT17), .Z(n878) );
  NAND2_X1 U560 ( .A1(G138), .A2(n878), .ZN(n516) );
  NAND2_X1 U561 ( .A1(n517), .A2(n516), .ZN(n522) );
  AND2_X1 U562 ( .A1(G2104), .A2(G2105), .ZN(n880) );
  NAND2_X1 U563 ( .A1(G114), .A2(n880), .ZN(n520) );
  NOR2_X1 U564 ( .A1(G2104), .A2(n518), .ZN(n881) );
  NAND2_X1 U565 ( .A1(G126), .A2(n881), .ZN(n519) );
  NAND2_X1 U566 ( .A1(n520), .A2(n519), .ZN(n521) );
  NOR2_X1 U567 ( .A1(n522), .A2(n521), .ZN(G164) );
  NAND2_X1 U568 ( .A1(n878), .A2(G137), .ZN(n525) );
  NAND2_X1 U569 ( .A1(G101), .A2(n886), .ZN(n523) );
  XOR2_X1 U570 ( .A(KEYINPUT23), .B(n523), .Z(n524) );
  NAND2_X1 U571 ( .A1(n525), .A2(n524), .ZN(n529) );
  NAND2_X1 U572 ( .A1(G113), .A2(n880), .ZN(n527) );
  NAND2_X1 U573 ( .A1(G125), .A2(n881), .ZN(n526) );
  NAND2_X1 U574 ( .A1(n527), .A2(n526), .ZN(n528) );
  NOR2_X1 U575 ( .A1(n529), .A2(n528), .ZN(G160) );
  XOR2_X1 U576 ( .A(KEYINPUT107), .B(G2435), .Z(n531) );
  XNOR2_X1 U577 ( .A(G2430), .B(G2438), .ZN(n530) );
  XNOR2_X1 U578 ( .A(n531), .B(n530), .ZN(n538) );
  XOR2_X1 U579 ( .A(G2446), .B(G2454), .Z(n533) );
  XNOR2_X1 U580 ( .A(G2451), .B(G2443), .ZN(n532) );
  XNOR2_X1 U581 ( .A(n533), .B(n532), .ZN(n534) );
  XOR2_X1 U582 ( .A(n534), .B(G2427), .Z(n536) );
  XNOR2_X1 U583 ( .A(G1341), .B(G1348), .ZN(n535) );
  XNOR2_X1 U584 ( .A(n536), .B(n535), .ZN(n537) );
  XNOR2_X1 U585 ( .A(n538), .B(n537), .ZN(n539) );
  AND2_X1 U586 ( .A1(n539), .A2(G14), .ZN(G401) );
  AND2_X1 U587 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U588 ( .A1(G123), .A2(n881), .ZN(n540) );
  XNOR2_X1 U589 ( .A(n540), .B(KEYINPUT18), .ZN(n547) );
  NAND2_X1 U590 ( .A1(G99), .A2(n886), .ZN(n542) );
  NAND2_X1 U591 ( .A1(G135), .A2(n878), .ZN(n541) );
  NAND2_X1 U592 ( .A1(n542), .A2(n541), .ZN(n545) );
  NAND2_X1 U593 ( .A1(n880), .A2(G111), .ZN(n543) );
  XOR2_X1 U594 ( .A(KEYINPUT80), .B(n543), .Z(n544) );
  NOR2_X1 U595 ( .A1(n545), .A2(n544), .ZN(n546) );
  NAND2_X1 U596 ( .A1(n547), .A2(n546), .ZN(n965) );
  XNOR2_X1 U597 ( .A(G2096), .B(n965), .ZN(n548) );
  OR2_X1 U598 ( .A1(G2100), .A2(n548), .ZN(G156) );
  INV_X1 U599 ( .A(G57), .ZN(G237) );
  INV_X1 U600 ( .A(G108), .ZN(G238) );
  INV_X1 U601 ( .A(G132), .ZN(G219) );
  INV_X1 U602 ( .A(G82), .ZN(G220) );
  XOR2_X1 U603 ( .A(G543), .B(KEYINPUT0), .Z(n639) );
  NAND2_X1 U604 ( .A1(n647), .A2(G52), .ZN(n552) );
  INV_X1 U605 ( .A(G651), .ZN(n553) );
  NOR2_X1 U606 ( .A1(G543), .A2(n553), .ZN(n550) );
  XNOR2_X1 U607 ( .A(KEYINPUT65), .B(KEYINPUT1), .ZN(n549) );
  XNOR2_X2 U608 ( .A(n550), .B(n549), .ZN(n646) );
  NAND2_X1 U609 ( .A1(n646), .A2(G64), .ZN(n551) );
  NAND2_X1 U610 ( .A1(n552), .A2(n551), .ZN(n559) );
  NOR2_X1 U611 ( .A1(G651), .A2(G543), .ZN(n651) );
  NAND2_X1 U612 ( .A1(G90), .A2(n651), .ZN(n555) );
  NAND2_X1 U613 ( .A1(G77), .A2(n652), .ZN(n554) );
  NAND2_X1 U614 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U615 ( .A(KEYINPUT67), .B(n556), .ZN(n557) );
  XNOR2_X1 U616 ( .A(KEYINPUT9), .B(n557), .ZN(n558) );
  NOR2_X1 U617 ( .A1(n559), .A2(n558), .ZN(G171) );
  INV_X1 U618 ( .A(G171), .ZN(G301) );
  NAND2_X1 U619 ( .A1(n646), .A2(G63), .ZN(n560) );
  XNOR2_X1 U620 ( .A(KEYINPUT77), .B(n560), .ZN(n563) );
  NAND2_X1 U621 ( .A1(n647), .A2(G51), .ZN(n561) );
  XOR2_X1 U622 ( .A(KEYINPUT78), .B(n561), .Z(n562) );
  NOR2_X1 U623 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U624 ( .A(KEYINPUT6), .B(n564), .ZN(n571) );
  XNOR2_X1 U625 ( .A(KEYINPUT76), .B(KEYINPUT5), .ZN(n569) );
  NAND2_X1 U626 ( .A1(n651), .A2(G89), .ZN(n565) );
  XNOR2_X1 U627 ( .A(n565), .B(KEYINPUT4), .ZN(n567) );
  NAND2_X1 U628 ( .A1(G76), .A2(n652), .ZN(n566) );
  NAND2_X1 U629 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U630 ( .A(n569), .B(n568), .ZN(n570) );
  NAND2_X1 U631 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U632 ( .A(n572), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U633 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U634 ( .A1(G7), .A2(G661), .ZN(n573) );
  XNOR2_X1 U635 ( .A(n573), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U636 ( .A(G223), .ZN(n830) );
  NAND2_X1 U637 ( .A1(n830), .A2(G567), .ZN(n574) );
  XOR2_X1 U638 ( .A(KEYINPUT11), .B(n574), .Z(G234) );
  NAND2_X1 U639 ( .A1(G56), .A2(n646), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n575), .B(KEYINPUT14), .ZN(n576) );
  XNOR2_X1 U641 ( .A(KEYINPUT69), .B(n576), .ZN(n584) );
  NAND2_X1 U642 ( .A1(n652), .A2(G68), .ZN(n577) );
  XNOR2_X1 U643 ( .A(KEYINPUT71), .B(n577), .ZN(n581) );
  XOR2_X1 U644 ( .A(KEYINPUT12), .B(KEYINPUT70), .Z(n579) );
  NAND2_X1 U645 ( .A1(G81), .A2(n651), .ZN(n578) );
  XNOR2_X1 U646 ( .A(n579), .B(n578), .ZN(n580) );
  NOR2_X1 U647 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U648 ( .A(KEYINPUT13), .B(n582), .ZN(n583) );
  NOR2_X1 U649 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U650 ( .A(n585), .B(KEYINPUT72), .ZN(n587) );
  NAND2_X1 U651 ( .A1(G43), .A2(n647), .ZN(n586) );
  NAND2_X1 U652 ( .A1(n587), .A2(n586), .ZN(n934) );
  INV_X1 U653 ( .A(G860), .ZN(n617) );
  OR2_X1 U654 ( .A1(n934), .A2(n617), .ZN(G153) );
  NAND2_X1 U655 ( .A1(G66), .A2(n646), .ZN(n588) );
  XNOR2_X1 U656 ( .A(n588), .B(KEYINPUT73), .ZN(n590) );
  AND2_X1 U657 ( .A1(n647), .A2(G54), .ZN(n589) );
  NOR2_X1 U658 ( .A1(n590), .A2(n589), .ZN(n594) );
  NAND2_X1 U659 ( .A1(G92), .A2(n651), .ZN(n592) );
  NAND2_X1 U660 ( .A1(G79), .A2(n652), .ZN(n591) );
  AND2_X1 U661 ( .A1(n592), .A2(n591), .ZN(n593) );
  AND2_X1 U662 ( .A1(n594), .A2(n593), .ZN(n595) );
  XNOR2_X1 U663 ( .A(n595), .B(KEYINPUT15), .ZN(n596) );
  XNOR2_X2 U664 ( .A(n596), .B(KEYINPUT74), .ZN(n948) );
  INV_X1 U665 ( .A(n948), .ZN(n615) );
  NOR2_X1 U666 ( .A1(G868), .A2(n615), .ZN(n597) );
  XNOR2_X1 U667 ( .A(n597), .B(KEYINPUT75), .ZN(n599) );
  NAND2_X1 U668 ( .A1(G868), .A2(G301), .ZN(n598) );
  NAND2_X1 U669 ( .A1(n599), .A2(n598), .ZN(G284) );
  NAND2_X1 U670 ( .A1(G65), .A2(n646), .ZN(n601) );
  NAND2_X1 U671 ( .A1(G53), .A2(n647), .ZN(n600) );
  NAND2_X1 U672 ( .A1(n601), .A2(n600), .ZN(n602) );
  XOR2_X1 U673 ( .A(KEYINPUT68), .B(n602), .Z(n606) );
  NAND2_X1 U674 ( .A1(G91), .A2(n651), .ZN(n604) );
  NAND2_X1 U675 ( .A1(G78), .A2(n652), .ZN(n603) );
  AND2_X1 U676 ( .A1(n604), .A2(n603), .ZN(n605) );
  NAND2_X1 U677 ( .A1(n606), .A2(n605), .ZN(G299) );
  INV_X1 U678 ( .A(G868), .ZN(n666) );
  NOR2_X1 U679 ( .A1(G286), .A2(n666), .ZN(n608) );
  NOR2_X1 U680 ( .A1(G868), .A2(G299), .ZN(n607) );
  NOR2_X1 U681 ( .A1(n608), .A2(n607), .ZN(G297) );
  NAND2_X1 U682 ( .A1(n617), .A2(G559), .ZN(n609) );
  NAND2_X1 U683 ( .A1(n609), .A2(n615), .ZN(n610) );
  XNOR2_X1 U684 ( .A(n610), .B(KEYINPUT16), .ZN(n611) );
  XOR2_X1 U685 ( .A(KEYINPUT79), .B(n611), .Z(G148) );
  NOR2_X1 U686 ( .A1(G868), .A2(n934), .ZN(n614) );
  NAND2_X1 U687 ( .A1(n615), .A2(G868), .ZN(n612) );
  NOR2_X1 U688 ( .A1(G559), .A2(n612), .ZN(n613) );
  NOR2_X1 U689 ( .A1(n614), .A2(n613), .ZN(G282) );
  NAND2_X1 U690 ( .A1(n615), .A2(G559), .ZN(n616) );
  XOR2_X1 U691 ( .A(n934), .B(n616), .Z(n664) );
  NAND2_X1 U692 ( .A1(n617), .A2(n664), .ZN(n625) );
  NAND2_X1 U693 ( .A1(G67), .A2(n646), .ZN(n619) );
  NAND2_X1 U694 ( .A1(G93), .A2(n651), .ZN(n618) );
  NAND2_X1 U695 ( .A1(n619), .A2(n618), .ZN(n622) );
  NAND2_X1 U696 ( .A1(G80), .A2(n652), .ZN(n620) );
  XNOR2_X1 U697 ( .A(KEYINPUT81), .B(n620), .ZN(n621) );
  NOR2_X1 U698 ( .A1(n622), .A2(n621), .ZN(n624) );
  NAND2_X1 U699 ( .A1(n647), .A2(G55), .ZN(n623) );
  NAND2_X1 U700 ( .A1(n624), .A2(n623), .ZN(n667) );
  XNOR2_X1 U701 ( .A(n625), .B(n667), .ZN(G145) );
  NAND2_X1 U702 ( .A1(G88), .A2(n651), .ZN(n627) );
  NAND2_X1 U703 ( .A1(G75), .A2(n652), .ZN(n626) );
  NAND2_X1 U704 ( .A1(n627), .A2(n626), .ZN(n631) );
  NAND2_X1 U705 ( .A1(G62), .A2(n646), .ZN(n629) );
  NAND2_X1 U706 ( .A1(G50), .A2(n647), .ZN(n628) );
  NAND2_X1 U707 ( .A1(n629), .A2(n628), .ZN(n630) );
  NOR2_X1 U708 ( .A1(n631), .A2(n630), .ZN(G166) );
  NAND2_X1 U709 ( .A1(G61), .A2(n646), .ZN(n633) );
  NAND2_X1 U710 ( .A1(G86), .A2(n651), .ZN(n632) );
  NAND2_X1 U711 ( .A1(n633), .A2(n632), .ZN(n636) );
  NAND2_X1 U712 ( .A1(n652), .A2(G73), .ZN(n634) );
  XOR2_X1 U713 ( .A(KEYINPUT2), .B(n634), .Z(n635) );
  NOR2_X1 U714 ( .A1(n636), .A2(n635), .ZN(n638) );
  NAND2_X1 U715 ( .A1(n647), .A2(G48), .ZN(n637) );
  NAND2_X1 U716 ( .A1(n638), .A2(n637), .ZN(G305) );
  NAND2_X1 U717 ( .A1(G74), .A2(G651), .ZN(n644) );
  NAND2_X1 U718 ( .A1(G49), .A2(n647), .ZN(n641) );
  NAND2_X1 U719 ( .A1(G87), .A2(n639), .ZN(n640) );
  NAND2_X1 U720 ( .A1(n641), .A2(n640), .ZN(n642) );
  NOR2_X1 U721 ( .A1(n646), .A2(n642), .ZN(n643) );
  NAND2_X1 U722 ( .A1(n644), .A2(n643), .ZN(n645) );
  XNOR2_X1 U723 ( .A(n645), .B(KEYINPUT82), .ZN(G288) );
  NAND2_X1 U724 ( .A1(G60), .A2(n646), .ZN(n649) );
  NAND2_X1 U725 ( .A1(G47), .A2(n647), .ZN(n648) );
  NAND2_X1 U726 ( .A1(n649), .A2(n648), .ZN(n650) );
  XOR2_X1 U727 ( .A(KEYINPUT66), .B(n650), .Z(n656) );
  NAND2_X1 U728 ( .A1(G85), .A2(n651), .ZN(n654) );
  NAND2_X1 U729 ( .A1(G72), .A2(n652), .ZN(n653) );
  AND2_X1 U730 ( .A1(n654), .A2(n653), .ZN(n655) );
  NAND2_X1 U731 ( .A1(n656), .A2(n655), .ZN(G290) );
  XOR2_X1 U732 ( .A(G305), .B(n667), .Z(n657) );
  XNOR2_X1 U733 ( .A(G166), .B(n657), .ZN(n661) );
  XOR2_X1 U734 ( .A(KEYINPUT84), .B(KEYINPUT83), .Z(n659) );
  XNOR2_X1 U735 ( .A(G288), .B(KEYINPUT19), .ZN(n658) );
  XNOR2_X1 U736 ( .A(n659), .B(n658), .ZN(n660) );
  XNOR2_X1 U737 ( .A(n661), .B(n660), .ZN(n662) );
  XNOR2_X1 U738 ( .A(n662), .B(G299), .ZN(n663) );
  XNOR2_X1 U739 ( .A(n663), .B(G290), .ZN(n836) );
  XNOR2_X1 U740 ( .A(n664), .B(n836), .ZN(n665) );
  NAND2_X1 U741 ( .A1(n665), .A2(G868), .ZN(n669) );
  NAND2_X1 U742 ( .A1(n667), .A2(n666), .ZN(n668) );
  NAND2_X1 U743 ( .A1(n669), .A2(n668), .ZN(G295) );
  NAND2_X1 U744 ( .A1(G2078), .A2(G2084), .ZN(n670) );
  XNOR2_X1 U745 ( .A(n670), .B(KEYINPUT85), .ZN(n671) );
  XNOR2_X1 U746 ( .A(n671), .B(KEYINPUT20), .ZN(n672) );
  NAND2_X1 U747 ( .A1(n672), .A2(G2090), .ZN(n673) );
  XNOR2_X1 U748 ( .A(KEYINPUT21), .B(n673), .ZN(n674) );
  NAND2_X1 U749 ( .A1(n674), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U750 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U751 ( .A1(G220), .A2(G219), .ZN(n675) );
  XNOR2_X1 U752 ( .A(KEYINPUT22), .B(n675), .ZN(n676) );
  NAND2_X1 U753 ( .A1(n676), .A2(G96), .ZN(n677) );
  NOR2_X1 U754 ( .A1(G218), .A2(n677), .ZN(n678) );
  XOR2_X1 U755 ( .A(KEYINPUT86), .B(n678), .Z(n835) );
  NAND2_X1 U756 ( .A1(n835), .A2(G2106), .ZN(n679) );
  XNOR2_X1 U757 ( .A(KEYINPUT87), .B(n679), .ZN(n686) );
  NAND2_X1 U758 ( .A1(G120), .A2(G69), .ZN(n680) );
  NOR2_X1 U759 ( .A1(G237), .A2(n680), .ZN(n681) );
  XOR2_X1 U760 ( .A(KEYINPUT88), .B(n681), .Z(n682) );
  NOR2_X1 U761 ( .A1(G238), .A2(n682), .ZN(n683) );
  XNOR2_X1 U762 ( .A(KEYINPUT89), .B(n683), .ZN(n834) );
  NAND2_X1 U763 ( .A1(G567), .A2(n834), .ZN(n684) );
  XOR2_X1 U764 ( .A(KEYINPUT90), .B(n684), .Z(n685) );
  NOR2_X1 U765 ( .A1(n686), .A2(n685), .ZN(G319) );
  INV_X1 U766 ( .A(G319), .ZN(n907) );
  NAND2_X1 U767 ( .A1(G483), .A2(G661), .ZN(n687) );
  NOR2_X1 U768 ( .A1(n907), .A2(n687), .ZN(n833) );
  NAND2_X1 U769 ( .A1(n833), .A2(G36), .ZN(G176) );
  XNOR2_X1 U770 ( .A(KEYINPUT91), .B(G166), .ZN(G303) );
  AND2_X1 U771 ( .A1(G160), .A2(G40), .ZN(n688) );
  NAND2_X1 U772 ( .A1(n777), .A2(n688), .ZN(n736) );
  NAND2_X1 U773 ( .A1(G8), .A2(n736), .ZN(n799) );
  NAND2_X1 U774 ( .A1(G1976), .A2(G288), .ZN(n941) );
  NOR2_X1 U775 ( .A1(G1976), .A2(G288), .ZN(n790) );
  NOR2_X1 U776 ( .A1(G1971), .A2(G303), .ZN(n689) );
  NOR2_X1 U777 ( .A1(n790), .A2(n689), .ZN(n942) );
  INV_X1 U778 ( .A(n942), .ZN(n752) );
  NAND2_X1 U779 ( .A1(n720), .A2(G2072), .ZN(n690) );
  XOR2_X1 U780 ( .A(KEYINPUT27), .B(n690), .Z(n692) );
  NAND2_X1 U781 ( .A1(G1956), .A2(n736), .ZN(n691) );
  NOR2_X1 U782 ( .A1(n712), .A2(G299), .ZN(n693) );
  XNOR2_X1 U783 ( .A(KEYINPUT97), .B(n693), .ZN(n711) );
  NAND2_X1 U784 ( .A1(n948), .A2(G2067), .ZN(n696) );
  NAND2_X1 U785 ( .A1(G1996), .A2(KEYINPUT26), .ZN(n694) );
  AND2_X1 U786 ( .A1(n694), .A2(n513), .ZN(n695) );
  NAND2_X1 U787 ( .A1(n696), .A2(n695), .ZN(n697) );
  AND2_X1 U788 ( .A1(n697), .A2(n720), .ZN(n698) );
  OR2_X1 U789 ( .A1(n698), .A2(n934), .ZN(n704) );
  AND2_X1 U790 ( .A1(G1348), .A2(n948), .ZN(n701) );
  INV_X1 U791 ( .A(G1341), .ZN(n699) );
  NAND2_X1 U792 ( .A1(KEYINPUT26), .A2(n699), .ZN(n700) );
  NOR2_X1 U793 ( .A1(n701), .A2(n700), .ZN(n702) );
  NOR2_X1 U794 ( .A1(n702), .A2(n720), .ZN(n703) );
  NOR2_X1 U795 ( .A1(n704), .A2(n703), .ZN(n709) );
  NAND2_X1 U796 ( .A1(G1348), .A2(n736), .ZN(n706) );
  NAND2_X1 U797 ( .A1(G2067), .A2(n720), .ZN(n705) );
  NAND2_X1 U798 ( .A1(n706), .A2(n705), .ZN(n707) );
  NOR2_X1 U799 ( .A1(n948), .A2(n707), .ZN(n708) );
  NOR2_X1 U800 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U801 ( .A1(n711), .A2(n710), .ZN(n716) );
  NAND2_X1 U802 ( .A1(n712), .A2(G299), .ZN(n713) );
  XNOR2_X1 U803 ( .A(n713), .B(KEYINPUT96), .ZN(n714) );
  XNOR2_X1 U804 ( .A(n714), .B(KEYINPUT28), .ZN(n715) );
  NAND2_X1 U805 ( .A1(n716), .A2(n715), .ZN(n719) );
  XOR2_X1 U806 ( .A(KEYINPUT29), .B(KEYINPUT98), .Z(n717) );
  XNOR2_X1 U807 ( .A(n719), .B(n718), .ZN(n724) );
  NAND2_X1 U808 ( .A1(G1961), .A2(n736), .ZN(n722) );
  XOR2_X1 U809 ( .A(KEYINPUT25), .B(G2078), .Z(n998) );
  NAND2_X1 U810 ( .A1(n720), .A2(n998), .ZN(n721) );
  NAND2_X1 U811 ( .A1(n722), .A2(n721), .ZN(n725) );
  NOR2_X1 U812 ( .A1(G301), .A2(n725), .ZN(n723) );
  NOR2_X1 U813 ( .A1(n724), .A2(n723), .ZN(n734) );
  NAND2_X1 U814 ( .A1(G301), .A2(n725), .ZN(n726) );
  XOR2_X1 U815 ( .A(KEYINPUT100), .B(n726), .Z(n731) );
  NOR2_X1 U816 ( .A1(G1966), .A2(n799), .ZN(n750) );
  NOR2_X1 U817 ( .A1(G2084), .A2(n736), .ZN(n747) );
  NOR2_X1 U818 ( .A1(n750), .A2(n747), .ZN(n727) );
  NAND2_X1 U819 ( .A1(G8), .A2(n727), .ZN(n728) );
  XNOR2_X1 U820 ( .A(KEYINPUT30), .B(n728), .ZN(n729) );
  NOR2_X1 U821 ( .A1(G168), .A2(n729), .ZN(n730) );
  NOR2_X1 U822 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U823 ( .A(n732), .B(KEYINPUT31), .ZN(n733) );
  NOR2_X1 U824 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U825 ( .A(n735), .B(KEYINPUT101), .ZN(n746) );
  NAND2_X1 U826 ( .A1(n746), .A2(G286), .ZN(n744) );
  INV_X1 U827 ( .A(G8), .ZN(n742) );
  NOR2_X1 U828 ( .A1(G2090), .A2(n736), .ZN(n737) );
  XNOR2_X1 U829 ( .A(n737), .B(KEYINPUT102), .ZN(n739) );
  NOR2_X1 U830 ( .A1(n799), .A2(G1971), .ZN(n738) );
  NOR2_X1 U831 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U832 ( .A1(n740), .A2(G303), .ZN(n741) );
  OR2_X1 U833 ( .A1(n742), .A2(n741), .ZN(n743) );
  AND2_X1 U834 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U835 ( .A1(G8), .A2(n747), .ZN(n748) );
  NAND2_X1 U836 ( .A1(n746), .A2(n748), .ZN(n749) );
  NOR2_X1 U837 ( .A1(n750), .A2(n749), .ZN(n751) );
  NOR2_X1 U838 ( .A1(n514), .A2(n751), .ZN(n803) );
  OR2_X1 U839 ( .A1(n752), .A2(n803), .ZN(n753) );
  NAND2_X1 U840 ( .A1(n941), .A2(n753), .ZN(n754) );
  XNOR2_X1 U841 ( .A(n755), .B(KEYINPUT64), .ZN(n756) );
  OR2_X1 U842 ( .A1(n756), .A2(KEYINPUT33), .ZN(n795) );
  XNOR2_X1 U843 ( .A(G1981), .B(KEYINPUT103), .ZN(n757) );
  XNOR2_X1 U844 ( .A(n757), .B(G305), .ZN(n935) );
  XOR2_X1 U845 ( .A(G1986), .B(G290), .Z(n952) );
  NAND2_X1 U846 ( .A1(G95), .A2(n886), .ZN(n759) );
  NAND2_X1 U847 ( .A1(G131), .A2(n878), .ZN(n758) );
  NAND2_X1 U848 ( .A1(n759), .A2(n758), .ZN(n764) );
  NAND2_X1 U849 ( .A1(G107), .A2(n880), .ZN(n761) );
  NAND2_X1 U850 ( .A1(G119), .A2(n881), .ZN(n760) );
  NAND2_X1 U851 ( .A1(n761), .A2(n760), .ZN(n762) );
  XOR2_X1 U852 ( .A(KEYINPUT93), .B(n762), .Z(n763) );
  NOR2_X1 U853 ( .A1(n764), .A2(n763), .ZN(n899) );
  INV_X1 U854 ( .A(G1991), .ZN(n996) );
  NOR2_X1 U855 ( .A1(n899), .A2(n996), .ZN(n775) );
  NAND2_X1 U856 ( .A1(n878), .A2(G141), .ZN(n765) );
  XNOR2_X1 U857 ( .A(KEYINPUT95), .B(n765), .ZN(n773) );
  NAND2_X1 U858 ( .A1(G117), .A2(n880), .ZN(n767) );
  NAND2_X1 U859 ( .A1(G129), .A2(n881), .ZN(n766) );
  NAND2_X1 U860 ( .A1(n767), .A2(n766), .ZN(n770) );
  NAND2_X1 U861 ( .A1(n886), .A2(G105), .ZN(n768) );
  XOR2_X1 U862 ( .A(KEYINPUT38), .B(n768), .Z(n769) );
  NOR2_X1 U863 ( .A1(n770), .A2(n769), .ZN(n771) );
  XOR2_X1 U864 ( .A(KEYINPUT94), .B(n771), .Z(n772) );
  NOR2_X1 U865 ( .A1(n773), .A2(n772), .ZN(n898) );
  INV_X1 U866 ( .A(G1996), .ZN(n993) );
  NOR2_X1 U867 ( .A1(n898), .A2(n993), .ZN(n774) );
  NOR2_X1 U868 ( .A1(n775), .A2(n774), .ZN(n970) );
  NAND2_X1 U869 ( .A1(n952), .A2(n970), .ZN(n778) );
  NAND2_X1 U870 ( .A1(G160), .A2(G40), .ZN(n776) );
  NOR2_X1 U871 ( .A1(n777), .A2(n776), .ZN(n822) );
  NAND2_X1 U872 ( .A1(n778), .A2(n822), .ZN(n789) );
  NAND2_X1 U873 ( .A1(n886), .A2(G104), .ZN(n779) );
  XNOR2_X1 U874 ( .A(n779), .B(KEYINPUT92), .ZN(n781) );
  NAND2_X1 U875 ( .A1(G140), .A2(n878), .ZN(n780) );
  NAND2_X1 U876 ( .A1(n781), .A2(n780), .ZN(n782) );
  XNOR2_X1 U877 ( .A(KEYINPUT34), .B(n782), .ZN(n787) );
  NAND2_X1 U878 ( .A1(G116), .A2(n880), .ZN(n784) );
  NAND2_X1 U879 ( .A1(G128), .A2(n881), .ZN(n783) );
  NAND2_X1 U880 ( .A1(n784), .A2(n783), .ZN(n785) );
  XOR2_X1 U881 ( .A(KEYINPUT35), .B(n785), .Z(n786) );
  NOR2_X1 U882 ( .A1(n787), .A2(n786), .ZN(n788) );
  XOR2_X1 U883 ( .A(KEYINPUT36), .B(n788), .Z(n902) );
  XOR2_X1 U884 ( .A(G2067), .B(KEYINPUT37), .Z(n820) );
  AND2_X1 U885 ( .A1(n902), .A2(n820), .ZN(n976) );
  NAND2_X1 U886 ( .A1(n976), .A2(n822), .ZN(n810) );
  AND2_X1 U887 ( .A1(n789), .A2(n810), .ZN(n796) );
  NAND2_X1 U888 ( .A1(n935), .A2(n796), .ZN(n793) );
  NAND2_X1 U889 ( .A1(n790), .A2(KEYINPUT33), .ZN(n791) );
  NOR2_X1 U890 ( .A1(n799), .A2(n791), .ZN(n792) );
  NOR2_X1 U891 ( .A1(n793), .A2(n792), .ZN(n794) );
  NAND2_X1 U892 ( .A1(n795), .A2(n794), .ZN(n828) );
  INV_X1 U893 ( .A(n796), .ZN(n809) );
  NOR2_X1 U894 ( .A1(G1981), .A2(G305), .ZN(n797) );
  XOR2_X1 U895 ( .A(n797), .B(KEYINPUT24), .Z(n798) );
  NOR2_X1 U896 ( .A1(n799), .A2(n798), .ZN(n807) );
  INV_X1 U897 ( .A(n799), .ZN(n805) );
  NOR2_X1 U898 ( .A1(G2090), .A2(G303), .ZN(n800) );
  NAND2_X1 U899 ( .A1(G8), .A2(n800), .ZN(n801) );
  XOR2_X1 U900 ( .A(KEYINPUT104), .B(n801), .Z(n802) );
  NOR2_X1 U901 ( .A1(n803), .A2(n802), .ZN(n804) );
  NOR2_X1 U902 ( .A1(n805), .A2(n804), .ZN(n806) );
  NOR2_X1 U903 ( .A1(n807), .A2(n806), .ZN(n808) );
  NOR2_X1 U904 ( .A1(n809), .A2(n808), .ZN(n826) );
  INV_X1 U905 ( .A(n810), .ZN(n819) );
  AND2_X1 U906 ( .A1(n993), .A2(n898), .ZN(n963) );
  INV_X1 U907 ( .A(n970), .ZN(n814) );
  NOR2_X1 U908 ( .A1(G1986), .A2(G290), .ZN(n811) );
  AND2_X1 U909 ( .A1(n996), .A2(n899), .ZN(n968) );
  NOR2_X1 U910 ( .A1(n811), .A2(n968), .ZN(n812) );
  XOR2_X1 U911 ( .A(KEYINPUT105), .B(n812), .Z(n813) );
  NOR2_X1 U912 ( .A1(n814), .A2(n813), .ZN(n815) );
  NOR2_X1 U913 ( .A1(n963), .A2(n815), .ZN(n816) );
  XNOR2_X1 U914 ( .A(KEYINPUT39), .B(n816), .ZN(n817) );
  NAND2_X1 U915 ( .A1(n817), .A2(n822), .ZN(n818) );
  OR2_X1 U916 ( .A1(n819), .A2(n818), .ZN(n824) );
  NOR2_X1 U917 ( .A1(n902), .A2(n820), .ZN(n821) );
  XNOR2_X1 U918 ( .A(KEYINPUT106), .B(n821), .ZN(n972) );
  NAND2_X1 U919 ( .A1(n972), .A2(n822), .ZN(n823) );
  NAND2_X1 U920 ( .A1(n824), .A2(n823), .ZN(n825) );
  NOR2_X1 U921 ( .A1(n826), .A2(n825), .ZN(n827) );
  NAND2_X1 U922 ( .A1(n828), .A2(n827), .ZN(n829) );
  XNOR2_X1 U923 ( .A(n829), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U924 ( .A1(G2106), .A2(n830), .ZN(G217) );
  AND2_X1 U925 ( .A1(G15), .A2(G2), .ZN(n831) );
  NAND2_X1 U926 ( .A1(G661), .A2(n831), .ZN(G259) );
  NAND2_X1 U927 ( .A1(G3), .A2(G1), .ZN(n832) );
  NAND2_X1 U928 ( .A1(n833), .A2(n832), .ZN(G188) );
  INV_X1 U930 ( .A(G120), .ZN(G236) );
  INV_X1 U931 ( .A(G96), .ZN(G221) );
  INV_X1 U932 ( .A(G69), .ZN(G235) );
  NOR2_X1 U933 ( .A1(n835), .A2(n834), .ZN(G325) );
  INV_X1 U934 ( .A(G325), .ZN(G261) );
  XOR2_X1 U935 ( .A(n836), .B(G286), .Z(n838) );
  XNOR2_X1 U936 ( .A(G171), .B(n948), .ZN(n837) );
  XNOR2_X1 U937 ( .A(n838), .B(n837), .ZN(n839) );
  XNOR2_X1 U938 ( .A(n839), .B(n934), .ZN(n840) );
  NOR2_X1 U939 ( .A1(G37), .A2(n840), .ZN(G397) );
  XOR2_X1 U940 ( .A(KEYINPUT109), .B(G1991), .Z(n842) );
  XNOR2_X1 U941 ( .A(G1996), .B(G1981), .ZN(n841) );
  XNOR2_X1 U942 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U943 ( .A(n843), .B(KEYINPUT41), .Z(n845) );
  XNOR2_X1 U944 ( .A(G1971), .B(G1986), .ZN(n844) );
  XNOR2_X1 U945 ( .A(n845), .B(n844), .ZN(n849) );
  XOR2_X1 U946 ( .A(G1976), .B(G1956), .Z(n847) );
  XNOR2_X1 U947 ( .A(G1966), .B(G1961), .ZN(n846) );
  XNOR2_X1 U948 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U949 ( .A(n849), .B(n848), .Z(n851) );
  XNOR2_X1 U950 ( .A(KEYINPUT110), .B(G2474), .ZN(n850) );
  XNOR2_X1 U951 ( .A(n851), .B(n850), .ZN(G229) );
  XOR2_X1 U952 ( .A(G2096), .B(KEYINPUT43), .Z(n853) );
  XNOR2_X1 U953 ( .A(G2090), .B(G2678), .ZN(n852) );
  XNOR2_X1 U954 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U955 ( .A(n854), .B(KEYINPUT108), .Z(n856) );
  XNOR2_X1 U956 ( .A(G2067), .B(G2072), .ZN(n855) );
  XNOR2_X1 U957 ( .A(n856), .B(n855), .ZN(n860) );
  XOR2_X1 U958 ( .A(KEYINPUT42), .B(G2100), .Z(n858) );
  XNOR2_X1 U959 ( .A(G2078), .B(G2084), .ZN(n857) );
  XNOR2_X1 U960 ( .A(n858), .B(n857), .ZN(n859) );
  XNOR2_X1 U961 ( .A(n860), .B(n859), .ZN(G227) );
  NAND2_X1 U962 ( .A1(G112), .A2(n880), .ZN(n862) );
  NAND2_X1 U963 ( .A1(G100), .A2(n886), .ZN(n861) );
  NAND2_X1 U964 ( .A1(n862), .A2(n861), .ZN(n863) );
  XNOR2_X1 U965 ( .A(n863), .B(KEYINPUT111), .ZN(n865) );
  NAND2_X1 U966 ( .A1(G136), .A2(n878), .ZN(n864) );
  NAND2_X1 U967 ( .A1(n865), .A2(n864), .ZN(n868) );
  NAND2_X1 U968 ( .A1(n881), .A2(G124), .ZN(n866) );
  XOR2_X1 U969 ( .A(KEYINPUT44), .B(n866), .Z(n867) );
  NOR2_X1 U970 ( .A1(n868), .A2(n867), .ZN(G162) );
  NAND2_X1 U971 ( .A1(G118), .A2(n880), .ZN(n870) );
  NAND2_X1 U972 ( .A1(G130), .A2(n881), .ZN(n869) );
  NAND2_X1 U973 ( .A1(n870), .A2(n869), .ZN(n871) );
  XNOR2_X1 U974 ( .A(KEYINPUT112), .B(n871), .ZN(n876) );
  NAND2_X1 U975 ( .A1(G106), .A2(n886), .ZN(n873) );
  NAND2_X1 U976 ( .A1(G142), .A2(n878), .ZN(n872) );
  NAND2_X1 U977 ( .A1(n873), .A2(n872), .ZN(n874) );
  XOR2_X1 U978 ( .A(n874), .B(KEYINPUT45), .Z(n875) );
  NOR2_X1 U979 ( .A1(n876), .A2(n875), .ZN(n877) );
  XNOR2_X1 U980 ( .A(n877), .B(n965), .ZN(n894) );
  XOR2_X1 U981 ( .A(KEYINPUT115), .B(KEYINPUT46), .Z(n892) );
  NAND2_X1 U982 ( .A1(n878), .A2(G139), .ZN(n879) );
  XNOR2_X1 U983 ( .A(KEYINPUT113), .B(n879), .ZN(n890) );
  NAND2_X1 U984 ( .A1(G115), .A2(n880), .ZN(n883) );
  NAND2_X1 U985 ( .A1(G127), .A2(n881), .ZN(n882) );
  NAND2_X1 U986 ( .A1(n883), .A2(n882), .ZN(n884) );
  XNOR2_X1 U987 ( .A(n884), .B(KEYINPUT114), .ZN(n885) );
  XNOR2_X1 U988 ( .A(n885), .B(KEYINPUT47), .ZN(n888) );
  NAND2_X1 U989 ( .A1(n886), .A2(G103), .ZN(n887) );
  NAND2_X1 U990 ( .A1(n888), .A2(n887), .ZN(n889) );
  NOR2_X1 U991 ( .A1(n890), .A2(n889), .ZN(n978) );
  XNOR2_X1 U992 ( .A(n978), .B(KEYINPUT48), .ZN(n891) );
  XNOR2_X1 U993 ( .A(n892), .B(n891), .ZN(n893) );
  XOR2_X1 U994 ( .A(n894), .B(n893), .Z(n896) );
  XNOR2_X1 U995 ( .A(G160), .B(G164), .ZN(n895) );
  XNOR2_X1 U996 ( .A(n896), .B(n895), .ZN(n897) );
  XOR2_X1 U997 ( .A(n897), .B(G162), .Z(n901) );
  XNOR2_X1 U998 ( .A(n899), .B(n898), .ZN(n900) );
  XNOR2_X1 U999 ( .A(n901), .B(n900), .ZN(n903) );
  XNOR2_X1 U1000 ( .A(n903), .B(n902), .ZN(n904) );
  NOR2_X1 U1001 ( .A1(G37), .A2(n904), .ZN(G395) );
  NOR2_X1 U1002 ( .A1(G229), .A2(G227), .ZN(n905) );
  XNOR2_X1 U1003 ( .A(KEYINPUT49), .B(n905), .ZN(n906) );
  NOR2_X1 U1004 ( .A1(G397), .A2(n906), .ZN(n911) );
  NOR2_X1 U1005 ( .A1(n907), .A2(G401), .ZN(n908) );
  XOR2_X1 U1006 ( .A(KEYINPUT116), .B(n908), .Z(n909) );
  NOR2_X1 U1007 ( .A1(G395), .A2(n909), .ZN(n910) );
  NAND2_X1 U1008 ( .A1(n911), .A2(n910), .ZN(G225) );
  INV_X1 U1009 ( .A(G225), .ZN(G308) );
  XNOR2_X1 U1010 ( .A(G1966), .B(G21), .ZN(n913) );
  XNOR2_X1 U1011 ( .A(G5), .B(G1961), .ZN(n912) );
  NOR2_X1 U1012 ( .A1(n913), .A2(n912), .ZN(n923) );
  XOR2_X1 U1013 ( .A(G1348), .B(KEYINPUT59), .Z(n914) );
  XNOR2_X1 U1014 ( .A(G4), .B(n914), .ZN(n916) );
  XNOR2_X1 U1015 ( .A(G20), .B(G1956), .ZN(n915) );
  NOR2_X1 U1016 ( .A1(n916), .A2(n915), .ZN(n920) );
  XNOR2_X1 U1017 ( .A(G1341), .B(G19), .ZN(n918) );
  XNOR2_X1 U1018 ( .A(G6), .B(G1981), .ZN(n917) );
  NOR2_X1 U1019 ( .A1(n918), .A2(n917), .ZN(n919) );
  NAND2_X1 U1020 ( .A1(n920), .A2(n919), .ZN(n921) );
  XOR2_X1 U1021 ( .A(KEYINPUT60), .B(n921), .Z(n922) );
  NAND2_X1 U1022 ( .A1(n923), .A2(n922), .ZN(n930) );
  XNOR2_X1 U1023 ( .A(G1971), .B(G22), .ZN(n925) );
  XNOR2_X1 U1024 ( .A(G23), .B(G1976), .ZN(n924) );
  NOR2_X1 U1025 ( .A1(n925), .A2(n924), .ZN(n927) );
  XOR2_X1 U1026 ( .A(G1986), .B(G24), .Z(n926) );
  NAND2_X1 U1027 ( .A1(n927), .A2(n926), .ZN(n928) );
  XNOR2_X1 U1028 ( .A(KEYINPUT58), .B(n928), .ZN(n929) );
  NOR2_X1 U1029 ( .A1(n930), .A2(n929), .ZN(n931) );
  XOR2_X1 U1030 ( .A(KEYINPUT61), .B(n931), .Z(n932) );
  NOR2_X1 U1031 ( .A1(G16), .A2(n932), .ZN(n933) );
  XNOR2_X1 U1032 ( .A(KEYINPUT125), .B(n933), .ZN(n960) );
  XNOR2_X1 U1033 ( .A(KEYINPUT56), .B(G16), .ZN(n958) );
  XNOR2_X1 U1034 ( .A(n934), .B(G1341), .ZN(n940) );
  XNOR2_X1 U1035 ( .A(G1966), .B(G168), .ZN(n936) );
  NAND2_X1 U1036 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1037 ( .A(n937), .B(KEYINPUT57), .ZN(n938) );
  XNOR2_X1 U1038 ( .A(KEYINPUT123), .B(n938), .ZN(n939) );
  NOR2_X1 U1039 ( .A1(n940), .A2(n939), .ZN(n956) );
  NAND2_X1 U1040 ( .A1(G303), .A2(G1971), .ZN(n946) );
  NAND2_X1 U1041 ( .A1(n942), .A2(n941), .ZN(n944) );
  XNOR2_X1 U1042 ( .A(G1956), .B(G299), .ZN(n943) );
  NOR2_X1 U1043 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1044 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1045 ( .A(n947), .B(KEYINPUT124), .ZN(n954) );
  XNOR2_X1 U1046 ( .A(G301), .B(G1961), .ZN(n950) );
  XNOR2_X1 U1047 ( .A(G1348), .B(n948), .ZN(n949) );
  NOR2_X1 U1048 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1049 ( .A1(n952), .A2(n951), .ZN(n953) );
  NOR2_X1 U1050 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1051 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1052 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1053 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1054 ( .A(n961), .B(KEYINPUT126), .ZN(n991) );
  INV_X1 U1055 ( .A(G29), .ZN(n988) );
  XOR2_X1 U1056 ( .A(G2090), .B(G162), .Z(n962) );
  NOR2_X1 U1057 ( .A1(n963), .A2(n962), .ZN(n964) );
  XOR2_X1 U1058 ( .A(KEYINPUT51), .B(n964), .Z(n974) );
  XNOR2_X1 U1059 ( .A(G160), .B(G2084), .ZN(n966) );
  NAND2_X1 U1060 ( .A1(n966), .A2(n965), .ZN(n967) );
  NOR2_X1 U1061 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1062 ( .A1(n970), .A2(n969), .ZN(n971) );
  NOR2_X1 U1063 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1064 ( .A1(n974), .A2(n973), .ZN(n975) );
  NOR2_X1 U1065 ( .A1(n976), .A2(n975), .ZN(n977) );
  XNOR2_X1 U1066 ( .A(KEYINPUT117), .B(n977), .ZN(n984) );
  XOR2_X1 U1067 ( .A(G2072), .B(n978), .Z(n980) );
  XOR2_X1 U1068 ( .A(G164), .B(G2078), .Z(n979) );
  NOR2_X1 U1069 ( .A1(n980), .A2(n979), .ZN(n981) );
  XOR2_X1 U1070 ( .A(KEYINPUT50), .B(n981), .Z(n982) );
  XNOR2_X1 U1071 ( .A(KEYINPUT118), .B(n982), .ZN(n983) );
  NOR2_X1 U1072 ( .A1(n984), .A2(n983), .ZN(n985) );
  XOR2_X1 U1073 ( .A(KEYINPUT52), .B(n985), .Z(n986) );
  NOR2_X1 U1074 ( .A1(KEYINPUT55), .A2(n986), .ZN(n987) );
  NOR2_X1 U1075 ( .A1(n988), .A2(n987), .ZN(n989) );
  XOR2_X1 U1076 ( .A(KEYINPUT119), .B(n989), .Z(n990) );
  NOR2_X1 U1077 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1078 ( .A1(G11), .A2(n992), .ZN(n1017) );
  XOR2_X1 U1079 ( .A(KEYINPUT121), .B(KEYINPUT55), .Z(n1013) );
  XNOR2_X1 U1080 ( .A(G2090), .B(G35), .ZN(n1008) );
  XOR2_X1 U1081 ( .A(G2072), .B(G33), .Z(n995) );
  XNOR2_X1 U1082 ( .A(n993), .B(G32), .ZN(n994) );
  NAND2_X1 U1083 ( .A1(n995), .A2(n994), .ZN(n1005) );
  XNOR2_X1 U1084 ( .A(G25), .B(n996), .ZN(n1003) );
  XOR2_X1 U1085 ( .A(G2067), .B(G26), .Z(n997) );
  NAND2_X1 U1086 ( .A1(n997), .A2(G28), .ZN(n1001) );
  XNOR2_X1 U1087 ( .A(G27), .B(n998), .ZN(n999) );
  XNOR2_X1 U1088 ( .A(KEYINPUT120), .B(n999), .ZN(n1000) );
  NOR2_X1 U1089 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1090 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NOR2_X1 U1091 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1092 ( .A(KEYINPUT53), .B(n1006), .ZN(n1007) );
  NOR2_X1 U1093 ( .A1(n1008), .A2(n1007), .ZN(n1011) );
  XOR2_X1 U1094 ( .A(G2084), .B(G34), .Z(n1009) );
  XNOR2_X1 U1095 ( .A(KEYINPUT54), .B(n1009), .ZN(n1010) );
  NAND2_X1 U1096 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1097 ( .A(n1013), .B(n1012), .ZN(n1014) );
  NOR2_X1 U1098 ( .A1(n1014), .A2(G29), .ZN(n1015) );
  XNOR2_X1 U1099 ( .A(KEYINPUT122), .B(n1015), .ZN(n1016) );
  NOR2_X1 U1100 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1101 ( .A(KEYINPUT62), .B(n1018), .ZN(G311) );
  INV_X1 U1102 ( .A(G311), .ZN(G150) );
endmodule

