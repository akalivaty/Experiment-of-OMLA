//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 1 1 1 1 0 0 0 1 0 1 1 1 1 1 1 0 1 1 1 1 1 1 1 0 0 0 0 1 0 0 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 1 0 1 0 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:38 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n734, new_n735, new_n736, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n767, new_n768, new_n769, new_n770, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n791, new_n792, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n819, new_n820, new_n821, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040;
  INV_X1    g000(.A(KEYINPUT6), .ZN(new_n187));
  NOR2_X1   g001(.A1(KEYINPUT2), .A2(G113), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT71), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  OAI21_X1  g004(.A(KEYINPUT71), .B1(KEYINPUT2), .B2(G113), .ZN(new_n191));
  AOI22_X1  g005(.A1(new_n190), .A2(new_n191), .B1(KEYINPUT2), .B2(G113), .ZN(new_n192));
  INV_X1    g006(.A(G119), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G116), .ZN(new_n194));
  INV_X1    g008(.A(G116), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G119), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n192), .A2(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(KEYINPUT72), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT72), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n192), .A2(new_n201), .A3(new_n198), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n200), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(new_n192), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(new_n197), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  AND2_X1   g020(.A1(KEYINPUT88), .A2(G104), .ZN(new_n207));
  NOR2_X1   g021(.A1(KEYINPUT88), .A2(G104), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G107), .ZN(new_n210));
  INV_X1    g024(.A(G104), .ZN(new_n211));
  NOR3_X1   g025(.A1(new_n211), .A2(KEYINPUT3), .A3(G107), .ZN(new_n212));
  INV_X1    g026(.A(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT88), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(new_n211), .ZN(new_n215));
  NAND2_X1  g029(.A1(KEYINPUT88), .A2(G104), .ZN(new_n216));
  AOI21_X1  g030(.A(G107), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT3), .ZN(new_n218));
  NOR3_X1   g032(.A1(new_n217), .A2(KEYINPUT89), .A3(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT89), .ZN(new_n220));
  INV_X1    g034(.A(G107), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n221), .B1(new_n207), .B2(new_n208), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n220), .B1(new_n222), .B2(KEYINPUT3), .ZN(new_n223));
  OAI211_X1 g037(.A(new_n210), .B(new_n213), .C1(new_n219), .C2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(G101), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n225), .A2(KEYINPUT4), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g041(.A(KEYINPUT89), .B1(new_n217), .B2(new_n218), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n222), .A2(new_n220), .A3(KEYINPUT3), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n212), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n225), .B1(new_n230), .B2(new_n210), .ZN(new_n231));
  AOI21_X1  g045(.A(G101), .B1(new_n209), .B2(G107), .ZN(new_n232));
  OAI211_X1 g046(.A(new_n213), .B(new_n232), .C1(new_n219), .C2(new_n223), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(KEYINPUT4), .ZN(new_n234));
  OAI211_X1 g048(.A(new_n206), .B(new_n227), .C1(new_n231), .C2(new_n234), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n221), .A2(G104), .ZN(new_n236));
  OAI21_X1  g050(.A(G101), .B1(new_n217), .B2(new_n236), .ZN(new_n237));
  AND2_X1   g051(.A1(new_n233), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT5), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n197), .A2(new_n239), .ZN(new_n240));
  OAI21_X1  g054(.A(G113), .B1(new_n194), .B2(KEYINPUT5), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n242), .B1(new_n200), .B2(new_n202), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n238), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n235), .A2(new_n244), .ZN(new_n245));
  XNOR2_X1  g059(.A(G110), .B(G122), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n187), .B1(new_n245), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n224), .A2(G101), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n249), .A2(KEYINPUT4), .A3(new_n233), .ZN(new_n250));
  AOI22_X1  g064(.A1(new_n203), .A2(new_n205), .B1(new_n224), .B2(new_n226), .ZN(new_n251));
  AOI22_X1  g065(.A1(new_n250), .A2(new_n251), .B1(new_n238), .B2(new_n243), .ZN(new_n252));
  AOI21_X1  g066(.A(KEYINPUT92), .B1(new_n252), .B2(new_n246), .ZN(new_n253));
  AND4_X1   g067(.A1(KEYINPUT92), .A2(new_n235), .A3(new_n244), .A4(new_n246), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n248), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n245), .A2(new_n187), .A3(new_n247), .ZN(new_n256));
  INV_X1    g070(.A(G146), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G143), .ZN(new_n258));
  INV_X1    g072(.A(G143), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G146), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  OAI21_X1  g075(.A(KEYINPUT1), .B1(new_n259), .B2(G146), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT69), .ZN(new_n263));
  OAI21_X1  g077(.A(G128), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  AOI21_X1  g078(.A(KEYINPUT69), .B1(new_n258), .B2(KEYINPUT1), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n261), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  XNOR2_X1  g080(.A(G143), .B(G146), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT1), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n267), .A2(new_n268), .A3(G128), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n266), .A2(new_n269), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n270), .A2(G125), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(G953), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(G224), .ZN(new_n274));
  AND2_X1   g088(.A1(KEYINPUT0), .A2(G128), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT64), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n275), .B1(new_n267), .B2(new_n276), .ZN(new_n277));
  NOR2_X1   g091(.A1(KEYINPUT0), .A2(G128), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n275), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n261), .A2(new_n279), .A3(KEYINPUT64), .ZN(new_n280));
  AND2_X1   g094(.A1(new_n277), .A2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(G125), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n272), .A2(new_n274), .A3(new_n284), .ZN(new_n285));
  OAI211_X1 g099(.A(G224), .B(new_n273), .C1(new_n271), .C2(new_n283), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n255), .A2(new_n256), .A3(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT92), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n289), .B1(new_n245), .B2(new_n247), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n252), .A2(KEYINPUT92), .A3(new_n246), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  XOR2_X1   g106(.A(new_n246), .B(KEYINPUT8), .Z(new_n293));
  OR2_X1    g107(.A1(new_n238), .A2(new_n243), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n293), .B1(new_n294), .B2(new_n244), .ZN(new_n295));
  AOI21_X1  g109(.A(KEYINPUT7), .B1(new_n273), .B2(G224), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n296), .B1(new_n285), .B2(new_n286), .ZN(new_n297));
  INV_X1    g111(.A(new_n296), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n298), .B1(new_n272), .B2(new_n284), .ZN(new_n299));
  NOR3_X1   g113(.A1(new_n295), .A2(new_n297), .A3(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(G902), .B1(new_n292), .B2(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(G210), .B1(G237), .B2(G902), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n288), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(KEYINPUT93), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT93), .ZN(new_n305));
  NAND4_X1  g119(.A1(new_n288), .A2(new_n301), .A3(new_n305), .A4(new_n302), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n288), .A2(new_n301), .ZN(new_n307));
  INV_X1    g121(.A(new_n302), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n304), .A2(new_n306), .A3(new_n309), .ZN(new_n310));
  OAI21_X1  g124(.A(G214), .B1(G237), .B2(G902), .ZN(new_n311));
  AND2_X1   g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  XOR2_X1   g126(.A(KEYINPUT9), .B(G234), .Z(new_n313));
  XNOR2_X1  g127(.A(new_n313), .B(KEYINPUT85), .ZN(new_n314));
  INV_X1    g128(.A(G902), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(G221), .ZN(new_n317));
  XOR2_X1   g131(.A(new_n317), .B(KEYINPUT86), .Z(new_n318));
  NAND2_X1  g132(.A1(new_n273), .A2(G227), .ZN(new_n319));
  XNOR2_X1  g133(.A(new_n319), .B(KEYINPUT87), .ZN(new_n320));
  XNOR2_X1  g134(.A(G110), .B(G140), .ZN(new_n321));
  XNOR2_X1  g135(.A(new_n320), .B(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT12), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n268), .B1(G143), .B2(new_n257), .ZN(new_n325));
  INV_X1    g139(.A(G128), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n261), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(new_n269), .ZN(new_n328));
  AND3_X1   g142(.A1(new_n233), .A2(new_n237), .A3(new_n328), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n270), .B1(new_n233), .B2(new_n237), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT91), .ZN(new_n331));
  NOR3_X1   g145(.A1(new_n329), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n233), .A2(new_n237), .ZN(new_n333));
  INV_X1    g147(.A(new_n270), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n333), .A2(new_n331), .A3(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(G137), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n336), .A2(G134), .ZN(new_n337));
  INV_X1    g151(.A(G134), .ZN(new_n338));
  OAI21_X1  g152(.A(KEYINPUT11), .B1(new_n338), .B2(G137), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT11), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n340), .A2(new_n336), .A3(G134), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n337), .B1(new_n339), .B2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(G131), .ZN(new_n343));
  AOI21_X1  g157(.A(KEYINPUT65), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(new_n337), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n340), .B1(G134), .B2(new_n336), .ZN(new_n346));
  NOR3_X1   g160(.A1(new_n338), .A2(KEYINPUT11), .A3(G137), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n345), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(G131), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n344), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n348), .A2(KEYINPUT65), .A3(G131), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n335), .A2(new_n353), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n324), .B1(new_n332), .B2(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n233), .A2(new_n237), .A3(new_n328), .ZN(new_n356));
  OAI211_X1 g170(.A(KEYINPUT91), .B(new_n356), .C1(new_n238), .C2(new_n270), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n357), .A2(KEYINPUT12), .A3(new_n353), .A4(new_n335), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n355), .A2(new_n358), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n326), .B1(new_n325), .B2(KEYINPUT69), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n262), .A2(new_n263), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n267), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(new_n269), .ZN(new_n363));
  OAI21_X1  g177(.A(KEYINPUT73), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT73), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n266), .A2(new_n365), .A3(new_n269), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n364), .A2(KEYINPUT10), .A3(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT10), .ZN(new_n369));
  AOI22_X1  g183(.A1(new_n368), .A2(new_n238), .B1(new_n369), .B2(new_n356), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n277), .A2(new_n280), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n371), .B1(new_n224), .B2(new_n226), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT90), .ZN(new_n373));
  OAI211_X1 g187(.A(new_n372), .B(new_n373), .C1(new_n231), .C2(new_n234), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n373), .B1(new_n250), .B2(new_n372), .ZN(new_n376));
  OAI211_X1 g190(.A(new_n352), .B(new_n370), .C1(new_n375), .C2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n359), .A2(new_n377), .ZN(new_n378));
  OAI22_X1  g192(.A1(new_n329), .A2(KEYINPUT10), .B1(new_n367), .B2(new_n333), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n372), .B1(new_n231), .B2(new_n234), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(KEYINPUT90), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n379), .B1(new_n381), .B2(new_n374), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n323), .B1(new_n382), .B2(new_n352), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n370), .B1(new_n375), .B2(new_n376), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(new_n353), .ZN(new_n385));
  AOI22_X1  g199(.A1(new_n323), .A2(new_n378), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  OAI21_X1  g200(.A(G469), .B1(new_n386), .B2(G902), .ZN(new_n387));
  INV_X1    g201(.A(G469), .ZN(new_n388));
  XOR2_X1   g202(.A(KEYINPUT79), .B(G902), .Z(new_n389));
  AOI21_X1  g203(.A(new_n322), .B1(new_n385), .B2(new_n377), .ZN(new_n390));
  AND3_X1   g204(.A1(new_n359), .A2(new_n322), .A3(new_n377), .ZN(new_n391));
  OAI211_X1 g205(.A(new_n388), .B(new_n389), .C1(new_n390), .C2(new_n391), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n318), .B1(new_n387), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n312), .A2(new_n393), .ZN(new_n394));
  XOR2_X1   g208(.A(G113), .B(G122), .Z(new_n395));
  XNOR2_X1  g209(.A(KEYINPUT96), .B(G104), .ZN(new_n396));
  XNOR2_X1  g210(.A(new_n395), .B(new_n396), .ZN(new_n397));
  XNOR2_X1  g211(.A(G125), .B(G140), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(KEYINPUT16), .ZN(new_n399));
  OR3_X1    g213(.A1(new_n282), .A2(KEYINPUT16), .A3(G140), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n399), .A2(G146), .A3(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT19), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n398), .A2(new_n403), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n398), .B(KEYINPUT83), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n404), .B1(new_n405), .B2(new_n403), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n402), .B1(new_n406), .B2(new_n257), .ZN(new_n407));
  INV_X1    g221(.A(G237), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n408), .A2(new_n273), .A3(G214), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n409), .B(new_n259), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(G131), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n409), .B(G143), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(new_n343), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(KEYINPUT95), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT95), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n411), .A2(new_n413), .A3(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n407), .A2(new_n415), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(KEYINPUT18), .A2(G131), .ZN(new_n419));
  XNOR2_X1  g233(.A(new_n410), .B(new_n419), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n398), .A2(new_n257), .ZN(new_n421));
  XOR2_X1   g235(.A(new_n421), .B(KEYINPUT94), .Z(new_n422));
  NAND2_X1  g236(.A1(new_n405), .A2(new_n257), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n420), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n397), .B1(new_n418), .B2(new_n425), .ZN(new_n426));
  XOR2_X1   g240(.A(new_n397), .B(KEYINPUT97), .Z(new_n427));
  INV_X1    g241(.A(KEYINPUT98), .ZN(new_n428));
  AOI21_X1  g242(.A(G146), .B1(new_n399), .B2(new_n400), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n428), .B1(new_n402), .B2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n429), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n431), .A2(KEYINPUT98), .A3(new_n401), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT17), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n411), .A2(new_n413), .A3(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n410), .A2(KEYINPUT17), .A3(G131), .ZN(new_n435));
  NAND4_X1  g249(.A1(new_n430), .A2(new_n432), .A3(new_n434), .A4(new_n435), .ZN(new_n436));
  AND3_X1   g250(.A1(new_n427), .A2(new_n436), .A3(new_n425), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n426), .A2(new_n437), .ZN(new_n438));
  NOR2_X1   g252(.A1(G475), .A2(G902), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  OAI21_X1  g254(.A(KEYINPUT20), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT20), .ZN(new_n442));
  OAI211_X1 g256(.A(new_n442), .B(new_n439), .C1(new_n426), .C2(new_n437), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n397), .B1(new_n436), .B2(new_n425), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n315), .B1(new_n437), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(G475), .ZN(new_n447));
  AND2_X1   g261(.A1(new_n444), .A2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(G122), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(G116), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n195), .A2(G122), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n221), .B1(new_n450), .B2(KEYINPUT14), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n453), .B(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT100), .ZN(new_n456));
  XNOR2_X1  g270(.A(G128), .B(G143), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(new_n338), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n457), .A2(new_n338), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n456), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(new_n460), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n462), .A2(KEYINPUT100), .A3(new_n458), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n455), .A2(new_n461), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(KEYINPUT101), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT101), .ZN(new_n466));
  NAND4_X1  g280(.A1(new_n455), .A2(new_n461), .A3(new_n463), .A4(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n314), .A2(G217), .A3(new_n273), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n259), .A2(KEYINPUT13), .A3(G128), .ZN(new_n471));
  OAI211_X1 g285(.A(new_n471), .B(KEYINPUT99), .C1(G128), .C2(new_n259), .ZN(new_n472));
  AOI21_X1  g286(.A(KEYINPUT13), .B1(new_n259), .B2(G128), .ZN(new_n473));
  OAI221_X1 g287(.A(G134), .B1(KEYINPUT99), .B2(new_n471), .C1(new_n472), .C2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n453), .A2(G107), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n452), .A2(new_n221), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n474), .A2(new_n458), .A3(new_n475), .A4(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n468), .A2(new_n470), .A3(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n470), .B1(new_n468), .B2(new_n477), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n389), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(G478), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n482), .A2(KEYINPUT15), .ZN(new_n483));
  OR2_X1    g297(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n481), .A2(new_n483), .ZN(new_n485));
  AND2_X1   g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT102), .ZN(new_n487));
  NAND2_X1  g301(.A1(G234), .A2(G237), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n488), .A2(G952), .A3(new_n273), .ZN(new_n489));
  INV_X1    g303(.A(new_n389), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n490), .A2(G953), .A3(new_n488), .ZN(new_n491));
  XNOR2_X1  g305(.A(KEYINPUT21), .B(G898), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n489), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  NAND4_X1  g308(.A1(new_n448), .A2(new_n486), .A3(new_n487), .A4(new_n494), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n444), .A2(new_n484), .A3(new_n485), .A4(new_n447), .ZN(new_n496));
  INV_X1    g310(.A(new_n494), .ZN(new_n497));
  OAI21_X1  g311(.A(KEYINPUT102), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n394), .B1(new_n495), .B2(new_n498), .ZN(new_n499));
  NOR2_X1   g313(.A1(G472), .A2(G902), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT32), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT76), .ZN(new_n504));
  OAI21_X1  g318(.A(KEYINPUT68), .B1(new_n336), .B2(G134), .ZN(new_n505));
  OAI21_X1  g319(.A(KEYINPUT67), .B1(new_n338), .B2(G137), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT68), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n507), .A2(new_n338), .A3(G137), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT67), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n509), .A2(new_n336), .A3(G134), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n505), .A2(new_n506), .A3(new_n508), .A4(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(G131), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n342), .A2(new_n343), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n364), .A2(new_n515), .A3(new_n366), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n350), .A2(new_n281), .A3(new_n351), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n516), .A2(KEYINPUT30), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(new_n206), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT30), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT66), .ZN(new_n521));
  AND2_X1   g335(.A1(new_n517), .A2(new_n521), .ZN(new_n522));
  NAND4_X1  g336(.A1(new_n350), .A2(new_n281), .A3(KEYINPUT66), .A4(new_n351), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n515), .A2(new_n270), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n520), .B1(new_n522), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(KEYINPUT70), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n517), .A2(new_n521), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n528), .A2(new_n524), .A3(new_n523), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT70), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n529), .A2(new_n530), .A3(new_n520), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n519), .B1(new_n527), .B2(new_n531), .ZN(new_n532));
  AOI22_X1  g346(.A1(new_n200), .A2(new_n202), .B1(new_n204), .B2(new_n197), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n516), .A2(new_n517), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(KEYINPUT74), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT74), .ZN(new_n536));
  NAND4_X1  g350(.A1(new_n516), .A2(new_n536), .A3(new_n517), .A4(new_n533), .ZN(new_n537));
  XOR2_X1   g351(.A(KEYINPUT75), .B(KEYINPUT27), .Z(new_n538));
  NAND3_X1  g352(.A1(new_n408), .A2(new_n273), .A3(G210), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n538), .B(new_n539), .ZN(new_n540));
  XNOR2_X1  g354(.A(KEYINPUT26), .B(G101), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n540), .B(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n535), .A2(new_n537), .A3(new_n542), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n504), .B1(new_n532), .B2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n519), .ZN(new_n545));
  AND3_X1   g359(.A1(new_n529), .A2(new_n530), .A3(new_n520), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n530), .B1(new_n529), .B2(new_n520), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n543), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n548), .A2(KEYINPUT76), .A3(new_n549), .ZN(new_n550));
  AND3_X1   g364(.A1(new_n544), .A2(KEYINPUT31), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n548), .A2(new_n549), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n529), .A2(new_n206), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n553), .A2(new_n535), .A3(new_n537), .ZN(new_n554));
  XOR2_X1   g368(.A(KEYINPUT77), .B(KEYINPUT28), .Z(new_n555));
  INV_X1    g369(.A(KEYINPUT28), .ZN(new_n556));
  AOI22_X1  g370(.A1(new_n554), .A2(new_n555), .B1(new_n556), .B2(new_n534), .ZN(new_n557));
  OAI22_X1  g371(.A1(new_n552), .A2(KEYINPUT31), .B1(new_n557), .B2(new_n542), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n503), .B1(new_n551), .B2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT80), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT31), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n527), .A2(new_n531), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n543), .B1(new_n563), .B2(new_n545), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n554), .A2(new_n555), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n534), .A2(new_n556), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n542), .ZN(new_n568));
  AOI22_X1  g382(.A1(new_n562), .A2(new_n564), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n544), .A2(new_n550), .A3(KEYINPUT31), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n571), .A2(KEYINPUT80), .A3(new_n503), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n561), .A2(new_n572), .ZN(new_n573));
  AND3_X1   g387(.A1(new_n266), .A2(new_n365), .A3(new_n269), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n365), .B1(new_n266), .B2(new_n269), .ZN(new_n575));
  NOR3_X1   g389(.A1(new_n574), .A2(new_n575), .A3(new_n514), .ZN(new_n576));
  INV_X1    g390(.A(new_n517), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n206), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n535), .A2(new_n537), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(KEYINPUT28), .ZN(new_n580));
  AND3_X1   g394(.A1(new_n534), .A2(KEYINPUT78), .A3(new_n556), .ZN(new_n581));
  AOI21_X1  g395(.A(KEYINPUT78), .B1(new_n534), .B2(new_n556), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(KEYINPUT29), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT29), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n557), .A2(new_n586), .ZN(new_n587));
  AND3_X1   g401(.A1(new_n585), .A2(new_n587), .A3(new_n542), .ZN(new_n588));
  AND2_X1   g402(.A1(new_n535), .A2(new_n537), .ZN(new_n589));
  NAND4_X1  g403(.A1(new_n548), .A2(new_n586), .A3(new_n589), .A4(new_n568), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(new_n389), .ZN(new_n591));
  OAI21_X1  g405(.A(G472), .B1(new_n588), .B2(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n501), .B1(new_n569), .B2(new_n570), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n592), .B1(KEYINPUT32), .B2(new_n593), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n573), .A2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(G217), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n596), .B1(new_n389), .B2(G234), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT25), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n193), .A2(G128), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n600), .A2(KEYINPUT81), .A3(KEYINPUT23), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n326), .A2(KEYINPUT82), .A3(G119), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n326), .A2(G119), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT82), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n601), .A2(new_n602), .A3(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(KEYINPUT81), .B1(new_n600), .B2(KEYINPUT23), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT23), .ZN(new_n608));
  OAI22_X1  g422(.A1(new_n606), .A2(new_n607), .B1(new_n608), .B2(new_n603), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(G110), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n603), .A2(new_n600), .ZN(new_n611));
  XNOR2_X1  g425(.A(KEYINPUT24), .B(G110), .ZN(new_n612));
  OAI221_X1 g426(.A(new_n610), .B1(new_n611), .B2(new_n612), .C1(new_n429), .C2(new_n402), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n611), .A2(new_n612), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n614), .B1(new_n609), .B2(G110), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n615), .A2(new_n401), .A3(new_n423), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n613), .A2(new_n616), .ZN(new_n617));
  XNOR2_X1  g431(.A(KEYINPUT22), .B(G137), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n273), .A2(G221), .A3(G234), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n618), .B(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n617), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n613), .A2(new_n616), .A3(new_n620), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n599), .B1(new_n624), .B2(new_n490), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n622), .A2(KEYINPUT25), .A3(new_n389), .A4(new_n623), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n598), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n597), .A2(G902), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n622), .A2(new_n629), .A3(new_n623), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  NOR3_X1   g445(.A1(new_n595), .A2(KEYINPUT84), .A3(new_n631), .ZN(new_n632));
  AOI21_X1  g446(.A(KEYINPUT80), .B1(new_n571), .B2(new_n503), .ZN(new_n633));
  INV_X1    g447(.A(new_n503), .ZN(new_n634));
  AOI211_X1 g448(.A(new_n560), .B(new_n634), .C1(new_n569), .C2(new_n570), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(G472), .ZN(new_n637));
  INV_X1    g451(.A(new_n591), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n585), .A2(new_n587), .A3(new_n542), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n637), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n571), .A2(new_n500), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n640), .B1(new_n641), .B2(new_n502), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n631), .B1(new_n636), .B2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT84), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n499), .B1(new_n632), .B2(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(KEYINPUT103), .B(G101), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G3));
  NAND2_X1  g462(.A1(new_n571), .A2(new_n389), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(G472), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT104), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n318), .ZN(new_n653));
  INV_X1    g467(.A(new_n377), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n381), .A2(new_n374), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n352), .B1(new_n655), .B2(new_n370), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n323), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n383), .A2(new_n359), .ZN(new_n658));
  AOI211_X1 g472(.A(G469), .B(new_n490), .C1(new_n657), .C2(new_n658), .ZN(new_n659));
  AOI22_X1  g473(.A1(new_n382), .A2(new_n352), .B1(new_n355), .B2(new_n358), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n377), .A2(new_n322), .ZN(new_n661));
  OAI22_X1  g475(.A1(new_n660), .A2(new_n322), .B1(new_n661), .B2(new_n656), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n388), .B1(new_n662), .B2(new_n315), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n653), .B1(new_n659), .B2(new_n663), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n664), .A2(new_n631), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n637), .B1(new_n571), .B2(new_n389), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(KEYINPUT104), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n652), .A2(new_n665), .A3(new_n641), .A4(new_n667), .ZN(new_n668));
  AND3_X1   g482(.A1(new_n288), .A2(new_n301), .A3(new_n302), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n302), .B1(new_n288), .B2(new_n301), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n311), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(KEYINPUT105), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT105), .ZN(new_n673));
  OAI211_X1 g487(.A(new_n673), .B(new_n311), .C1(new_n669), .C2(new_n670), .ZN(new_n674));
  INV_X1    g488(.A(new_n480), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(new_n478), .ZN(new_n676));
  AOI21_X1  g490(.A(G478), .B1(new_n676), .B2(new_n389), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(KEYINPUT33), .ZN(new_n678));
  OR3_X1    g492(.A1(new_n479), .A2(KEYINPUT33), .A3(new_n480), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n490), .A2(new_n482), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n677), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n448), .A2(new_n682), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n672), .A2(new_n674), .A3(new_n494), .A4(new_n683), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n668), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(KEYINPUT34), .B(G104), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n685), .B(new_n686), .ZN(G6));
  NAND2_X1  g501(.A1(new_n444), .A2(new_n447), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n486), .A2(new_n688), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n672), .A2(new_n674), .A3(new_n494), .A4(new_n689), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n668), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(KEYINPUT35), .B(G107), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(G9));
  NOR2_X1   g507(.A1(new_n621), .A2(KEYINPUT36), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n617), .B(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(new_n629), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n627), .A2(new_n697), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n698), .B1(new_n495), .B2(new_n498), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n312), .A2(new_n393), .A3(new_n699), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n652), .A2(new_n641), .A3(new_n667), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(KEYINPUT37), .B(G110), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n702), .B(new_n703), .ZN(G12));
  AND3_X1   g518(.A1(new_n672), .A2(new_n393), .A3(new_n674), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n641), .A2(new_n502), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n706), .A2(new_n561), .A3(new_n592), .A4(new_n572), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n489), .B(KEYINPUT106), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n708), .B1(new_n491), .B2(G900), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n689), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n710), .A2(new_n698), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n705), .A2(new_n707), .A3(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G128), .ZN(G30));
  XNOR2_X1  g527(.A(new_n709), .B(KEYINPUT39), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n393), .A2(new_n714), .ZN(new_n715));
  OR2_X1    g529(.A1(new_n715), .A2(KEYINPUT40), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n310), .B(KEYINPUT38), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n448), .A2(new_n486), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n718), .A2(new_n311), .A3(new_n698), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n719), .B1(new_n715), .B2(KEYINPUT40), .ZN(new_n720));
  AND3_X1   g534(.A1(new_n716), .A2(new_n717), .A3(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n579), .A2(new_n568), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n544), .A2(new_n550), .A3(new_n722), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n637), .B1(new_n723), .B2(new_n315), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n724), .B1(new_n641), .B2(new_n502), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n636), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(KEYINPUT107), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT107), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n636), .A2(new_n728), .A3(new_n725), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  AND2_X1   g544(.A1(new_n721), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(new_n259), .ZN(G45));
  INV_X1    g546(.A(new_n683), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n709), .B1(new_n627), .B2(new_n697), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n705), .A2(new_n707), .A3(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G146), .ZN(G48));
  INV_X1    g551(.A(new_n631), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n389), .B1(new_n390), .B2(new_n391), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(G469), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n738), .A2(new_n740), .A3(new_n317), .A4(new_n392), .ZN(new_n741));
  INV_X1    g555(.A(new_n741), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n742), .B1(new_n573), .B2(new_n594), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n743), .A2(new_n684), .ZN(new_n744));
  XOR2_X1   g558(.A(KEYINPUT41), .B(G113), .Z(new_n745));
  XNOR2_X1  g559(.A(new_n744), .B(new_n745), .ZN(G15));
  NOR2_X1   g560(.A1(new_n743), .A2(new_n690), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(new_n195), .ZN(G18));
  NAND2_X1  g562(.A1(new_n740), .A2(new_n392), .ZN(new_n749));
  INV_X1    g563(.A(new_n317), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n751), .A2(new_n674), .A3(new_n672), .ZN(new_n752));
  INV_X1    g566(.A(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n753), .A2(new_n707), .A3(new_n699), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G119), .ZN(G21));
  AND4_X1   g569(.A1(new_n494), .A2(new_n740), .A3(new_n317), .A4(new_n392), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n756), .A2(new_n672), .A3(new_n674), .A4(new_n718), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT108), .ZN(new_n758));
  AOI22_X1  g572(.A1(new_n564), .A2(new_n562), .B1(new_n584), .B2(new_n568), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n570), .A2(new_n759), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n758), .B1(new_n760), .B2(new_n500), .ZN(new_n761));
  INV_X1    g575(.A(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n760), .A2(new_n758), .A3(new_n500), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n762), .A2(new_n650), .A3(new_n738), .A4(new_n763), .ZN(new_n764));
  OR2_X1    g578(.A1(new_n757), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G122), .ZN(G24));
  AND2_X1   g580(.A1(new_n672), .A2(new_n674), .ZN(new_n767));
  AOI211_X1 g581(.A(KEYINPUT108), .B(new_n501), .C1(new_n570), .C2(new_n759), .ZN(new_n768));
  NOR3_X1   g582(.A1(new_n666), .A2(new_n761), .A3(new_n768), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n767), .A2(new_n769), .A3(new_n735), .A4(new_n751), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G125), .ZN(G27));
  OAI211_X1 g585(.A(new_n592), .B(new_n559), .C1(KEYINPUT32), .C2(new_n593), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(new_n738), .ZN(new_n773));
  AND3_X1   g587(.A1(new_n304), .A2(new_n306), .A3(new_n309), .ZN(new_n774));
  INV_X1    g588(.A(new_n709), .ZN(new_n775));
  NOR3_X1   g589(.A1(new_n448), .A2(new_n682), .A3(new_n775), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n750), .B1(new_n387), .B2(new_n392), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n774), .A2(new_n311), .A3(new_n776), .A4(new_n777), .ZN(new_n778));
  OAI21_X1  g592(.A(KEYINPUT42), .B1(new_n773), .B2(new_n778), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n304), .A2(new_n309), .A3(new_n311), .A4(new_n306), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n317), .B1(new_n659), .B2(new_n663), .ZN(new_n781));
  INV_X1    g595(.A(new_n682), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n782), .A2(new_n688), .A3(new_n709), .ZN(new_n783));
  NOR3_X1   g597(.A1(new_n780), .A2(new_n781), .A3(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT42), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n784), .A2(new_n707), .A3(new_n785), .A4(new_n738), .ZN(new_n786));
  AND3_X1   g600(.A1(new_n779), .A2(new_n786), .A3(KEYINPUT109), .ZN(new_n787));
  AOI21_X1  g601(.A(KEYINPUT109), .B1(new_n779), .B2(new_n786), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G131), .ZN(G33));
  NOR3_X1   g604(.A1(new_n780), .A2(new_n781), .A3(new_n710), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n791), .A2(new_n707), .A3(new_n738), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G134), .ZN(G36));
  AOI21_X1  g607(.A(KEYINPUT43), .B1(new_n448), .B2(KEYINPUT110), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n794), .B1(new_n682), .B2(new_n688), .ZN(new_n795));
  OAI211_X1 g609(.A(new_n782), .B(new_n448), .C1(KEYINPUT110), .C2(KEYINPUT43), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n698), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n701), .A2(new_n797), .ZN(new_n798));
  OR2_X1    g612(.A1(new_n798), .A2(KEYINPUT44), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n701), .A2(KEYINPUT44), .A3(new_n797), .ZN(new_n800));
  INV_X1    g614(.A(new_n780), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n800), .A2(KEYINPUT111), .A3(new_n801), .ZN(new_n802));
  OR2_X1    g616(.A1(new_n386), .A2(KEYINPUT45), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n386), .A2(KEYINPUT45), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n803), .A2(G469), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(G469), .A2(G902), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT46), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n809), .A2(new_n392), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n807), .A2(new_n808), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n317), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(new_n714), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n799), .A2(new_n802), .A3(new_n814), .ZN(new_n815));
  AOI21_X1  g629(.A(KEYINPUT111), .B1(new_n800), .B2(new_n801), .ZN(new_n816));
  OR2_X1    g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(G137), .ZN(G39));
  XNOR2_X1  g632(.A(new_n812), .B(KEYINPUT47), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n595), .A2(new_n631), .A3(new_n776), .A4(new_n801), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  XOR2_X1   g635(.A(new_n821), .B(G140), .Z(G42));
  INV_X1    g636(.A(KEYINPUT53), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT112), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n743), .B1(new_n684), .B2(new_n690), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n699), .B1(new_n573), .B2(new_n594), .ZN(new_n826));
  OAI22_X1  g640(.A1(new_n826), .A2(new_n752), .B1(new_n757), .B2(new_n764), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n824), .B1(new_n825), .B2(new_n827), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n741), .B1(new_n636), .B2(new_n642), .ZN(new_n829));
  AND3_X1   g643(.A1(new_n672), .A2(new_n674), .A3(new_n494), .ZN(new_n830));
  OAI211_X1 g644(.A(new_n829), .B(new_n830), .C1(new_n683), .C2(new_n689), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n831), .A2(new_n754), .A3(new_n765), .A4(KEYINPUT112), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n828), .A2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(new_n689), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n497), .B1(new_n733), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n312), .A2(new_n835), .ZN(new_n836));
  OAI22_X1  g650(.A1(new_n668), .A2(new_n836), .B1(new_n700), .B2(new_n701), .ZN(new_n837));
  XNOR2_X1  g651(.A(new_n643), .B(new_n644), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n837), .B1(new_n838), .B2(new_n499), .ZN(new_n839));
  INV_X1    g653(.A(new_n698), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n784), .A2(new_n769), .A3(new_n840), .ZN(new_n841));
  OR2_X1    g655(.A1(new_n734), .A2(new_n496), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n780), .A2(new_n664), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n843), .A2(new_n707), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n792), .A2(new_n841), .A3(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n845), .A2(KEYINPUT113), .ZN(new_n846));
  AOI22_X1  g660(.A1(new_n643), .A2(new_n791), .B1(new_n843), .B2(new_n707), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT113), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n847), .A2(new_n848), .A3(new_n841), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n846), .A2(new_n849), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n833), .A2(new_n789), .A3(new_n839), .A4(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT52), .ZN(new_n852));
  OAI211_X1 g666(.A(new_n705), .B(new_n707), .C1(new_n711), .C2(new_n735), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(new_n770), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n781), .A2(new_n840), .A3(new_n775), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n855), .A2(new_n674), .A3(new_n672), .A4(new_n718), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n856), .B1(new_n729), .B2(new_n727), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n852), .B1(new_n854), .B2(new_n857), .ZN(new_n858));
  AND3_X1   g672(.A1(new_n672), .A2(new_n674), .A3(new_n718), .ZN(new_n859));
  AND3_X1   g673(.A1(new_n636), .A2(new_n728), .A3(new_n725), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n728), .B1(new_n636), .B2(new_n725), .ZN(new_n861));
  OAI211_X1 g675(.A(new_n859), .B(new_n855), .C1(new_n860), .C2(new_n861), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n862), .A2(new_n853), .A3(KEYINPUT52), .A4(new_n770), .ZN(new_n863));
  AND2_X1   g677(.A1(new_n858), .A2(new_n863), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n823), .B1(new_n851), .B2(new_n864), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n825), .A2(new_n827), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n779), .A2(new_n786), .A3(KEYINPUT53), .ZN(new_n867));
  INV_X1    g681(.A(new_n668), .ZN(new_n868));
  INV_X1    g682(.A(new_n836), .ZN(new_n869));
  INV_X1    g683(.A(new_n701), .ZN(new_n870));
  AND3_X1   g684(.A1(new_n312), .A2(new_n393), .A3(new_n699), .ZN(new_n871));
  AOI22_X1  g685(.A1(new_n868), .A2(new_n869), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n866), .A2(new_n646), .A3(new_n867), .A4(new_n872), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n848), .B1(new_n847), .B2(new_n841), .ZN(new_n874));
  AND4_X1   g688(.A1(new_n848), .A2(new_n792), .A3(new_n841), .A4(new_n844), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n873), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n862), .A2(new_n853), .A3(new_n770), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT114), .ZN(new_n879));
  AOI22_X1  g693(.A1(new_n858), .A2(new_n863), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n878), .A2(new_n879), .A3(KEYINPUT52), .ZN(new_n881));
  INV_X1    g695(.A(new_n881), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n877), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT54), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n865), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  OR2_X1    g699(.A1(new_n885), .A2(KEYINPUT115), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n885), .A2(KEYINPUT115), .ZN(new_n887));
  OAI21_X1  g701(.A(KEYINPUT53), .B1(new_n851), .B2(new_n864), .ZN(new_n888));
  OR2_X1    g702(.A1(new_n851), .A2(KEYINPUT53), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n880), .A2(new_n882), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n888), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  OAI211_X1 g705(.A(new_n886), .B(new_n887), .C1(new_n884), .C2(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n795), .A2(new_n796), .ZN(new_n893));
  INV_X1    g707(.A(new_n708), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n751), .A2(new_n801), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(new_n773), .ZN(new_n898));
  AND4_X1   g712(.A1(KEYINPUT118), .A2(new_n897), .A3(KEYINPUT48), .A4(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n897), .A2(new_n898), .ZN(new_n900));
  XOR2_X1   g714(.A(KEYINPUT118), .B(KEYINPUT48), .Z(new_n901));
  AOI21_X1  g715(.A(new_n899), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n273), .A2(G952), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n895), .A2(new_n764), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n903), .B1(new_n904), .B2(new_n753), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n896), .A2(new_n489), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n727), .A2(new_n906), .A3(new_n738), .A4(new_n729), .ZN(new_n907));
  OAI211_X1 g721(.A(new_n902), .B(new_n905), .C1(new_n733), .C2(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n897), .A2(new_n840), .A3(new_n769), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n448), .A2(new_n682), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n909), .B1(new_n907), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n819), .B1(new_n653), .B2(new_n749), .ZN(new_n912));
  NOR3_X1   g726(.A1(new_n895), .A2(new_n764), .A3(new_n780), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n911), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NOR4_X1   g728(.A1(new_n717), .A2(new_n311), .A3(new_n750), .A4(new_n749), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(new_n904), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT50), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  XOR2_X1   g732(.A(new_n918), .B(KEYINPUT117), .Z(new_n919));
  NAND2_X1  g733(.A1(new_n916), .A2(new_n917), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n920), .B(KEYINPUT116), .Z(new_n921));
  OAI21_X1  g735(.A(new_n914), .B1(new_n919), .B2(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT51), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n908), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n924), .B1(new_n923), .B2(new_n922), .ZN(new_n925));
  OAI22_X1  g739(.A1(new_n892), .A2(new_n925), .B1(G952), .B2(G953), .ZN(new_n926));
  OR2_X1    g740(.A1(new_n749), .A2(KEYINPUT49), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n749), .A2(KEYINPUT49), .ZN(new_n928));
  AND4_X1   g742(.A1(new_n448), .A2(new_n782), .A3(new_n311), .A4(new_n653), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n927), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  OR4_X1    g744(.A1(new_n631), .A2(new_n730), .A3(new_n717), .A4(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n926), .A2(new_n931), .ZN(G75));
  NOR2_X1   g746(.A1(new_n273), .A2(G952), .ZN(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n389), .B1(new_n865), .B2(new_n883), .ZN(new_n935));
  AOI21_X1  g749(.A(KEYINPUT56), .B1(new_n935), .B2(new_n308), .ZN(new_n936));
  AND2_X1   g750(.A1(new_n255), .A2(new_n256), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(new_n287), .ZN(new_n938));
  XNOR2_X1  g752(.A(KEYINPUT119), .B(KEYINPUT55), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n938), .B(new_n939), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n934), .B1(new_n936), .B2(new_n940), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n941), .B1(new_n936), .B2(new_n940), .ZN(G51));
  INV_X1    g756(.A(KEYINPUT120), .ZN(new_n943));
  AOI211_X1 g757(.A(new_n389), .B(new_n805), .C1(new_n865), .C2(new_n883), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n806), .B(KEYINPUT57), .Z(new_n945));
  AND3_X1   g759(.A1(new_n865), .A2(new_n883), .A3(new_n884), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n884), .B1(new_n865), .B2(new_n883), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n945), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n390), .A2(new_n391), .ZN(new_n949));
  INV_X1    g763(.A(new_n949), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n944), .B1(new_n948), .B2(new_n950), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n943), .B1(new_n951), .B2(new_n933), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n865), .A2(new_n883), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n953), .A2(KEYINPUT54), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(new_n885), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n949), .B1(new_n955), .B2(new_n945), .ZN(new_n956));
  OAI211_X1 g770(.A(KEYINPUT120), .B(new_n934), .C1(new_n956), .C2(new_n944), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n952), .A2(new_n957), .ZN(G54));
  NAND2_X1  g772(.A1(KEYINPUT58), .A2(G475), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n959), .B(KEYINPUT121), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n935), .A2(new_n960), .ZN(new_n961));
  AND2_X1   g775(.A1(new_n961), .A2(new_n438), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n961), .A2(new_n438), .ZN(new_n963));
  NOR3_X1   g777(.A1(new_n962), .A2(new_n963), .A3(new_n933), .ZN(G60));
  NAND2_X1  g778(.A1(G478), .A2(G902), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n965), .B(KEYINPUT59), .Z(new_n966));
  INV_X1    g780(.A(new_n966), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n955), .A2(new_n680), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n968), .A2(new_n934), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n892), .A2(new_n967), .ZN(new_n970));
  INV_X1    g784(.A(new_n680), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n969), .B1(new_n970), .B2(new_n971), .ZN(G63));
  NAND2_X1  g786(.A1(G217), .A2(G902), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n973), .B(KEYINPUT60), .Z(new_n974));
  NAND2_X1  g788(.A1(new_n953), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n975), .A2(new_n624), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n953), .A2(new_n695), .A3(new_n974), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n976), .A2(new_n934), .A3(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(KEYINPUT122), .ZN(new_n979));
  AND3_X1   g793(.A1(new_n978), .A2(new_n979), .A3(KEYINPUT61), .ZN(new_n980));
  AOI21_X1  g794(.A(KEYINPUT61), .B1(new_n978), .B2(new_n979), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n980), .A2(new_n981), .ZN(G66));
  AOI21_X1  g796(.A(new_n273), .B1(new_n493), .B2(G224), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n833), .A2(new_n839), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n983), .B1(new_n984), .B2(new_n273), .ZN(new_n985));
  INV_X1    g799(.A(G898), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n937), .B1(new_n986), .B2(G953), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n987), .B(KEYINPUT123), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n985), .B(new_n988), .ZN(G69));
  NOR2_X1   g803(.A1(new_n731), .A2(new_n854), .ZN(new_n990));
  INV_X1    g804(.A(KEYINPUT62), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n992), .B1(new_n819), .B2(new_n820), .ZN(new_n993));
  INV_X1    g807(.A(new_n993), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n990), .A2(new_n991), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n995), .A2(KEYINPUT124), .ZN(new_n996));
  INV_X1    g810(.A(new_n996), .ZN(new_n997));
  NOR2_X1   g811(.A1(new_n995), .A2(KEYINPUT124), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n994), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  INV_X1    g813(.A(KEYINPUT125), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n715), .B1(new_n733), .B2(new_n834), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n838), .A2(new_n801), .A3(new_n1001), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n1000), .B1(new_n817), .B2(new_n1002), .ZN(new_n1003));
  OAI211_X1 g817(.A(new_n1000), .B(new_n1002), .C1(new_n815), .C2(new_n816), .ZN(new_n1004));
  INV_X1    g818(.A(new_n1004), .ZN(new_n1005));
  NOR2_X1   g819(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g820(.A(KEYINPUT126), .B1(new_n999), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n817), .A2(new_n1002), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1008), .A2(KEYINPUT125), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1009), .A2(new_n1004), .ZN(new_n1010));
  INV_X1    g824(.A(KEYINPUT126), .ZN(new_n1011));
  OR2_X1    g825(.A1(new_n995), .A2(KEYINPUT124), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n993), .B1(new_n1012), .B2(new_n996), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n1010), .A2(new_n1011), .A3(new_n1013), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1007), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n563), .A2(new_n518), .ZN(new_n1016));
  XOR2_X1   g830(.A(new_n1016), .B(new_n406), .Z(new_n1017));
  INV_X1    g831(.A(new_n1017), .ZN(new_n1018));
  NAND3_X1  g832(.A1(new_n1015), .A2(new_n273), .A3(new_n1018), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n1017), .B1(G227), .B2(new_n273), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1020), .A2(G900), .ZN(new_n1021));
  NOR2_X1   g835(.A1(new_n1017), .A2(G227), .ZN(new_n1022));
  OAI21_X1  g836(.A(G953), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g837(.A1(new_n814), .A2(new_n859), .A3(new_n898), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1024), .A2(new_n792), .ZN(new_n1025));
  NOR3_X1   g839(.A1(new_n821), .A2(new_n1025), .A3(new_n854), .ZN(new_n1026));
  NAND3_X1  g840(.A1(new_n1026), .A2(new_n789), .A3(new_n817), .ZN(new_n1027));
  OAI211_X1 g841(.A(new_n1019), .B(new_n1023), .C1(new_n1020), .C2(new_n1027), .ZN(G72));
  NAND2_X1  g842(.A1(G472), .A2(G902), .ZN(new_n1029));
  XOR2_X1   g843(.A(new_n1029), .B(KEYINPUT63), .Z(new_n1030));
  OAI21_X1  g844(.A(new_n1030), .B1(new_n1027), .B2(new_n984), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n548), .A2(new_n589), .ZN(new_n1032));
  NOR2_X1   g846(.A1(new_n1032), .A2(new_n542), .ZN(new_n1033));
  AOI21_X1  g847(.A(new_n933), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g848(.A1(new_n1032), .A2(new_n568), .ZN(new_n1035));
  NAND3_X1  g849(.A1(new_n1035), .A2(new_n544), .A3(new_n550), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n1036), .A2(new_n1030), .ZN(new_n1037));
  OAI21_X1  g851(.A(new_n1034), .B1(new_n891), .B2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g852(.A(new_n1030), .B1(new_n1015), .B2(new_n984), .ZN(new_n1039));
  AOI21_X1  g853(.A(new_n568), .B1(new_n548), .B2(new_n589), .ZN(new_n1040));
  AOI21_X1  g854(.A(new_n1038), .B1(new_n1039), .B2(new_n1040), .ZN(G57));
endmodule


