//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 0 0 1 0 1 1 0 0 0 0 0 1 1 0 0 1 0 1 0 0 0 0 0 0 1 0 0 0 0 1 0 0 0 1 0 1 0 0 0 1 0 0 1 1 1 0 0 0 0 1 1 0 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:47 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1282, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1348, new_n1349, new_n1350, new_n1351, new_n1352, new_n1353,
    new_n1354;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G68), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  AOI22_X1  g0005(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n206), .B(KEYINPUT65), .ZN(new_n207));
  INV_X1    g0007(.A(G68), .ZN(new_n208));
  INV_X1    g0008(.A(G238), .ZN(new_n209));
  INV_X1    g0009(.A(G87), .ZN(new_n210));
  INV_X1    g0010(.A(G250), .ZN(new_n211));
  OAI22_X1  g0011(.A1(new_n208), .A2(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  AOI21_X1  g0012(.A(new_n212), .B1(G58), .B2(G232), .ZN(new_n213));
  XNOR2_X1  g0013(.A(KEYINPUT66), .B(G244), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(G77), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G97), .A2(G257), .B1(G107), .B2(G264), .ZN(new_n217));
  NAND4_X1  g0017(.A1(new_n207), .A2(new_n213), .A3(new_n216), .A4(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G20), .ZN(new_n219));
  AND2_X1   g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(KEYINPUT1), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT67), .ZN(new_n223));
  OAI21_X1  g0023(.A(G50), .B1(G58), .B2(G68), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT64), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  INV_X1    g0026(.A(G20), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n225), .A2(new_n228), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n219), .A2(G13), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n230), .B(G250), .C1(G257), .C2(G264), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT0), .ZN(new_n232));
  OAI211_X1 g0032(.A(new_n229), .B(new_n232), .C1(new_n220), .C2(new_n221), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n223), .A2(new_n233), .ZN(G361));
  XOR2_X1   g0034(.A(G238), .B(G244), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XOR2_X1   g0036(.A(KEYINPUT2), .B(G226), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G264), .B(G270), .Z(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G107), .B(G116), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(KEYINPUT69), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G87), .B(G97), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G68), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(KEYINPUT68), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G50), .B(G58), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n246), .B(new_n250), .ZN(G351));
  NOR2_X1   g0051(.A1(G20), .A2(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(G50), .ZN(new_n253));
  INV_X1    g0053(.A(G77), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n227), .A2(G33), .ZN(new_n255));
  OAI221_X1 g0055(.A(new_n253), .B1(new_n227), .B2(G68), .C1(new_n254), .C2(new_n255), .ZN(new_n256));
  NAND3_X1  g0056(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(new_n226), .ZN(new_n258));
  AND2_X1   g0058(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G1), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(G20), .ZN(new_n261));
  XNOR2_X1  g0061(.A(new_n261), .B(KEYINPUT73), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n260), .A2(G13), .A3(G20), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n264), .A2(new_n258), .ZN(new_n265));
  AND2_X1   g0065(.A1(new_n262), .A2(new_n265), .ZN(new_n266));
  AOI22_X1  g0066(.A1(new_n259), .A2(KEYINPUT11), .B1(new_n266), .B2(G68), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT75), .ZN(new_n268));
  AOI21_X1  g0068(.A(KEYINPUT11), .B1(new_n256), .B2(new_n258), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n263), .A2(G68), .ZN(new_n270));
  XNOR2_X1  g0070(.A(new_n270), .B(KEYINPUT12), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  AND3_X1   g0072(.A1(new_n267), .A2(new_n268), .A3(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n268), .B1(new_n267), .B2(new_n272), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT13), .ZN(new_n277));
  AND2_X1   g0077(.A1(KEYINPUT3), .A2(G33), .ZN(new_n278));
  NOR2_X1   g0078(.A1(KEYINPUT3), .A2(G33), .ZN(new_n279));
  OAI211_X1 g0079(.A(G232), .B(G1698), .C1(new_n278), .C2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(G33), .A2(G97), .ZN(new_n281));
  OR2_X1    g0081(.A1(KEYINPUT71), .A2(G1698), .ZN(new_n282));
  NAND2_X1  g0082(.A1(KEYINPUT71), .A2(G1698), .ZN(new_n283));
  OAI211_X1 g0083(.A(new_n282), .B(new_n283), .C1(new_n278), .C2(new_n279), .ZN(new_n284));
  INV_X1    g0084(.A(G226), .ZN(new_n285));
  OAI211_X1 g0085(.A(new_n280), .B(new_n281), .C1(new_n284), .C2(new_n285), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n226), .B1(G33), .B2(G41), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n260), .B1(G41), .B2(G45), .ZN(new_n289));
  INV_X1    g0089(.A(G274), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(G33), .A2(G41), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n293), .A2(G1), .A3(G13), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT70), .ZN(new_n295));
  AND3_X1   g0095(.A1(new_n294), .A2(new_n295), .A3(new_n289), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n295), .B1(new_n294), .B2(new_n289), .ZN(new_n297));
  OAI21_X1  g0097(.A(G238), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  AND4_X1   g0098(.A1(new_n277), .A2(new_n288), .A3(new_n292), .A4(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n294), .A2(new_n289), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(KEYINPUT70), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n294), .A2(new_n295), .A3(new_n289), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n291), .B1(new_n303), .B2(G238), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n277), .B1(new_n304), .B2(new_n288), .ZN(new_n305));
  OAI21_X1  g0105(.A(G200), .B1(new_n299), .B2(new_n305), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n299), .A2(new_n305), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(G190), .ZN(new_n308));
  AND3_X1   g0108(.A1(new_n276), .A2(new_n306), .A3(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT76), .ZN(new_n310));
  AND2_X1   g0110(.A1(new_n286), .A2(new_n287), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n298), .A2(new_n292), .ZN(new_n312));
  OAI21_X1  g0112(.A(KEYINPUT13), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n304), .A2(new_n277), .A3(new_n288), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n313), .A2(G179), .A3(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(G169), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n316), .B1(new_n313), .B2(new_n314), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT14), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n315), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  AOI211_X1 g0119(.A(KEYINPUT14), .B(new_n316), .C1(new_n313), .C2(new_n314), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n310), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  OAI21_X1  g0121(.A(G169), .B1(new_n299), .B2(new_n305), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(KEYINPUT14), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n317), .A2(new_n318), .ZN(new_n324));
  NAND4_X1  g0124(.A1(new_n323), .A2(new_n324), .A3(KEYINPUT76), .A4(new_n315), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n321), .A2(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n309), .B1(new_n326), .B2(new_n275), .ZN(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  XNOR2_X1  g0128(.A(KEYINPUT8), .B(G58), .ZN(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n330), .A2(new_n264), .ZN(new_n331));
  INV_X1    g0131(.A(new_n266), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n331), .B1(new_n332), .B2(new_n330), .ZN(new_n333));
  INV_X1    g0133(.A(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT16), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n202), .A2(new_n208), .ZN(new_n336));
  NOR2_X1   g0136(.A1(G58), .A2(G68), .ZN(new_n337));
  OAI21_X1  g0137(.A(G20), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n252), .A2(G159), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  OR2_X1    g0140(.A1(KEYINPUT3), .A2(G33), .ZN(new_n341));
  NAND2_X1  g0141(.A1(KEYINPUT3), .A2(G33), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n341), .A2(new_n227), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(KEYINPUT7), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT7), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n341), .A2(new_n345), .A3(new_n227), .A4(new_n342), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n344), .A2(G68), .A3(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT77), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND4_X1  g0149(.A1(new_n344), .A2(KEYINPUT77), .A3(G68), .A4(new_n346), .ZN(new_n350));
  AOI211_X1 g0150(.A(new_n335), .B(new_n340), .C1(new_n349), .C2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n340), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(new_n347), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(new_n335), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(new_n258), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n334), .B1(new_n351), .B2(new_n355), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n278), .A2(new_n279), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n282), .A2(G223), .A3(new_n283), .ZN(new_n358));
  NAND2_X1  g0158(.A1(G226), .A2(G1698), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n357), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(G33), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n361), .A2(new_n210), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n287), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n300), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n291), .B1(new_n364), .B2(G232), .ZN(new_n365));
  AND2_X1   g0165(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(G179), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n367), .B1(new_n316), .B2(new_n366), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n356), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(KEYINPUT18), .ZN(new_n370));
  INV_X1    g0170(.A(G200), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n371), .B1(new_n363), .B2(new_n365), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n372), .B1(G190), .B2(new_n366), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n373), .B(new_n334), .C1(new_n351), .C2(new_n355), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT17), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n340), .B1(new_n349), .B2(new_n350), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(KEYINPUT16), .ZN(new_n378));
  INV_X1    g0178(.A(new_n258), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n379), .B1(new_n353), .B2(new_n335), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n333), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n381), .A2(KEYINPUT17), .A3(new_n373), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT18), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n356), .A2(new_n368), .A3(new_n383), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n370), .A2(new_n376), .A3(new_n382), .A4(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n341), .A2(new_n342), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(G1698), .ZN(new_n388));
  INV_X1    g0188(.A(G223), .ZN(new_n389));
  OAI22_X1  g0189(.A1(new_n388), .A2(new_n389), .B1(new_n254), .B2(new_n387), .ZN(new_n390));
  AND2_X1   g0190(.A1(KEYINPUT71), .A2(G1698), .ZN(new_n391));
  NOR2_X1   g0191(.A1(KEYINPUT71), .A2(G1698), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  AND3_X1   g0193(.A1(new_n387), .A2(new_n393), .A3(G222), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n287), .B1(new_n390), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n303), .A2(G226), .ZN(new_n396));
  AND3_X1   g0196(.A1(new_n395), .A2(new_n292), .A3(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(G179), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  OAI21_X1  g0199(.A(G20), .B1(new_n203), .B2(G68), .ZN(new_n400));
  INV_X1    g0200(.A(G150), .ZN(new_n401));
  INV_X1    g0201(.A(new_n252), .ZN(new_n402));
  OAI221_X1 g0202(.A(new_n400), .B1(new_n401), .B2(new_n402), .C1(new_n255), .C2(new_n329), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(new_n258), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(KEYINPUT72), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n263), .A2(G50), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n406), .B1(new_n266), .B2(G50), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT72), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n403), .A2(new_n408), .A3(new_n258), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n405), .A2(new_n407), .A3(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n395), .A2(new_n292), .A3(new_n396), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(new_n316), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n399), .A2(new_n410), .A3(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT74), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT9), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n410), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n415), .A2(new_n416), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n405), .A2(new_n407), .A3(new_n418), .A4(new_n409), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n395), .A2(G190), .A3(new_n292), .A4(new_n396), .ZN(new_n421));
  OAI221_X1 g0221(.A(new_n421), .B1(KEYINPUT74), .B2(KEYINPUT9), .C1(new_n397), .C2(new_n371), .ZN(new_n422));
  OAI21_X1  g0222(.A(KEYINPUT10), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  XNOR2_X1  g0223(.A(new_n410), .B(new_n418), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n397), .A2(new_n371), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n421), .B1(KEYINPUT74), .B2(KEYINPUT9), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT10), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n424), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n414), .B1(new_n423), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n266), .A2(G77), .ZN(new_n431));
  XNOR2_X1  g0231(.A(KEYINPUT15), .B(G87), .ZN(new_n432));
  OAI22_X1  g0232(.A1(new_n432), .A2(new_n255), .B1(new_n227), .B2(new_n254), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n329), .A2(new_n402), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n258), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n431), .B(new_n435), .C1(G77), .C2(new_n263), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n387), .A2(new_n393), .A3(G232), .ZN(new_n437));
  INV_X1    g0237(.A(G107), .ZN(new_n438));
  OAI221_X1 g0238(.A(new_n437), .B1(new_n438), .B2(new_n387), .C1(new_n209), .C2(new_n388), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(new_n287), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n303), .A2(new_n215), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n440), .A2(new_n292), .A3(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n436), .B1(new_n443), .B2(G190), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n444), .B1(new_n371), .B2(new_n443), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n442), .A2(new_n316), .ZN(new_n446));
  AND2_X1   g0246(.A1(new_n446), .A2(new_n436), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n443), .A2(new_n398), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n386), .A2(new_n430), .A3(new_n445), .A4(new_n449), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n328), .A2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT23), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n452), .B1(new_n227), .B2(G107), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n438), .A2(KEYINPUT23), .A3(G20), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(G33), .A2(G116), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n455), .B1(G20), .B2(new_n456), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n227), .B(G87), .C1(new_n278), .C2(new_n279), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(KEYINPUT22), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT22), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n387), .A2(new_n460), .A3(new_n227), .A4(G87), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n457), .B1(new_n459), .B2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT84), .ZN(new_n463));
  NOR3_X1   g0263(.A1(new_n462), .A2(new_n463), .A3(KEYINPUT24), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n464), .A2(new_n379), .ZN(new_n465));
  AND2_X1   g0265(.A1(new_n459), .A2(new_n461), .ZN(new_n466));
  OAI21_X1  g0266(.A(KEYINPUT84), .B1(new_n466), .B2(new_n457), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n462), .A2(new_n463), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n467), .A2(new_n468), .A3(KEYINPUT24), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n465), .A2(new_n469), .ZN(new_n470));
  OR3_X1    g0270(.A1(new_n361), .A2(KEYINPUT78), .A3(G1), .ZN(new_n471));
  OAI21_X1  g0271(.A(KEYINPUT78), .B1(new_n361), .B2(G1), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n379), .A2(new_n471), .A3(new_n263), .A4(new_n472), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n473), .A2(new_n438), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT25), .ZN(new_n475));
  AOI211_X1 g0275(.A(G107), .B(new_n263), .C1(KEYINPUT85), .C2(new_n475), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n475), .A2(KEYINPUT85), .ZN(new_n477));
  OR2_X1    g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n476), .A2(new_n477), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n474), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n470), .A2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(G190), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT87), .ZN(new_n483));
  OAI211_X1 g0283(.A(G257), .B(G1698), .C1(new_n278), .C2(new_n279), .ZN(new_n484));
  NAND2_X1  g0284(.A1(G33), .A2(G294), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n484), .B(new_n485), .C1(new_n284), .C2(new_n211), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT86), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n294), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n387), .A2(new_n393), .A3(G250), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n489), .A2(KEYINPUT86), .A3(new_n484), .A4(new_n485), .ZN(new_n490));
  INV_X1    g0290(.A(G45), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n491), .A2(G1), .ZN(new_n492));
  XNOR2_X1  g0292(.A(KEYINPUT5), .B(G41), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n287), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  AOI22_X1  g0294(.A1(new_n488), .A2(new_n490), .B1(G264), .B2(new_n494), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n493), .A2(G274), .A3(new_n294), .A4(new_n492), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n483), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n486), .A2(new_n487), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n498), .A2(new_n287), .A3(new_n490), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n494), .A2(G264), .ZN(new_n500));
  AND4_X1   g0300(.A1(new_n483), .A2(new_n499), .A3(new_n496), .A4(new_n500), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n482), .B1(new_n497), .B2(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n499), .A2(new_n496), .A3(new_n500), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(new_n371), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n481), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(new_n480), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n506), .B1(new_n465), .B2(new_n469), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n503), .A2(KEYINPUT87), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n495), .A2(new_n483), .A3(new_n496), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n508), .A2(new_n509), .A3(G169), .ZN(new_n510));
  INV_X1    g0310(.A(new_n503), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(G179), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n507), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n505), .A2(new_n513), .ZN(new_n514));
  AND3_X1   g0314(.A1(new_n344), .A2(G107), .A3(new_n346), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n402), .A2(new_n254), .ZN(new_n516));
  INV_X1    g0316(.A(new_n516), .ZN(new_n517));
  AND3_X1   g0317(.A1(new_n438), .A2(KEYINPUT6), .A3(G97), .ZN(new_n518));
  XNOR2_X1  g0318(.A(G97), .B(G107), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT6), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n517), .B1(new_n521), .B2(new_n227), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n258), .B1(new_n515), .B2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(G97), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n264), .A2(new_n524), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n525), .B1(new_n473), .B2(new_n524), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n523), .A2(new_n527), .ZN(new_n528));
  AND2_X1   g0328(.A1(KEYINPUT5), .A2(G41), .ZN(new_n529));
  NOR2_X1   g0329(.A1(KEYINPUT5), .A2(G41), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n492), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(new_n294), .ZN(new_n532));
  INV_X1    g0332(.A(G257), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n496), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT4), .ZN(new_n535));
  INV_X1    g0335(.A(G244), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n535), .B1(new_n284), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(G33), .A2(G283), .ZN(new_n538));
  INV_X1    g0338(.A(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(G1698), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n540), .B1(new_n341), .B2(new_n342), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n539), .B1(new_n541), .B2(G250), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n387), .A2(new_n393), .A3(KEYINPUT4), .A4(G244), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n537), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n534), .B1(new_n544), .B2(new_n287), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n545), .A2(new_n316), .ZN(new_n546));
  AOI211_X1 g0346(.A(new_n398), .B(new_n534), .C1(new_n544), .C2(new_n287), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n528), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  OAI211_X1 g0348(.A(G250), .B(G1698), .C1(new_n278), .C2(new_n279), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n538), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n387), .A2(new_n393), .A3(G244), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n550), .B1(new_n535), .B2(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n294), .B1(new_n552), .B2(new_n543), .ZN(new_n553));
  OAI211_X1 g0353(.A(KEYINPUT80), .B(G200), .C1(new_n553), .C2(new_n534), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT80), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n555), .B1(new_n545), .B2(new_n371), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n523), .A2(KEYINPUT79), .A3(new_n527), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT79), .ZN(new_n559));
  AND2_X1   g0359(.A1(G97), .A2(G107), .ZN(new_n560));
  NOR2_X1   g0360(.A1(G97), .A2(G107), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n520), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n438), .A2(KEYINPUT6), .A3(G97), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n516), .B1(new_n564), .B2(G20), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n344), .A2(G107), .A3(new_n346), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n379), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n559), .B1(new_n567), .B2(new_n526), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n544), .A2(new_n287), .ZN(new_n569));
  INV_X1    g0369(.A(new_n534), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n569), .A2(new_n570), .A3(G190), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n558), .A2(new_n568), .A3(new_n571), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n548), .B1(new_n557), .B2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT19), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n227), .B1(new_n281), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n561), .A2(new_n210), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n227), .B(G68), .C1(new_n278), .C2(new_n279), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n574), .B1(new_n255), .B2(new_n524), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  AOI22_X1  g0380(.A1(new_n580), .A2(new_n258), .B1(new_n264), .B2(new_n432), .ZN(new_n581));
  AND2_X1   g0381(.A1(new_n471), .A2(new_n472), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n582), .A2(G87), .A3(new_n265), .ZN(new_n583));
  AND2_X1   g0383(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n260), .A2(G45), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(G250), .ZN(new_n586));
  OAI22_X1  g0386(.A1(new_n287), .A2(new_n586), .B1(new_n290), .B2(new_n585), .ZN(new_n587));
  OAI211_X1 g0387(.A(G244), .B(G1698), .C1(new_n278), .C2(new_n279), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n456), .B(new_n588), .C1(new_n284), .C2(new_n209), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n587), .B1(new_n589), .B2(new_n287), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(G190), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n584), .B(new_n591), .C1(new_n371), .C2(new_n590), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n580), .A2(new_n258), .ZN(new_n593));
  INV_X1    g0393(.A(new_n432), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n582), .A2(new_n265), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n432), .A2(new_n264), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n593), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT81), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  AND2_X1   g0399(.A1(new_n588), .A2(new_n456), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n387), .A2(new_n393), .A3(G238), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n294), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n316), .B1(new_n602), .B2(new_n587), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n581), .A2(KEYINPUT81), .A3(new_n595), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n590), .A2(new_n398), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n599), .A2(new_n603), .A3(new_n604), .A4(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n592), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g0407(.A(KEYINPUT82), .B1(new_n573), .B2(new_n607), .ZN(new_n608));
  AOI21_X1  g0408(.A(KEYINPUT79), .B1(new_n523), .B2(new_n527), .ZN(new_n609));
  NOR3_X1   g0409(.A1(new_n567), .A2(new_n559), .A3(new_n526), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n611), .A2(new_n571), .A3(new_n556), .A4(new_n554), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT82), .ZN(new_n613));
  AND2_X1   g0413(.A1(new_n592), .A2(new_n606), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n612), .A2(new_n613), .A3(new_n548), .A4(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n608), .A2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT21), .ZN(new_n617));
  OAI211_X1 g0417(.A(G264), .B(G1698), .C1(new_n278), .C2(new_n279), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n341), .A2(G303), .A3(new_n342), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n618), .B(new_n619), .C1(new_n284), .C2(new_n533), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(new_n287), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n531), .A2(G270), .A3(new_n294), .ZN(new_n622));
  AND2_X1   g0422(.A1(new_n622), .A2(new_n496), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(G169), .ZN(new_n625));
  INV_X1    g0425(.A(G116), .ZN(new_n626));
  AOI22_X1  g0426(.A1(new_n257), .A2(new_n226), .B1(G20), .B2(new_n626), .ZN(new_n627));
  OAI211_X1 g0427(.A(new_n538), .B(new_n227), .C1(G33), .C2(new_n524), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g0429(.A(new_n629), .B(KEYINPUT20), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n264), .A2(new_n626), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n631), .B1(new_n473), .B2(new_n626), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n617), .B1(new_n625), .B2(new_n633), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n624), .A2(KEYINPUT21), .A3(G169), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n621), .A2(new_n623), .A3(G179), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n633), .ZN(new_n638));
  AOI21_X1  g0438(.A(KEYINPUT83), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT83), .ZN(new_n640));
  AOI211_X1 g0440(.A(new_n640), .B(new_n633), .C1(new_n635), .C2(new_n636), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n634), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n624), .A2(new_n482), .ZN(new_n643));
  AOI211_X1 g0443(.A(new_n638), .B(new_n643), .C1(G200), .C2(new_n624), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  AND4_X1   g0445(.A1(new_n451), .A2(new_n514), .A3(new_n616), .A4(new_n645), .ZN(G372));
  NOR3_X1   g0446(.A1(new_n420), .A2(new_n422), .A3(KEYINPUT10), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n428), .B1(new_n424), .B2(new_n427), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n376), .A2(new_n382), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n309), .A2(new_n449), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n276), .B1(new_n321), .B2(new_n325), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n651), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n370), .A2(new_n384), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n649), .B1(new_n657), .B2(KEYINPUT89), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT89), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n654), .A2(new_n659), .A3(new_n656), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n414), .B1(new_n658), .B2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n451), .ZN(new_n662));
  OAI21_X1  g0462(.A(KEYINPUT88), .B1(new_n590), .B2(G169), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT88), .ZN(new_n664));
  OAI211_X1 g0464(.A(new_n664), .B(new_n316), .C1(new_n602), .C2(new_n587), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n663), .A2(new_n665), .A3(new_n597), .A4(new_n605), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(new_n592), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n573), .A2(new_n667), .ZN(new_n668));
  AOI21_X1  g0468(.A(G190), .B1(new_n508), .B2(new_n509), .ZN(new_n669));
  INV_X1    g0469(.A(new_n504), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n507), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n637), .A2(new_n638), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(new_n634), .ZN(new_n673));
  OAI211_X1 g0473(.A(new_n668), .B(new_n671), .C1(new_n513), .C2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n569), .A2(new_n570), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(G169), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n545), .A2(G179), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n678), .A2(new_n528), .A3(new_n592), .A4(new_n606), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(KEYINPUT26), .ZN(new_n680));
  AND2_X1   g0480(.A1(new_n666), .A2(new_n592), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT26), .ZN(new_n682));
  AOI22_X1  g0482(.A1(new_n676), .A2(new_n677), .B1(new_n558), .B2(new_n568), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n681), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  AND3_X1   g0484(.A1(new_n680), .A2(new_n684), .A3(new_n666), .ZN(new_n685));
  AND2_X1   g0485(.A1(new_n674), .A2(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n661), .B1(new_n662), .B2(new_n686), .ZN(G369));
  XNOR2_X1  g0487(.A(KEYINPUT92), .B(G330), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n260), .A2(new_n227), .A3(G13), .ZN(new_n689));
  XNOR2_X1  g0489(.A(new_n689), .B(KEYINPUT90), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT27), .ZN(new_n691));
  OR2_X1    g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n690), .A2(new_n691), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n692), .A2(new_n693), .A3(G213), .ZN(new_n694));
  INV_X1    g0494(.A(G343), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(new_n638), .ZN(new_n697));
  XOR2_X1   g0497(.A(new_n697), .B(KEYINPUT91), .Z(new_n698));
  NAND2_X1  g0498(.A1(new_n645), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n673), .ZN(new_n700));
  OR2_X1    g0500(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n688), .B1(new_n699), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n510), .A2(new_n512), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(new_n481), .ZN(new_n704));
  INV_X1    g0504(.A(new_n696), .ZN(new_n705));
  OAI211_X1 g0505(.A(new_n704), .B(new_n671), .C1(new_n507), .C2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n513), .A2(new_n696), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n702), .A2(new_n708), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n704), .A2(new_n671), .A3(new_n642), .A4(new_n705), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n513), .A2(new_n705), .ZN(new_n711));
  AOI21_X1  g0511(.A(KEYINPUT93), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n710), .A2(KEYINPUT93), .A3(new_n711), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n709), .B1(new_n712), .B2(new_n714), .ZN(new_n715));
  XOR2_X1   g0515(.A(new_n715), .B(KEYINPUT94), .Z(G399));
  NOR2_X1   g0516(.A1(new_n576), .A2(G116), .ZN(new_n717));
  INV_X1    g0517(.A(G41), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n230), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n717), .A2(G1), .A3(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n225), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n720), .B1(new_n721), .B2(new_n719), .ZN(new_n722));
  XOR2_X1   g0522(.A(new_n722), .B(KEYINPUT28), .Z(new_n723));
  OAI211_X1 g0523(.A(new_n668), .B(new_n671), .C1(new_n642), .C2(new_n513), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n666), .B1(new_n679), .B2(KEYINPUT26), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n682), .B1(new_n681), .B2(new_n683), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n696), .B1(new_n724), .B2(new_n727), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n728), .A2(KEYINPUT96), .A3(KEYINPUT29), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n696), .B1(new_n674), .B2(new_n685), .ZN(new_n731));
  OR2_X1    g0531(.A1(new_n731), .A2(KEYINPUT29), .ZN(new_n732));
  AOI21_X1  g0532(.A(KEYINPUT96), .B1(new_n728), .B2(KEYINPUT29), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n730), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n616), .A2(new_n514), .A3(new_n645), .A4(new_n705), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n545), .B1(new_n495), .B2(new_n496), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n590), .A2(G179), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT95), .ZN(new_n738));
  AND3_X1   g0538(.A1(new_n737), .A2(new_n738), .A3(new_n624), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n738), .B1(new_n737), .B2(new_n624), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n736), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n636), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n495), .A2(new_n742), .A3(new_n545), .A4(new_n590), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT30), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  AND2_X1   g0545(.A1(new_n545), .A2(new_n590), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n746), .A2(KEYINPUT30), .A3(new_n495), .A4(new_n742), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n741), .A2(new_n745), .A3(new_n747), .ZN(new_n748));
  AND3_X1   g0548(.A1(new_n748), .A2(KEYINPUT31), .A3(new_n696), .ZN(new_n749));
  AOI21_X1  g0549(.A(KEYINPUT31), .B1(new_n748), .B2(new_n696), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n688), .B1(new_n735), .B2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n734), .A2(new_n753), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n723), .B1(new_n754), .B2(new_n260), .ZN(new_n755));
  XNOR2_X1  g0555(.A(new_n755), .B(KEYINPUT97), .ZN(G364));
  AND2_X1   g0556(.A1(new_n227), .A2(G13), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n260), .B1(new_n757), .B2(G45), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n719), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n702), .A2(new_n761), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n699), .A2(new_n701), .A3(new_n688), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(G13), .A2(G33), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(G20), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n699), .A2(new_n701), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n387), .A2(new_n230), .ZN(new_n769));
  INV_X1    g0569(.A(G355), .ZN(new_n770));
  OAI22_X1  g0570(.A1(new_n769), .A2(new_n770), .B1(G116), .B2(new_n230), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n250), .A2(G45), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n357), .A2(new_n230), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n773), .B1(new_n225), .B2(new_n491), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n771), .B1(new_n772), .B2(new_n774), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n226), .B1(G20), .B2(new_n316), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n767), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n761), .B1(new_n775), .B2(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(G179), .A2(G200), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n227), .B1(new_n780), .B2(G190), .ZN(new_n781));
  XOR2_X1   g0581(.A(new_n781), .B(KEYINPUT101), .Z(new_n782));
  OR2_X1    g0582(.A1(new_n782), .A2(KEYINPUT102), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n782), .A2(KEYINPUT102), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(G97), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n227), .A2(new_n482), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n398), .A2(new_n371), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n227), .A2(G190), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  OAI22_X1  g0592(.A1(new_n790), .A2(new_n201), .B1(new_n792), .B2(new_n208), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n791), .A2(new_n780), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(G159), .ZN(new_n796));
  XNOR2_X1  g0596(.A(new_n796), .B(KEYINPUT32), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n371), .A2(G179), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n791), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  AOI211_X1 g0600(.A(new_n793), .B(new_n797), .C1(G107), .C2(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n788), .A2(new_n798), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n357), .B1(new_n803), .B2(G87), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n804), .A2(KEYINPUT100), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n398), .A2(G200), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n791), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(KEYINPUT99), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n807), .A2(KEYINPUT99), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n805), .B1(new_n812), .B2(G77), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n788), .A2(new_n806), .ZN(new_n814));
  XNOR2_X1  g0614(.A(new_n814), .B(KEYINPUT98), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  AOI22_X1  g0616(.A1(new_n816), .A2(G58), .B1(KEYINPUT100), .B2(new_n804), .ZN(new_n817));
  NAND4_X1  g0617(.A1(new_n787), .A2(new_n801), .A3(new_n813), .A4(new_n817), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n802), .B(KEYINPUT103), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n812), .A2(G311), .B1(G303), .B2(new_n819), .ZN(new_n820));
  XOR2_X1   g0620(.A(KEYINPUT33), .B(G317), .Z(new_n821));
  INV_X1    g0621(.A(G322), .ZN(new_n822));
  OAI22_X1  g0622(.A1(new_n821), .A2(new_n792), .B1(new_n814), .B2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(G326), .ZN(new_n824));
  INV_X1    g0624(.A(G329), .ZN(new_n825));
  OAI22_X1  g0625(.A1(new_n790), .A2(new_n824), .B1(new_n794), .B2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(G283), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n357), .B1(new_n799), .B2(new_n827), .ZN(new_n828));
  NOR3_X1   g0628(.A1(new_n823), .A2(new_n826), .A3(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(G294), .ZN(new_n830));
  OAI211_X1 g0630(.A(new_n820), .B(new_n829), .C1(new_n830), .C2(new_n782), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n818), .A2(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n779), .B1(new_n832), .B2(new_n776), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n768), .A2(new_n833), .ZN(new_n834));
  AND2_X1   g0634(.A1(new_n764), .A2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(G396));
  NAND2_X1  g0636(.A1(new_n696), .A2(new_n436), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n445), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n838), .A2(new_n449), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n447), .A2(new_n448), .A3(new_n705), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  XNOR2_X1  g0642(.A(new_n731), .B(new_n842), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n761), .B1(new_n843), .B2(new_n753), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n844), .B1(new_n753), .B2(new_n843), .ZN(new_n845));
  INV_X1    g0645(.A(G303), .ZN(new_n846));
  OAI22_X1  g0646(.A1(new_n790), .A2(new_n846), .B1(new_n792), .B2(new_n827), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n847), .B1(new_n812), .B2(G116), .ZN(new_n848));
  OR2_X1    g0648(.A1(new_n848), .A2(KEYINPUT106), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n848), .A2(KEYINPUT106), .ZN(new_n850));
  INV_X1    g0650(.A(G311), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n357), .B1(new_n794), .B2(new_n851), .ZN(new_n852));
  OAI22_X1  g0652(.A1(new_n814), .A2(new_n830), .B1(new_n799), .B2(new_n210), .ZN(new_n853));
  AOI211_X1 g0653(.A(new_n852), .B(new_n853), .C1(new_n819), .C2(G107), .ZN(new_n854));
  AND4_X1   g0654(.A1(new_n787), .A2(new_n849), .A3(new_n850), .A4(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n790), .ZN(new_n856));
  INV_X1    g0656(.A(new_n792), .ZN(new_n857));
  AOI22_X1  g0657(.A1(G137), .A2(new_n856), .B1(new_n857), .B2(G150), .ZN(new_n858));
  INV_X1    g0658(.A(G143), .ZN(new_n859));
  INV_X1    g0659(.A(G159), .ZN(new_n860));
  OAI221_X1 g0660(.A(new_n858), .B1(new_n815), .B2(new_n859), .C1(new_n811), .C2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT34), .ZN(new_n862));
  AND2_X1   g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n861), .A2(new_n862), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n819), .A2(G50), .ZN(new_n865));
  INV_X1    g0665(.A(G132), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n387), .B1(new_n794), .B2(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n867), .B1(G68), .B2(new_n800), .ZN(new_n868));
  OAI211_X1 g0668(.A(new_n865), .B(new_n868), .C1(new_n202), .C2(new_n782), .ZN(new_n869));
  NOR3_X1   g0669(.A1(new_n863), .A2(new_n864), .A3(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n776), .B1(new_n855), .B2(new_n870), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n776), .A2(new_n765), .ZN(new_n872));
  XOR2_X1   g0672(.A(new_n872), .B(KEYINPUT104), .Z(new_n873));
  OAI21_X1  g0673(.A(new_n761), .B1(new_n873), .B2(G77), .ZN(new_n874));
  XNOR2_X1  g0674(.A(new_n874), .B(KEYINPUT105), .ZN(new_n875));
  OAI211_X1 g0675(.A(new_n871), .B(new_n875), .C1(new_n842), .C2(new_n766), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n845), .A2(new_n876), .ZN(G384));
  OR2_X1    g0677(.A1(new_n564), .A2(KEYINPUT35), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n564), .A2(KEYINPUT35), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n878), .A2(new_n879), .A3(G116), .A4(new_n228), .ZN(new_n880));
  XOR2_X1   g0680(.A(new_n880), .B(KEYINPUT36), .Z(new_n881));
  OAI211_X1 g0681(.A(new_n225), .B(G77), .C1(new_n202), .C2(new_n208), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n208), .A2(G50), .ZN(new_n883));
  XNOR2_X1  g0683(.A(new_n883), .B(KEYINPUT107), .ZN(new_n884));
  AOI211_X1 g0684(.A(new_n260), .B(G13), .C1(new_n882), .C2(new_n884), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n881), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g0686(.A1(KEYINPUT109), .A2(KEYINPUT16), .ZN(new_n887));
  AND2_X1   g0687(.A1(new_n349), .A2(new_n350), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n887), .B1(new_n888), .B2(new_n340), .ZN(new_n889));
  INV_X1    g0689(.A(new_n887), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n379), .B1(new_n377), .B2(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n333), .B1(new_n889), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n374), .B1(new_n892), .B2(new_n694), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n889), .A2(new_n891), .ZN(new_n894));
  OR2_X1    g0694(.A1(new_n366), .A2(new_n316), .ZN(new_n895));
  AOI22_X1  g0695(.A1(new_n894), .A2(new_n334), .B1(new_n895), .B2(new_n367), .ZN(new_n896));
  OAI21_X1  g0696(.A(KEYINPUT37), .B1(new_n893), .B2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(new_n694), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n356), .A2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT37), .ZN(new_n900));
  NAND4_X1  g0700(.A1(new_n369), .A2(new_n899), .A3(new_n374), .A4(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n897), .A2(new_n901), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n892), .A2(new_n694), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n385), .A2(new_n903), .ZN(new_n904));
  AND3_X1   g0704(.A1(new_n902), .A2(KEYINPUT38), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(KEYINPUT38), .B1(new_n902), .B2(new_n904), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT39), .ZN(new_n907));
  NOR3_X1   g0707(.A1(new_n905), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(new_n899), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n385), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n369), .A2(new_n899), .A3(new_n374), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(KEYINPUT37), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n901), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n910), .A2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT38), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n902), .A2(KEYINPUT38), .A3(new_n904), .ZN(new_n917));
  AOI21_X1  g0717(.A(KEYINPUT39), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n908), .A2(new_n918), .ZN(new_n919));
  AOI22_X1  g0719(.A1(new_n322), .A2(KEYINPUT14), .B1(new_n307), .B2(G179), .ZN(new_n920));
  AOI21_X1  g0720(.A(KEYINPUT76), .B1(new_n920), .B2(new_n324), .ZN(new_n921));
  NOR3_X1   g0721(.A1(new_n319), .A2(new_n310), .A3(new_n320), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n275), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n923), .A2(new_n696), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n919), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n276), .A2(new_n705), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n326), .A2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT108), .ZN(new_n928));
  INV_X1    g0728(.A(new_n926), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n928), .B1(new_n327), .B2(new_n929), .ZN(new_n930));
  NOR4_X1   g0730(.A1(new_n653), .A2(KEYINPUT108), .A3(new_n309), .A4(new_n926), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n927), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n731), .A2(new_n842), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(new_n840), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n932), .B(new_n934), .C1(new_n905), .C2(new_n906), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n655), .A2(new_n694), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n925), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n657), .A2(KEYINPUT89), .ZN(new_n938));
  INV_X1    g0738(.A(new_n649), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n938), .A2(new_n939), .A3(new_n660), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(new_n413), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n724), .A2(new_n727), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n942), .A2(KEYINPUT29), .A3(new_n705), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT96), .ZN(new_n944));
  OAI211_X1 g0744(.A(new_n943), .B(new_n944), .C1(KEYINPUT29), .C2(new_n731), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n662), .B1(new_n945), .B2(new_n729), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n941), .A2(new_n946), .ZN(new_n947));
  XOR2_X1   g0747(.A(new_n937), .B(new_n947), .Z(new_n948));
  NAND2_X1  g0748(.A1(new_n916), .A2(new_n917), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n841), .B1(new_n735), .B2(new_n751), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n932), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(KEYINPUT40), .ZN(new_n952));
  INV_X1    g0752(.A(new_n906), .ZN(new_n953));
  AOI21_X1  g0753(.A(KEYINPUT40), .B1(new_n953), .B2(new_n917), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n954), .A2(new_n932), .A3(new_n950), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n952), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n735), .A2(new_n751), .ZN(new_n957));
  AND2_X1   g0757(.A1(new_n451), .A2(new_n957), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n956), .B(new_n958), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n948), .B1(new_n959), .B2(new_n688), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n960), .B1(new_n260), .B2(new_n757), .ZN(new_n961));
  NOR3_X1   g0761(.A1(new_n948), .A2(new_n959), .A3(new_n688), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n886), .B1(new_n961), .B2(new_n962), .ZN(G367));
  OAI221_X1 g0763(.A(new_n777), .B1(new_n230), .B2(new_n432), .C1(new_n241), .C2(new_n773), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n964), .A2(new_n761), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n819), .A2(KEYINPUT46), .A3(G116), .ZN(new_n966));
  OAI221_X1 g0766(.A(new_n966), .B1(new_n827), .B2(new_n811), .C1(new_n846), .C2(new_n815), .ZN(new_n967));
  AOI22_X1  g0767(.A1(new_n856), .A2(G311), .B1(new_n800), .B2(G97), .ZN(new_n968));
  INV_X1    g0768(.A(G317), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n968), .B1(new_n969), .B2(new_n794), .ZN(new_n970));
  AOI21_X1  g0770(.A(KEYINPUT46), .B1(new_n803), .B2(G116), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n357), .B1(new_n792), .B2(new_n830), .ZN(new_n972));
  NOR3_X1   g0772(.A1(new_n970), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n973), .B1(new_n438), .B2(new_n782), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n785), .A2(new_n208), .ZN(new_n975));
  AOI22_X1  g0775(.A1(G58), .A2(new_n803), .B1(new_n795), .B2(G137), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(KEYINPUT113), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n387), .B1(new_n790), .B2(new_n859), .ZN(new_n978));
  OAI22_X1  g0778(.A1(new_n792), .A2(new_n860), .B1(new_n799), .B2(new_n254), .ZN(new_n979));
  INV_X1    g0779(.A(new_n814), .ZN(new_n980));
  AOI211_X1 g0780(.A(new_n978), .B(new_n979), .C1(G150), .C2(new_n980), .ZN(new_n981));
  OAI211_X1 g0781(.A(new_n977), .B(new_n981), .C1(new_n201), .C2(new_n811), .ZN(new_n982));
  OAI22_X1  g0782(.A1(new_n967), .A2(new_n974), .B1(new_n975), .B2(new_n982), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(KEYINPUT47), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n965), .B1(new_n984), .B2(new_n776), .ZN(new_n985));
  OR2_X1    g0785(.A1(new_n705), .A2(new_n584), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n681), .A2(new_n986), .ZN(new_n987));
  OAI211_X1 g0787(.A(new_n987), .B(new_n767), .C1(new_n666), .C2(new_n986), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n985), .A2(new_n988), .ZN(new_n989));
  OAI211_X1 g0789(.A(new_n612), .B(new_n548), .C1(new_n611), .C2(new_n705), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n683), .A2(new_n696), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n992), .B1(new_n714), .B2(new_n712), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT45), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  OAI211_X1 g0795(.A(KEYINPUT45), .B(new_n992), .C1(new_n714), .C2(new_n712), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n710), .A2(new_n711), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT93), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n992), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n1000), .A2(new_n713), .A3(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT44), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND4_X1  g0804(.A1(new_n1000), .A2(KEYINPUT44), .A3(new_n713), .A4(new_n1001), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n997), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n709), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1008), .A2(KEYINPUT111), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1007), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n642), .A2(new_n705), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n706), .A2(new_n707), .A3(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1013), .A2(new_n710), .ZN(new_n1014));
  XOR2_X1   g0814(.A(new_n1014), .B(new_n702), .Z(new_n1015));
  NAND2_X1  g0815(.A1(new_n945), .A2(new_n729), .ZN(new_n1016));
  NOR3_X1   g0816(.A1(new_n1015), .A2(new_n1016), .A3(new_n752), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n997), .A2(new_n1006), .A3(new_n1009), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1011), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n754), .ZN(new_n1020));
  AND2_X1   g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n719), .B(KEYINPUT41), .ZN(new_n1022));
  OAI21_X1  g0822(.A(KEYINPUT112), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1022), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT112), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n759), .B1(new_n1023), .B2(new_n1026), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n709), .A2(new_n1001), .ZN(new_n1028));
  OR2_X1    g0828(.A1(new_n1001), .A2(new_n710), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n548), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n1029), .A2(KEYINPUT42), .B1(new_n1030), .B2(new_n705), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n711), .A2(KEYINPUT42), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n998), .A2(new_n992), .A3(new_n1032), .ZN(new_n1033));
  AND2_X1   g0833(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n987), .B1(new_n666), .B2(new_n986), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n1035), .A2(KEYINPUT43), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1034), .A2(new_n1036), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT110), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n1038), .ZN(new_n1039));
  XOR2_X1   g0839(.A(new_n1035), .B(KEYINPUT43), .Z(new_n1040));
  INV_X1    g0840(.A(new_n1040), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n1034), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n1042), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1028), .B1(new_n1039), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1028), .ZN(new_n1045));
  NOR3_X1   g0845(.A1(new_n1038), .A2(new_n1045), .A3(new_n1042), .ZN(new_n1046));
  OR2_X1    g0846(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n989), .B1(new_n1027), .B2(new_n1047), .ZN(G387));
  INV_X1    g0848(.A(new_n1017), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n754), .A2(new_n1015), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1049), .A2(new_n760), .A3(new_n1050), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n769), .A2(new_n717), .B1(G107), .B2(new_n230), .ZN(new_n1052));
  OR2_X1    g0852(.A1(new_n238), .A2(new_n491), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n717), .ZN(new_n1054));
  AOI211_X1 g0854(.A(G45), .B(new_n1054), .C1(G68), .C2(G77), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n329), .A2(G50), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT50), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n773), .B1(new_n1055), .B2(new_n1057), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1052), .B1(new_n1053), .B2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n761), .B1(new_n1059), .B2(new_n778), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n786), .A2(new_n594), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n330), .A2(new_n857), .B1(new_n795), .B2(G150), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1062), .B1(new_n860), .B2(new_n790), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n357), .B1(new_n800), .B2(G97), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n1064), .B1(new_n201), .B2(new_n814), .C1(new_n254), .C2(new_n802), .ZN(new_n1065));
  AOI211_X1 g0865(.A(new_n1063), .B(new_n1065), .C1(G68), .C2(new_n812), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1061), .A2(new_n1066), .ZN(new_n1067));
  XOR2_X1   g0867(.A(new_n1067), .B(KEYINPUT114), .Z(new_n1068));
  NAND2_X1  g0868(.A1(new_n803), .A2(G294), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(G322), .A2(new_n856), .B1(new_n857), .B2(G311), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n1070), .B1(new_n815), .B2(new_n969), .C1(new_n811), .C2(new_n846), .ZN(new_n1071));
  INV_X1    g0871(.A(KEYINPUT48), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n1069), .B1(new_n827), .B2(new_n782), .C1(new_n1071), .C2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1073), .B1(new_n1072), .B2(new_n1071), .ZN(new_n1074));
  XOR2_X1   g0874(.A(KEYINPUT115), .B(KEYINPUT49), .Z(new_n1075));
  XNOR2_X1  g0875(.A(new_n1074), .B(new_n1075), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n357), .B1(new_n794), .B2(new_n824), .C1(new_n626), .C2(new_n799), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1068), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1060), .B1(new_n1078), .B2(new_n776), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n767), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1079), .B1(new_n708), .B2(new_n1080), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n1051), .B(new_n1081), .C1(new_n758), .C2(new_n1015), .ZN(G393));
  NOR2_X1   g0882(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n709), .B1(new_n997), .B2(new_n1006), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  OAI21_X1  g0885(.A(KEYINPUT116), .B1(new_n1085), .B2(new_n1017), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT116), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n1049), .B(new_n1087), .C1(new_n1083), .C2(new_n1084), .ZN(new_n1088));
  NAND4_X1  g0888(.A1(new_n1086), .A2(new_n760), .A3(new_n1019), .A4(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1001), .A2(new_n767), .ZN(new_n1090));
  AND3_X1   g0890(.A1(new_n246), .A2(new_n230), .A3(new_n357), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n777), .B1(new_n524), .B2(new_n230), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n761), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n785), .A2(new_n254), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n387), .B1(new_n799), .B2(new_n210), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n792), .A2(new_n201), .B1(new_n794), .B2(new_n859), .ZN(new_n1096));
  AOI211_X1 g0896(.A(new_n1095), .B(new_n1096), .C1(G68), .C2(new_n803), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n812), .A2(new_n330), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(G150), .A2(new_n856), .B1(new_n980), .B2(G159), .ZN(new_n1099));
  OR2_X1    g0899(.A1(new_n1099), .A2(KEYINPUT51), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1099), .A2(KEYINPUT51), .ZN(new_n1101));
  NAND4_X1  g0901(.A1(new_n1097), .A2(new_n1098), .A3(new_n1100), .A4(new_n1101), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n790), .A2(new_n969), .B1(new_n814), .B2(new_n851), .ZN(new_n1103));
  XNOR2_X1  g0903(.A(new_n1103), .B(KEYINPUT52), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1104), .B1(new_n830), .B2(new_n811), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n802), .A2(new_n827), .B1(new_n794), .B2(new_n822), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1106), .B1(G303), .B2(new_n857), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n387), .B1(new_n800), .B2(G107), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n1107), .B(new_n1108), .C1(new_n626), .C2(new_n782), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n1094), .A2(new_n1102), .B1(new_n1105), .B2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1093), .B1(new_n1110), .B2(new_n776), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n1085), .A2(new_n759), .B1(new_n1090), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1089), .A2(new_n1112), .ZN(G390));
  INV_X1    g0913(.A(new_n927), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n309), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n923), .A2(new_n1115), .A3(new_n929), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(KEYINPUT108), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n327), .A2(new_n928), .A3(new_n929), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1114), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n950), .A2(G330), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  AOI211_X1 g0921(.A(new_n688), .B(new_n841), .C1(new_n735), .C2(new_n751), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n932), .A2(new_n1122), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n934), .B1(new_n1121), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n728), .A2(new_n839), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1125), .A2(new_n840), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1126), .B1(new_n932), .B2(new_n1122), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1124), .A2(new_n1129), .ZN(new_n1130));
  AND3_X1   g0930(.A1(new_n451), .A2(G330), .A3(new_n957), .ZN(new_n1131));
  NOR3_X1   g0931(.A1(new_n941), .A2(new_n946), .A3(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n924), .B1(new_n916), .B2(new_n917), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n840), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1135), .B1(new_n728), .B2(new_n839), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1134), .B1(new_n1119), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n932), .A2(new_n1122), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n924), .B1(new_n932), .B2(new_n934), .ZN(new_n1139));
  OAI211_X1 g0939(.A(new_n1137), .B(new_n1138), .C1(new_n1139), .C2(new_n919), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n924), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1135), .B1(new_n731), .B2(new_n842), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1141), .B1(new_n1119), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n949), .A2(new_n907), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n953), .A2(KEYINPUT39), .A3(new_n917), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n932), .A2(new_n1126), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(new_n1143), .A2(new_n1146), .B1(new_n1147), .B2(new_n1134), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n932), .A2(G330), .A3(new_n950), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1140), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1133), .A2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1137), .B1(new_n1139), .B2(new_n919), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1152), .A2(new_n1121), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n1153), .A2(new_n1130), .A3(new_n1132), .A4(new_n1140), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1151), .A2(new_n760), .A3(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1153), .A2(new_n759), .A3(new_n1140), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n761), .B1(new_n873), .B2(new_n330), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n857), .A2(G137), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(KEYINPUT54), .B(G143), .ZN(new_n1159));
  OAI221_X1 g0959(.A(new_n1158), .B1(new_n811), .B2(new_n1159), .C1(new_n785), .C2(new_n860), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(new_n1160), .B(KEYINPUT117), .ZN(new_n1161));
  INV_X1    g0961(.A(G128), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n802), .A2(new_n401), .ZN(new_n1163));
  INV_X1    g0963(.A(KEYINPUT53), .ZN(new_n1164));
  OAI221_X1 g0964(.A(new_n387), .B1(new_n1162), .B2(new_n790), .C1(new_n1163), .C2(new_n1164), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(G132), .A2(new_n980), .B1(new_n795), .B2(G125), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1166), .B1(new_n201), .B2(new_n799), .ZN(new_n1167));
  AOI211_X1 g0967(.A(new_n1165), .B(new_n1167), .C1(new_n1164), .C2(new_n1163), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1161), .A2(new_n1168), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n814), .A2(new_n626), .B1(new_n799), .B2(new_n208), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(G283), .A2(new_n856), .B1(new_n857), .B2(G107), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1171), .B1(new_n830), .B2(new_n794), .ZN(new_n1172));
  AOI211_X1 g0972(.A(new_n1170), .B(new_n1172), .C1(G97), .C2(new_n812), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n387), .B1(new_n819), .B2(G87), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(new_n1174), .B(KEYINPUT118), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n1173), .B(new_n1175), .C1(new_n254), .C2(new_n785), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(new_n1176), .B(KEYINPUT119), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1169), .A2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1157), .B1(new_n1178), .B2(new_n776), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1179), .B1(new_n919), .B2(new_n766), .ZN(new_n1180));
  AND2_X1   g0980(.A1(new_n1156), .A2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1155), .A2(new_n1181), .ZN(G378));
  INV_X1    g0982(.A(new_n937), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n413), .B1(new_n647), .B2(new_n648), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n410), .A2(new_n898), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT122), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(new_n1185), .B(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1184), .A2(new_n1187), .ZN(new_n1188));
  XOR2_X1   g0988(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1189));
  INV_X1    g0989(.A(new_n1187), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n430), .A2(new_n1190), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1188), .A2(new_n1189), .A3(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1189), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n430), .A2(new_n1190), .ZN(new_n1194));
  AOI211_X1 g0994(.A(new_n414), .B(new_n1187), .C1(new_n423), .C2(new_n429), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1193), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(new_n956), .A2(G330), .B1(new_n1192), .B2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(G330), .ZN(new_n1198));
  AND3_X1   g0998(.A1(new_n1196), .A2(new_n1192), .A3(KEYINPUT123), .ZN(new_n1199));
  AOI21_X1  g0999(.A(KEYINPUT123), .B1(new_n1196), .B2(new_n1192), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  AOI211_X1 g1001(.A(new_n1198), .B(new_n1201), .C1(new_n952), .C2(new_n955), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1183), .B1(new_n1197), .B2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1196), .A2(new_n1192), .ZN(new_n1204));
  AND2_X1   g1004(.A1(new_n932), .A2(new_n950), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(new_n1205), .A2(new_n954), .B1(new_n951), .B2(KEYINPUT40), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1204), .B1(new_n1206), .B2(new_n1198), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1201), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n956), .A2(G330), .A3(new_n1208), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1207), .A2(new_n1209), .A3(new_n937), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n758), .B1(new_n1203), .B2(new_n1210), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n201), .B1(new_n278), .B2(G41), .ZN(new_n1212));
  XNOR2_X1  g1012(.A(new_n1212), .B(KEYINPUT120), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(G97), .A2(new_n857), .B1(new_n795), .B2(G283), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1214), .B1(new_n626), .B2(new_n790), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n718), .B(new_n357), .C1(new_n802), .C2(new_n254), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n814), .A2(new_n438), .B1(new_n799), .B2(new_n202), .ZN(new_n1217));
  NOR3_X1   g1017(.A1(new_n1215), .A2(new_n1216), .A3(new_n1217), .ZN(new_n1218));
  OAI221_X1 g1018(.A(new_n1218), .B1(new_n432), .B2(new_n811), .C1(new_n785), .C2(new_n208), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT58), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1213), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1221));
  AOI211_X1 g1021(.A(G33), .B(G41), .C1(new_n795), .C2(G124), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n802), .A2(new_n1159), .ZN(new_n1223));
  XNOR2_X1  g1023(.A(new_n1223), .B(KEYINPUT121), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(G125), .A2(new_n856), .B1(new_n857), .B2(G132), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1225), .B1(new_n1162), .B2(new_n814), .ZN(new_n1226));
  AOI211_X1 g1026(.A(new_n1224), .B(new_n1226), .C1(G137), .C2(new_n812), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1227), .B1(new_n401), .B2(new_n785), .ZN(new_n1228));
  OAI221_X1 g1028(.A(new_n1222), .B1(new_n860), .B2(new_n799), .C1(new_n1228), .C2(KEYINPUT59), .ZN(new_n1229));
  AND2_X1   g1029(.A1(new_n1228), .A2(KEYINPUT59), .ZN(new_n1230));
  OAI221_X1 g1030(.A(new_n1221), .B1(new_n1220), .B2(new_n1219), .C1(new_n1229), .C2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1231), .A2(new_n776), .ZN(new_n1232));
  OAI211_X1 g1032(.A(new_n1232), .B(new_n761), .C1(G50), .C2(new_n873), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1233), .B1(new_n1208), .B2(new_n765), .ZN(new_n1234));
  OR2_X1    g1034(.A1(new_n1211), .A2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1203), .A2(new_n1210), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1119), .B1(new_n753), .B2(new_n841), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1237), .A2(new_n1149), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n1238), .A2(new_n934), .B1(new_n1128), .B2(new_n1127), .ZN(new_n1239));
  OAI211_X1 g1039(.A(KEYINPUT124), .B(new_n1132), .C1(new_n1150), .C2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(KEYINPUT124), .B1(new_n1154), .B2(new_n1132), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1236), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT57), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1132), .B1(new_n1150), .B2(new_n1239), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT124), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1248), .A2(new_n1240), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1244), .B1(new_n1203), .B2(new_n1210), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n719), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1235), .B1(new_n1245), .B2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(G375));
  INV_X1    g1053(.A(new_n1022), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1131), .ZN(new_n1255));
  OAI211_X1 g1055(.A(new_n661), .B(new_n1255), .C1(new_n734), .C2(new_n662), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1256), .A2(new_n1124), .A3(new_n1129), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1133), .A2(new_n1254), .A3(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1119), .A2(new_n765), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n761), .B1(new_n873), .B2(G68), .ZN(new_n1260));
  AOI22_X1  g1060(.A1(new_n856), .A2(G294), .B1(new_n795), .B2(G303), .ZN(new_n1261));
  OAI221_X1 g1061(.A(new_n1261), .B1(new_n626), .B2(new_n792), .C1(new_n827), .C2(new_n814), .ZN(new_n1262));
  AOI211_X1 g1062(.A(new_n387), .B(new_n1262), .C1(G77), .C2(new_n800), .ZN(new_n1263));
  AOI22_X1  g1063(.A1(new_n812), .A2(G107), .B1(G97), .B2(new_n819), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1263), .A2(new_n1061), .A3(new_n1264), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n785), .A2(new_n201), .ZN(new_n1266));
  AOI22_X1  g1066(.A1(new_n812), .A2(G150), .B1(new_n816), .B2(G137), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n387), .B1(new_n799), .B2(new_n202), .ZN(new_n1268));
  OAI22_X1  g1068(.A1(new_n790), .A2(new_n866), .B1(new_n792), .B2(new_n1159), .ZN(new_n1269));
  AOI211_X1 g1069(.A(new_n1268), .B(new_n1269), .C1(G128), .C2(new_n795), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n819), .A2(G159), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1267), .A2(new_n1270), .A3(new_n1271), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1265), .B1(new_n1266), .B2(new_n1272), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1260), .B1(new_n1273), .B2(new_n776), .ZN(new_n1274));
  AOI22_X1  g1074(.A1(new_n1130), .A2(new_n759), .B1(new_n1259), .B2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1258), .A2(new_n1275), .ZN(G381));
  INV_X1    g1076(.A(G387), .ZN(new_n1277));
  OR2_X1    g1077(.A1(G393), .A2(G396), .ZN(new_n1278));
  NOR4_X1   g1078(.A1(G390), .A2(new_n1278), .A3(G384), .A4(G381), .ZN(new_n1279));
  INV_X1    g1079(.A(G378), .ZN(new_n1280));
  NAND4_X1  g1080(.A1(new_n1277), .A2(new_n1279), .A3(new_n1252), .A4(new_n1280), .ZN(G407));
  NAND2_X1  g1081(.A1(new_n1252), .A2(new_n1280), .ZN(new_n1282));
  OAI211_X1 g1082(.A(G407), .B(G213), .C1(G343), .C2(new_n1282), .ZN(G409));
  XNOR2_X1  g1083(.A(G393), .B(new_n835), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n989), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1287));
  AOI211_X1 g1087(.A(KEYINPUT112), .B(new_n1022), .C1(new_n1019), .C2(new_n1020), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n758), .B1(new_n1287), .B2(new_n1288), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1290));
  AOI221_X4 g1090(.A(new_n1286), .B1(new_n1089), .B2(new_n1112), .C1(new_n1289), .C2(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1292));
  AOI21_X1  g1092(.A(G390), .B1(new_n1292), .B2(new_n989), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1285), .B1(new_n1291), .B2(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(G390), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(G387), .A2(new_n1295), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1292), .A2(new_n989), .A3(G390), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1296), .A2(new_n1284), .A3(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1294), .A2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT127), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1294), .A2(new_n1298), .A3(KEYINPUT127), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  AND2_X1   g1103(.A1(new_n695), .A2(G213), .ZN(new_n1304));
  NOR3_X1   g1104(.A1(G378), .A2(new_n1211), .A3(new_n1234), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1249), .A2(new_n1254), .A3(new_n1236), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1304), .B1(new_n1305), .B2(new_n1306), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n719), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT60), .ZN(new_n1309));
  AOI211_X1 g1109(.A(KEYINPUT125), .B(new_n1309), .C1(new_n1239), .C2(new_n1256), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT125), .ZN(new_n1311));
  AOI21_X1  g1111(.A(KEYINPUT60), .B1(new_n1257), .B2(new_n1311), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1308), .B1(new_n1310), .B2(new_n1312), .ZN(new_n1313));
  AND3_X1   g1113(.A1(new_n1313), .A2(G384), .A3(new_n1275), .ZN(new_n1314));
  AOI21_X1  g1114(.A(G384), .B1(new_n1313), .B2(new_n1275), .ZN(new_n1315));
  NOR2_X1   g1115(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1316));
  OAI211_X1 g1116(.A(new_n1307), .B(new_n1316), .C1(new_n1252), .C2(new_n1280), .ZN(new_n1317));
  OR2_X1    g1117(.A1(new_n1317), .A2(KEYINPUT62), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1307), .B1(new_n1252), .B2(new_n1280), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1304), .A2(G2897), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1320), .ZN(new_n1321));
  NOR3_X1   g1121(.A1(new_n1314), .A2(new_n1315), .A3(new_n1321), .ZN(new_n1322));
  INV_X1    g1122(.A(G384), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1308), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1257), .A2(new_n1311), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1325), .A2(new_n1309), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1257), .A2(new_n1311), .A3(KEYINPUT60), .ZN(new_n1327));
  AOI21_X1  g1127(.A(new_n1324), .B1(new_n1326), .B2(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1275), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1323), .B1(new_n1328), .B2(new_n1329), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1313), .A2(G384), .A3(new_n1275), .ZN(new_n1331));
  AOI21_X1  g1131(.A(new_n1320), .B1(new_n1330), .B2(new_n1331), .ZN(new_n1332));
  NOR2_X1   g1132(.A1(new_n1322), .A2(new_n1332), .ZN(new_n1333));
  AOI21_X1  g1133(.A(KEYINPUT61), .B1(new_n1319), .B2(new_n1333), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1317), .A2(KEYINPUT62), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1318), .A2(new_n1334), .A3(new_n1335), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1303), .A2(new_n1336), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT63), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1317), .A2(new_n1338), .ZN(new_n1339));
  AND2_X1   g1139(.A1(new_n1334), .A2(new_n1339), .ZN(new_n1340));
  OAI211_X1 g1140(.A(new_n1294), .B(new_n1298), .C1(new_n1317), .C2(new_n1338), .ZN(new_n1341));
  INV_X1    g1141(.A(new_n1341), .ZN(new_n1342));
  AOI21_X1  g1142(.A(KEYINPUT126), .B1(new_n1340), .B2(new_n1342), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1334), .A2(new_n1339), .ZN(new_n1344));
  INV_X1    g1144(.A(KEYINPUT126), .ZN(new_n1345));
  NOR3_X1   g1145(.A1(new_n1344), .A2(new_n1341), .A3(new_n1345), .ZN(new_n1346));
  OAI21_X1  g1146(.A(new_n1337), .B1(new_n1343), .B2(new_n1346), .ZN(G405));
  NAND2_X1  g1147(.A1(G375), .A2(G378), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1348), .A2(new_n1282), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1349), .A2(new_n1316), .ZN(new_n1350));
  OAI211_X1 g1150(.A(new_n1348), .B(new_n1282), .C1(new_n1315), .C2(new_n1314), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1350), .A2(new_n1351), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1303), .A2(new_n1352), .ZN(new_n1353));
  NAND4_X1  g1153(.A1(new_n1301), .A2(new_n1350), .A3(new_n1302), .A4(new_n1351), .ZN(new_n1354));
  AND2_X1   g1154(.A1(new_n1353), .A2(new_n1354), .ZN(G402));
endmodule


