//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 1 0 1 1 1 0 0 1 0 0 0 1 0 1 0 0 1 0 0 1 1 0 0 0 0 1 0 1 0 1 1 1 0 1 1 0 1 0 1 0 0 1 0 0 0 0 1 0 0 0 1 0 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:17 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n613, new_n614, new_n615, new_n616, new_n617,
    new_n618, new_n619, new_n620, new_n621, new_n622, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n663,
    new_n664, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n708, new_n709, new_n710,
    new_n711, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n869, new_n870,
    new_n871, new_n872, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G146), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G143), .ZN(new_n190));
  INV_X1    g004(.A(G143), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G146), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n190), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G128), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n189), .A2(G143), .ZN(new_n195));
  AOI22_X1  g009(.A1(new_n193), .A2(new_n194), .B1(KEYINPUT1), .B2(new_n195), .ZN(new_n196));
  XNOR2_X1  g010(.A(G143), .B(G146), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT1), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n197), .A2(new_n198), .A3(G128), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n196), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G125), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n193), .A2(new_n194), .ZN(new_n204));
  AOI22_X1  g018(.A1(new_n190), .A2(new_n192), .B1(KEYINPUT0), .B2(G128), .ZN(new_n205));
  OAI21_X1  g019(.A(KEYINPUT0), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(G128), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(new_n208), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n203), .B1(new_n209), .B2(new_n202), .ZN(new_n210));
  INV_X1    g024(.A(G224), .ZN(new_n211));
  OAI21_X1  g025(.A(KEYINPUT7), .B1(new_n211), .B2(G953), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  XOR2_X1   g027(.A(new_n213), .B(KEYINPUT85), .Z(new_n214));
  INV_X1    g028(.A(G101), .ZN(new_n215));
  INV_X1    g029(.A(G107), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G104), .ZN(new_n217));
  INV_X1    g031(.A(G104), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G107), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n215), .B1(new_n217), .B2(new_n219), .ZN(new_n220));
  XNOR2_X1  g034(.A(new_n220), .B(KEYINPUT78), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n216), .A2(G104), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n222), .A2(G101), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n218), .A2(G107), .ZN(new_n224));
  AOI21_X1  g038(.A(KEYINPUT3), .B1(new_n224), .B2(KEYINPUT76), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n216), .A2(KEYINPUT76), .A3(KEYINPUT3), .A4(G104), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n223), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n221), .A2(new_n228), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n229), .A2(KEYINPUT84), .ZN(new_n230));
  XNOR2_X1  g044(.A(G116), .B(G119), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(KEYINPUT5), .ZN(new_n232));
  INV_X1    g046(.A(G116), .ZN(new_n233));
  NOR3_X1   g047(.A1(new_n233), .A2(KEYINPUT5), .A3(G119), .ZN(new_n234));
  INV_X1    g048(.A(G113), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  XOR2_X1   g050(.A(KEYINPUT2), .B(G113), .Z(new_n237));
  AOI22_X1  g051(.A1(new_n232), .A2(new_n236), .B1(new_n237), .B2(new_n231), .ZN(new_n238));
  XOR2_X1   g052(.A(new_n230), .B(new_n238), .Z(new_n239));
  XNOR2_X1  g053(.A(G110), .B(G122), .ZN(new_n240));
  XOR2_X1   g054(.A(new_n240), .B(KEYINPUT8), .Z(new_n241));
  OAI22_X1  g055(.A1(new_n239), .A2(new_n241), .B1(new_n210), .B2(new_n212), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n214), .A2(new_n242), .ZN(new_n243));
  AND3_X1   g057(.A1(new_n221), .A2(new_n228), .A3(new_n238), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT77), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n228), .A2(KEYINPUT4), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n216), .A2(KEYINPUT76), .A3(G104), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT3), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n222), .B1(new_n249), .B2(new_n226), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n250), .A2(new_n215), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n245), .B1(new_n246), .B2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n249), .A2(new_n226), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n253), .B1(new_n254), .B2(new_n223), .ZN(new_n255));
  OAI211_X1 g069(.A(new_n255), .B(KEYINPUT77), .C1(new_n215), .C2(new_n250), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n252), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n251), .A2(new_n253), .ZN(new_n258));
  XNOR2_X1  g072(.A(new_n237), .B(new_n231), .ZN(new_n259));
  AND2_X1   g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n244), .B1(new_n257), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(new_n240), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n243), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(G902), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  OAI21_X1  g080(.A(KEYINPUT81), .B1(new_n261), .B2(new_n240), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT6), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n268), .B1(new_n261), .B2(new_n240), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT81), .ZN(new_n270));
  INV_X1    g084(.A(new_n240), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n258), .A2(new_n259), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n272), .B1(new_n252), .B2(new_n256), .ZN(new_n273));
  OAI211_X1 g087(.A(new_n270), .B(new_n271), .C1(new_n273), .C2(new_n244), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n267), .A2(new_n269), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(KEYINPUT82), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT82), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n267), .A2(new_n269), .A3(new_n277), .A4(new_n274), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n261), .A2(new_n240), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(new_n268), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n211), .A2(G953), .ZN(new_n282));
  XNOR2_X1  g096(.A(new_n210), .B(new_n282), .ZN(new_n283));
  AND4_X1   g097(.A1(KEYINPUT83), .A2(new_n279), .A3(new_n281), .A4(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(new_n281), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n285), .B1(new_n276), .B2(new_n278), .ZN(new_n286));
  AOI21_X1  g100(.A(KEYINPUT83), .B1(new_n286), .B2(new_n283), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n266), .B1(new_n284), .B2(new_n287), .ZN(new_n288));
  OAI21_X1  g102(.A(G210), .B1(G237), .B2(G902), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  OAI211_X1 g105(.A(new_n266), .B(new_n289), .C1(new_n284), .C2(new_n287), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n188), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(G953), .ZN(new_n294));
  AND2_X1   g108(.A1(new_n294), .A2(G952), .ZN(new_n295));
  NAND2_X1  g109(.A1(G234), .A2(G237), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n296), .A2(G902), .A3(G953), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  XNOR2_X1  g114(.A(KEYINPUT21), .B(G898), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n298), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  NOR2_X1   g117(.A1(G475), .A2(G902), .ZN(new_n304));
  XNOR2_X1  g118(.A(G125), .B(G140), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(KEYINPUT73), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT73), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n307), .A2(new_n202), .A3(G140), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT19), .ZN(new_n310));
  OAI21_X1  g124(.A(KEYINPUT86), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT86), .ZN(new_n312));
  NAND4_X1  g126(.A1(new_n306), .A2(new_n312), .A3(KEYINPUT19), .A4(new_n308), .ZN(new_n313));
  OR2_X1    g127(.A1(new_n305), .A2(KEYINPUT74), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n305), .A2(KEYINPUT74), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n314), .A2(new_n315), .A3(new_n310), .ZN(new_n316));
  NAND4_X1  g130(.A1(new_n311), .A2(new_n189), .A3(new_n313), .A4(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT16), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n318), .B1(new_n202), .B2(G140), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n319), .B1(new_n309), .B2(new_n318), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(G146), .ZN(new_n321));
  NOR2_X1   g135(.A1(G237), .A2(G953), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n322), .A2(G143), .A3(G214), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  AOI21_X1  g138(.A(G143), .B1(new_n322), .B2(G214), .ZN(new_n325));
  OAI21_X1  g139(.A(G131), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(new_n325), .ZN(new_n327));
  INV_X1    g141(.A(G131), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n327), .A2(new_n328), .A3(new_n323), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n326), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n317), .A2(new_n321), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n327), .A2(new_n323), .ZN(new_n332));
  NAND2_X1  g146(.A1(KEYINPUT18), .A2(G131), .ZN(new_n333));
  XNOR2_X1  g147(.A(new_n332), .B(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n314), .A2(new_n189), .A3(new_n315), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n335), .B1(new_n189), .B2(new_n309), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n331), .A2(new_n337), .ZN(new_n338));
  XNOR2_X1  g152(.A(G113), .B(G122), .ZN(new_n339));
  XNOR2_X1  g153(.A(KEYINPUT87), .B(G104), .ZN(new_n340));
  XOR2_X1   g154(.A(new_n339), .B(new_n340), .Z(new_n341));
  NAND2_X1  g155(.A1(new_n338), .A2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(new_n341), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT17), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n326), .A2(new_n329), .A3(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT88), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n345), .B(new_n346), .ZN(new_n347));
  OAI211_X1 g161(.A(new_n189), .B(new_n319), .C1(new_n309), .C2(new_n318), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n332), .A2(KEYINPUT17), .A3(G131), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n321), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  OAI211_X1 g164(.A(new_n343), .B(new_n337), .C1(new_n347), .C2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT89), .ZN(new_n352));
  AND3_X1   g166(.A1(new_n342), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n352), .B1(new_n342), .B2(new_n351), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n304), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(KEYINPUT20), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n342), .A2(new_n351), .ZN(new_n357));
  NOR3_X1   g171(.A1(KEYINPUT20), .A2(G475), .A3(G902), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n356), .A2(new_n359), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n337), .B1(new_n347), .B2(new_n350), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(new_n341), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(new_n351), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(new_n264), .ZN(new_n364));
  AND2_X1   g178(.A1(new_n364), .A2(G475), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n360), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g181(.A(KEYINPUT13), .B1(new_n191), .B2(G128), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT91), .ZN(new_n369));
  XNOR2_X1  g183(.A(new_n368), .B(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT92), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n371), .B1(new_n191), .B2(G128), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n194), .A2(KEYINPUT92), .A3(G143), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n191), .A2(KEYINPUT13), .A3(G128), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(KEYINPUT93), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT93), .ZN(new_n377));
  NAND4_X1  g191(.A1(new_n377), .A2(new_n191), .A3(KEYINPUT13), .A4(G128), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n374), .A2(new_n376), .A3(new_n378), .ZN(new_n379));
  OAI21_X1  g193(.A(G134), .B1(new_n370), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n233), .A2(G122), .ZN(new_n381));
  INV_X1    g195(.A(G122), .ZN(new_n382));
  AND3_X1   g196(.A1(new_n382), .A2(KEYINPUT90), .A3(G116), .ZN(new_n383));
  AOI21_X1  g197(.A(KEYINPUT90), .B1(new_n382), .B2(G116), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n381), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  AOI22_X1  g199(.A1(new_n372), .A2(new_n373), .B1(G128), .B2(new_n191), .ZN(new_n386));
  INV_X1    g200(.A(G134), .ZN(new_n387));
  AOI22_X1  g201(.A1(new_n385), .A2(new_n216), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  OAI211_X1 g202(.A(new_n380), .B(new_n388), .C1(new_n216), .C2(new_n385), .ZN(new_n389));
  OAI21_X1  g203(.A(KEYINPUT14), .B1(new_n383), .B2(new_n384), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n385), .A2(new_n390), .A3(G107), .ZN(new_n391));
  OAI221_X1 g205(.A(new_n381), .B1(KEYINPUT14), .B2(new_n216), .C1(new_n383), .C2(new_n384), .ZN(new_n392));
  AND2_X1   g206(.A1(new_n386), .A2(new_n387), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n386), .A2(new_n387), .ZN(new_n394));
  OAI211_X1 g208(.A(new_n391), .B(new_n392), .C1(new_n393), .C2(new_n394), .ZN(new_n395));
  XNOR2_X1  g209(.A(KEYINPUT9), .B(G234), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n397), .A2(G217), .A3(new_n294), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n389), .A2(new_n395), .A3(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n399), .B1(new_n389), .B2(new_n395), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n264), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  OR2_X1    g217(.A1(new_n403), .A2(KEYINPUT94), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(KEYINPUT94), .ZN(new_n405));
  INV_X1    g219(.A(G478), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n406), .A2(KEYINPUT15), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n404), .A2(new_n405), .A3(new_n407), .ZN(new_n408));
  OAI211_X1 g222(.A(new_n403), .B(KEYINPUT94), .C1(KEYINPUT15), .C2(new_n406), .ZN(new_n409));
  AND2_X1   g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n367), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n293), .A2(new_n303), .A3(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(G137), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n413), .B1(KEYINPUT11), .B2(G134), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT11), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n414), .B1(new_n415), .B2(new_n387), .ZN(new_n416));
  XNOR2_X1  g230(.A(KEYINPUT64), .B(G137), .ZN(new_n417));
  AND2_X1   g231(.A1(KEYINPUT11), .A2(G134), .ZN(new_n418));
  AOI21_X1  g232(.A(KEYINPUT65), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n413), .A2(KEYINPUT64), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT64), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(G137), .ZN(new_n422));
  AND4_X1   g236(.A1(KEYINPUT65), .A2(new_n420), .A3(new_n422), .A4(new_n418), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n416), .B1(new_n419), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(G131), .ZN(new_n425));
  OAI211_X1 g239(.A(new_n328), .B(new_n416), .C1(new_n419), .C2(new_n423), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(new_n209), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n417), .A2(new_n387), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n328), .B1(G134), .B2(G137), .ZN(new_n430));
  AOI22_X1  g244(.A1(new_n196), .A2(new_n199), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(new_n426), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n428), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(new_n259), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n208), .B1(new_n425), .B2(new_n426), .ZN(new_n435));
  INV_X1    g249(.A(new_n432), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n259), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n434), .A2(new_n439), .A3(KEYINPUT69), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT69), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n433), .A2(new_n441), .A3(new_n259), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n440), .A2(KEYINPUT28), .A3(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT28), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n438), .B1(new_n437), .B2(KEYINPUT68), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT68), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n433), .A2(new_n446), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n444), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n322), .A2(G210), .ZN(new_n449));
  XOR2_X1   g263(.A(new_n449), .B(KEYINPUT27), .Z(new_n450));
  XNOR2_X1  g264(.A(KEYINPUT26), .B(G101), .ZN(new_n451));
  XOR2_X1   g265(.A(new_n450), .B(new_n451), .Z(new_n452));
  NAND4_X1  g266(.A1(new_n443), .A2(new_n448), .A3(KEYINPUT29), .A4(new_n452), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n453), .B(KEYINPUT70), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT29), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n428), .A2(KEYINPUT30), .A3(new_n432), .ZN(new_n456));
  AND3_X1   g270(.A1(new_n431), .A2(new_n426), .A3(KEYINPUT66), .ZN(new_n457));
  AOI21_X1  g271(.A(KEYINPUT66), .B1(new_n431), .B2(new_n426), .ZN(new_n458));
  NOR3_X1   g272(.A1(new_n435), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  OAI211_X1 g273(.A(new_n456), .B(new_n259), .C1(new_n459), .C2(KEYINPUT30), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(new_n439), .ZN(new_n461));
  INV_X1    g275(.A(new_n452), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n439), .B1(new_n438), .B2(new_n459), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(KEYINPUT28), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(new_n448), .ZN(new_n466));
  OAI211_X1 g280(.A(new_n455), .B(new_n463), .C1(new_n466), .C2(new_n462), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(new_n264), .ZN(new_n468));
  OAI21_X1  g282(.A(G472), .B1(new_n454), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n466), .A2(new_n462), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT31), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n460), .A2(new_n439), .A3(new_n452), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT67), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND4_X1  g288(.A1(new_n460), .A2(KEYINPUT67), .A3(new_n439), .A4(new_n452), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n471), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  AND2_X1   g290(.A1(new_n472), .A2(new_n471), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n470), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT32), .ZN(new_n479));
  NOR2_X1   g293(.A1(G472), .A2(G902), .ZN(new_n480));
  AND3_X1   g294(.A1(new_n478), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n479), .B1(new_n478), .B2(new_n480), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n469), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(G234), .ZN(new_n484));
  OAI21_X1  g298(.A(G217), .B1(new_n484), .B2(G902), .ZN(new_n485));
  XNOR2_X1  g299(.A(new_n485), .B(KEYINPUT71), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT23), .ZN(new_n488));
  INV_X1    g302(.A(G119), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n488), .B1(new_n489), .B2(G128), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n194), .A2(KEYINPUT23), .A3(G119), .ZN(new_n491));
  OAI211_X1 g305(.A(new_n490), .B(new_n491), .C1(G119), .C2(new_n194), .ZN(new_n492));
  XNOR2_X1  g306(.A(KEYINPUT24), .B(G110), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  XNOR2_X1  g308(.A(G119), .B(G128), .ZN(new_n495));
  OAI22_X1  g309(.A1(new_n492), .A2(G110), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n321), .A2(new_n335), .A3(new_n496), .ZN(new_n497));
  AND2_X1   g311(.A1(new_n321), .A2(new_n348), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n492), .A2(G110), .ZN(new_n499));
  XNOR2_X1  g313(.A(new_n499), .B(KEYINPUT72), .ZN(new_n500));
  INV_X1    g314(.A(new_n495), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n500), .B1(new_n501), .B2(new_n493), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n497), .B1(new_n498), .B2(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n294), .A2(G221), .A3(G234), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n504), .B(KEYINPUT75), .ZN(new_n505));
  XNOR2_X1  g319(.A(KEYINPUT22), .B(G137), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n505), .B(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  OR2_X1    g322(.A1(new_n503), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n503), .A2(new_n508), .ZN(new_n510));
  AOI21_X1  g324(.A(G902), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT25), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n487), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n503), .B(new_n507), .ZN(new_n514));
  NOR3_X1   g328(.A1(new_n514), .A2(KEYINPUT25), .A3(G902), .ZN(new_n515));
  OR2_X1    g329(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  OR3_X1    g330(.A1(new_n514), .A2(G902), .A3(new_n487), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  OAI21_X1  g333(.A(G221), .B1(new_n396), .B2(G902), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(G469), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n522), .A2(new_n264), .ZN(new_n523));
  XNOR2_X1  g337(.A(G110), .B(G140), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n294), .A2(G227), .ZN(new_n525));
  XOR2_X1   g339(.A(new_n524), .B(new_n525), .Z(new_n526));
  NAND3_X1  g340(.A1(new_n257), .A2(new_n258), .A3(new_n209), .ZN(new_n527));
  AND2_X1   g341(.A1(new_n221), .A2(new_n228), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT10), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n201), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n199), .A2(KEYINPUT79), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT79), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n197), .A2(new_n532), .A3(new_n198), .A4(G128), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n531), .A2(new_n196), .A3(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n534), .A2(new_n228), .A3(new_n221), .ZN(new_n535));
  AOI22_X1  g349(.A1(new_n528), .A2(new_n530), .B1(new_n535), .B2(new_n529), .ZN(new_n536));
  INV_X1    g350(.A(new_n427), .ZN(new_n537));
  AND3_X1   g351(.A1(new_n527), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n537), .B1(new_n527), .B2(new_n536), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n526), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n200), .B1(new_n221), .B2(new_n228), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n535), .B1(new_n541), .B2(KEYINPUT80), .ZN(new_n542));
  AND3_X1   g356(.A1(new_n229), .A2(KEYINPUT80), .A3(new_n201), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n427), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(KEYINPUT12), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n527), .A2(new_n536), .A3(new_n537), .ZN(new_n546));
  INV_X1    g360(.A(new_n526), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT12), .ZN(new_n548));
  OAI211_X1 g362(.A(new_n548), .B(new_n427), .C1(new_n542), .C2(new_n543), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n545), .A2(new_n546), .A3(new_n547), .A4(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(G902), .B1(new_n540), .B2(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n523), .B1(new_n551), .B2(new_n522), .ZN(new_n552));
  OR3_X1    g366(.A1(new_n538), .A2(new_n539), .A3(new_n526), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n545), .A2(new_n546), .A3(new_n549), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(new_n526), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n553), .A2(new_n555), .A3(G469), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n521), .B1(new_n552), .B2(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n483), .A2(new_n519), .A3(new_n557), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n412), .A2(new_n558), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n559), .B(new_n215), .ZN(G3));
  NAND2_X1  g374(.A1(new_n293), .A2(new_n303), .ZN(new_n561));
  OAI21_X1  g375(.A(KEYINPUT33), .B1(new_n401), .B2(new_n402), .ZN(new_n562));
  INV_X1    g376(.A(new_n402), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT33), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n563), .A2(new_n564), .A3(new_n400), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n562), .A2(new_n565), .A3(G478), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n406), .A2(new_n264), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n569), .B1(new_n403), .B2(G478), .ZN(new_n570));
  OAI21_X1  g384(.A(KEYINPUT95), .B1(new_n567), .B2(new_n570), .ZN(new_n571));
  OR2_X1    g385(.A1(new_n403), .A2(G478), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT95), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n572), .A2(new_n573), .A3(new_n566), .A4(new_n569), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n367), .A2(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(KEYINPUT96), .B1(new_n561), .B2(new_n576), .ZN(new_n577));
  AOI211_X1 g391(.A(new_n188), .B(new_n302), .C1(new_n291), .C2(new_n292), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT96), .ZN(new_n579));
  INV_X1    g393(.A(new_n576), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n478), .A2(new_n480), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(G472), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n584), .B1(new_n478), .B2(new_n264), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n586), .A2(new_n519), .A3(new_n557), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n577), .A2(new_n581), .A3(new_n588), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n589), .B(G104), .ZN(new_n590));
  XNOR2_X1  g404(.A(KEYINPUT97), .B(KEYINPUT34), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n590), .B(new_n591), .ZN(G6));
  NOR2_X1   g406(.A1(new_n353), .A2(new_n354), .ZN(new_n593));
  INV_X1    g407(.A(new_n358), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n356), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(new_n366), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n408), .A2(new_n409), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n293), .A2(new_n303), .A3(new_n598), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n599), .A2(new_n587), .ZN(new_n600));
  XNOR2_X1  g414(.A(KEYINPUT35), .B(G107), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n600), .B(new_n601), .ZN(G9));
  NOR2_X1   g416(.A1(new_n507), .A2(KEYINPUT36), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n503), .B(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n604), .A2(new_n264), .A3(new_n486), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n605), .B1(new_n513), .B2(new_n515), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n557), .A2(new_n606), .ZN(new_n607));
  NOR3_X1   g421(.A1(new_n583), .A2(new_n607), .A3(new_n585), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n293), .A2(new_n303), .A3(new_n411), .A4(new_n608), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n609), .B(KEYINPUT98), .ZN(new_n610));
  XOR2_X1   g424(.A(KEYINPUT37), .B(G110), .Z(new_n611));
  XNOR2_X1  g425(.A(new_n610), .B(new_n611), .ZN(G12));
  NAND2_X1  g426(.A1(new_n582), .A2(KEYINPUT32), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n478), .A2(new_n479), .A3(new_n480), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n607), .B1(new_n615), .B2(new_n469), .ZN(new_n616));
  XOR2_X1   g430(.A(KEYINPUT99), .B(G900), .Z(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(new_n300), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(new_n297), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NOR3_X1   g434(.A1(new_n596), .A2(new_n597), .A3(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n616), .A2(new_n293), .A3(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(G128), .ZN(G30));
  NAND2_X1  g437(.A1(new_n291), .A2(new_n292), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(KEYINPUT38), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n474), .A2(new_n475), .ZN(new_n626));
  AND2_X1   g440(.A1(new_n440), .A2(new_n442), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n626), .B1(new_n462), .B2(new_n627), .ZN(new_n628));
  OAI21_X1  g442(.A(G472), .B1(new_n628), .B2(G902), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n615), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n619), .B(KEYINPUT39), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n557), .A2(new_n631), .ZN(new_n632));
  XOR2_X1   g446(.A(new_n632), .B(KEYINPUT40), .Z(new_n633));
  AOI22_X1  g447(.A1(new_n355), .A2(KEYINPUT20), .B1(new_n357), .B2(new_n358), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n634), .A2(new_n365), .ZN(new_n635));
  NOR4_X1   g449(.A1(new_n635), .A2(new_n606), .A3(new_n188), .A4(new_n597), .ZN(new_n636));
  AND4_X1   g450(.A1(new_n625), .A2(new_n630), .A3(new_n633), .A4(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(new_n191), .ZN(G45));
  OAI211_X1 g452(.A(new_n575), .B(new_n619), .C1(new_n634), .C2(new_n365), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n279), .A2(new_n281), .A3(new_n283), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT83), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n286), .A2(KEYINPUT83), .A3(new_n283), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n289), .B1(new_n645), .B2(new_n266), .ZN(new_n646));
  AOI211_X1 g460(.A(new_n290), .B(new_n265), .C1(new_n643), .C2(new_n644), .ZN(new_n647));
  OAI211_X1 g461(.A(new_n187), .B(new_n640), .C1(new_n646), .C2(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(KEYINPUT100), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT100), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n624), .A2(new_n650), .A3(new_n187), .A4(new_n640), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n649), .A2(new_n616), .A3(new_n651), .ZN(new_n652));
  XOR2_X1   g466(.A(KEYINPUT101), .B(G146), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G48));
  AOI21_X1  g468(.A(new_n518), .B1(new_n615), .B2(new_n469), .ZN(new_n655));
  OR2_X1    g469(.A1(new_n551), .A2(new_n522), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n551), .A2(new_n522), .ZN(new_n657));
  AND2_X1   g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  AND2_X1   g472(.A1(new_n658), .A2(new_n520), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n577), .A2(new_n655), .A3(new_n581), .A4(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(KEYINPUT41), .B(G113), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G15));
  NAND3_X1  g476(.A1(new_n483), .A2(new_n519), .A3(new_n659), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n599), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(new_n233), .ZN(G18));
  INV_X1    g479(.A(new_n606), .ZN(new_n666));
  NOR4_X1   g480(.A1(new_n666), .A2(new_n367), .A3(new_n302), .A4(new_n410), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n293), .A2(new_n483), .A3(new_n659), .A4(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(G119), .ZN(G21));
  AND2_X1   g483(.A1(new_n443), .A2(new_n448), .ZN(new_n670));
  OAI22_X1  g484(.A1(new_n476), .A2(new_n477), .B1(new_n452), .B2(new_n670), .ZN(new_n671));
  AND2_X1   g485(.A1(new_n671), .A2(new_n480), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n656), .A2(new_n303), .A3(new_n520), .A4(new_n657), .ZN(new_n673));
  NOR4_X1   g487(.A1(new_n672), .A2(new_n585), .A3(new_n518), .A4(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n367), .A2(new_n410), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT102), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n674), .A2(new_n293), .A3(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G122), .ZN(G24));
  AND3_X1   g493(.A1(new_n624), .A2(new_n187), .A3(new_n659), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT103), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n639), .B(new_n681), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n672), .A2(new_n585), .ZN(new_n683));
  AND3_X1   g497(.A1(new_n682), .A2(new_n606), .A3(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n680), .A2(new_n684), .ZN(new_n685));
  XOR2_X1   g499(.A(KEYINPUT104), .B(G125), .Z(new_n686));
  XNOR2_X1  g500(.A(new_n685), .B(new_n686), .ZN(G27));
  INV_X1    g501(.A(KEYINPUT105), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n555), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n554), .A2(KEYINPUT105), .A3(new_n526), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n689), .A2(G469), .A3(new_n553), .A4(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n552), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT106), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n691), .A2(new_n552), .A3(KEYINPUT106), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n521), .A2(new_n188), .ZN(new_n697));
  AND4_X1   g511(.A1(new_n291), .A2(new_n292), .A3(new_n696), .A4(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n698), .A2(new_n655), .A3(new_n682), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT42), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n483), .A2(new_n519), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n291), .A2(new_n696), .A3(new_n292), .A4(new_n697), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n704), .A2(KEYINPUT42), .A3(new_n682), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n701), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G131), .ZN(G33));
  INV_X1    g521(.A(KEYINPUT107), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n708), .B1(new_n704), .B2(new_n621), .ZN(new_n709));
  AND4_X1   g523(.A1(new_n708), .A2(new_n698), .A3(new_n655), .A4(new_n621), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(new_n387), .ZN(G36));
  NOR2_X1   g526(.A1(new_n586), .A2(new_n666), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n635), .A2(new_n575), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n714), .A2(KEYINPUT110), .A3(KEYINPUT43), .ZN(new_n715));
  INV_X1    g529(.A(new_n715), .ZN(new_n716));
  AOI21_X1  g530(.A(KEYINPUT43), .B1(new_n714), .B2(KEYINPUT110), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT111), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NOR3_X1   g534(.A1(new_n716), .A2(KEYINPUT111), .A3(new_n717), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n713), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT44), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  OAI211_X1 g538(.A(KEYINPUT44), .B(new_n713), .C1(new_n720), .C2(new_n721), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n624), .A2(new_n188), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n724), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT112), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n724), .A2(new_n725), .A3(KEYINPUT112), .A4(new_n726), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT45), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n556), .B1(new_n731), .B2(new_n522), .ZN(new_n732));
  OR2_X1    g546(.A1(new_n732), .A2(KEYINPUT108), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n689), .A2(KEYINPUT45), .A3(new_n553), .A4(new_n690), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n732), .A2(KEYINPUT108), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n733), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(new_n523), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT46), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n736), .A2(KEYINPUT46), .A3(new_n737), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n740), .A2(new_n657), .A3(new_n741), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n742), .A2(new_n520), .A3(new_n631), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(KEYINPUT109), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n729), .A2(new_n730), .A3(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G137), .ZN(G39));
  INV_X1    g560(.A(KEYINPUT47), .ZN(new_n747));
  INV_X1    g561(.A(new_n742), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n747), .B1(new_n748), .B2(new_n521), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n742), .A2(KEYINPUT47), .A3(new_n520), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(new_n726), .ZN(new_n752));
  NOR4_X1   g566(.A1(new_n752), .A2(new_n483), .A3(new_n519), .A4(new_n639), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G140), .ZN(G42));
  XOR2_X1   g569(.A(new_n658), .B(KEYINPUT49), .Z(new_n756));
  OR4_X1    g570(.A1(new_n188), .A2(new_n756), .A3(new_n521), .A4(new_n714), .ZN(new_n757));
  OR4_X1    g571(.A1(new_n518), .A2(new_n757), .A3(new_n625), .A4(new_n630), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT54), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT53), .ZN(new_n760));
  OAI211_X1 g574(.A(new_n668), .B(new_n678), .C1(new_n412), .C2(new_n558), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n609), .B1(new_n599), .B2(new_n663), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT113), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n293), .A2(new_n764), .A3(new_n303), .A4(new_n580), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n410), .A2(KEYINPUT114), .ZN(new_n766));
  AND3_X1   g580(.A1(new_n408), .A2(KEYINPUT114), .A3(new_n409), .ZN(new_n767));
  OR2_X1    g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n768), .A2(new_n367), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n293), .A2(new_n303), .A3(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n765), .A2(new_n770), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n764), .B1(new_n578), .B2(new_n580), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n588), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n763), .A2(new_n660), .A3(new_n773), .A4(new_n706), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n768), .A2(new_n366), .A3(new_n595), .A4(new_n619), .ZN(new_n775));
  NOR3_X1   g589(.A1(new_n624), .A2(new_n775), .A3(new_n188), .ZN(new_n776));
  AOI22_X1  g590(.A1(new_n776), .A2(new_n616), .B1(new_n684), .B2(new_n698), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n777), .B1(new_n709), .B2(new_n710), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT115), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  OAI211_X1 g594(.A(new_n777), .B(KEYINPUT115), .C1(new_n709), .C2(new_n710), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n774), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  AND2_X1   g596(.A1(new_n619), .A2(KEYINPUT116), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n619), .A2(KEYINPUT116), .ZN(new_n784));
  NOR3_X1   g598(.A1(new_n783), .A2(new_n784), .A3(new_n521), .ZN(new_n785));
  AND3_X1   g599(.A1(new_n696), .A2(new_n666), .A3(new_n785), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n293), .A2(new_n786), .A3(new_n630), .A4(new_n677), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n652), .A2(new_n622), .A3(new_n685), .A4(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT118), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT52), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n791), .A2(KEYINPUT117), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  OAI211_X1 g607(.A(new_n788), .B(new_n789), .C1(KEYINPUT117), .C2(new_n791), .ZN(new_n794));
  OAI21_X1  g608(.A(KEYINPUT117), .B1(new_n788), .B2(new_n791), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n793), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n760), .B1(new_n782), .B2(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(new_n774), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n780), .A2(new_n781), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n685), .A2(new_n622), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n800), .A2(KEYINPUT52), .A3(new_n652), .A4(new_n787), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n788), .A2(new_n791), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  AND4_X1   g617(.A1(new_n760), .A2(new_n798), .A3(new_n799), .A4(new_n803), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n759), .B1(new_n797), .B2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT119), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n798), .A2(new_n799), .A3(new_n803), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(KEYINPUT53), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n782), .A2(new_n760), .A3(new_n796), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n808), .A2(new_n809), .A3(KEYINPUT54), .ZN(new_n810));
  AND3_X1   g624(.A1(new_n805), .A2(new_n806), .A3(new_n810), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n806), .B1(new_n805), .B2(new_n810), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n718), .A2(new_n298), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n291), .A2(new_n292), .A3(new_n658), .A4(new_n697), .ZN(new_n814));
  NOR3_X1   g628(.A1(new_n813), .A2(new_n702), .A3(new_n814), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(KEYINPUT48), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n683), .A2(new_n519), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n813), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(new_n680), .ZN(new_n819));
  OR4_X1    g633(.A1(new_n297), .A2(new_n814), .A3(new_n630), .A4(new_n518), .ZN(new_n820));
  OAI211_X1 g634(.A(new_n819), .B(new_n295), .C1(new_n820), .C2(new_n576), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n816), .A2(new_n821), .ZN(new_n822));
  XOR2_X1   g636(.A(new_n822), .B(KEYINPUT121), .Z(new_n823));
  NOR2_X1   g637(.A1(new_n813), .A2(new_n814), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n824), .A2(new_n606), .A3(new_n683), .ZN(new_n825));
  XOR2_X1   g639(.A(new_n825), .B(KEYINPUT120), .Z(new_n826));
  INV_X1    g640(.A(new_n625), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n827), .A2(new_n818), .A3(new_n188), .A4(new_n659), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT50), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n828), .B(new_n829), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n820), .A2(new_n367), .A3(new_n575), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n658), .A2(new_n521), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n749), .A2(new_n750), .A3(new_n832), .ZN(new_n833));
  NOR3_X1   g647(.A1(new_n752), .A2(new_n813), .A3(new_n817), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n831), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n826), .A2(new_n830), .A3(new_n835), .ZN(new_n836));
  AND2_X1   g650(.A1(new_n836), .A2(KEYINPUT51), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n836), .A2(KEYINPUT51), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n823), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n811), .A2(new_n812), .A3(new_n839), .ZN(new_n840));
  NOR2_X1   g654(.A1(G952), .A2(G953), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n758), .B1(new_n840), .B2(new_n841), .ZN(G75));
  NOR2_X1   g656(.A1(new_n294), .A2(G952), .ZN(new_n843));
  INV_X1    g657(.A(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n782), .A2(new_n796), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n845), .A2(KEYINPUT53), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n782), .A2(new_n760), .A3(new_n803), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n846), .A2(G210), .A3(G902), .A4(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT56), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  XOR2_X1   g664(.A(new_n286), .B(new_n283), .Z(new_n851));
  XOR2_X1   g665(.A(new_n851), .B(KEYINPUT55), .Z(new_n852));
  OAI21_X1  g666(.A(new_n844), .B1(new_n850), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g667(.A(KEYINPUT122), .B1(new_n850), .B2(new_n852), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT122), .ZN(new_n855));
  INV_X1    g669(.A(new_n852), .ZN(new_n856));
  AOI211_X1 g670(.A(new_n855), .B(new_n856), .C1(new_n848), .C2(new_n849), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n853), .A2(new_n854), .A3(new_n857), .ZN(G51));
  XNOR2_X1  g672(.A(new_n523), .B(KEYINPUT57), .ZN(new_n859));
  INV_X1    g673(.A(new_n805), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n797), .A2(new_n804), .A3(new_n759), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n859), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n540), .A2(new_n550), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n797), .A2(new_n804), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n865), .A2(G902), .ZN(new_n866));
  OR2_X1    g680(.A1(new_n866), .A2(new_n736), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n843), .B1(new_n864), .B2(new_n867), .ZN(G54));
  NAND2_X1  g682(.A1(KEYINPUT58), .A2(G475), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n593), .B1(new_n866), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(new_n844), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n866), .A2(new_n593), .A3(new_n869), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n871), .A2(new_n872), .ZN(G60));
  AND2_X1   g687(.A1(new_n562), .A2(new_n565), .ZN(new_n874));
  XNOR2_X1  g688(.A(KEYINPUT123), .B(KEYINPUT59), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n569), .B(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(new_n876), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n878), .B1(new_n860), .B2(new_n861), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(new_n844), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n876), .B1(new_n811), .B2(new_n812), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n880), .B1(new_n881), .B2(new_n874), .ZN(G63));
  NAND2_X1  g696(.A1(G217), .A2(G902), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n883), .B(KEYINPUT60), .ZN(new_n884));
  INV_X1    g698(.A(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n865), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n886), .A2(new_n514), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n865), .A2(new_n604), .A3(new_n885), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n887), .A2(new_n844), .A3(new_n888), .ZN(new_n889));
  XNOR2_X1  g703(.A(KEYINPUT124), .B(KEYINPUT61), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n887), .A2(new_n844), .A3(new_n888), .A4(new_n890), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n892), .A2(new_n893), .ZN(G66));
  OAI21_X1  g708(.A(G953), .B1(new_n301), .B2(new_n211), .ZN(new_n895));
  XOR2_X1   g709(.A(new_n895), .B(KEYINPUT125), .Z(new_n896));
  NAND3_X1  g710(.A1(new_n763), .A2(new_n660), .A3(new_n773), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n896), .B1(new_n897), .B2(new_n294), .ZN(new_n898));
  INV_X1    g712(.A(G898), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n286), .B1(new_n899), .B2(G953), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n898), .B(new_n900), .ZN(G69));
  NAND3_X1  g715(.A1(new_n652), .A2(new_n622), .A3(new_n685), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n637), .A2(new_n902), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(KEYINPUT62), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n769), .A2(new_n580), .ZN(new_n905));
  OR4_X1    g719(.A1(new_n702), .A2(new_n752), .A3(new_n632), .A4(new_n905), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n904), .A2(new_n745), .A3(new_n754), .A4(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(new_n294), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n456), .B1(new_n459), .B2(KEYINPUT30), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n311), .A2(new_n313), .A3(new_n316), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n909), .B(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n908), .A2(new_n912), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n294), .A2(G900), .ZN(new_n914));
  AND3_X1   g728(.A1(new_n655), .A2(new_n293), .A3(new_n677), .ZN(new_n915));
  AOI22_X1  g729(.A1(new_n744), .A2(new_n915), .B1(new_n701), .B2(new_n705), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n711), .A2(new_n902), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n745), .A2(new_n916), .A3(new_n754), .A4(new_n917), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n912), .A2(G953), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n914), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n294), .B1(G227), .B2(G900), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(KEYINPUT126), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n913), .A2(new_n920), .A3(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT127), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n913), .A2(KEYINPUT127), .A3(new_n920), .A4(new_n922), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n913), .A2(new_n920), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(new_n921), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n925), .A2(new_n926), .A3(new_n928), .ZN(G72));
  NAND2_X1  g743(.A1(G472), .A2(G902), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n930), .B(KEYINPUT63), .Z(new_n931));
  OAI21_X1  g745(.A(new_n931), .B1(new_n907), .B2(new_n897), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n932), .A2(new_n452), .A3(new_n461), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n931), .B1(new_n918), .B2(new_n897), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n461), .A2(new_n452), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n843), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n474), .A2(new_n475), .A3(new_n463), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n808), .A2(new_n809), .A3(new_n931), .A4(new_n937), .ZN(new_n938));
  AND3_X1   g752(.A1(new_n933), .A2(new_n936), .A3(new_n938), .ZN(G57));
endmodule


