//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 0 0 1 0 1 0 1 1 1 0 1 0 0 1 1 0 1 0 1 1 0 0 1 1 1 0 1 1 0 1 0 0 0 0 1 0 1 0 0 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:40 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n778, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n804, new_n805, new_n806, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n849, new_n851, new_n853, new_n854, new_n855, new_n856, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n935, new_n936, new_n937, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n946, new_n947, new_n948,
    new_n949, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n982, new_n983, new_n984, new_n985;
  INV_X1    g000(.A(KEYINPUT89), .ZN(new_n202));
  INV_X1    g001(.A(G50gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(G43gat), .ZN(new_n204));
  INV_X1    g003(.A(G43gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G50gat), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n204), .A2(new_n206), .A3(KEYINPUT15), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n204), .A2(new_n206), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT15), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(G29gat), .A2(G36gat), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n211), .B(KEYINPUT88), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT14), .ZN(new_n213));
  INV_X1    g012(.A(G29gat), .ZN(new_n214));
  INV_X1    g013(.A(G36gat), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n213), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  OAI21_X1  g015(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  AND4_X1   g017(.A1(new_n207), .A2(new_n210), .A3(new_n212), .A4(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n216), .A2(KEYINPUT87), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT87), .ZN(new_n221));
  NAND4_X1  g020(.A1(new_n221), .A2(new_n213), .A3(new_n214), .A4(new_n215), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n220), .A2(new_n222), .A3(new_n217), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n207), .B1(new_n223), .B2(new_n212), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n202), .B1(new_n219), .B2(new_n224), .ZN(new_n225));
  NAND4_X1  g024(.A1(new_n210), .A2(new_n212), .A3(new_n207), .A4(new_n218), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT88), .ZN(new_n227));
  XNOR2_X1  g026(.A(new_n211), .B(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(new_n217), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n229), .B1(KEYINPUT87), .B2(new_n216), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n228), .B1(new_n230), .B2(new_n222), .ZN(new_n231));
  OAI211_X1 g030(.A(KEYINPUT89), .B(new_n226), .C1(new_n231), .C2(new_n207), .ZN(new_n232));
  XNOR2_X1  g031(.A(KEYINPUT90), .B(KEYINPUT17), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n225), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  OAI211_X1 g033(.A(KEYINPUT17), .B(new_n226), .C1(new_n231), .C2(new_n207), .ZN(new_n235));
  XNOR2_X1  g034(.A(G15gat), .B(G22gat), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT16), .ZN(new_n237));
  AOI21_X1  g036(.A(G1gat), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT91), .ZN(new_n240));
  INV_X1    g039(.A(G8gat), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n236), .A2(new_n240), .A3(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n241), .B1(new_n236), .B2(new_n240), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n239), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n244), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n246), .A2(new_n238), .A3(new_n242), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n245), .A2(new_n247), .A3(KEYINPUT92), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT92), .ZN(new_n249));
  NOR3_X1   g048(.A1(new_n239), .A2(new_n243), .A3(new_n244), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n238), .B1(new_n246), .B2(new_n242), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n249), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND4_X1  g051(.A1(new_n234), .A2(new_n235), .A3(new_n248), .A4(new_n252), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n250), .A2(new_n251), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n254), .A2(new_n225), .A3(new_n232), .ZN(new_n255));
  NAND2_X1  g054(.A1(G229gat), .A2(G233gat), .ZN(new_n256));
  NAND4_X1  g055(.A1(new_n253), .A2(KEYINPUT18), .A3(new_n255), .A4(new_n256), .ZN(new_n257));
  XOR2_X1   g056(.A(new_n256), .B(KEYINPUT13), .Z(new_n258));
  INV_X1    g057(.A(new_n255), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n254), .B1(new_n225), .B2(new_n232), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n258), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  AND2_X1   g060(.A1(new_n257), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n234), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n252), .A2(new_n235), .A3(new_n248), .ZN(new_n264));
  OAI211_X1 g063(.A(new_n255), .B(new_n256), .C1(new_n263), .C2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT18), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT93), .ZN(new_n268));
  XNOR2_X1  g067(.A(G113gat), .B(G141gat), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n269), .B(G197gat), .ZN(new_n270));
  XOR2_X1   g069(.A(KEYINPUT11), .B(G169gat), .Z(new_n271));
  XNOR2_X1  g070(.A(new_n270), .B(new_n271), .ZN(new_n272));
  XOR2_X1   g071(.A(new_n272), .B(KEYINPUT12), .Z(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  OAI211_X1 g073(.A(new_n262), .B(new_n267), .C1(new_n268), .C2(new_n274), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n257), .A2(new_n268), .A3(new_n261), .ZN(new_n276));
  AND2_X1   g075(.A1(new_n265), .A2(new_n266), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n257), .A2(new_n261), .ZN(new_n278));
  OAI211_X1 g077(.A(new_n276), .B(new_n273), .C1(new_n277), .C2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n275), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  XOR2_X1   g080(.A(G1gat), .B(G29gat), .Z(new_n282));
  XNOR2_X1  g081(.A(new_n282), .B(KEYINPUT80), .ZN(new_n283));
  XOR2_X1   g082(.A(G57gat), .B(G85gat), .Z(new_n284));
  XNOR2_X1  g083(.A(new_n283), .B(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n286));
  XOR2_X1   g085(.A(new_n285), .B(new_n286), .Z(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(G225gat), .A2(G233gat), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(G113gat), .ZN(new_n291));
  INV_X1    g090(.A(G120gat), .ZN(new_n292));
  AOI21_X1  g091(.A(KEYINPUT1), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n293), .B1(new_n291), .B2(new_n292), .ZN(new_n294));
  XNOR2_X1  g093(.A(G127gat), .B(G134gat), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT69), .ZN(new_n298));
  XOR2_X1   g097(.A(KEYINPUT68), .B(KEYINPUT1), .Z(new_n299));
  NAND2_X1  g098(.A1(new_n291), .A2(new_n292), .ZN(new_n300));
  AND3_X1   g099(.A1(new_n299), .A2(new_n295), .A3(new_n300), .ZN(new_n301));
  XNOR2_X1  g100(.A(KEYINPUT67), .B(G120gat), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n302), .A2(new_n291), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n298), .B1(new_n301), .B2(new_n304), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n299), .A2(new_n295), .A3(new_n300), .ZN(new_n306));
  NOR3_X1   g105(.A1(new_n306), .A2(KEYINPUT69), .A3(new_n303), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n297), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  XNOR2_X1  g107(.A(G141gat), .B(G148gat), .ZN(new_n309));
  AOI21_X1  g108(.A(KEYINPUT2), .B1(new_n309), .B2(KEYINPUT77), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n310), .B1(KEYINPUT77), .B2(new_n309), .ZN(new_n311));
  XOR2_X1   g110(.A(G155gat), .B(G162gat), .Z(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  XNOR2_X1  g112(.A(KEYINPUT78), .B(G155gat), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(G162gat), .ZN(new_n316));
  OAI21_X1  g115(.A(KEYINPUT2), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n312), .A2(new_n309), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n313), .A2(new_n319), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n308), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n301), .A2(new_n298), .A3(new_n304), .ZN(new_n322));
  OAI21_X1  g121(.A(KEYINPUT69), .B1(new_n306), .B2(new_n303), .ZN(new_n323));
  AOI22_X1  g122(.A1(new_n322), .A2(new_n323), .B1(new_n296), .B2(new_n294), .ZN(new_n324));
  AOI22_X1  g123(.A1(new_n311), .A2(new_n312), .B1(new_n317), .B2(new_n318), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n290), .B1(new_n321), .B2(new_n326), .ZN(new_n327));
  OAI21_X1  g126(.A(KEYINPUT4), .B1(new_n308), .B2(new_n320), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT4), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n324), .A2(new_n329), .A3(new_n325), .ZN(new_n330));
  AND2_X1   g129(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n320), .A2(KEYINPUT3), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT3), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n325), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n332), .A2(new_n308), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(new_n289), .ZN(new_n336));
  OAI211_X1 g135(.A(KEYINPUT5), .B(new_n327), .C1(new_n331), .C2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT81), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n328), .A2(new_n338), .A3(new_n330), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n321), .A2(KEYINPUT81), .A3(new_n329), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n290), .A2(KEYINPUT5), .ZN(new_n341));
  NAND4_X1  g140(.A1(new_n339), .A2(new_n340), .A3(new_n335), .A4(new_n341), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n288), .B1(new_n337), .B2(new_n342), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n339), .A2(new_n335), .A3(new_n340), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(new_n290), .ZN(new_n345));
  OR2_X1    g144(.A1(new_n345), .A2(KEYINPUT39), .ZN(new_n346));
  OR2_X1    g145(.A1(new_n321), .A2(new_n326), .ZN(new_n347));
  OAI211_X1 g146(.A(new_n345), .B(KEYINPUT39), .C1(new_n290), .C2(new_n347), .ZN(new_n348));
  AND3_X1   g147(.A1(new_n346), .A2(new_n348), .A3(new_n288), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n343), .B1(new_n349), .B2(KEYINPUT40), .ZN(new_n350));
  NAND2_X1  g149(.A1(G169gat), .A2(G176gat), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT26), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(G169gat), .ZN(new_n354));
  INV_X1    g153(.A(G176gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT66), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n353), .A2(KEYINPUT66), .A3(new_n356), .ZN(new_n360));
  OAI211_X1 g159(.A(new_n359), .B(new_n360), .C1(KEYINPUT26), .C2(new_n356), .ZN(new_n361));
  XNOR2_X1  g160(.A(KEYINPUT27), .B(G183gat), .ZN(new_n362));
  INV_X1    g161(.A(G190gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT28), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(KEYINPUT65), .ZN(new_n366));
  OR2_X1    g165(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  AOI22_X1  g166(.A1(new_n364), .A2(new_n366), .B1(G183gat), .B2(G190gat), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n361), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT23), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n356), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n354), .A2(new_n355), .A3(KEYINPUT23), .ZN(new_n372));
  AND3_X1   g171(.A1(new_n371), .A2(new_n351), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(G183gat), .A2(G190gat), .ZN(new_n374));
  OAI211_X1 g173(.A(new_n373), .B(new_n374), .C1(KEYINPUT64), .C2(KEYINPUT25), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n371), .A2(new_n351), .A3(new_n372), .ZN(new_n376));
  OAI21_X1  g175(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n371), .A2(KEYINPUT64), .A3(new_n351), .A4(new_n372), .ZN(new_n379));
  NAND4_X1  g178(.A1(new_n371), .A2(new_n351), .A3(new_n374), .A4(new_n372), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT25), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n379), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  AND3_X1   g181(.A1(new_n375), .A2(new_n378), .A3(new_n382), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n378), .B1(new_n375), .B2(new_n382), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n369), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT29), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(G226gat), .A2(G233gat), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  XOR2_X1   g188(.A(KEYINPUT74), .B(G197gat), .Z(new_n390));
  INV_X1    g189(.A(G204gat), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  XNOR2_X1  g191(.A(KEYINPUT74), .B(G197gat), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(G204gat), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(G211gat), .A2(G218gat), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT22), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n395), .A2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT75), .ZN(new_n400));
  INV_X1    g199(.A(new_n396), .ZN(new_n401));
  NOR2_X1   g200(.A1(G211gat), .A2(G218gat), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n399), .A2(new_n400), .A3(new_n404), .ZN(new_n405));
  AOI22_X1  g204(.A1(new_n392), .A2(new_n394), .B1(new_n397), .B2(new_n396), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n403), .B1(new_n406), .B2(KEYINPUT75), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n385), .A2(G226gat), .A3(G233gat), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n389), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT76), .ZN(new_n412));
  NAND4_X1  g211(.A1(new_n385), .A2(new_n412), .A3(G226gat), .A4(G233gat), .ZN(new_n413));
  AND3_X1   g212(.A1(new_n361), .A2(new_n367), .A3(new_n368), .ZN(new_n414));
  AND3_X1   g213(.A1(new_n379), .A2(new_n380), .A3(new_n381), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n380), .B1(new_n381), .B2(new_n379), .ZN(new_n416));
  OAI22_X1  g215(.A1(new_n415), .A2(new_n416), .B1(new_n376), .B2(new_n377), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n375), .A2(new_n378), .A3(new_n382), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n414), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  OAI21_X1  g218(.A(KEYINPUT76), .B1(new_n419), .B2(new_n388), .ZN(new_n420));
  AOI22_X1  g219(.A1(new_n413), .A2(new_n420), .B1(new_n387), .B2(new_n388), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n411), .B1(new_n421), .B2(new_n409), .ZN(new_n422));
  XNOR2_X1  g221(.A(G8gat), .B(G36gat), .ZN(new_n423));
  XNOR2_X1  g222(.A(G64gat), .B(G92gat), .ZN(new_n424));
  XOR2_X1   g223(.A(new_n423), .B(new_n424), .Z(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n422), .A2(new_n426), .ZN(new_n427));
  OAI211_X1 g226(.A(new_n411), .B(new_n425), .C1(new_n421), .C2(new_n409), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n427), .A2(KEYINPUT30), .A3(new_n428), .ZN(new_n429));
  OR3_X1    g228(.A1(new_n422), .A2(KEYINPUT30), .A3(new_n426), .ZN(new_n430));
  AND2_X1   g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  OAI211_X1 g230(.A(new_n350), .B(new_n431), .C1(KEYINPUT40), .C2(new_n349), .ZN(new_n432));
  NAND2_X1  g231(.A1(G228gat), .A2(G233gat), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n333), .B1(new_n408), .B2(KEYINPUT29), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n433), .B1(new_n434), .B2(new_n320), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT83), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n334), .A2(new_n386), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n436), .B1(new_n437), .B2(new_n408), .ZN(new_n438));
  AOI21_X1  g237(.A(KEYINPUT29), .B1(new_n325), .B2(new_n333), .ZN(new_n439));
  NOR3_X1   g238(.A1(new_n409), .A2(new_n439), .A3(KEYINPUT83), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n435), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  XOR2_X1   g240(.A(new_n433), .B(KEYINPUT82), .Z(new_n442));
  AOI21_X1  g241(.A(KEYINPUT29), .B1(new_n399), .B2(new_n404), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n443), .B1(new_n404), .B2(new_n399), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n325), .B1(new_n444), .B2(new_n333), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n409), .A2(new_n439), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n442), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n441), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(G22gat), .ZN(new_n449));
  INV_X1    g248(.A(G22gat), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n441), .A2(new_n450), .A3(new_n447), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  XNOR2_X1  g251(.A(G78gat), .B(G106gat), .ZN(new_n453));
  XNOR2_X1  g252(.A(KEYINPUT31), .B(G50gat), .ZN(new_n454));
  XNOR2_X1  g253(.A(new_n453), .B(new_n454), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n450), .B1(new_n441), .B2(new_n447), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n455), .B1(new_n456), .B2(KEYINPUT84), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n452), .A2(new_n457), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n449), .A2(KEYINPUT84), .A3(new_n451), .A4(new_n455), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n426), .B1(new_n422), .B2(KEYINPUT37), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT38), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n421), .A2(new_n408), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n389), .A2(new_n408), .A3(new_n410), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(KEYINPUT37), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n462), .B1(new_n463), .B2(new_n465), .ZN(new_n466));
  OR3_X1    g265(.A1(new_n461), .A2(new_n466), .A3(KEYINPUT85), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n337), .A2(new_n342), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(new_n287), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT6), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n337), .A2(new_n288), .A3(new_n342), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n469), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n343), .A2(KEYINPUT6), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(KEYINPUT86), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT86), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n473), .A2(new_n476), .ZN(new_n477));
  OAI21_X1  g276(.A(KEYINPUT85), .B1(new_n461), .B2(new_n466), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n467), .A2(new_n475), .A3(new_n477), .A4(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n461), .B1(KEYINPUT37), .B2(new_n422), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n428), .B1(new_n480), .B2(new_n462), .ZN(new_n481));
  OAI211_X1 g280(.A(new_n432), .B(new_n460), .C1(new_n479), .C2(new_n481), .ZN(new_n482));
  AOI22_X1  g281(.A1(new_n429), .A2(new_n430), .B1(new_n472), .B2(new_n473), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n483), .A2(new_n460), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT36), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT32), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n385), .A2(new_n324), .ZN(new_n487));
  OAI211_X1 g286(.A(new_n308), .B(new_n369), .C1(new_n383), .C2(new_n384), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(G227gat), .ZN(new_n491));
  INV_X1    g290(.A(G233gat), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n486), .B1(new_n490), .B2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT34), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT72), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n493), .B1(new_n489), .B2(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n487), .A2(KEYINPUT72), .A3(new_n488), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n495), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n493), .A2(KEYINPUT34), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n419), .A2(new_n308), .ZN(new_n501));
  INV_X1    g300(.A(new_n488), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(KEYINPUT73), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT73), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n489), .A2(new_n505), .A3(new_n500), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n494), .B1(new_n499), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n490), .A2(new_n493), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT33), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  XOR2_X1   g310(.A(G15gat), .B(G43gat), .Z(new_n512));
  XNOR2_X1  g311(.A(KEYINPUT70), .B(KEYINPUT71), .ZN(new_n513));
  XNOR2_X1  g312(.A(new_n512), .B(new_n513), .ZN(new_n514));
  XNOR2_X1  g313(.A(G71gat), .B(G99gat), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n514), .B(new_n515), .ZN(new_n516));
  AND2_X1   g315(.A1(new_n511), .A2(new_n516), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n496), .B1(new_n501), .B2(new_n502), .ZN(new_n518));
  INV_X1    g317(.A(new_n493), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n518), .A2(new_n519), .A3(new_n498), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(KEYINPUT34), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n509), .A2(KEYINPUT32), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n505), .B1(new_n489), .B2(new_n500), .ZN(new_n523));
  INV_X1    g322(.A(new_n500), .ZN(new_n524));
  AOI211_X1 g323(.A(KEYINPUT73), .B(new_n524), .C1(new_n487), .C2(new_n488), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n521), .A2(new_n522), .A3(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n508), .A2(new_n517), .A3(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(new_n528), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n517), .B1(new_n508), .B2(new_n527), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n485), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n508), .A2(new_n527), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n511), .A2(new_n516), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n534), .A2(KEYINPUT36), .A3(new_n528), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n484), .B1(new_n531), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n482), .A2(new_n536), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n529), .A2(new_n530), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n475), .A2(new_n477), .ZN(new_n539));
  AOI21_X1  g338(.A(KEYINPUT35), .B1(new_n429), .B2(new_n430), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n538), .A2(new_n539), .A3(new_n460), .A4(new_n540), .ZN(new_n541));
  NAND4_X1  g340(.A1(new_n483), .A2(new_n534), .A3(new_n460), .A4(new_n528), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(KEYINPUT35), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n281), .B1(new_n537), .B2(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(G57gat), .B(G64gat), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  OR2_X1    g346(.A1(G71gat), .A2(G78gat), .ZN(new_n548));
  NAND2_X1  g347(.A1(G71gat), .A2(G78gat), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT9), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n547), .A2(new_n550), .A3(new_n552), .ZN(new_n553));
  OAI211_X1 g352(.A(new_n549), .B(new_n548), .C1(new_n546), .C2(new_n551), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n254), .B1(KEYINPUT21), .B2(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n557), .B(KEYINPUT94), .ZN(new_n558));
  XNOR2_X1  g357(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n559));
  XOR2_X1   g358(.A(new_n559), .B(G155gat), .Z(new_n560));
  XNOR2_X1  g359(.A(new_n558), .B(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT21), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n555), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(G231gat), .A2(G233gat), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n563), .B(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(G127gat), .ZN(new_n566));
  XOR2_X1   g365(.A(G183gat), .B(G211gat), .Z(new_n567));
  XNOR2_X1  g366(.A(new_n566), .B(new_n567), .ZN(new_n568));
  XOR2_X1   g367(.A(new_n561), .B(new_n568), .Z(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  AND2_X1   g369(.A1(G232gat), .A2(G233gat), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n571), .A2(KEYINPUT41), .ZN(new_n572));
  XNOR2_X1  g371(.A(G134gat), .B(G162gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n572), .B(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n225), .A2(new_n232), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT96), .ZN(new_n578));
  AND2_X1   g377(.A1(G99gat), .A2(G106gat), .ZN(new_n579));
  NOR2_X1   g378(.A1(G99gat), .A2(G106gat), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  AND2_X1   g381(.A1(G85gat), .A2(G92gat), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT95), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n585), .A2(KEYINPUT7), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT7), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n587), .A2(KEYINPUT95), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n584), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n587), .A2(KEYINPUT95), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n585), .A2(KEYINPUT7), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n590), .A2(new_n591), .A3(new_n583), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(G99gat), .A2(G106gat), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n594), .A2(KEYINPUT8), .ZN(new_n595));
  OR2_X1    g394(.A1(G85gat), .A2(G92gat), .ZN(new_n596));
  AND2_X1   g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n582), .B1(new_n593), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n595), .A2(new_n596), .ZN(new_n599));
  AOI211_X1 g398(.A(new_n581), .B(new_n599), .C1(new_n589), .C2(new_n592), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n578), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  AND3_X1   g400(.A1(new_n590), .A2(new_n591), .A3(new_n583), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n583), .B1(new_n590), .B2(new_n591), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n597), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n604), .A2(new_n581), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n593), .A2(new_n582), .A3(new_n597), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n605), .A2(new_n606), .A3(KEYINPUT96), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n601), .A2(new_n607), .ZN(new_n608));
  AOI22_X1  g407(.A1(new_n577), .A2(new_n608), .B1(KEYINPUT41), .B2(new_n571), .ZN(new_n609));
  XOR2_X1   g408(.A(G190gat), .B(G218gat), .Z(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  NAND4_X1  g410(.A1(new_n234), .A2(new_n235), .A3(new_n607), .A4(new_n601), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n609), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n611), .B1(new_n609), .B2(new_n612), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n575), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n615), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n617), .A2(new_n574), .A3(new_n613), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n570), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n556), .B1(new_n598), .B2(new_n600), .ZN(new_n621));
  NAND2_X1  g420(.A1(G230gat), .A2(G233gat), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n605), .A2(new_n606), .A3(new_n555), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n621), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(G120gat), .B(G148gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(G176gat), .B(G204gat), .ZN(new_n627));
  XOR2_X1   g426(.A(new_n626), .B(new_n627), .Z(new_n628));
  INV_X1    g427(.A(KEYINPUT10), .ZN(new_n629));
  AND3_X1   g428(.A1(new_n605), .A2(new_n555), .A3(new_n606), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n555), .B1(new_n605), .B2(new_n606), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n629), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n555), .A2(new_n629), .ZN(new_n633));
  AND3_X1   g432(.A1(new_n605), .A2(KEYINPUT96), .A3(new_n606), .ZN(new_n634));
  AOI21_X1  g433(.A(KEYINPUT96), .B1(new_n605), .B2(new_n606), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n633), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n632), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT97), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n623), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n632), .A2(new_n636), .A3(KEYINPUT97), .ZN(new_n640));
  AOI21_X1  g439(.A(KEYINPUT98), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  AOI21_X1  g440(.A(KEYINPUT10), .B1(new_n621), .B2(new_n624), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n556), .A2(KEYINPUT10), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n643), .B1(new_n601), .B2(new_n607), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n638), .B1(new_n642), .B2(new_n644), .ZN(new_n645));
  NAND4_X1  g444(.A1(new_n645), .A2(new_n640), .A3(KEYINPUT98), .A4(new_n622), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  OAI211_X1 g446(.A(new_n625), .B(new_n628), .C1(new_n641), .C2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT100), .ZN(new_n649));
  XOR2_X1   g448(.A(new_n622), .B(KEYINPUT99), .Z(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n637), .A2(new_n651), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n628), .B1(new_n652), .B2(new_n625), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n648), .A2(new_n649), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n625), .A2(new_n628), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n645), .A2(new_n640), .A3(new_n622), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT98), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n656), .B1(new_n659), .B2(new_n646), .ZN(new_n660));
  OAI21_X1  g459(.A(KEYINPUT100), .B1(new_n660), .B2(new_n653), .ZN(new_n661));
  AND2_X1   g460(.A1(new_n655), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n620), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n545), .A2(new_n663), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n664), .A2(new_n474), .ZN(new_n665));
  XOR2_X1   g464(.A(new_n665), .B(G1gat), .Z(G1324gat));
  INV_X1    g465(.A(new_n431), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g467(.A(KEYINPUT16), .B(G8gat), .Z(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n670), .B1(new_n241), .B2(new_n668), .ZN(new_n671));
  MUX2_X1   g470(.A(new_n670), .B(new_n671), .S(KEYINPUT42), .Z(G1325gat));
  INV_X1    g471(.A(KEYINPUT101), .ZN(new_n673));
  NOR3_X1   g472(.A1(new_n529), .A2(new_n530), .A3(new_n485), .ZN(new_n674));
  AOI21_X1  g473(.A(KEYINPUT36), .B1(new_n534), .B2(new_n528), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n673), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n531), .A2(KEYINPUT101), .A3(new_n535), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  OAI21_X1  g477(.A(G15gat), .B1(new_n664), .B2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n538), .ZN(new_n680));
  OR2_X1    g479(.A1(new_n680), .A2(G15gat), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n679), .B1(new_n664), .B2(new_n681), .ZN(G1326gat));
  INV_X1    g481(.A(new_n460), .ZN(new_n683));
  AND2_X1   g482(.A1(new_n545), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(new_n663), .ZN(new_n685));
  XNOR2_X1  g484(.A(KEYINPUT43), .B(G22gat), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n685), .B(new_n686), .ZN(G1327gat));
  INV_X1    g486(.A(new_n662), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n688), .A2(new_n569), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n689), .A2(new_n619), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n474), .A2(G29gat), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n545), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(KEYINPUT45), .ZN(new_n693));
  AND3_X1   g492(.A1(new_n541), .A2(new_n543), .A3(KEYINPUT102), .ZN(new_n694));
  AOI21_X1  g493(.A(KEYINPUT102), .B1(new_n541), .B2(new_n543), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n537), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n619), .ZN(new_n697));
  AOI21_X1  g496(.A(KEYINPUT44), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT44), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n619), .A2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n701), .B1(new_n537), .B2(new_n544), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n689), .A2(new_n281), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  NOR4_X1   g503(.A1(new_n698), .A2(new_n474), .A3(new_n702), .A4(new_n704), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n693), .B1(new_n705), .B2(new_n214), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT103), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n706), .B(new_n707), .ZN(G1328gat));
  AND2_X1   g507(.A1(new_n545), .A2(new_n690), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n709), .A2(new_n215), .A3(new_n431), .ZN(new_n710));
  AND2_X1   g509(.A1(KEYINPUT104), .A2(KEYINPUT46), .ZN(new_n711));
  NOR2_X1   g510(.A1(KEYINPUT104), .A2(KEYINPUT46), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n710), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT102), .ZN(new_n714));
  AND2_X1   g513(.A1(new_n542), .A2(KEYINPUT35), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n476), .B1(new_n472), .B2(new_n473), .ZN(new_n716));
  INV_X1    g515(.A(new_n477), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n540), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n534), .A2(new_n460), .A3(new_n528), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n714), .B1(new_n715), .B2(new_n720), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n541), .A2(new_n543), .A3(KEYINPUT102), .ZN(new_n722));
  AOI22_X1  g521(.A1(new_n721), .A2(new_n722), .B1(new_n482), .B2(new_n536), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n699), .B1(new_n723), .B2(new_n619), .ZN(new_n724));
  INV_X1    g523(.A(new_n702), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NOR3_X1   g525(.A1(new_n726), .A2(new_n667), .A3(new_n704), .ZN(new_n727));
  OAI221_X1 g526(.A(new_n713), .B1(new_n711), .B2(new_n710), .C1(new_n727), .C2(new_n215), .ZN(G1329gat));
  NOR2_X1   g527(.A1(new_n680), .A2(G43gat), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n545), .A2(new_n690), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(KEYINPUT47), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n674), .A2(new_n675), .ZN(new_n732));
  NAND4_X1  g531(.A1(new_n724), .A2(new_n732), .A3(new_n725), .A4(new_n703), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n731), .B1(new_n733), .B2(G43gat), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT106), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  AOI211_X1 g535(.A(KEYINPUT106), .B(new_n731), .C1(new_n733), .C2(G43gat), .ZN(new_n737));
  INV_X1    g536(.A(new_n678), .ZN(new_n738));
  NAND4_X1  g537(.A1(new_n724), .A2(new_n738), .A3(new_n725), .A4(new_n703), .ZN(new_n739));
  AOI22_X1  g538(.A1(new_n739), .A2(G43gat), .B1(new_n709), .B2(new_n729), .ZN(new_n740));
  XOR2_X1   g539(.A(KEYINPUT105), .B(KEYINPUT47), .Z(new_n741));
  OAI22_X1  g540(.A1(new_n736), .A2(new_n737), .B1(new_n740), .B2(new_n741), .ZN(G1330gat));
  NOR3_X1   g541(.A1(new_n689), .A2(G50gat), .A3(new_n619), .ZN(new_n743));
  AND2_X1   g542(.A1(new_n684), .A2(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(new_n744), .ZN(new_n745));
  NOR4_X1   g544(.A1(new_n698), .A2(new_n460), .A3(new_n702), .A4(new_n704), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n745), .B1(new_n746), .B2(new_n203), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT107), .ZN(new_n748));
  AOI21_X1  g547(.A(KEYINPUT48), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n724), .A2(new_n683), .A3(new_n725), .A4(new_n703), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n744), .B1(new_n750), .B2(G50gat), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT48), .ZN(new_n752));
  NOR3_X1   g551(.A1(new_n751), .A2(KEYINPUT107), .A3(new_n752), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n749), .A2(new_n753), .ZN(G1331gat));
  NOR3_X1   g553(.A1(new_n620), .A2(new_n280), .A3(new_n688), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n696), .A2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT108), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n696), .A2(KEYINPUT108), .A3(new_n755), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n760), .A2(new_n474), .ZN(new_n761));
  XOR2_X1   g560(.A(KEYINPUT109), .B(G57gat), .Z(new_n762));
  XNOR2_X1  g561(.A(new_n761), .B(new_n762), .ZN(G1332gat));
  AOI21_X1  g562(.A(new_n667), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n758), .A2(new_n759), .A3(new_n764), .ZN(new_n765));
  NOR2_X1   g564(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(KEYINPUT110), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(KEYINPUT111), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n765), .B(new_n768), .ZN(G1333gat));
  OAI21_X1  g568(.A(G71gat), .B1(new_n760), .B2(new_n678), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n680), .A2(G71gat), .ZN(new_n771));
  INV_X1    g570(.A(new_n771), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n770), .B1(new_n760), .B2(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT50), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  OAI211_X1 g574(.A(new_n770), .B(KEYINPUT50), .C1(new_n760), .C2(new_n772), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(G1334gat));
  NOR2_X1   g576(.A1(new_n760), .A2(new_n460), .ZN(new_n778));
  XOR2_X1   g577(.A(new_n778), .B(G78gat), .Z(G1335gat));
  NAND2_X1  g578(.A1(new_n569), .A2(new_n281), .ZN(new_n780));
  XOR2_X1   g579(.A(new_n780), .B(KEYINPUT112), .Z(new_n781));
  NAND3_X1  g580(.A1(new_n696), .A2(new_n697), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(KEYINPUT51), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT51), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n696), .A2(new_n784), .A3(new_n697), .A4(new_n781), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n783), .A2(new_n662), .A3(new_n785), .ZN(new_n786));
  OR2_X1    g585(.A1(new_n786), .A2(new_n474), .ZN(new_n787));
  INV_X1    g586(.A(G85gat), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n781), .A2(new_n662), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n726), .A2(new_n789), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n474), .A2(new_n788), .ZN(new_n791));
  AOI22_X1  g590(.A1(new_n787), .A2(new_n788), .B1(new_n790), .B2(new_n791), .ZN(G1336gat));
  OR2_X1    g591(.A1(KEYINPUT113), .A2(KEYINPUT52), .ZN(new_n793));
  INV_X1    g592(.A(new_n789), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n724), .A2(new_n431), .A3(new_n725), .A4(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(G92gat), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n667), .A2(G92gat), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n783), .A2(new_n662), .A3(new_n785), .A4(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(KEYINPUT113), .A2(KEYINPUT52), .ZN(new_n799));
  AND4_X1   g598(.A1(new_n793), .A2(new_n796), .A3(new_n798), .A4(new_n799), .ZN(new_n800));
  AOI22_X1  g599(.A1(new_n795), .A2(G92gat), .B1(KEYINPUT113), .B2(KEYINPUT52), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n793), .B1(new_n801), .B2(new_n798), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n800), .A2(new_n802), .ZN(G1337gat));
  OR2_X1    g602(.A1(new_n786), .A2(new_n680), .ZN(new_n804));
  INV_X1    g603(.A(G99gat), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n678), .A2(new_n805), .ZN(new_n806));
  AOI22_X1  g605(.A1(new_n804), .A2(new_n805), .B1(new_n790), .B2(new_n806), .ZN(G1338gat));
  INV_X1    g606(.A(KEYINPUT53), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n460), .A2(G106gat), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n783), .A2(new_n662), .A3(new_n785), .A4(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT114), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n808), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NOR4_X1   g611(.A1(new_n698), .A2(new_n460), .A3(new_n702), .A4(new_n789), .ZN(new_n813));
  INV_X1    g612(.A(G106gat), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n810), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n812), .A2(new_n815), .ZN(new_n816));
  OAI221_X1 g615(.A(new_n810), .B1(new_n811), .B2(new_n808), .C1(new_n813), .C2(new_n814), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(G1339gat));
  OAI21_X1  g617(.A(KEYINPUT54), .B1(new_n637), .B2(new_n651), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n820), .B1(new_n641), .B2(new_n647), .ZN(new_n821));
  INV_X1    g620(.A(new_n628), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n822), .B1(new_n652), .B2(KEYINPUT54), .ZN(new_n823));
  INV_X1    g622(.A(new_n823), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n821), .A2(KEYINPUT55), .A3(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT55), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n819), .B1(new_n659), .B2(new_n646), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n826), .B1(new_n827), .B2(new_n823), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n825), .A2(new_n828), .A3(new_n280), .A4(new_n648), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n267), .A2(new_n261), .A3(new_n257), .A4(new_n274), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n256), .B1(new_n253), .B2(new_n255), .ZN(new_n831));
  NOR3_X1   g630(.A1(new_n259), .A2(new_n260), .A3(new_n258), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n272), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n830), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n655), .A2(new_n661), .A3(new_n834), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n697), .B1(new_n829), .B2(new_n835), .ZN(new_n836));
  AND4_X1   g635(.A1(new_n618), .A2(new_n616), .A3(new_n833), .A4(new_n830), .ZN(new_n837));
  AND4_X1   g636(.A1(new_n648), .A2(new_n837), .A3(new_n825), .A4(new_n828), .ZN(new_n838));
  NOR3_X1   g637(.A1(new_n836), .A2(new_n838), .A3(KEYINPUT115), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  OAI21_X1  g639(.A(KEYINPUT115), .B1(new_n836), .B2(new_n838), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n840), .A2(new_n569), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n663), .A2(new_n281), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n719), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n431), .A2(new_n474), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n846), .A2(new_n281), .ZN(new_n847));
  XNOR2_X1  g646(.A(new_n847), .B(new_n291), .ZN(G1340gat));
  NOR2_X1   g647(.A1(new_n846), .A2(new_n688), .ZN(new_n849));
  MUX2_X1   g648(.A(G120gat), .B(new_n302), .S(new_n849), .Z(G1341gat));
  NOR2_X1   g649(.A1(new_n846), .A2(new_n569), .ZN(new_n851));
  XOR2_X1   g650(.A(new_n851), .B(G127gat), .Z(G1342gat));
  NOR2_X1   g651(.A1(new_n474), .A2(G134gat), .ZN(new_n853));
  NAND4_X1  g652(.A1(new_n844), .A2(new_n667), .A3(new_n697), .A4(new_n853), .ZN(new_n854));
  XOR2_X1   g653(.A(new_n854), .B(KEYINPUT56), .Z(new_n855));
  OAI21_X1  g654(.A(G134gat), .B1(new_n846), .B2(new_n619), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(G1343gat));
  INV_X1    g656(.A(G141gat), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n845), .B1(new_n674), .B2(new_n675), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT117), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n821), .A2(KEYINPUT116), .A3(new_n824), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT116), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n862), .B1(new_n827), .B2(new_n823), .ZN(new_n863));
  AND3_X1   g662(.A1(new_n861), .A2(new_n863), .A3(new_n826), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n825), .A2(new_n280), .A3(new_n648), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n835), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n838), .B1(new_n866), .B2(new_n619), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n860), .B1(new_n867), .B2(new_n570), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n861), .A2(new_n863), .A3(new_n826), .ZN(new_n869));
  NAND4_X1  g668(.A1(new_n869), .A2(new_n280), .A3(new_n648), .A4(new_n825), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n697), .B1(new_n870), .B2(new_n835), .ZN(new_n871));
  OAI211_X1 g670(.A(KEYINPUT117), .B(new_n569), .C1(new_n871), .C2(new_n838), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n868), .A2(new_n843), .A3(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT57), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n460), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n841), .A2(new_n569), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n843), .B1(new_n877), .B2(new_n839), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(new_n683), .ZN(new_n879));
  AOI22_X1  g678(.A1(new_n876), .A2(KEYINPUT118), .B1(new_n879), .B2(new_n874), .ZN(new_n880));
  INV_X1    g679(.A(new_n875), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n569), .B1(new_n871), .B2(new_n838), .ZN(new_n882));
  AOI22_X1  g681(.A1(new_n882), .A2(new_n860), .B1(new_n281), .B2(new_n663), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n881), .B1(new_n883), .B2(new_n872), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT118), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n859), .B1(new_n880), .B2(new_n886), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n858), .B1(new_n887), .B2(new_n280), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n678), .A2(new_n683), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT119), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n460), .B1(new_n676), .B2(new_n677), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n474), .B1(new_n892), .B2(KEYINPUT119), .ZN(new_n893));
  NAND4_X1  g692(.A1(new_n891), .A2(new_n893), .A3(new_n667), .A4(new_n878), .ZN(new_n894));
  NOR3_X1   g693(.A1(new_n894), .A2(G141gat), .A3(new_n281), .ZN(new_n895));
  OAI21_X1  g694(.A(KEYINPUT58), .B1(new_n888), .B2(new_n895), .ZN(new_n896));
  INV_X1    g695(.A(new_n859), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n879), .A2(new_n874), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n898), .B1(new_n884), .B2(new_n885), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n876), .A2(KEYINPUT118), .ZN(new_n900));
  OAI211_X1 g699(.A(new_n280), .B(new_n897), .C1(new_n899), .C2(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(G141gat), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT58), .ZN(new_n903));
  INV_X1    g702(.A(new_n895), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n896), .A2(new_n905), .ZN(G1344gat));
  NOR3_X1   g705(.A1(new_n894), .A2(G148gat), .A3(new_n688), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT120), .ZN(new_n908));
  XNOR2_X1  g707(.A(new_n907), .B(new_n908), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT59), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(G148gat), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n911), .B1(new_n887), .B2(new_n662), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n882), .A2(new_n843), .ZN(new_n913));
  AOI21_X1  g712(.A(KEYINPUT57), .B1(new_n913), .B2(new_n683), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n881), .B1(new_n842), .B2(new_n843), .ZN(new_n915));
  OR2_X1    g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n688), .B1(new_n859), .B2(KEYINPUT121), .ZN(new_n917));
  OAI211_X1 g716(.A(new_n916), .B(new_n917), .C1(KEYINPUT121), .C2(new_n859), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n910), .B1(new_n918), .B2(G148gat), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n909), .B1(new_n912), .B2(new_n919), .ZN(G1345gat));
  AND3_X1   g719(.A1(new_n891), .A2(new_n893), .A3(new_n878), .ZN(new_n921));
  NAND4_X1  g720(.A1(new_n921), .A2(KEYINPUT122), .A3(new_n667), .A4(new_n570), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT122), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n923), .B1(new_n894), .B2(new_n569), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(new_n315), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT123), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n887), .A2(new_n314), .A3(new_n570), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n926), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n314), .B1(new_n922), .B2(new_n924), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n570), .A2(new_n314), .ZN(new_n931));
  AOI211_X1 g730(.A(new_n859), .B(new_n931), .C1(new_n880), .C2(new_n886), .ZN(new_n932));
  OAI21_X1  g731(.A(KEYINPUT123), .B1(new_n930), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n929), .A2(new_n933), .ZN(G1346gat));
  NAND4_X1  g733(.A1(new_n921), .A2(new_n316), .A3(new_n667), .A4(new_n697), .ZN(new_n935));
  XNOR2_X1  g734(.A(new_n935), .B(KEYINPUT124), .ZN(new_n936));
  AND2_X1   g735(.A1(new_n887), .A2(new_n697), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n936), .B1(new_n316), .B2(new_n937), .ZN(G1347gat));
  NAND2_X1  g737(.A1(new_n431), .A2(new_n474), .ZN(new_n939));
  INV_X1    g738(.A(new_n939), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n844), .A2(new_n940), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n941), .A2(new_n281), .ZN(new_n942));
  XNOR2_X1  g741(.A(new_n942), .B(new_n354), .ZN(G1348gat));
  NOR2_X1   g742(.A1(new_n941), .A2(new_n688), .ZN(new_n944));
  XNOR2_X1  g743(.A(new_n944), .B(new_n355), .ZN(G1349gat));
  NAND3_X1  g744(.A1(new_n844), .A2(new_n570), .A3(new_n940), .ZN(new_n946));
  INV_X1    g745(.A(G183gat), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n948), .B1(new_n362), .B2(new_n946), .ZN(new_n949));
  XOR2_X1   g748(.A(new_n949), .B(KEYINPUT60), .Z(G1350gat));
  NAND3_X1  g749(.A1(new_n844), .A2(new_n697), .A3(new_n940), .ZN(new_n951));
  OR2_X1    g750(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(KEYINPUT125), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT125), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n951), .A2(new_n955), .A3(new_n952), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  AND2_X1   g756(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n958));
  XNOR2_X1  g757(.A(new_n957), .B(new_n958), .ZN(G1351gat));
  NOR2_X1   g758(.A1(new_n738), .A2(new_n939), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n916), .A2(new_n280), .A3(new_n960), .ZN(new_n961));
  AND3_X1   g760(.A1(new_n878), .A2(new_n892), .A3(new_n940), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n281), .A2(G197gat), .ZN(new_n963));
  AOI22_X1  g762(.A1(new_n961), .A2(G197gat), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  XNOR2_X1  g763(.A(new_n964), .B(KEYINPUT126), .ZN(G1352gat));
  NAND3_X1  g764(.A1(new_n962), .A2(new_n391), .A3(new_n662), .ZN(new_n966));
  XOR2_X1   g765(.A(new_n966), .B(KEYINPUT62), .Z(new_n967));
  AND2_X1   g766(.A1(new_n916), .A2(new_n960), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n968), .A2(new_n662), .ZN(new_n969));
  INV_X1    g768(.A(new_n969), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n967), .B1(new_n970), .B2(new_n391), .ZN(G1353gat));
  INV_X1    g770(.A(G211gat), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n962), .A2(new_n972), .A3(new_n570), .ZN(new_n973));
  OAI211_X1 g772(.A(new_n570), .B(new_n960), .C1(new_n914), .C2(new_n915), .ZN(new_n974));
  AND3_X1   g773(.A1(new_n974), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n975));
  AOI21_X1  g774(.A(KEYINPUT63), .B1(new_n974), .B2(G211gat), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n973), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n977), .A2(KEYINPUT127), .ZN(new_n978));
  INV_X1    g777(.A(KEYINPUT127), .ZN(new_n979));
  OAI211_X1 g778(.A(new_n979), .B(new_n973), .C1(new_n975), .C2(new_n976), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n978), .A2(new_n980), .ZN(G1354gat));
  INV_X1    g780(.A(G218gat), .ZN(new_n982));
  NAND3_X1  g781(.A1(new_n962), .A2(new_n982), .A3(new_n697), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n968), .A2(new_n697), .ZN(new_n984));
  INV_X1    g783(.A(new_n984), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n983), .B1(new_n985), .B2(new_n982), .ZN(G1355gat));
endmodule


