//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 1 0 1 1 0 1 1 0 1 0 1 1 1 0 1 0 0 1 0 1 1 1 1 1 0 0 1 1 1 0 0 1 0 1 1 0 1 1 1 1 0 0 0 0 0 0 1 0 0 0 0 1 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:00 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n670, new_n671, new_n672, new_n673, new_n674, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n696, new_n697, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n712, new_n713, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n744, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n924, new_n925, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G469), .ZN(new_n190));
  INV_X1    g004(.A(G902), .ZN(new_n191));
  INV_X1    g005(.A(G104), .ZN(new_n192));
  OAI21_X1  g006(.A(KEYINPUT3), .B1(new_n192), .B2(G107), .ZN(new_n193));
  AOI21_X1  g007(.A(G101), .B1(new_n192), .B2(G107), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT3), .ZN(new_n195));
  INV_X1    g009(.A(G107), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n195), .A2(new_n196), .A3(G104), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n193), .A2(new_n194), .A3(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(KEYINPUT81), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT81), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n193), .A2(new_n194), .A3(new_n197), .A4(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n199), .A2(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n196), .A2(G104), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n192), .A2(G107), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G101), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n202), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT84), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G143), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n210), .A2(KEYINPUT1), .A3(G146), .ZN(new_n211));
  INV_X1    g025(.A(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G146), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G143), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n210), .A2(G146), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G128), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n212), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  XNOR2_X1  g032(.A(G143), .B(G146), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT1), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n219), .A2(new_n220), .A3(G128), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n218), .A2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT10), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  AOI22_X1  g039(.A1(new_n199), .A2(new_n201), .B1(G101), .B2(new_n205), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(KEYINPUT84), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n209), .A2(new_n225), .A3(new_n227), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n193), .A2(new_n197), .A3(new_n204), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT4), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n229), .A2(new_n230), .A3(G101), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(KEYINPUT82), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT82), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n229), .A2(new_n233), .A3(new_n230), .A4(G101), .ZN(new_n234));
  AND2_X1   g048(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT66), .ZN(new_n236));
  AND2_X1   g050(.A1(KEYINPUT0), .A2(G128), .ZN(new_n237));
  NOR2_X1   g051(.A1(KEYINPUT0), .A2(G128), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT64), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n216), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n219), .A2(new_n237), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n240), .B1(new_n216), .B2(new_n239), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n236), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  XNOR2_X1  g059(.A(KEYINPUT0), .B(G128), .ZN(new_n246));
  OAI21_X1  g060(.A(KEYINPUT64), .B1(new_n219), .B2(new_n246), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n247), .A2(new_n241), .A3(KEYINPUT66), .A4(new_n242), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n230), .B1(new_n229), .B2(G101), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n202), .A2(new_n249), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n235), .A2(new_n245), .A3(new_n248), .A4(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT11), .ZN(new_n252));
  INV_X1    g066(.A(G134), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n252), .B1(new_n253), .B2(G137), .ZN(new_n254));
  INV_X1    g068(.A(G137), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n255), .A2(KEYINPUT11), .A3(G134), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n253), .A2(G137), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n254), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(G131), .ZN(new_n259));
  INV_X1    g073(.A(G131), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n254), .A2(new_n256), .A3(new_n260), .A4(new_n257), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(KEYINPUT67), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT67), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n259), .A2(new_n264), .A3(new_n261), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n211), .B1(new_n219), .B2(G128), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(KEYINPUT83), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT83), .ZN(new_n269));
  OAI211_X1 g083(.A(new_n269), .B(new_n211), .C1(new_n219), .C2(G128), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n268), .A2(new_n221), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(new_n226), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(new_n224), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n228), .A2(new_n251), .A3(new_n266), .A4(new_n273), .ZN(new_n274));
  XNOR2_X1  g088(.A(G110), .B(G140), .ZN(new_n275));
  INV_X1    g089(.A(G953), .ZN(new_n276));
  AND2_X1   g090(.A1(new_n276), .A2(G227), .ZN(new_n277));
  XNOR2_X1  g091(.A(new_n275), .B(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n274), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n207), .A2(new_n223), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(new_n272), .ZN(new_n282));
  INV_X1    g096(.A(new_n266), .ZN(new_n283));
  AOI21_X1  g097(.A(KEYINPUT12), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(KEYINPUT85), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT85), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n266), .B1(new_n281), .B2(new_n272), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n286), .B1(new_n287), .B2(KEYINPUT12), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n285), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n282), .A2(KEYINPUT12), .A3(new_n262), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n280), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n228), .A2(new_n251), .A3(new_n273), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(new_n283), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n279), .B1(new_n293), .B2(new_n274), .ZN(new_n294));
  OAI211_X1 g108(.A(new_n190), .B(new_n191), .C1(new_n291), .C2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(KEYINPUT86), .ZN(new_n296));
  AND2_X1   g110(.A1(new_n293), .A2(new_n274), .ZN(new_n297));
  INV_X1    g111(.A(new_n290), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n298), .B1(new_n285), .B2(new_n288), .ZN(new_n299));
  OAI22_X1  g113(.A1(new_n297), .A2(new_n279), .B1(new_n299), .B2(new_n280), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT86), .ZN(new_n301));
  NAND4_X1  g115(.A1(new_n300), .A2(new_n301), .A3(new_n190), .A4(new_n191), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n296), .A2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(new_n288), .ZN(new_n304));
  NOR3_X1   g118(.A1(new_n287), .A2(new_n286), .A3(KEYINPUT12), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n290), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n279), .B1(new_n306), .B2(new_n274), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n280), .B1(new_n283), .B2(new_n292), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n191), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(G469), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n189), .B1(new_n303), .B2(new_n310), .ZN(new_n311));
  OAI21_X1  g125(.A(G214), .B1(G237), .B2(G902), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(G119), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(G116), .ZN(new_n315));
  INV_X1    g129(.A(G116), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(G119), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  XNOR2_X1  g133(.A(KEYINPUT2), .B(G113), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n318), .A2(new_n320), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n250), .A2(new_n324), .A3(new_n232), .A4(new_n234), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(KEYINPUT87), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n319), .A2(KEYINPUT5), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n315), .A2(KEYINPUT5), .ZN(new_n328));
  INV_X1    g142(.A(G113), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  AOI22_X1  g144(.A1(new_n327), .A2(new_n330), .B1(new_n321), .B2(new_n319), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n209), .A2(new_n227), .A3(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT87), .ZN(new_n333));
  NAND4_X1  g147(.A1(new_n235), .A2(new_n333), .A3(new_n324), .A4(new_n250), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n326), .A2(new_n332), .A3(new_n334), .ZN(new_n335));
  XNOR2_X1  g149(.A(G110), .B(G122), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  NAND4_X1  g152(.A1(new_n326), .A2(new_n332), .A3(new_n334), .A4(new_n336), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n338), .A2(KEYINPUT6), .A3(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n247), .A2(new_n242), .A3(new_n241), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(G125), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n342), .B1(G125), .B2(new_n222), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n276), .A2(G224), .ZN(new_n344));
  XOR2_X1   g158(.A(new_n343), .B(new_n344), .Z(new_n345));
  INV_X1    g159(.A(KEYINPUT6), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n335), .A2(new_n346), .A3(new_n337), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n340), .A2(new_n345), .A3(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT90), .ZN(new_n349));
  XOR2_X1   g163(.A(new_n336), .B(KEYINPUT8), .Z(new_n350));
  INV_X1    g164(.A(KEYINPUT88), .ZN(new_n351));
  OAI21_X1  g165(.A(KEYINPUT89), .B1(new_n207), .B2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT89), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n331), .B1(new_n226), .B2(new_n353), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n350), .B1(new_n352), .B2(new_n354), .ZN(new_n355));
  OAI211_X1 g169(.A(KEYINPUT89), .B(new_n331), .C1(new_n207), .C2(new_n351), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n343), .A2(KEYINPUT7), .A3(new_n344), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n344), .A2(KEYINPUT7), .ZN(new_n358));
  OAI211_X1 g172(.A(new_n342), .B(new_n358), .C1(G125), .C2(new_n222), .ZN(new_n359));
  AOI22_X1  g173(.A1(new_n355), .A2(new_n356), .B1(new_n357), .B2(new_n359), .ZN(new_n360));
  AOI211_X1 g174(.A(new_n349), .B(G902), .C1(new_n360), .C2(new_n339), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n355), .A2(new_n356), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n357), .A2(new_n359), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n339), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(KEYINPUT90), .B1(new_n364), .B2(new_n191), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n348), .B1(new_n361), .B2(new_n365), .ZN(new_n366));
  OAI21_X1  g180(.A(G210), .B1(G237), .B2(G902), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n366), .A2(KEYINPUT91), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(KEYINPUT91), .ZN(new_n370));
  OAI211_X1 g184(.A(new_n348), .B(new_n370), .C1(new_n361), .C2(new_n365), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n313), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  AND2_X1   g186(.A1(new_n311), .A2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT71), .ZN(new_n374));
  NOR2_X1   g188(.A1(G237), .A2(G953), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(G210), .ZN(new_n376));
  XNOR2_X1  g190(.A(new_n376), .B(KEYINPUT27), .ZN(new_n377));
  XNOR2_X1  g191(.A(KEYINPUT26), .B(G101), .ZN(new_n378));
  XNOR2_X1  g192(.A(new_n377), .B(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  NAND4_X1  g194(.A1(new_n245), .A2(new_n263), .A3(new_n265), .A4(new_n248), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n253), .A2(G137), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n255), .A2(G134), .ZN(new_n383));
  OAI21_X1  g197(.A(G131), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n261), .A2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT68), .ZN(new_n386));
  AOI22_X1  g200(.A1(new_n385), .A2(new_n386), .B1(new_n218), .B2(new_n221), .ZN(new_n387));
  AND2_X1   g201(.A1(new_n261), .A2(new_n384), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(KEYINPUT68), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n324), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  AOI21_X1  g204(.A(KEYINPUT28), .B1(new_n381), .B2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  AND3_X1   g206(.A1(new_n381), .A2(KEYINPUT69), .A3(new_n390), .ZN(new_n393));
  AOI21_X1  g207(.A(KEYINPUT69), .B1(new_n381), .B2(new_n390), .ZN(new_n394));
  INV_X1    g208(.A(new_n324), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n341), .A2(KEYINPUT65), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT65), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n247), .A2(new_n241), .A3(new_n397), .A4(new_n242), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n396), .A2(new_n398), .A3(new_n262), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n222), .A2(new_n388), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n395), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NOR3_X1   g215(.A1(new_n393), .A2(new_n394), .A3(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT28), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n392), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT31), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n387), .A2(new_n389), .ZN(new_n406));
  AND3_X1   g220(.A1(new_n381), .A2(KEYINPUT30), .A3(new_n406), .ZN(new_n407));
  AOI21_X1  g221(.A(KEYINPUT30), .B1(new_n399), .B2(new_n400), .ZN(new_n408));
  NOR3_X1   g222(.A1(new_n407), .A2(new_n395), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n381), .A2(new_n390), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT69), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n381), .A2(new_n390), .A3(KEYINPUT69), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n412), .A2(new_n413), .A3(new_n379), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n405), .B1(new_n409), .B2(new_n414), .ZN(new_n415));
  NOR3_X1   g229(.A1(new_n393), .A2(new_n394), .A3(new_n380), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n381), .A2(KEYINPUT30), .A3(new_n406), .ZN(new_n417));
  AOI22_X1  g231(.A1(new_n341), .A2(KEYINPUT65), .B1(new_n261), .B2(new_n259), .ZN(new_n418));
  AOI22_X1  g232(.A1(new_n418), .A2(new_n398), .B1(new_n222), .B2(new_n388), .ZN(new_n419));
  OAI211_X1 g233(.A(new_n417), .B(new_n324), .C1(new_n419), .C2(KEYINPUT30), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n416), .A2(KEYINPUT31), .A3(new_n420), .ZN(new_n421));
  AOI22_X1  g235(.A1(new_n380), .A2(new_n404), .B1(new_n415), .B2(new_n421), .ZN(new_n422));
  NOR2_X1   g236(.A1(G472), .A2(G902), .ZN(new_n423));
  XNOR2_X1  g237(.A(new_n423), .B(KEYINPUT70), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n374), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT32), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n393), .A2(new_n394), .ZN(new_n427));
  AND4_X1   g241(.A1(KEYINPUT31), .A2(new_n427), .A3(new_n420), .A4(new_n379), .ZN(new_n428));
  AOI21_X1  g242(.A(KEYINPUT31), .B1(new_n416), .B2(new_n420), .ZN(new_n429));
  INV_X1    g243(.A(new_n401), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n430), .A2(new_n412), .A3(new_n413), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n391), .B1(new_n431), .B2(KEYINPUT28), .ZN(new_n432));
  OAI22_X1  g246(.A1(new_n428), .A2(new_n429), .B1(new_n432), .B2(new_n379), .ZN(new_n433));
  INV_X1    g247(.A(new_n424), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n433), .A2(KEYINPUT71), .A3(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n425), .A2(new_n426), .A3(new_n435), .ZN(new_n436));
  NOR3_X1   g250(.A1(new_n422), .A2(new_n426), .A3(new_n424), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT75), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n427), .A2(new_n420), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(new_n380), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT72), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT29), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n440), .A2(KEYINPUT72), .A3(new_n380), .ZN(new_n445));
  OAI211_X1 g259(.A(new_n379), .B(new_n392), .C1(new_n402), .C2(new_n403), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n443), .A2(new_n444), .A3(new_n445), .A4(new_n446), .ZN(new_n447));
  XNOR2_X1  g261(.A(new_n391), .B(KEYINPUT74), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n381), .A2(new_n406), .ZN(new_n449));
  AOI21_X1  g263(.A(KEYINPUT73), .B1(new_n449), .B2(new_n324), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT73), .ZN(new_n451));
  AOI211_X1 g265(.A(new_n451), .B(new_n395), .C1(new_n381), .C2(new_n406), .ZN(new_n452));
  OAI211_X1 g266(.A(new_n412), .B(new_n413), .C1(new_n450), .C2(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n448), .B1(new_n453), .B2(KEYINPUT28), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n380), .A2(new_n444), .ZN(new_n455));
  AOI21_X1  g269(.A(G902), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n447), .A2(new_n456), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n439), .B1(new_n457), .B2(G472), .ZN(new_n458));
  INV_X1    g272(.A(G472), .ZN(new_n459));
  AOI211_X1 g273(.A(KEYINPUT75), .B(new_n459), .C1(new_n447), .C2(new_n456), .ZN(new_n460));
  OAI211_X1 g274(.A(new_n436), .B(new_n438), .C1(new_n458), .C2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n217), .A2(G119), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT23), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n462), .B1(KEYINPUT76), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n314), .A2(G128), .ZN(new_n465));
  XNOR2_X1  g279(.A(KEYINPUT76), .B(KEYINPUT23), .ZN(new_n466));
  OAI211_X1 g280(.A(new_n464), .B(new_n465), .C1(new_n466), .C2(new_n462), .ZN(new_n467));
  AND2_X1   g281(.A1(new_n462), .A2(new_n465), .ZN(new_n468));
  XOR2_X1   g282(.A(KEYINPUT24), .B(G110), .Z(new_n469));
  OAI22_X1  g283(.A1(new_n467), .A2(G110), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(KEYINPUT77), .A2(G125), .ZN(new_n471));
  INV_X1    g285(.A(G140), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(KEYINPUT77), .A2(G125), .A3(G140), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n473), .A2(KEYINPUT16), .A3(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT16), .ZN(new_n476));
  INV_X1    g290(.A(G125), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n476), .B1(new_n477), .B2(G140), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n213), .B1(new_n475), .B2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  XNOR2_X1  g294(.A(G125), .B(G140), .ZN(new_n481));
  AOI21_X1  g295(.A(KEYINPUT78), .B1(new_n481), .B2(new_n213), .ZN(new_n482));
  AND3_X1   g296(.A1(new_n481), .A2(KEYINPUT78), .A3(new_n213), .ZN(new_n483));
  OAI211_X1 g297(.A(new_n470), .B(new_n480), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n467), .A2(G110), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n468), .A2(new_n469), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n475), .A2(new_n478), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n487), .A2(G146), .ZN(new_n488));
  OAI211_X1 g302(.A(new_n485), .B(new_n486), .C1(new_n488), .C2(new_n479), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n484), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n276), .A2(G221), .A3(G234), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n491), .B(KEYINPUT79), .ZN(new_n492));
  XNOR2_X1  g306(.A(KEYINPUT22), .B(G137), .ZN(new_n493));
  XNOR2_X1  g307(.A(new_n492), .B(new_n493), .ZN(new_n494));
  XNOR2_X1  g308(.A(new_n490), .B(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT80), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT25), .ZN(new_n497));
  AOI21_X1  g311(.A(G902), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n495), .A2(new_n498), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n496), .A2(new_n497), .ZN(new_n500));
  OR2_X1    g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(G234), .ZN(new_n502));
  OAI21_X1  g316(.A(G217), .B1(new_n502), .B2(G902), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n503), .B1(new_n499), .B2(new_n500), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n501), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(G902), .B1(new_n502), .B2(G217), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n495), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  NOR2_X1   g323(.A1(G475), .A2(G902), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(G237), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n512), .A2(new_n276), .A3(G214), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n513), .A2(KEYINPUT92), .A3(new_n210), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n210), .A2(KEYINPUT92), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n515), .A2(G214), .A3(new_n375), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(G131), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n514), .A2(new_n260), .A3(new_n516), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n479), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n473), .A2(new_n474), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT93), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n473), .A2(KEYINPUT93), .A3(new_n474), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n523), .A2(new_n524), .A3(KEYINPUT19), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT19), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n481), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n525), .A2(new_n213), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n520), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n523), .A2(new_n524), .A3(G146), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n530), .B1(new_n482), .B2(new_n483), .ZN(new_n531));
  NAND2_X1  g345(.A1(KEYINPUT18), .A2(G131), .ZN(new_n532));
  AND3_X1   g346(.A1(new_n514), .A2(new_n532), .A3(new_n516), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n532), .B1(new_n514), .B2(new_n516), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n531), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n529), .A2(new_n536), .ZN(new_n537));
  XOR2_X1   g351(.A(G113), .B(G122), .Z(new_n538));
  XOR2_X1   g352(.A(KEYINPUT94), .B(G104), .Z(new_n539));
  XOR2_X1   g353(.A(new_n538), .B(new_n539), .Z(new_n540));
  NAND2_X1  g354(.A1(new_n537), .A2(new_n540), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n488), .A2(new_n479), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT17), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n518), .A2(new_n543), .A3(new_n519), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n517), .A2(KEYINPUT17), .A3(G131), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n542), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(new_n540), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n546), .A2(new_n547), .A3(new_n536), .ZN(new_n548));
  AOI211_X1 g362(.A(KEYINPUT20), .B(new_n511), .C1(new_n541), .C2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT20), .ZN(new_n550));
  AOI22_X1  g364(.A1(new_n520), .A2(new_n528), .B1(new_n531), .B2(new_n535), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n548), .B1(new_n547), .B2(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n550), .B1(new_n552), .B2(new_n510), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n549), .A2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(G475), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n546), .A2(new_n536), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT95), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n556), .A2(new_n557), .A3(new_n540), .ZN(new_n558));
  AND2_X1   g372(.A1(new_n558), .A2(new_n191), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n556), .A2(new_n540), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n560), .A2(KEYINPUT95), .A3(new_n548), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n555), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n554), .A2(new_n562), .ZN(new_n563));
  XNOR2_X1  g377(.A(G128), .B(G143), .ZN(new_n564));
  XNOR2_X1  g378(.A(KEYINPUT96), .B(KEYINPUT13), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n210), .A2(G128), .ZN(new_n567));
  OAI211_X1 g381(.A(new_n566), .B(G134), .C1(new_n567), .C2(new_n565), .ZN(new_n568));
  XNOR2_X1  g382(.A(G116), .B(G122), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n569), .B(new_n196), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n564), .A2(new_n253), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n568), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n564), .B(new_n253), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n316), .A2(KEYINPUT14), .A3(G122), .ZN(new_n574));
  INV_X1    g388(.A(new_n569), .ZN(new_n575));
  OAI211_X1 g389(.A(G107), .B(new_n574), .C1(new_n575), .C2(KEYINPUT14), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n569), .A2(new_n196), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n573), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(G217), .ZN(new_n579));
  NOR3_X1   g393(.A1(new_n187), .A2(new_n579), .A3(G953), .ZN(new_n580));
  AND3_X1   g394(.A1(new_n572), .A2(new_n578), .A3(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n580), .B1(new_n572), .B2(new_n578), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n191), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(G478), .ZN(new_n584));
  OR2_X1    g398(.A1(new_n584), .A2(KEYINPUT15), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n583), .B(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n563), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(G234), .A2(G237), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n588), .A2(G952), .A3(new_n276), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n588), .A2(G902), .A3(G953), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n590), .B(KEYINPUT97), .ZN(new_n591));
  XNOR2_X1  g405(.A(KEYINPUT21), .B(G898), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n589), .B1(new_n591), .B2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n587), .A2(new_n595), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n373), .A2(new_n461), .A3(new_n509), .A4(new_n596), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n597), .B(G101), .ZN(G3));
  NAND2_X1  g412(.A1(new_n303), .A2(new_n310), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(new_n188), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n404), .A2(new_n380), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n415), .A2(new_n421), .ZN(new_n602));
  AOI211_X1 g416(.A(new_n374), .B(new_n424), .C1(new_n601), .C2(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(KEYINPUT71), .B1(new_n433), .B2(new_n434), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  OAI21_X1  g419(.A(G472), .B1(new_n422), .B2(G902), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n600), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n366), .A2(new_n367), .ZN(new_n609));
  OAI211_X1 g423(.A(new_n348), .B(new_n368), .C1(new_n361), .C2(new_n365), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n609), .A2(new_n312), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n583), .A2(new_n584), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT33), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n581), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n572), .A2(new_n578), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n580), .B(KEYINPUT98), .ZN(new_n616));
  AND3_X1   g430(.A1(new_n615), .A2(KEYINPUT99), .A3(new_n616), .ZN(new_n617));
  AOI21_X1  g431(.A(KEYINPUT99), .B1(new_n615), .B2(new_n616), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n614), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n613), .B1(new_n581), .B2(new_n582), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n191), .A2(G478), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n612), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n623), .B1(new_n554), .B2(new_n562), .ZN(new_n624));
  NOR4_X1   g438(.A1(new_n611), .A2(new_n508), .A3(new_n595), .A4(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n608), .A2(new_n625), .ZN(new_n626));
  XOR2_X1   g440(.A(KEYINPUT34), .B(G104), .Z(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(G6));
  NOR3_X1   g442(.A1(new_n554), .A2(new_n562), .A3(new_n586), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  NOR4_X1   g444(.A1(new_n611), .A2(new_n508), .A3(new_n595), .A4(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n608), .A2(new_n631), .ZN(new_n632));
  XOR2_X1   g446(.A(KEYINPUT35), .B(G107), .Z(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G9));
  INV_X1    g448(.A(new_n494), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n635), .A2(KEYINPUT36), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(new_n490), .ZN(new_n637));
  AOI22_X1  g451(.A1(new_n501), .A2(new_n504), .B1(new_n506), .B2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n596), .A2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n373), .A2(new_n605), .A3(new_n606), .A4(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT37), .B(G110), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G12));
  AOI21_X1  g458(.A(new_n313), .B1(new_n366), .B2(new_n367), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n645), .A2(new_n639), .A3(new_n610), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n589), .B(KEYINPUT100), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n647), .B1(new_n591), .B2(G900), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n629), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n461), .A2(new_n311), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(G128), .ZN(G30));
  XNOR2_X1  g466(.A(new_n648), .B(KEYINPUT39), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n311), .A2(new_n653), .ZN(new_n654));
  XOR2_X1   g468(.A(new_n654), .B(KEYINPUT40), .Z(new_n655));
  NAND2_X1  g469(.A1(new_n369), .A2(new_n371), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(KEYINPUT38), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  AOI22_X1  g472(.A1(new_n453), .A2(new_n380), .B1(new_n420), .B2(new_n416), .ZN(new_n659));
  OAI21_X1  g473(.A(G472), .B1(new_n659), .B2(G902), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n436), .A2(new_n438), .A3(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(new_n554), .ZN(new_n663));
  INV_X1    g477(.A(new_n562), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n586), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n638), .A2(new_n665), .A3(new_n312), .ZN(new_n666));
  NOR3_X1   g480(.A1(new_n658), .A2(new_n662), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n655), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(G143), .ZN(G45));
  OAI211_X1 g483(.A(new_n623), .B(new_n648), .C1(new_n554), .C2(new_n562), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n646), .A2(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n458), .A2(new_n460), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n436), .A2(new_n438), .ZN(new_n673));
  OAI211_X1 g487(.A(new_n311), .B(new_n671), .C1(new_n672), .C2(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G146), .ZN(G48));
  OAI21_X1  g489(.A(new_n625), .B1(new_n672), .B2(new_n673), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n300), .A2(new_n191), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(G469), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n303), .A2(new_n188), .A3(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT101), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  AOI22_X1  g495(.A1(new_n296), .A2(new_n302), .B1(G469), .B2(new_n677), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n682), .A2(KEYINPUT101), .A3(new_n188), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  OAI21_X1  g498(.A(KEYINPUT102), .B1(new_n676), .B2(new_n684), .ZN(new_n685));
  AND4_X1   g499(.A1(KEYINPUT101), .A2(new_n303), .A3(new_n188), .A4(new_n678), .ZN(new_n686));
  AOI21_X1  g500(.A(KEYINPUT101), .B1(new_n682), .B2(new_n188), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT102), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n688), .A2(new_n689), .A3(new_n461), .A4(new_n625), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n685), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(KEYINPUT41), .B(G113), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(G15));
  NAND4_X1  g507(.A1(new_n461), .A2(new_n631), .A3(new_n681), .A4(new_n683), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G116), .ZN(G18));
  NOR2_X1   g509(.A1(new_n679), .A2(new_n611), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n461), .A2(new_n641), .A3(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G119), .ZN(G21));
  NAND4_X1  g512(.A1(new_n609), .A2(new_n312), .A3(new_n610), .A4(new_n665), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(KEYINPUT104), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT104), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n645), .A2(new_n701), .A3(new_n610), .A4(new_n665), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(KEYINPUT103), .B(G472), .ZN(new_n704));
  OAI21_X1  g518(.A(new_n704), .B1(new_n422), .B2(G902), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n602), .B1(new_n454), .B2(new_n379), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(new_n434), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n509), .A2(new_n705), .A3(new_n707), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n708), .A2(new_n595), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n703), .A2(new_n681), .A3(new_n709), .A4(new_n683), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G122), .ZN(G24));
  NAND3_X1  g525(.A1(new_n705), .A2(new_n639), .A3(new_n707), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n670), .B(KEYINPUT105), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n696), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G125), .ZN(G27));
  AOI22_X1  g530(.A1(new_n296), .A2(new_n302), .B1(new_n309), .B2(G469), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n369), .A2(new_n312), .A3(new_n371), .ZN(new_n718));
  NOR3_X1   g532(.A1(new_n717), .A2(new_n718), .A3(new_n189), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n713), .A2(KEYINPUT42), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n461), .A2(new_n509), .A3(new_n719), .A4(new_n720), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n426), .B1(new_n422), .B2(new_n424), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n438), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n446), .A2(new_n444), .ZN(new_n724));
  AOI21_X1  g538(.A(KEYINPUT72), .B1(new_n440), .B2(new_n380), .ZN(new_n725));
  AOI211_X1 g539(.A(new_n442), .B(new_n379), .C1(new_n427), .C2(new_n420), .ZN(new_n726));
  NOR3_X1   g540(.A1(new_n724), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n453), .A2(KEYINPUT28), .ZN(new_n728));
  INV_X1    g542(.A(new_n448), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n728), .A2(new_n729), .A3(new_n455), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(new_n191), .ZN(new_n731));
  OAI21_X1  g545(.A(G472), .B1(new_n727), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(KEYINPUT75), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n457), .A2(new_n439), .A3(G472), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n723), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT105), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n670), .B(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(new_n718), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n311), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  NOR3_X1   g553(.A1(new_n735), .A2(new_n739), .A3(new_n508), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT42), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n721), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(new_n260), .ZN(G33));
  INV_X1    g557(.A(new_n649), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n461), .A2(new_n509), .A3(new_n719), .A4(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G134), .ZN(G36));
  NAND2_X1  g560(.A1(new_n563), .A2(new_n623), .ZN(new_n747));
  XOR2_X1   g561(.A(new_n747), .B(KEYINPUT43), .Z(new_n748));
  NAND3_X1  g562(.A1(new_n607), .A2(new_n748), .A3(new_n639), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT44), .ZN(new_n750));
  OR2_X1    g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n749), .A2(new_n750), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n751), .A2(new_n738), .A3(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT107), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n751), .A2(KEYINPUT107), .A3(new_n738), .A4(new_n752), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT45), .ZN(new_n758));
  OR3_X1    g572(.A1(new_n307), .A2(new_n758), .A3(new_n308), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n758), .B1(new_n307), .B2(new_n308), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n759), .A2(G469), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(G469), .A2(G902), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT46), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(new_n303), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n763), .A2(new_n764), .ZN(new_n767));
  OAI211_X1 g581(.A(new_n188), .B(new_n653), .C1(new_n766), .C2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT106), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n768), .B(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n757), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G137), .ZN(G39));
  OAI21_X1  g586(.A(new_n188), .B1(new_n766), .B2(new_n767), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT47), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NOR4_X1   g589(.A1(new_n461), .A2(new_n509), .A3(new_n670), .A4(new_n718), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G140), .ZN(G42));
  NAND4_X1  g592(.A1(new_n682), .A2(new_n188), .A3(new_n610), .A4(new_n645), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n737), .A2(new_n639), .A3(new_n707), .A4(new_n705), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n733), .A2(new_n734), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n437), .B1(new_n605), .B2(new_n426), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n600), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n781), .B1(new_n784), .B2(new_n650), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT110), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n638), .A2(new_n648), .ZN(new_n787));
  INV_X1    g601(.A(new_n787), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n786), .B1(new_n311), .B2(new_n788), .ZN(new_n789));
  NOR4_X1   g603(.A1(new_n717), .A2(KEYINPUT110), .A3(new_n189), .A4(new_n787), .ZN(new_n790));
  OAI211_X1 g604(.A(new_n661), .B(new_n703), .C1(new_n789), .C2(new_n790), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n785), .A2(KEYINPUT52), .A3(new_n674), .A4(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT111), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n651), .A2(new_n674), .A3(new_n715), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n703), .A2(new_n661), .ZN(new_n796));
  OAI21_X1  g610(.A(KEYINPUT110), .B1(new_n600), .B2(new_n787), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n311), .A2(new_n786), .A3(new_n788), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n796), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n795), .A2(new_n799), .ZN(new_n800));
  XOR2_X1   g614(.A(KEYINPUT112), .B(KEYINPUT52), .Z(new_n801));
  OR3_X1    g615(.A1(new_n800), .A2(KEYINPUT113), .A3(new_n801), .ZN(new_n802));
  OAI21_X1  g616(.A(KEYINPUT113), .B1(new_n800), .B2(new_n801), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n794), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  AND3_X1   g618(.A1(new_n694), .A2(new_n697), .A3(new_n710), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n691), .A2(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT109), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n630), .A2(new_n624), .ZN(new_n809));
  AND4_X1   g623(.A1(new_n509), .A2(new_n372), .A3(new_n594), .A4(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n608), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n597), .A2(new_n642), .A3(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(new_n648), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n638), .A2(new_n587), .A3(new_n813), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n714), .B1(new_n461), .B2(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(new_n719), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n745), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n742), .A2(new_n812), .A3(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n691), .A2(new_n805), .A3(KEYINPUT109), .ZN(new_n819));
  AND3_X1   g633(.A1(new_n808), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT53), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n804), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT52), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n823), .B1(new_n795), .B2(new_n799), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n824), .A2(new_n792), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n808), .A2(new_n818), .A3(new_n825), .A4(new_n819), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(KEYINPUT53), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n822), .A2(new_n827), .ZN(new_n828));
  AND4_X1   g642(.A1(KEYINPUT53), .A2(new_n818), .A3(new_n691), .A4(new_n805), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n804), .A2(new_n829), .ZN(new_n830));
  AND3_X1   g644(.A1(new_n826), .A2(KEYINPUT114), .A3(new_n821), .ZN(new_n831));
  AOI21_X1  g645(.A(KEYINPUT114), .B1(new_n826), .B2(new_n821), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n830), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT54), .ZN(new_n834));
  MUX2_X1   g648(.A(new_n828), .B(new_n833), .S(new_n834), .Z(new_n835));
  INV_X1    g649(.A(new_n679), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(new_n738), .ZN(new_n837));
  INV_X1    g651(.A(new_n647), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n748), .A2(new_n838), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n837), .A2(new_n839), .A3(new_n712), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n839), .A2(new_n708), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n841), .A2(new_n313), .A3(new_n658), .A4(new_n836), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n842), .B(KEYINPUT50), .ZN(new_n843));
  NOR4_X1   g657(.A1(new_n837), .A2(new_n508), .A3(new_n589), .A4(new_n661), .ZN(new_n844));
  NOR3_X1   g658(.A1(new_n623), .A2(new_n554), .A3(new_n562), .ZN(new_n845));
  AOI211_X1 g659(.A(new_n840), .B(new_n843), .C1(new_n844), .C2(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n841), .A2(new_n738), .ZN(new_n847));
  XOR2_X1   g661(.A(new_n847), .B(KEYINPUT115), .Z(new_n848));
  INV_X1    g662(.A(new_n682), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n849), .A2(new_n188), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n848), .B1(new_n775), .B2(new_n850), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n846), .A2(KEYINPUT51), .A3(new_n851), .ZN(new_n852));
  AOI21_X1  g666(.A(KEYINPUT51), .B1(new_n846), .B2(new_n851), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n276), .A2(G952), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n841), .A2(new_n696), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n854), .B1(new_n855), .B2(KEYINPUT116), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n856), .B1(KEYINPUT116), .B2(new_n855), .ZN(new_n857));
  INV_X1    g671(.A(new_n624), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n857), .B1(new_n858), .B2(new_n844), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n509), .B1(new_n672), .B2(new_n723), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n860), .A2(new_n839), .A3(new_n837), .ZN(new_n861));
  XOR2_X1   g675(.A(new_n861), .B(KEYINPUT48), .Z(new_n862));
  NAND2_X1  g676(.A1(new_n859), .A2(new_n862), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n852), .A2(new_n853), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n835), .A2(new_n864), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n865), .B1(G952), .B2(G953), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n849), .A2(KEYINPUT49), .ZN(new_n867));
  XOR2_X1   g681(.A(new_n867), .B(KEYINPUT108), .Z(new_n868));
  NAND3_X1  g682(.A1(new_n509), .A2(new_n312), .A3(new_n188), .ZN(new_n869));
  AOI211_X1 g683(.A(new_n747), .B(new_n869), .C1(new_n849), .C2(KEYINPUT49), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n868), .A2(new_n658), .A3(new_n662), .A4(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n866), .A2(new_n871), .ZN(G75));
  NOR2_X1   g686(.A1(new_n276), .A2(G952), .ZN(new_n873));
  INV_X1    g687(.A(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n826), .A2(new_n821), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT114), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n826), .A2(KEYINPUT114), .A3(new_n821), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n191), .B1(new_n879), .B2(new_n830), .ZN(new_n880));
  AOI21_X1  g694(.A(KEYINPUT56), .B1(new_n880), .B2(G210), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n340), .A2(new_n347), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n882), .B(new_n345), .ZN(new_n883));
  XNOR2_X1  g697(.A(KEYINPUT117), .B(KEYINPUT55), .ZN(new_n884));
  XOR2_X1   g698(.A(new_n883), .B(new_n884), .Z(new_n885));
  OAI21_X1  g699(.A(new_n874), .B1(new_n881), .B2(new_n885), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n886), .B1(new_n881), .B2(new_n885), .ZN(G51));
  AOI21_X1  g701(.A(new_n834), .B1(new_n879), .B2(new_n830), .ZN(new_n888));
  OAI211_X1 g702(.A(new_n830), .B(new_n834), .C1(new_n831), .C2(new_n832), .ZN(new_n889));
  INV_X1    g703(.A(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  XOR2_X1   g705(.A(new_n762), .B(KEYINPUT118), .Z(new_n892));
  XNOR2_X1  g706(.A(new_n892), .B(KEYINPUT57), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n300), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n761), .B(KEYINPUT119), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n880), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n873), .B1(new_n894), .B2(new_n896), .ZN(G54));
  NAND2_X1  g711(.A1(KEYINPUT58), .A2(G475), .ZN(new_n898));
  XOR2_X1   g712(.A(new_n898), .B(KEYINPUT120), .Z(new_n899));
  NAND2_X1  g713(.A1(new_n880), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n900), .B1(new_n548), .B2(new_n541), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n552), .B1(new_n880), .B2(new_n899), .ZN(new_n902));
  NOR3_X1   g716(.A1(new_n901), .A2(new_n873), .A3(new_n902), .ZN(G60));
  NAND2_X1  g717(.A1(G478), .A2(G902), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n904), .B(KEYINPUT59), .Z(new_n905));
  NOR2_X1   g719(.A1(new_n621), .A2(new_n905), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n906), .B1(new_n888), .B2(new_n890), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT121), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n907), .A2(new_n908), .A3(new_n874), .ZN(new_n909));
  INV_X1    g723(.A(new_n906), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n833), .A2(KEYINPUT54), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n910), .B1(new_n911), .B2(new_n889), .ZN(new_n912));
  OAI21_X1  g726(.A(KEYINPUT121), .B1(new_n912), .B2(new_n873), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n621), .B1(new_n835), .B2(new_n905), .ZN(new_n914));
  AND3_X1   g728(.A1(new_n909), .A2(new_n913), .A3(new_n914), .ZN(G63));
  NAND2_X1  g729(.A1(G217), .A2(G902), .ZN(new_n916));
  XOR2_X1   g730(.A(new_n916), .B(KEYINPUT60), .Z(new_n917));
  NAND3_X1  g731(.A1(new_n833), .A2(new_n637), .A3(new_n917), .ZN(new_n918));
  AND2_X1   g732(.A1(new_n833), .A2(new_n917), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n495), .B(KEYINPUT122), .ZN(new_n920));
  OAI211_X1 g734(.A(new_n874), .B(new_n918), .C1(new_n919), .C2(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT61), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n921), .B(new_n922), .ZN(G66));
  AOI21_X1  g737(.A(new_n276), .B1(new_n593), .B2(G224), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n808), .A2(new_n819), .ZN(new_n925));
  OR2_X1    g739(.A1(new_n925), .A2(new_n812), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n924), .B1(new_n926), .B2(new_n276), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n882), .B1(G898), .B2(new_n276), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n927), .B(new_n928), .Z(G69));
  NOR2_X1   g743(.A1(new_n407), .A2(new_n408), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n525), .A2(new_n527), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n930), .B(new_n931), .Z(new_n932));
  AOI21_X1  g746(.A(new_n508), .B1(new_n782), .B2(new_n783), .ZN(new_n933));
  AOI211_X1 g747(.A(new_n718), .B(new_n654), .C1(new_n624), .C2(new_n630), .ZN(new_n934));
  AOI22_X1  g748(.A1(new_n775), .A2(new_n776), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(new_n668), .ZN(new_n936));
  OAI21_X1  g750(.A(KEYINPUT62), .B1(new_n936), .B2(new_n795), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT62), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n668), .A2(new_n938), .A3(new_n674), .A4(new_n785), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n935), .A2(new_n771), .A3(new_n937), .A4(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n932), .B1(new_n940), .B2(new_n276), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n860), .B1(new_n702), .B2(new_n700), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n770), .B1(new_n757), .B2(new_n942), .ZN(new_n943));
  OAI211_X1 g757(.A(new_n721), .B(new_n745), .C1(new_n740), .C2(new_n741), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n944), .A2(new_n795), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n943), .A2(new_n777), .A3(new_n945), .ZN(new_n946));
  OR2_X1    g760(.A1(new_n946), .A2(G953), .ZN(new_n947));
  NAND2_X1  g761(.A1(G900), .A2(G953), .ZN(new_n948));
  AND2_X1   g762(.A1(new_n932), .A2(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n941), .B1(new_n947), .B2(new_n949), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n276), .B1(G227), .B2(G900), .ZN(new_n951));
  XOR2_X1   g765(.A(new_n950), .B(new_n951), .Z(G72));
  NAND2_X1  g766(.A1(G472), .A2(G902), .ZN(new_n953));
  XOR2_X1   g767(.A(new_n953), .B(KEYINPUT63), .Z(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(KEYINPUT123), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n955), .B1(new_n926), .B2(new_n940), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n440), .B(KEYINPUT124), .ZN(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n958), .A2(new_n380), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n873), .B1(new_n956), .B2(new_n959), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n955), .B1(new_n926), .B2(new_n946), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n961), .A2(new_n380), .A3(new_n958), .ZN(new_n962));
  AND2_X1   g776(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  AND2_X1   g777(.A1(new_n822), .A2(new_n827), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT126), .ZN(new_n965));
  INV_X1    g779(.A(new_n954), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n725), .A2(new_n726), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n416), .A2(new_n420), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n966), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n969), .B(KEYINPUT125), .Z(new_n970));
  AND3_X1   g784(.A1(new_n964), .A2(new_n965), .A3(new_n970), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n965), .B1(new_n964), .B2(new_n970), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n963), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n973), .A2(KEYINPUT127), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT127), .ZN(new_n975));
  OAI211_X1 g789(.A(new_n963), .B(new_n975), .C1(new_n971), .C2(new_n972), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n974), .A2(new_n976), .ZN(G57));
endmodule


