//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 1 0 1 0 1 0 0 0 0 0 1 1 0 0 1 0 1 1 0 1 1 0 0 0 1 0 1 1 0 0 0 0 1 1 0 0 1 0 0 1 0 1 1 0 1 0 1 1 0 1 1 1 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:47 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1241, new_n1242, new_n1243,
    new_n1244, new_n1245, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311,
    new_n1312, new_n1313;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  AOI22_X1  g0003(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n204));
  INV_X1    g0004(.A(G68), .ZN(new_n205));
  INV_X1    g0005(.A(G238), .ZN(new_n206));
  INV_X1    g0006(.A(G87), .ZN(new_n207));
  INV_X1    g0007(.A(G250), .ZN(new_n208));
  OAI221_X1 g0008(.A(new_n204), .B1(new_n205), .B2(new_n206), .C1(new_n207), .C2(new_n208), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  OAI21_X1  g0012(.A(new_n203), .B1(new_n209), .B2(new_n212), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT65), .ZN(new_n214));
  INV_X1    g0014(.A(KEYINPUT1), .ZN(new_n215));
  OR2_X1    g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n214), .A2(new_n215), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n203), .A2(G13), .ZN(new_n218));
  OAI211_X1 g0018(.A(new_n218), .B(G250), .C1(G257), .C2(G264), .ZN(new_n219));
  XNOR2_X1  g0019(.A(KEYINPUT64), .B(KEYINPUT0), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n219), .B(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G13), .ZN(new_n222));
  INV_X1    g0022(.A(G20), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(G50), .B1(G58), .B2(G68), .ZN(new_n225));
  INV_X1    g0025(.A(new_n225), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n221), .B1(new_n224), .B2(new_n226), .ZN(new_n227));
  AND3_X1   g0027(.A1(new_n216), .A2(new_n217), .A3(new_n227), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  INV_X1    g0029(.A(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(KEYINPUT2), .B(G226), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT66), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G107), .B(G116), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G50), .B(G68), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G58), .B(G77), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n241), .B(new_n244), .Z(G351));
  AOI21_X1  g0045(.A(new_n222), .B1(G33), .B2(G41), .ZN(new_n246));
  INV_X1    g0046(.A(G274), .ZN(new_n247));
  NOR2_X1   g0047(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(G41), .ZN(new_n249));
  INV_X1    g0049(.A(G45), .ZN(new_n250));
  AOI21_X1  g0050(.A(G1), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(KEYINPUT67), .B(G1), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n249), .A2(new_n250), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(new_n246), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G226), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n252), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  XNOR2_X1  g0059(.A(KEYINPUT3), .B(G33), .ZN(new_n260));
  INV_X1    g0060(.A(G1698), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n260), .A2(G222), .A3(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G77), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n260), .A2(G1698), .ZN(new_n264));
  INV_X1    g0064(.A(G223), .ZN(new_n265));
  OAI221_X1 g0065(.A(new_n262), .B1(new_n263), .B2(new_n260), .C1(new_n264), .C2(new_n265), .ZN(new_n266));
  OR2_X1    g0066(.A1(new_n266), .A2(KEYINPUT68), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n256), .B1(new_n266), .B2(KEYINPUT68), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n259), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G190), .ZN(new_n270));
  NAND3_X1  g0070(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(new_n222), .ZN(new_n272));
  XNOR2_X1  g0072(.A(KEYINPUT8), .B(G58), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n223), .A2(G33), .ZN(new_n274));
  INV_X1    g0074(.A(G150), .ZN(new_n275));
  NOR2_X1   g0075(.A1(G20), .A2(G33), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  OAI22_X1  g0077(.A1(new_n273), .A2(new_n274), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  NOR2_X1   g0078(.A1(G58), .A2(G68), .ZN(new_n279));
  INV_X1    g0079(.A(G50), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n223), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n272), .B1(new_n278), .B2(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n272), .B1(new_n253), .B2(G20), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G50), .ZN(new_n284));
  INV_X1    g0084(.A(G1), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(KEYINPUT67), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT67), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(G1), .ZN(new_n288));
  NAND4_X1  g0088(.A1(new_n286), .A2(new_n288), .A3(G13), .A4(G20), .ZN(new_n289));
  OAI211_X1 g0089(.A(new_n282), .B(new_n284), .C1(G50), .C2(new_n289), .ZN(new_n290));
  XNOR2_X1  g0090(.A(new_n290), .B(KEYINPUT9), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n270), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G200), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n269), .A2(new_n293), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n295), .A2(KEYINPUT69), .A3(KEYINPUT10), .ZN(new_n296));
  NAND2_X1  g0096(.A1(KEYINPUT69), .A2(KEYINPUT10), .ZN(new_n297));
  OR2_X1    g0097(.A1(KEYINPUT69), .A2(KEYINPUT10), .ZN(new_n298));
  OAI211_X1 g0098(.A(new_n297), .B(new_n298), .C1(new_n292), .C2(new_n294), .ZN(new_n299));
  INV_X1    g0099(.A(G179), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n269), .A2(new_n300), .ZN(new_n301));
  OAI211_X1 g0101(.A(new_n301), .B(new_n290), .C1(G169), .C2(new_n269), .ZN(new_n302));
  AND2_X1   g0102(.A1(new_n248), .A2(new_n251), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n246), .B1(new_n253), .B2(new_n254), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n303), .B1(G244), .B2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(G107), .ZN(new_n306));
  OAI22_X1  g0106(.A1(new_n264), .A2(new_n206), .B1(new_n306), .B2(new_n260), .ZN(new_n307));
  INV_X1    g0107(.A(G33), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(KEYINPUT3), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT3), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(G33), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  NOR3_X1   g0112(.A1(new_n312), .A2(new_n230), .A3(G1698), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n246), .B1(new_n307), .B2(new_n313), .ZN(new_n314));
  AND2_X1   g0114(.A1(new_n305), .A2(new_n314), .ZN(new_n315));
  OR2_X1    g0115(.A1(new_n315), .A2(G169), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(new_n300), .ZN(new_n317));
  OAI22_X1  g0117(.A1(new_n273), .A2(new_n277), .B1(new_n223), .B2(new_n263), .ZN(new_n318));
  XNOR2_X1  g0118(.A(KEYINPUT15), .B(G87), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n319), .A2(new_n274), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n272), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n283), .A2(G77), .ZN(new_n322));
  OAI211_X1 g0122(.A(new_n321), .B(new_n322), .C1(G77), .C2(new_n289), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n316), .A2(new_n317), .A3(new_n323), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n323), .B1(new_n315), .B2(G190), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n325), .B1(new_n293), .B2(new_n315), .ZN(new_n326));
  AND2_X1   g0126(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  NAND4_X1  g0127(.A1(new_n296), .A2(new_n299), .A3(new_n302), .A4(new_n327), .ZN(new_n328));
  XNOR2_X1  g0128(.A(new_n328), .B(KEYINPUT70), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n289), .A2(new_n273), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n330), .B1(new_n283), .B2(new_n273), .ZN(new_n331));
  XNOR2_X1  g0131(.A(new_n331), .B(KEYINPUT75), .ZN(new_n332));
  INV_X1    g0132(.A(new_n272), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT7), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n334), .A2(G20), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  AND2_X1   g0136(.A1(KEYINPUT73), .A2(KEYINPUT3), .ZN(new_n337));
  NOR2_X1   g0137(.A1(KEYINPUT73), .A2(KEYINPUT3), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n308), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n336), .B1(new_n339), .B2(new_n311), .ZN(new_n340));
  AOI21_X1  g0140(.A(KEYINPUT7), .B1(new_n312), .B2(new_n223), .ZN(new_n341));
  OAI21_X1  g0141(.A(G68), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(G58), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n343), .A2(new_n205), .ZN(new_n344));
  OAI21_X1  g0144(.A(G20), .B1(new_n344), .B2(new_n279), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n276), .A2(G159), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n342), .A2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT16), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n333), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NOR2_X1   g0151(.A1(KEYINPUT74), .A2(KEYINPUT7), .ZN(new_n352));
  NOR3_X1   g0152(.A1(new_n337), .A2(new_n338), .A3(new_n308), .ZN(new_n353));
  INV_X1    g0153(.A(new_n309), .ZN(new_n354));
  OAI211_X1 g0154(.A(new_n223), .B(new_n352), .C1(new_n353), .C2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(G68), .ZN(new_n356));
  XNOR2_X1  g0156(.A(KEYINPUT74), .B(KEYINPUT7), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT73), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(new_n310), .ZN(new_n359));
  NAND2_X1  g0159(.A1(KEYINPUT73), .A2(KEYINPUT3), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n359), .A2(G33), .A3(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(new_n309), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n357), .B1(new_n362), .B2(new_n223), .ZN(new_n363));
  OAI211_X1 g0163(.A(KEYINPUT16), .B(new_n348), .C1(new_n356), .C2(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n332), .B1(new_n351), .B2(new_n364), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n252), .B1(new_n257), .B2(new_n230), .ZN(new_n366));
  NOR2_X1   g0166(.A1(G223), .A2(G1698), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n367), .B1(new_n258), .B2(G1698), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n368), .A2(new_n361), .A3(new_n309), .ZN(new_n369));
  NAND2_X1  g0169(.A1(G33), .A2(G87), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n256), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n293), .B1(new_n366), .B2(new_n371), .ZN(new_n372));
  AOI22_X1  g0172(.A1(new_n304), .A2(G232), .B1(new_n248), .B2(new_n251), .ZN(new_n373));
  INV_X1    g0173(.A(G190), .ZN(new_n374));
  AND2_X1   g0174(.A1(new_n369), .A2(new_n370), .ZN(new_n375));
  OAI211_X1 g0175(.A(new_n373), .B(new_n374), .C1(new_n375), .C2(new_n256), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n372), .A2(new_n376), .ZN(new_n377));
  AOI21_X1  g0177(.A(KEYINPUT17), .B1(new_n365), .B2(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(G33), .B1(new_n359), .B2(new_n360), .ZN(new_n379));
  INV_X1    g0179(.A(new_n311), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n335), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n334), .B1(new_n260), .B2(G20), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n205), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n350), .B1(new_n383), .B2(new_n347), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n364), .A2(new_n384), .A3(new_n272), .ZN(new_n385));
  XOR2_X1   g0185(.A(new_n331), .B(KEYINPUT75), .Z(new_n386));
  NAND3_X1  g0186(.A1(new_n385), .A2(new_n377), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(KEYINPUT76), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT76), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n365), .A2(new_n389), .A3(new_n377), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n378), .B1(new_n391), .B2(KEYINPUT17), .ZN(new_n392));
  OAI21_X1  g0192(.A(G169), .B1(new_n366), .B2(new_n371), .ZN(new_n393));
  OAI211_X1 g0193(.A(new_n373), .B(G179), .C1(new_n375), .C2(new_n256), .ZN(new_n394));
  AOI22_X1  g0194(.A1(new_n385), .A2(new_n386), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT18), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n393), .A2(new_n394), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  OAI21_X1  g0199(.A(KEYINPUT18), .B1(new_n365), .B2(new_n399), .ZN(new_n400));
  AND2_X1   g0200(.A1(new_n397), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n392), .A2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(KEYINPUT77), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n329), .A2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT13), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n303), .B1(G238), .B2(new_n304), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n260), .A2(G232), .A3(G1698), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n260), .A2(G226), .A3(new_n261), .ZN(new_n409));
  NAND2_X1  g0209(.A1(G33), .A2(G97), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n408), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(new_n246), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n406), .B1(new_n407), .B2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n407), .A2(new_n406), .A3(new_n412), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT72), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT14), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n416), .A2(new_n417), .A3(new_n418), .A4(G169), .ZN(new_n419));
  INV_X1    g0219(.A(new_n415), .ZN(new_n420));
  OAI211_X1 g0220(.A(new_n417), .B(G169), .C1(new_n420), .C2(new_n413), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(KEYINPUT14), .ZN(new_n422));
  OR2_X1    g0222(.A1(new_n413), .A2(KEYINPUT71), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n413), .A2(KEYINPUT71), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n423), .A2(G179), .A3(new_n424), .A4(new_n415), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n419), .A2(new_n422), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n205), .A2(G20), .ZN(new_n427));
  OAI221_X1 g0227(.A(new_n427), .B1(new_n274), .B2(new_n263), .C1(new_n277), .C2(new_n280), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(new_n272), .ZN(new_n429));
  XNOR2_X1  g0229(.A(new_n429), .B(KEYINPUT11), .ZN(new_n430));
  INV_X1    g0230(.A(new_n289), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(new_n205), .ZN(new_n432));
  XNOR2_X1  g0232(.A(new_n432), .B(KEYINPUT12), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n283), .A2(G68), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n430), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n426), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n435), .B1(new_n416), .B2(G200), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n423), .A2(G190), .A3(new_n424), .A4(new_n415), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  OAI211_X1 g0239(.A(new_n436), .B(new_n439), .C1(new_n403), .C2(KEYINPUT77), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n405), .A2(new_n440), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n260), .A2(KEYINPUT4), .A3(G244), .A4(new_n261), .ZN(new_n442));
  NAND2_X1  g0242(.A1(G33), .A2(G283), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n260), .A2(G250), .A3(G1698), .ZN(new_n444));
  AND3_X1   g0244(.A1(new_n442), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n361), .A2(G244), .A3(new_n261), .A4(new_n309), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT4), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n445), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(new_n246), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n286), .A2(new_n288), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n451), .A2(new_n250), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT78), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT5), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n453), .B1(new_n454), .B2(G41), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n249), .A2(KEYINPUT78), .A3(KEYINPUT5), .ZN(new_n456));
  AOI22_X1  g0256(.A1(new_n455), .A2(new_n456), .B1(new_n454), .B2(G41), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n248), .A2(new_n452), .A3(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n246), .B1(new_n452), .B2(new_n457), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n459), .B1(G257), .B2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT79), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n450), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n460), .A2(G257), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(new_n458), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n256), .B1(new_n445), .B2(new_n448), .ZN(new_n466));
  OAI21_X1  g0266(.A(KEYINPUT79), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n463), .A2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(G169), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n465), .A2(new_n466), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(new_n300), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n306), .A2(KEYINPUT6), .A3(G97), .ZN(new_n473));
  INV_X1    g0273(.A(G97), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n474), .A2(new_n306), .ZN(new_n475));
  NOR2_X1   g0275(.A1(G97), .A2(G107), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n473), .B1(new_n477), .B2(KEYINPUT6), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n478), .A2(G20), .B1(G77), .B2(new_n276), .ZN(new_n479));
  OAI21_X1  g0279(.A(G107), .B1(new_n340), .B2(new_n341), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n333), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT80), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n289), .A2(G97), .ZN(new_n484));
  OAI211_X1 g0284(.A(new_n289), .B(new_n333), .C1(new_n308), .C2(new_n451), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n484), .B1(new_n486), .B2(G97), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n482), .A2(new_n483), .A3(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(new_n487), .ZN(new_n489));
  OAI21_X1  g0289(.A(KEYINPUT80), .B1(new_n489), .B2(new_n481), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n470), .A2(new_n472), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n482), .A2(new_n487), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  OAI21_X1  g0294(.A(G200), .B1(new_n465), .B2(new_n466), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n494), .B(new_n495), .C1(new_n468), .C2(new_n374), .ZN(new_n496));
  INV_X1    g0296(.A(new_n319), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n497), .A2(new_n289), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n337), .A2(new_n338), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n354), .B1(new_n499), .B2(G33), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n500), .A2(new_n223), .A3(G68), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT19), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n502), .B1(new_n274), .B2(new_n474), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n223), .B1(new_n410), .B2(new_n502), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n476), .A2(new_n207), .ZN(new_n505));
  AOI22_X1  g0305(.A1(new_n503), .A2(KEYINPUT82), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n501), .B(new_n506), .C1(KEYINPUT82), .C2(new_n503), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n498), .B1(new_n507), .B2(new_n272), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n508), .B1(new_n319), .B2(new_n485), .ZN(new_n509));
  INV_X1    g0309(.A(new_n452), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n246), .B1(new_n510), .B2(new_n208), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n452), .A2(new_n247), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n261), .A2(G238), .ZN(new_n514));
  INV_X1    g0314(.A(G116), .ZN(new_n515));
  OAI22_X1  g0315(.A1(new_n362), .A2(new_n514), .B1(new_n308), .B2(new_n515), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n361), .A2(G244), .A3(G1698), .A4(new_n309), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT81), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n500), .A2(KEYINPUT81), .A3(G244), .A4(G1698), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n516), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n513), .B1(new_n521), .B2(new_n256), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(new_n469), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n509), .B(new_n523), .C1(G179), .C2(new_n522), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n522), .A2(G200), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n485), .A2(new_n207), .ZN(new_n526));
  AOI211_X1 g0326(.A(new_n498), .B(new_n526), .C1(new_n507), .C2(new_n272), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n525), .B(new_n527), .C1(new_n374), .C2(new_n522), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n492), .A2(new_n496), .A3(new_n524), .A4(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT21), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n460), .A2(G270), .ZN(new_n532));
  MUX2_X1   g0332(.A(G257), .B(G264), .S(G1698), .Z(new_n533));
  AOI22_X1  g0333(.A1(new_n500), .A2(new_n533), .B1(G303), .B2(new_n312), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n532), .B(new_n458), .C1(new_n256), .C2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(new_n535), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n443), .B(new_n223), .C1(G33), .C2(new_n474), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n537), .B(new_n272), .C1(new_n223), .C2(G116), .ZN(new_n538));
  XNOR2_X1  g0338(.A(new_n538), .B(KEYINPUT20), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n431), .A2(new_n515), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n540), .B1(new_n485), .B2(new_n515), .ZN(new_n541));
  OAI21_X1  g0341(.A(G169), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n531), .B1(new_n536), .B2(new_n542), .ZN(new_n543));
  OR2_X1    g0343(.A1(new_n539), .A2(new_n541), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n536), .A2(new_n544), .A3(G179), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n544), .A2(new_n535), .A3(KEYINPUT21), .A4(G169), .ZN(new_n546));
  AND3_X1   g0346(.A1(new_n543), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n535), .A2(G200), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT83), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n539), .A2(new_n541), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n551), .B1(new_n374), .B2(new_n535), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n549), .B1(new_n548), .B2(new_n550), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n547), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n460), .A2(G264), .ZN(new_n555));
  MUX2_X1   g0355(.A(G250), .B(G257), .S(G1698), .Z(new_n556));
  AOI22_X1  g0356(.A1(new_n500), .A2(new_n556), .B1(G33), .B2(G294), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n555), .B(new_n458), .C1(new_n256), .C2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(new_n469), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n559), .B1(G179), .B2(new_n558), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT24), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n500), .A2(new_n223), .A3(G87), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(KEYINPUT22), .ZN(new_n563));
  XOR2_X1   g0363(.A(KEYINPUT84), .B(KEYINPUT22), .Z(new_n564));
  NOR4_X1   g0364(.A1(new_n564), .A2(new_n312), .A3(G20), .A4(new_n207), .ZN(new_n565));
  INV_X1    g0365(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n563), .A2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT23), .ZN(new_n568));
  OAI22_X1  g0368(.A1(KEYINPUT85), .A2(new_n568), .B1(new_n223), .B2(G107), .ZN(new_n569));
  AND2_X1   g0369(.A1(new_n568), .A2(KEYINPUT85), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT86), .ZN(new_n571));
  OR3_X1    g0371(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n571), .B1(new_n569), .B2(new_n570), .ZN(new_n573));
  NOR3_X1   g0373(.A1(new_n308), .A2(new_n515), .A3(G20), .ZN(new_n574));
  NOR3_X1   g0374(.A1(new_n223), .A2(KEYINPUT23), .A3(G107), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n572), .A2(new_n573), .A3(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n561), .B1(new_n567), .B2(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n565), .B1(KEYINPUT22), .B2(new_n562), .ZN(new_n580));
  NOR3_X1   g0380(.A1(new_n580), .A2(KEYINPUT24), .A3(new_n577), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n272), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT25), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n583), .B1(new_n289), .B2(G107), .ZN(new_n584));
  INV_X1    g0384(.A(new_n584), .ZN(new_n585));
  NOR3_X1   g0385(.A1(new_n289), .A2(new_n583), .A3(G107), .ZN(new_n586));
  OAI22_X1  g0386(.A1(new_n585), .A2(new_n586), .B1(new_n306), .B2(new_n485), .ZN(new_n587));
  INV_X1    g0387(.A(new_n587), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n560), .B1(new_n582), .B2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(new_n558), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(G190), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n558), .A2(G200), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n582), .A2(new_n588), .A3(new_n591), .A4(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  NOR3_X1   g0394(.A1(new_n554), .A2(new_n589), .A3(new_n594), .ZN(new_n595));
  AND3_X1   g0395(.A1(new_n441), .A2(new_n530), .A3(new_n595), .ZN(G372));
  NAND3_X1  g0396(.A1(new_n543), .A2(new_n546), .A3(new_n545), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n593), .B1(new_n589), .B2(new_n597), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n524), .B1(new_n529), .B2(new_n598), .ZN(new_n599));
  AND2_X1   g0399(.A1(new_n524), .A2(new_n528), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT26), .ZN(new_n601));
  AOI22_X1  g0401(.A1(new_n468), .A2(new_n469), .B1(new_n300), .B2(new_n471), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n600), .A2(new_n601), .A3(new_n602), .A4(new_n493), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n602), .A2(new_n491), .A3(new_n524), .A4(new_n528), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(KEYINPUT26), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n441), .B1(new_n599), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n296), .A2(new_n299), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT88), .ZN(new_n609));
  XNOR2_X1  g0409(.A(new_n608), .B(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(new_n439), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n436), .B1(new_n611), .B2(new_n324), .ZN(new_n612));
  AND2_X1   g0412(.A1(new_n612), .A2(new_n392), .ZN(new_n613));
  AND3_X1   g0413(.A1(new_n397), .A2(KEYINPUT87), .A3(new_n400), .ZN(new_n614));
  AOI21_X1  g0414(.A(KEYINPUT87), .B1(new_n397), .B2(new_n400), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(new_n616), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n610), .B1(new_n613), .B2(new_n617), .ZN(new_n618));
  AND2_X1   g0418(.A1(new_n618), .A2(new_n302), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n607), .A2(new_n619), .ZN(G369));
  INV_X1    g0420(.A(KEYINPUT91), .ZN(new_n621));
  INV_X1    g0421(.A(G13), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n622), .A2(G20), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n253), .A2(new_n623), .ZN(new_n624));
  OR2_X1    g0424(.A1(new_n624), .A2(KEYINPUT27), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(KEYINPUT27), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n625), .A2(G213), .A3(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(G343), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n544), .A2(new_n629), .ZN(new_n630));
  OAI211_X1 g0430(.A(new_n547), .B(new_n630), .C1(new_n552), .C2(new_n553), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT89), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n597), .A2(new_n544), .A3(new_n629), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n631), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n632), .B1(new_n631), .B2(new_n633), .ZN(new_n636));
  OAI21_X1  g0436(.A(G330), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n590), .A2(new_n300), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n567), .A2(new_n561), .A3(new_n578), .ZN(new_n639));
  OAI21_X1  g0439(.A(KEYINPUT24), .B1(new_n580), .B2(new_n577), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n333), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  OAI211_X1 g0441(.A(new_n559), .B(new_n638), .C1(new_n641), .C2(new_n587), .ZN(new_n642));
  INV_X1    g0442(.A(new_n629), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n629), .B1(new_n641), .B2(new_n587), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n642), .A2(new_n593), .A3(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT90), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n642), .A2(new_n593), .A3(KEYINPUT90), .A4(new_n645), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n644), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n621), .B1(new_n637), .B2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(G330), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n631), .A2(new_n633), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(KEYINPUT89), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n652), .B1(new_n654), .B2(new_n634), .ZN(new_n655));
  INV_X1    g0455(.A(new_n650), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n655), .A2(KEYINPUT91), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n651), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n589), .A2(new_n643), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n547), .A2(new_n629), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n648), .A2(new_n649), .A3(new_n660), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n658), .A2(new_n659), .A3(new_n661), .ZN(G399));
  INV_X1    g0462(.A(new_n218), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n663), .A2(G41), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n505), .A2(G116), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n665), .A2(G1), .A3(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n667), .B1(new_n225), .B2(new_n665), .ZN(new_n668));
  XNOR2_X1  g0468(.A(new_n668), .B(KEYINPUT28), .ZN(new_n669));
  INV_X1    g0469(.A(new_n599), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT94), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n604), .A2(new_n671), .A3(new_n601), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n600), .A2(new_n602), .A3(new_n493), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n672), .B1(new_n673), .B2(new_n601), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n671), .B1(new_n604), .B2(new_n601), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n670), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n676), .A2(KEYINPUT29), .A3(new_n643), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n643), .B1(new_n606), .B2(new_n599), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT29), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  AND2_X1   g0481(.A1(new_n500), .A2(new_n533), .ZN(new_n682));
  INV_X1    g0482(.A(G303), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n260), .A2(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n246), .B1(new_n682), .B2(new_n684), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n685), .A2(G179), .A3(new_n458), .A4(new_n532), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n555), .B1(new_n256), .B2(new_n557), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n522), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n688), .A2(new_n689), .A3(new_n467), .A4(new_n463), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT30), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n558), .A2(new_n535), .A3(new_n300), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n692), .A2(new_n471), .ZN(new_n693));
  AOI22_X1  g0493(.A1(new_n690), .A2(new_n691), .B1(new_n522), .B2(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(KEYINPUT92), .B1(new_n690), .B2(new_n691), .ZN(new_n695));
  INV_X1    g0495(.A(new_n468), .ZN(new_n696));
  NOR3_X1   g0496(.A1(new_n522), .A2(new_n686), .A3(new_n687), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT92), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n696), .A2(new_n697), .A3(new_n698), .A4(KEYINPUT30), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n694), .A2(new_n695), .A3(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(new_n629), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT31), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT93), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n701), .A2(KEYINPUT93), .A3(new_n702), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n700), .A2(KEYINPUT31), .A3(new_n629), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n595), .A2(new_n530), .A3(new_n643), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n705), .A2(new_n706), .A3(new_n707), .A4(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(G330), .ZN(new_n710));
  AND2_X1   g0510(.A1(new_n681), .A2(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n669), .B1(new_n711), .B2(G1), .ZN(G364));
  OAI21_X1  g0512(.A(G20), .B1(KEYINPUT95), .B2(G169), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(KEYINPUT95), .A2(G169), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n222), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(G20), .A2(G179), .ZN(new_n718));
  NOR3_X1   g0518(.A1(new_n718), .A2(G190), .A3(G200), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NOR3_X1   g0520(.A1(new_n718), .A2(new_n374), .A3(G200), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  OAI221_X1 g0522(.A(new_n260), .B1(new_n720), .B2(new_n263), .C1(new_n343), .C2(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n223), .A2(G179), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n724), .A2(new_n374), .A3(G200), .ZN(new_n725));
  INV_X1    g0525(.A(new_n718), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n726), .A2(G190), .A3(G200), .ZN(new_n727));
  OAI22_X1  g0527(.A1(new_n725), .A2(new_n306), .B1(new_n727), .B2(new_n280), .ZN(new_n728));
  NOR3_X1   g0528(.A1(new_n374), .A2(G179), .A3(G200), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(new_n223), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n726), .A2(new_n374), .A3(G200), .ZN(new_n731));
  OAI22_X1  g0531(.A1(new_n730), .A2(new_n474), .B1(new_n731), .B2(new_n205), .ZN(new_n732));
  NOR3_X1   g0532(.A1(new_n723), .A2(new_n728), .A3(new_n732), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n724), .A2(G190), .A3(G200), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n734), .A2(new_n207), .ZN(new_n735));
  NOR2_X1   g0535(.A1(G190), .A2(G200), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n724), .A2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(G159), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n735), .B1(new_n739), .B2(KEYINPUT32), .ZN(new_n740));
  OAI211_X1 g0540(.A(new_n733), .B(new_n740), .C1(KEYINPUT32), .C2(new_n739), .ZN(new_n741));
  INV_X1    g0541(.A(G322), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n722), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(G311), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n312), .B1(new_n720), .B2(new_n744), .ZN(new_n745));
  AOI211_X1 g0545(.A(new_n743), .B(new_n745), .C1(G329), .C2(new_n738), .ZN(new_n746));
  INV_X1    g0546(.A(new_n727), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(G326), .ZN(new_n748));
  INV_X1    g0548(.A(new_n734), .ZN(new_n749));
  INV_X1    g0549(.A(new_n731), .ZN(new_n750));
  XNOR2_X1  g0550(.A(KEYINPUT33), .B(G317), .ZN(new_n751));
  AOI22_X1  g0551(.A1(G303), .A2(new_n749), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n730), .ZN(new_n753));
  INV_X1    g0553(.A(new_n725), .ZN(new_n754));
  AOI22_X1  g0554(.A1(new_n753), .A2(G294), .B1(new_n754), .B2(G283), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n746), .A2(new_n748), .A3(new_n752), .A4(new_n755), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n717), .B1(new_n741), .B2(new_n756), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n285), .B1(new_n623), .B2(G45), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n664), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n663), .A2(new_n312), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(G355), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n762), .B1(G116), .B2(new_n218), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n500), .A2(new_n663), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n765), .B1(new_n250), .B2(new_n226), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n244), .A2(G45), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n763), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(G13), .A2(G33), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(G20), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n716), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n760), .B1(new_n768), .B2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n757), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n654), .A2(new_n634), .ZN(new_n776));
  INV_X1    g0576(.A(new_n771), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n775), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n760), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n637), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n776), .A2(G330), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n778), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  AND2_X1   g0582(.A1(new_n782), .A2(KEYINPUT96), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n782), .A2(KEYINPUT96), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(G396));
  NAND2_X1  g0586(.A1(new_n629), .A2(new_n323), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n326), .A2(new_n787), .ZN(new_n788));
  AND2_X1   g0588(.A1(new_n788), .A2(new_n324), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n324), .A2(new_n629), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n678), .A2(new_n792), .ZN(new_n793));
  OAI211_X1 g0593(.A(new_n643), .B(new_n791), .C1(new_n606), .C2(new_n599), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  OR2_X1    g0595(.A1(new_n710), .A2(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n760), .B1(new_n710), .B2(new_n795), .ZN(new_n797));
  AND2_X1   g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(G283), .ZN(new_n799));
  OAI22_X1  g0599(.A1(new_n734), .A2(new_n306), .B1(new_n731), .B2(new_n799), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n800), .B1(G87), .B2(new_n754), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n260), .B1(new_n719), .B2(G116), .ZN(new_n802));
  AOI22_X1  g0602(.A1(new_n738), .A2(G311), .B1(G294), .B2(new_n721), .ZN(new_n803));
  AOI22_X1  g0603(.A1(new_n753), .A2(G97), .B1(new_n747), .B2(G303), .ZN(new_n804));
  NAND4_X1  g0604(.A1(new_n801), .A2(new_n802), .A3(new_n803), .A4(new_n804), .ZN(new_n805));
  AOI22_X1  g0605(.A1(G143), .A2(new_n721), .B1(new_n719), .B2(G159), .ZN(new_n806));
  INV_X1    g0606(.A(G137), .ZN(new_n807));
  OAI221_X1 g0607(.A(new_n806), .B1(new_n807), .B2(new_n727), .C1(new_n275), .C2(new_n731), .ZN(new_n808));
  XNOR2_X1  g0608(.A(new_n808), .B(KEYINPUT34), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(KEYINPUT97), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n725), .A2(new_n205), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n811), .B1(G58), .B2(new_n753), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n812), .B1(new_n280), .B2(new_n734), .ZN(new_n813));
  AOI211_X1 g0613(.A(new_n362), .B(new_n813), .C1(G132), .C2(new_n738), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n810), .A2(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n809), .A2(KEYINPUT97), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n805), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(new_n716), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n716), .A2(new_n769), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n779), .B1(new_n819), .B2(new_n263), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n821), .B1(new_n769), .B2(new_n792), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n798), .A2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(G384));
  NOR2_X1   g0624(.A1(new_n253), .A2(new_n623), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n617), .A2(new_n627), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n385), .A2(new_n386), .ZN(new_n827));
  AOI21_X1  g0627(.A(KEYINPUT37), .B1(new_n827), .B2(new_n398), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n627), .B1(new_n385), .B2(new_n386), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  NAND4_X1  g0630(.A1(new_n828), .A2(new_n388), .A3(new_n830), .A4(new_n390), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n831), .A2(KEYINPUT101), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n389), .B1(new_n365), .B2(new_n377), .ZN(new_n833));
  AND4_X1   g0633(.A1(new_n389), .A2(new_n385), .A3(new_n386), .A4(new_n377), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NOR3_X1   g0635(.A1(new_n395), .A2(new_n829), .A3(KEYINPUT37), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT101), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n835), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n832), .A2(new_n838), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n348), .B1(new_n356), .B2(new_n363), .ZN(new_n840));
  NOR2_X1   g0640(.A1(KEYINPUT100), .A2(KEYINPUT16), .ZN(new_n841));
  AND2_X1   g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n272), .B1(new_n840), .B2(new_n841), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n331), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n627), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n844), .B1(new_n398), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n835), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n847), .A2(KEYINPUT37), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n839), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n844), .A2(new_n845), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n850), .B1(new_n392), .B2(new_n401), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n849), .A2(new_n852), .A3(KEYINPUT38), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT38), .ZN(new_n854));
  AOI22_X1  g0654(.A1(new_n832), .A2(new_n838), .B1(new_n847), .B2(KEYINPUT37), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n854), .B1(new_n855), .B2(new_n851), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n853), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n435), .A2(new_n629), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n436), .A2(new_n439), .A3(new_n858), .ZN(new_n859));
  OAI211_X1 g0659(.A(new_n435), .B(new_n629), .C1(new_n611), .C2(new_n426), .ZN(new_n860));
  AND2_X1   g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n790), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n861), .B1(new_n794), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n857), .B1(new_n863), .B2(KEYINPUT99), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT99), .ZN(new_n865));
  AOI211_X1 g0665(.A(new_n865), .B(new_n861), .C1(new_n862), .C2(new_n794), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n826), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n853), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n868), .A2(KEYINPUT39), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n831), .A2(KEYINPUT101), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n837), .B1(new_n835), .B2(new_n836), .ZN(new_n871));
  OAI21_X1  g0671(.A(KEYINPUT103), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT103), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n832), .A2(new_n838), .A3(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT37), .ZN(new_n875));
  OAI21_X1  g0675(.A(KEYINPUT87), .B1(new_n365), .B2(new_n399), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT87), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n827), .A2(new_n877), .A3(new_n398), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n365), .A2(KEYINPUT102), .A3(new_n377), .ZN(new_n879));
  AND3_X1   g0679(.A1(new_n876), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT102), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n829), .B1(new_n881), .B2(new_n387), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n875), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n872), .A2(new_n874), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n830), .B1(new_n616), .B2(new_n392), .ZN(new_n886));
  INV_X1    g0686(.A(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(KEYINPUT104), .B1(new_n888), .B2(new_n854), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT104), .ZN(new_n890));
  AOI211_X1 g0690(.A(new_n890), .B(KEYINPUT38), .C1(new_n885), .C2(new_n887), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n869), .B1(new_n889), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n857), .A2(KEYINPUT39), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n436), .A2(new_n629), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n867), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n441), .A2(new_n680), .A3(new_n677), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(new_n619), .ZN(new_n898));
  XOR2_X1   g0698(.A(new_n896), .B(new_n898), .Z(new_n899));
  NOR2_X1   g0699(.A1(new_n861), .A2(new_n792), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT105), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n707), .A2(new_n901), .ZN(new_n902));
  NAND4_X1  g0702(.A1(new_n700), .A2(KEYINPUT105), .A3(KEYINPUT31), .A4(new_n629), .ZN(new_n903));
  NAND4_X1  g0703(.A1(new_n902), .A2(new_n708), .A3(new_n703), .A4(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n900), .A2(KEYINPUT40), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n883), .B1(new_n839), .B2(KEYINPUT103), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n886), .B1(new_n906), .B2(new_n874), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n890), .B1(new_n907), .B2(KEYINPUT38), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n888), .A2(KEYINPUT104), .A3(new_n854), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n905), .B1(new_n910), .B2(new_n853), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT40), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n900), .A2(new_n857), .A3(new_n904), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n911), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  AND2_X1   g0714(.A1(new_n441), .A2(new_n904), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n652), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n916), .B1(new_n914), .B2(new_n915), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n825), .B1(new_n899), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n918), .B1(new_n899), .B2(new_n917), .ZN(new_n919));
  OR2_X1    g0719(.A1(new_n478), .A2(KEYINPUT35), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n478), .A2(KEYINPUT35), .ZN(new_n921));
  NAND4_X1  g0721(.A1(new_n920), .A2(G116), .A3(new_n224), .A4(new_n921), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n922), .B(KEYINPUT36), .ZN(new_n923));
  NOR3_X1   g0723(.A1(new_n344), .A2(new_n225), .A3(new_n263), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT98), .ZN(new_n925));
  AOI22_X1  g0725(.A1(new_n924), .A2(new_n925), .B1(new_n280), .B2(G68), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n926), .B1(new_n925), .B2(new_n924), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n927), .A2(new_n622), .A3(new_n451), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n919), .A2(new_n923), .A3(new_n928), .ZN(new_n929));
  XOR2_X1   g0729(.A(new_n929), .B(KEYINPUT106), .Z(G367));
  INV_X1    g0730(.A(new_n661), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n493), .A2(new_n629), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n602), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n492), .A2(new_n496), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n933), .B1(new_n934), .B2(new_n932), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n931), .A2(new_n935), .ZN(new_n936));
  OR2_X1    g0736(.A1(new_n936), .A2(KEYINPUT42), .ZN(new_n937));
  INV_X1    g0737(.A(new_n935), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n492), .B1(new_n938), .B2(new_n642), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(new_n643), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n936), .A2(KEYINPUT42), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n937), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  OR2_X1    g0742(.A1(new_n527), .A2(new_n643), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n600), .A2(new_n943), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n524), .A2(new_n943), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT43), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n946), .A2(KEYINPUT43), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n942), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n658), .A2(new_n938), .ZN(new_n952));
  AND2_X1   g0752(.A1(new_n941), .A2(new_n940), .ZN(new_n953));
  NAND4_X1  g0753(.A1(new_n953), .A2(new_n948), .A3(new_n947), .A4(new_n937), .ZN(new_n954));
  AND3_X1   g0754(.A1(new_n951), .A2(new_n952), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n952), .B1(new_n951), .B2(new_n954), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  XOR2_X1   g0757(.A(new_n664), .B(KEYINPUT41), .Z(new_n958));
  NAND2_X1  g0758(.A1(new_n661), .A2(new_n659), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(new_n938), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT44), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n959), .A2(KEYINPUT44), .A3(new_n938), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT45), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(new_n959), .B2(new_n938), .ZN(new_n966));
  NAND4_X1  g0766(.A1(new_n661), .A2(KEYINPUT45), .A3(new_n659), .A4(new_n935), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n964), .A2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(new_n658), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT107), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n969), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  AOI22_X1  g0772(.A1(new_n962), .A2(new_n963), .B1(new_n966), .B2(new_n967), .ZN(new_n973));
  OAI21_X1  g0773(.A(KEYINPUT107), .B1(new_n973), .B2(new_n658), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n650), .B1(new_n547), .B2(new_n629), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n637), .A2(new_n975), .A3(new_n661), .ZN(new_n976));
  AOI211_X1 g0776(.A(new_n644), .B(new_n660), .C1(new_n648), .C2(new_n649), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n655), .B1(new_n977), .B2(new_n931), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  AND3_X1   g0779(.A1(new_n681), .A2(new_n710), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n973), .A2(new_n658), .ZN(new_n981));
  NAND4_X1  g0781(.A1(new_n972), .A2(new_n974), .A3(new_n980), .A4(new_n981), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n958), .B1(new_n982), .B2(new_n711), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n957), .B1(new_n983), .B2(new_n759), .ZN(new_n984));
  OAI221_X1 g0784(.A(new_n772), .B1(new_n218), .B2(new_n319), .C1(new_n765), .C2(new_n236), .ZN(new_n985));
  AND2_X1   g0785(.A1(new_n985), .A2(new_n760), .ZN(new_n986));
  INV_X1    g0786(.A(G159), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n734), .A2(new_n343), .B1(new_n731), .B2(new_n987), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n988), .B1(G68), .B2(new_n753), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n312), .B1(new_n738), .B2(G137), .ZN(new_n990));
  AOI22_X1  g0790(.A1(G50), .A2(new_n719), .B1(new_n721), .B2(G150), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n725), .A2(new_n263), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n992), .B1(G143), .B2(new_n747), .ZN(new_n993));
  NAND4_X1  g0793(.A1(new_n989), .A2(new_n990), .A3(new_n991), .A4(new_n993), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n730), .A2(new_n306), .B1(new_n720), .B2(new_n799), .ZN(new_n995));
  OR2_X1    g0795(.A1(new_n995), .A2(KEYINPUT108), .ZN(new_n996));
  INV_X1    g0796(.A(G294), .ZN(new_n997));
  OAI22_X1  g0797(.A1(new_n997), .A2(new_n731), .B1(new_n727), .B2(new_n744), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n998), .B1(G97), .B2(new_n754), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n995), .A2(KEYINPUT108), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n996), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(new_n738), .A2(G317), .B1(G303), .B2(new_n721), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n749), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT46), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1004), .B1(new_n734), .B2(new_n515), .ZN(new_n1005));
  NAND4_X1  g0805(.A1(new_n1002), .A2(new_n1003), .A3(new_n362), .A4(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n994), .B1(new_n1001), .B2(new_n1006), .ZN(new_n1007));
  XOR2_X1   g0807(.A(new_n1007), .B(KEYINPUT47), .Z(new_n1008));
  OAI221_X1 g0808(.A(new_n986), .B1(new_n717), .B2(new_n1008), .C1(new_n946), .C2(new_n777), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n984), .A2(new_n1009), .ZN(G387));
  INV_X1    g0810(.A(new_n666), .ZN(new_n1011));
  AOI211_X1 g0811(.A(G45), .B(new_n1011), .C1(G68), .C2(G77), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n273), .A2(G50), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1013), .B(KEYINPUT50), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n765), .B1(new_n1012), .B2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1015), .B1(new_n233), .B2(new_n250), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n1011), .A2(new_n761), .B1(new_n306), .B2(new_n663), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n1018), .A2(KEYINPUT109), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1018), .A2(KEYINPUT109), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1020), .A2(new_n772), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n722), .A2(new_n280), .B1(new_n720), .B2(new_n205), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1022), .B1(G150), .B2(new_n738), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n730), .A2(new_n319), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1024), .B1(G159), .B2(new_n747), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n273), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(G77), .A2(new_n749), .B1(new_n750), .B2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n362), .B1(G97), .B2(new_n754), .ZN(new_n1028));
  NAND4_X1  g0828(.A1(new_n1023), .A2(new_n1025), .A3(new_n1027), .A4(new_n1028), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(G303), .A2(new_n719), .B1(new_n721), .B2(G317), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n1030), .B1(new_n744), .B2(new_n731), .C1(new_n742), .C2(new_n727), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT48), .ZN(new_n1032));
  AND2_X1   g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1034));
  OAI22_X1  g0834(.A1(new_n730), .A2(new_n799), .B1(new_n734), .B2(new_n997), .ZN(new_n1035));
  NOR3_X1   g0835(.A1(new_n1033), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1036), .A2(KEYINPUT49), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n754), .A2(G116), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n500), .B1(G326), .B2(new_n738), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1037), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n1036), .A2(KEYINPUT49), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1029), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  XOR2_X1   g0842(.A(new_n1042), .B(KEYINPUT110), .Z(new_n1043));
  OAI221_X1 g0843(.A(new_n760), .B1(new_n1019), .B2(new_n1021), .C1(new_n1043), .C2(new_n717), .ZN(new_n1044));
  XOR2_X1   g0844(.A(new_n1044), .B(KEYINPUT111), .Z(new_n1045));
  NAND2_X1  g0845(.A1(new_n650), .A2(new_n771), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n1045), .A2(new_n1046), .B1(new_n759), .B2(new_n979), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n711), .A2(new_n979), .ZN(new_n1048));
  OR2_X1    g0848(.A1(new_n980), .A2(new_n665), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1047), .B1(new_n1048), .B2(new_n1049), .ZN(G393));
  XNOR2_X1  g0850(.A(new_n970), .B(new_n973), .ZN(new_n1051));
  OAI211_X1 g0851(.A(new_n982), .B(new_n664), .C1(new_n1051), .C2(new_n980), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n938), .A2(new_n771), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n312), .B1(new_n737), .B2(new_n742), .C1(new_n306), .C2(new_n725), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(G283), .B2(new_n749), .ZN(new_n1055));
  XOR2_X1   g0855(.A(new_n1055), .B(KEYINPUT112), .Z(new_n1056));
  AOI22_X1  g0856(.A1(new_n747), .A2(G317), .B1(G311), .B2(new_n721), .ZN(new_n1057));
  XOR2_X1   g0857(.A(new_n1057), .B(KEYINPUT52), .Z(new_n1058));
  OAI22_X1  g0858(.A1(new_n730), .A2(new_n515), .B1(new_n720), .B2(new_n997), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1059), .B1(G303), .B2(new_n750), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n1056), .A2(new_n1058), .A3(new_n1060), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n722), .A2(new_n987), .B1(new_n727), .B2(new_n275), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1062), .B(KEYINPUT51), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(G143), .A2(new_n738), .B1(new_n1026), .B2(new_n719), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n730), .A2(new_n263), .B1(new_n731), .B2(new_n280), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n205), .A2(new_n734), .B1(new_n725), .B2(new_n207), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NAND4_X1  g0867(.A1(new_n1063), .A2(new_n500), .A3(new_n1064), .A4(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n717), .B1(new_n1061), .B2(new_n1068), .ZN(new_n1069));
  OR2_X1    g0869(.A1(new_n241), .A2(new_n765), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n773), .B1(G97), .B2(new_n663), .ZN(new_n1071));
  AOI211_X1 g0871(.A(new_n779), .B(new_n1069), .C1(new_n1070), .C2(new_n1071), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n1051), .A2(new_n759), .B1(new_n1053), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1052), .A2(new_n1073), .ZN(G390));
  NAND2_X1  g0874(.A1(new_n904), .A2(G330), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n441), .A2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n897), .A2(new_n1077), .A3(new_n619), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1078), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n709), .A2(G330), .A3(new_n791), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1080), .A2(new_n861), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1076), .A2(new_n900), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n1081), .A2(new_n1082), .B1(new_n862), .B2(new_n794), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n861), .B1(new_n1075), .B2(new_n792), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n789), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n676), .A2(new_n643), .A3(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1086), .A2(new_n862), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n861), .ZN(new_n1089));
  NAND4_X1  g0889(.A1(new_n709), .A2(G330), .A3(new_n1089), .A4(new_n791), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1084), .A2(new_n1088), .A3(new_n1090), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1091), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1079), .B1(new_n1083), .B2(new_n1092), .ZN(new_n1093));
  OR2_X1    g0893(.A1(new_n863), .A2(new_n895), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n892), .A2(new_n893), .A3(new_n1094), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n853), .B1(new_n889), .B2(new_n891), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n895), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1096), .A2(new_n1097), .A3(new_n1098), .ZN(new_n1099));
  AND3_X1   g0899(.A1(new_n1095), .A2(new_n1099), .A3(new_n1090), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1082), .B1(new_n1095), .B2(new_n1099), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1093), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1095), .A2(new_n1099), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1082), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n794), .A2(new_n862), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1078), .B1(new_n1108), .B2(new_n1091), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1095), .A2(new_n1099), .A3(new_n1090), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1105), .A2(new_n1109), .A3(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1102), .A2(new_n1111), .A3(new_n664), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n894), .A2(new_n770), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(KEYINPUT54), .B(G143), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n720), .A2(new_n1114), .B1(new_n731), .B2(new_n807), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n1115), .A2(KEYINPUT113), .B1(G159), .B2(new_n753), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1116), .B1(KEYINPUT113), .B2(new_n1115), .ZN(new_n1117));
  XOR2_X1   g0917(.A(new_n1117), .B(KEYINPUT114), .Z(new_n1118));
  NAND2_X1  g0918(.A1(new_n749), .A2(G150), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(new_n1119), .B(KEYINPUT53), .ZN(new_n1120));
  INV_X1    g0920(.A(G125), .ZN(new_n1121));
  INV_X1    g0921(.A(G132), .ZN(new_n1122));
  OAI221_X1 g0922(.A(new_n260), .B1(new_n737), .B2(new_n1121), .C1(new_n722), .C2(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(G128), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n725), .A2(new_n280), .B1(new_n727), .B2(new_n1124), .ZN(new_n1125));
  OR3_X1    g0925(.A1(new_n1120), .A2(new_n1123), .A3(new_n1125), .ZN(new_n1126));
  OAI22_X1  g0926(.A1(new_n730), .A2(new_n263), .B1(new_n722), .B2(new_n515), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(new_n1127), .B(KEYINPUT115), .ZN(new_n1128));
  OAI221_X1 g0928(.A(new_n312), .B1(new_n737), .B2(new_n997), .C1(new_n720), .C2(new_n474), .ZN(new_n1129));
  OAI22_X1  g0929(.A1(new_n306), .A2(new_n731), .B1(new_n727), .B2(new_n799), .ZN(new_n1130));
  OR4_X1    g0930(.A1(new_n735), .A2(new_n1129), .A3(new_n811), .A4(new_n1130), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n1118), .A2(new_n1126), .B1(new_n1128), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT116), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n717), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1134), .B1(new_n1133), .B2(new_n1132), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n779), .B1(new_n819), .B2(new_n273), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n1113), .A2(new_n1137), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1138), .B1(new_n1139), .B2(new_n759), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1112), .A2(new_n1140), .ZN(G378));
  NAND2_X1  g0941(.A1(new_n1108), .A2(new_n1091), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1078), .B1(new_n1139), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n610), .A2(new_n302), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n290), .A2(new_n845), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1144), .A2(new_n1146), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n608), .A2(new_n609), .ZN(new_n1148));
  AOI21_X1  g0948(.A(KEYINPUT88), .B1(new_n296), .B2(new_n299), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n302), .B(new_n1145), .C1(new_n1148), .C2(new_n1149), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1147), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1151), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1145), .B1(new_n610), .B2(new_n302), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1150), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1153), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1152), .A2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n652), .B1(new_n913), .B2(new_n912), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n868), .B1(new_n908), .B2(new_n909), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n1157), .B(new_n1158), .C1(new_n1159), .C2(new_n905), .ZN(new_n1160));
  AND2_X1   g0960(.A1(new_n1152), .A2(new_n1156), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n913), .A2(new_n912), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1162), .A2(G330), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1161), .B1(new_n911), .B2(new_n1163), .ZN(new_n1164));
  AND3_X1   g0964(.A1(new_n896), .A2(new_n1160), .A3(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n894), .A2(new_n895), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n867), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n1164), .A2(new_n1160), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  OAI21_X1  g0968(.A(KEYINPUT57), .B1(new_n1165), .B2(new_n1168), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n664), .B1(new_n1143), .B2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1111), .A2(new_n1079), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1164), .A2(new_n1160), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n896), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n896), .A2(new_n1164), .A3(new_n1160), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(KEYINPUT57), .B1(new_n1171), .B2(new_n1176), .ZN(new_n1177));
  OR2_X1    g0977(.A1(new_n1170), .A2(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1114), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n749), .A2(new_n1179), .B1(G128), .B2(new_n721), .ZN(new_n1180));
  XOR2_X1   g0980(.A(new_n1180), .B(KEYINPUT119), .Z(new_n1181));
  OAI22_X1  g0981(.A1(new_n720), .A2(new_n807), .B1(new_n727), .B2(new_n1121), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n730), .A2(new_n275), .B1(new_n731), .B2(new_n1122), .ZN(new_n1183));
  OR3_X1    g0983(.A1(new_n1181), .A2(new_n1182), .A3(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1184), .A2(KEYINPUT59), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(G33), .A2(G41), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(new_n1186), .B(KEYINPUT117), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1187), .B1(G124), .B2(new_n738), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n1185), .B(new_n1188), .C1(new_n987), .C2(new_n725), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n1184), .A2(KEYINPUT59), .ZN(new_n1190));
  INV_X1    g0990(.A(KEYINPUT58), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n722), .A2(new_n306), .B1(new_n737), .B2(new_n799), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1192), .B1(new_n497), .B2(new_n719), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n725), .A2(new_n343), .B1(new_n727), .B2(new_n515), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(G97), .B2(new_n750), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n500), .A2(G41), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(new_n753), .A2(G68), .B1(new_n749), .B2(G77), .ZN(new_n1197));
  NAND4_X1  g0997(.A1(new_n1193), .A2(new_n1195), .A3(new_n1196), .A4(new_n1197), .ZN(new_n1198));
  OAI22_X1  g0998(.A1(new_n1189), .A2(new_n1190), .B1(new_n1191), .B2(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1187), .ZN(new_n1200));
  NOR3_X1   g1000(.A1(new_n1196), .A2(G50), .A3(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1201), .B1(new_n1198), .B2(new_n1191), .ZN(new_n1202));
  XOR2_X1   g1002(.A(new_n1202), .B(KEYINPUT118), .Z(new_n1203));
  OAI21_X1  g1003(.A(new_n716), .B1(new_n1199), .B2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n779), .B1(new_n819), .B2(new_n280), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n1204), .B(new_n1205), .C1(new_n1157), .C2(new_n770), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1207), .B1(new_n1176), .B2(new_n759), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1178), .A2(new_n1208), .ZN(G375));
  NAND2_X1  g1009(.A1(new_n1142), .A2(new_n759), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n861), .A2(new_n769), .ZN(new_n1211));
  XNOR2_X1  g1011(.A(new_n1211), .B(KEYINPUT121), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n779), .B1(new_n819), .B2(new_n205), .ZN(new_n1213));
  OAI22_X1  g1013(.A1(new_n734), .A2(new_n474), .B1(new_n737), .B2(new_n683), .ZN(new_n1214));
  XOR2_X1   g1014(.A(new_n1214), .B(KEYINPUT122), .Z(new_n1215));
  INV_X1    g1015(.A(new_n1215), .ZN(new_n1216));
  OAI221_X1 g1016(.A(new_n312), .B1(new_n720), .B2(new_n306), .C1(new_n799), .C2(new_n722), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n515), .A2(new_n731), .B1(new_n727), .B2(new_n997), .ZN(new_n1218));
  NOR4_X1   g1018(.A1(new_n1217), .A2(new_n1218), .A3(new_n992), .A4(new_n1024), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n722), .A2(new_n807), .B1(new_n720), .B2(new_n275), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n500), .B1(new_n343), .B2(new_n725), .ZN(new_n1221));
  AOI211_X1 g1021(.A(new_n1220), .B(new_n1221), .C1(G128), .C2(new_n738), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n731), .A2(new_n1114), .ZN(new_n1223));
  OAI22_X1  g1023(.A1(new_n730), .A2(new_n280), .B1(new_n727), .B2(new_n1122), .ZN(new_n1224));
  AOI211_X1 g1024(.A(new_n1223), .B(new_n1224), .C1(G159), .C2(new_n749), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(new_n1216), .A2(new_n1219), .B1(new_n1222), .B2(new_n1225), .ZN(new_n1226));
  OAI211_X1 g1026(.A(new_n1212), .B(new_n1213), .C1(new_n717), .C2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1210), .A2(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1108), .A2(new_n1078), .A3(new_n1091), .ZN(new_n1230));
  XOR2_X1   g1030(.A(new_n958), .B(KEYINPUT120), .Z(new_n1231));
  NAND3_X1  g1031(.A1(new_n1093), .A2(new_n1230), .A3(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1229), .A2(new_n1232), .ZN(G381));
  AND2_X1   g1033(.A1(new_n1178), .A2(new_n1208), .ZN(new_n1234));
  INV_X1    g1034(.A(G378), .ZN(new_n1235));
  INV_X1    g1035(.A(G390), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(new_n823), .ZN(new_n1237));
  OAI211_X1 g1037(.A(new_n1047), .B(new_n785), .C1(new_n1048), .C2(new_n1049), .ZN(new_n1238));
  NOR4_X1   g1038(.A1(G381), .A2(new_n1237), .A3(G387), .A4(new_n1238), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1234), .A2(new_n1235), .A3(new_n1239), .ZN(G407));
  NAND2_X1  g1040(.A1(new_n628), .A2(G213), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1234), .A2(new_n1235), .A3(new_n1242), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(G407), .A2(new_n1243), .A3(G213), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT123), .ZN(new_n1245));
  XNOR2_X1  g1045(.A(new_n1244), .B(new_n1245), .ZN(G409));
  NAND2_X1  g1046(.A1(new_n1093), .A2(KEYINPUT60), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(new_n1230), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1108), .A2(KEYINPUT60), .A3(new_n1078), .A4(new_n1091), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1249), .A2(new_n664), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1248), .A2(new_n1251), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1252), .A2(G384), .A3(new_n1229), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1250), .B1(new_n1247), .B2(new_n1230), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n823), .B1(new_n1254), .B2(new_n1228), .ZN(new_n1255));
  AND2_X1   g1055(.A1(new_n1242), .A2(G2897), .ZN(new_n1256));
  AND3_X1   g1056(.A1(new_n1253), .A2(new_n1255), .A3(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1256), .B1(new_n1253), .B2(new_n1255), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  OAI21_X1  g1059(.A(KEYINPUT124), .B1(new_n1165), .B2(new_n1168), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT124), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1174), .A2(new_n1261), .A3(new_n1175), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1260), .A2(new_n1262), .A3(new_n759), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1171), .A2(new_n1176), .A3(new_n1231), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1263), .A2(new_n1264), .A3(new_n1206), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(new_n1235), .ZN(new_n1266));
  OAI211_X1 g1066(.A(G378), .B(new_n1208), .C1(new_n1170), .C2(new_n1177), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1242), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1259), .B1(new_n1268), .B2(KEYINPUT125), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1270), .A2(new_n1241), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT125), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1269), .A2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1253), .A2(new_n1255), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1268), .A2(KEYINPUT63), .A3(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT61), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(G393), .A2(G396), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1279), .A2(new_n1238), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1280), .A2(KEYINPUT126), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT126), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1279), .A2(new_n1238), .A3(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1281), .A2(new_n1283), .ZN(new_n1284));
  AOI21_X1  g1084(.A(G390), .B1(new_n984), .B2(new_n1009), .ZN(new_n1285));
  AND3_X1   g1085(.A1(new_n984), .A2(new_n1009), .A3(G390), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT127), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1285), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n984), .A2(new_n1009), .A3(G390), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1289), .A2(KEYINPUT127), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1284), .B1(new_n1288), .B2(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1285), .ZN(new_n1292));
  AND3_X1   g1092(.A1(new_n1292), .A2(new_n1289), .A3(new_n1280), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1278), .B1(new_n1291), .B2(new_n1293), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1270), .A2(new_n1241), .A3(new_n1276), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT63), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1294), .B1(new_n1295), .B2(new_n1296), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1274), .A2(new_n1277), .A3(new_n1297), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n1295), .A2(KEYINPUT62), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1278), .B1(new_n1268), .B2(new_n1259), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT62), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1301), .B1(new_n1268), .B2(new_n1276), .ZN(new_n1302));
  NOR3_X1   g1102(.A1(new_n1299), .A2(new_n1300), .A3(new_n1302), .ZN(new_n1303));
  NOR2_X1   g1103(.A1(new_n1291), .A2(new_n1293), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1304), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1298), .B1(new_n1303), .B2(new_n1305), .ZN(G405));
  AOI21_X1  g1106(.A(G378), .B1(new_n1178), .B2(new_n1208), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1307), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1308), .A2(new_n1267), .A3(new_n1275), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1267), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1276), .B1(new_n1307), .B2(new_n1310), .ZN(new_n1311));
  AND3_X1   g1111(.A1(new_n1309), .A2(new_n1304), .A3(new_n1311), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1304), .B1(new_n1309), .B2(new_n1311), .ZN(new_n1313));
  NOR2_X1   g1113(.A1(new_n1312), .A2(new_n1313), .ZN(G402));
endmodule


