

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760;

  NOR2_X1 U363 ( .A1(n597), .A2(n343), .ZN(n650) );
  OR2_X1 U364 ( .A1(n608), .A2(n607), .ZN(n610) );
  AND2_X1 U365 ( .A1(n443), .A2(n355), .ZN(n441) );
  OR2_X1 U366 ( .A1(n677), .A2(n678), .ZN(n567) );
  XNOR2_X1 U367 ( .A(n684), .B(KEYINPUT6), .ZN(n608) );
  XNOR2_X1 U368 ( .A(n412), .B(KEYINPUT1), .ZN(n677) );
  INV_X1 U369 ( .A(n684), .ZN(n404) );
  NAND2_X1 U370 ( .A1(n406), .A2(n664), .ZN(n612) );
  XNOR2_X1 U371 ( .A(n436), .B(n733), .ZN(n702) );
  XNOR2_X1 U372 ( .A(n515), .B(G134), .ZN(n411) );
  NAND2_X1 U373 ( .A1(n387), .A2(n386), .ZN(n744) );
  NAND2_X1 U374 ( .A1(n361), .A2(n549), .ZN(n368) );
  XNOR2_X1 U375 ( .A(n524), .B(n391), .ZN(n361) );
  XNOR2_X2 U376 ( .A(n341), .B(KEYINPUT65), .ZN(n629) );
  NAND2_X2 U377 ( .A1(n433), .A2(n477), .ZN(n341) );
  XNOR2_X2 U378 ( .A(n342), .B(KEYINPUT33), .ZN(n662) );
  NAND2_X2 U379 ( .A1(n555), .A2(n554), .ZN(n342) );
  XNOR2_X2 U380 ( .A(n411), .B(n526), .ZN(n743) );
  NAND2_X2 U381 ( .A1(n428), .A2(n427), .ZN(n425) );
  XNOR2_X1 U382 ( .A(n481), .B(G110), .ZN(n734) );
  NOR2_X1 U383 ( .A1(n404), .A2(n607), .ZN(n423) );
  INV_X1 U384 ( .A(G953), .ZN(n752) );
  NOR2_X2 U385 ( .A1(n613), .A2(n612), .ZN(n614) );
  XNOR2_X2 U386 ( .A(n616), .B(n615), .ZN(n628) );
  XNOR2_X2 U387 ( .A(n612), .B(n493), .ZN(n598) );
  XNOR2_X2 U388 ( .A(G104), .B(G107), .ZN(n481) );
  XNOR2_X2 U389 ( .A(KEYINPUT42), .B(n595), .ZN(n758) );
  XNOR2_X2 U390 ( .A(n455), .B(n454), .ZN(n515) );
  XNOR2_X1 U391 ( .A(n543), .B(n437), .ZN(n709) );
  NOR2_X1 U392 ( .A1(n667), .A2(n666), .ZN(n432) );
  NOR2_X1 U393 ( .A1(G902), .A2(n709), .ZN(n530) );
  INV_X1 U394 ( .A(G469), .ZN(n527) );
  INV_X1 U395 ( .A(KEYINPUT28), .ZN(n422) );
  NOR2_X1 U396 ( .A1(n757), .A2(n644), .ZN(n558) );
  AND2_X1 U397 ( .A1(n566), .A2(n344), .ZN(n644) );
  XNOR2_X1 U398 ( .A(n407), .B(KEYINPUT98), .ZN(n640) );
  XNOR2_X1 U399 ( .A(n368), .B(n551), .ZN(n757) );
  XNOR2_X1 U400 ( .A(n432), .B(n431), .ZN(n689) );
  NOR2_X1 U401 ( .A1(n594), .A2(n412), .ZN(n596) );
  XNOR2_X1 U402 ( .A(n423), .B(n422), .ZN(n594) );
  XNOR2_X1 U403 ( .A(n606), .B(KEYINPUT107), .ZN(n637) );
  NAND2_X2 U404 ( .A1(n394), .A2(n392), .ZN(n406) );
  AND2_X1 U405 ( .A1(n396), .A2(n395), .ZN(n394) );
  INV_X1 U406 ( .A(n440), .ZN(n343) );
  XNOR2_X1 U407 ( .A(n545), .B(n472), .ZN(n390) );
  XNOR2_X2 U408 ( .A(n580), .B(n475), .ZN(n479) );
  NOR2_X2 U409 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X2 U410 ( .A(n743), .B(n457), .ZN(n543) );
  INV_X1 U411 ( .A(KEYINPUT67), .ZN(n459) );
  XNOR2_X1 U412 ( .A(n449), .B(n448), .ZN(n666) );
  INV_X1 U413 ( .A(KEYINPUT104), .ZN(n448) );
  NOR2_X1 U414 ( .A1(n561), .A2(n560), .ZN(n449) );
  XNOR2_X1 U415 ( .A(n542), .B(n352), .ZN(n733) );
  NAND2_X1 U416 ( .A1(n470), .A2(n469), .ZN(n468) );
  NAND2_X1 U417 ( .A1(KEYINPUT0), .A2(KEYINPUT89), .ZN(n470) );
  NAND2_X1 U418 ( .A1(n471), .A2(n499), .ZN(n469) );
  INV_X1 U419 ( .A(G143), .ZN(n454) );
  XNOR2_X1 U420 ( .A(n473), .B(n483), .ZN(n542) );
  XNOR2_X1 U421 ( .A(n484), .B(n482), .ZN(n473) );
  XNOR2_X1 U422 ( .A(KEYINPUT74), .B(KEYINPUT90), .ZN(n484) );
  XNOR2_X1 U423 ( .A(n511), .B(n510), .ZN(n560) );
  INV_X1 U424 ( .A(KEYINPUT95), .ZN(n559) );
  XNOR2_X1 U425 ( .A(n500), .B(KEYINPUT10), .ZN(n532) );
  XNOR2_X1 U426 ( .A(n734), .B(KEYINPUT76), .ZN(n472) );
  XNOR2_X1 U427 ( .A(n430), .B(KEYINPUT86), .ZN(n413) );
  NAND2_X1 U428 ( .A1(n749), .A2(KEYINPUT2), .ZN(n430) );
  INV_X1 U429 ( .A(KEYINPUT22), .ZN(n391) );
  NAND2_X1 U430 ( .A1(n345), .A2(n490), .ZN(n395) );
  XNOR2_X1 U431 ( .A(n402), .B(n421), .ZN(n401) );
  INV_X1 U432 ( .A(G137), .ZN(n421) );
  NAND2_X1 U433 ( .A1(n544), .A2(G210), .ZN(n402) );
  XNOR2_X1 U434 ( .A(n400), .B(KEYINPUT97), .ZN(n399) );
  INV_X1 U435 ( .A(KEYINPUT5), .ZN(n400) );
  AND2_X1 U436 ( .A1(n752), .A2(n403), .ZN(n544) );
  INV_X1 U437 ( .A(G237), .ZN(n403) );
  XNOR2_X1 U438 ( .A(G131), .B(KEYINPUT70), .ZN(n526) );
  INV_X1 U439 ( .A(KEYINPUT91), .ZN(n485) );
  NOR2_X1 U440 ( .A1(n383), .A2(n382), .ZN(n381) );
  NOR2_X1 U441 ( .A1(n760), .A2(n623), .ZN(n627) );
  XNOR2_X1 U442 ( .A(n533), .B(n373), .ZN(n372) );
  XNOR2_X1 U443 ( .A(n374), .B(KEYINPUT75), .ZN(n373) );
  INV_X1 U444 ( .A(KEYINPUT23), .ZN(n374) );
  XNOR2_X1 U445 ( .A(n532), .B(n531), .ZN(n742) );
  XNOR2_X1 U446 ( .A(n516), .B(G116), .ZN(n453) );
  XOR2_X1 U447 ( .A(KEYINPUT7), .B(G107), .Z(n516) );
  INV_X1 U448 ( .A(G146), .ZN(n457) );
  INV_X1 U449 ( .A(KEYINPUT45), .ZN(n475) );
  XNOR2_X1 U450 ( .A(n429), .B(KEYINPUT39), .ZN(n622) );
  XNOR2_X1 U451 ( .A(n369), .B(KEYINPUT106), .ZN(n548) );
  OR2_X1 U452 ( .A1(n438), .A2(n675), .ZN(n369) );
  NAND2_X1 U453 ( .A1(n440), .A2(n444), .ZN(n439) );
  NOR2_X1 U454 ( .A1(n445), .A2(n359), .ZN(n444) );
  XNOR2_X1 U455 ( .A(n541), .B(n461), .ZN(n460) );
  OR2_X1 U456 ( .A1(n724), .A2(G902), .ZN(n462) );
  INV_X1 U457 ( .A(KEYINPUT81), .ZN(n461) );
  XNOR2_X1 U458 ( .A(n520), .B(n450), .ZN(n561) );
  XNOR2_X1 U459 ( .A(n519), .B(G478), .ZN(n450) );
  AND2_X1 U460 ( .A1(n361), .A2(n438), .ZN(n566) );
  XNOR2_X1 U461 ( .A(n506), .B(n434), .ZN(n508) );
  INV_X1 U462 ( .A(G475), .ZN(n366) );
  XNOR2_X1 U463 ( .A(n390), .B(n489), .ZN(n436) );
  INV_X1 U464 ( .A(G210), .ZN(n367) );
  NOR2_X1 U465 ( .A1(G952), .A2(n414), .ZN(n726) );
  NAND2_X1 U466 ( .A1(n379), .A2(n378), .ZN(n375) );
  NOR2_X1 U467 ( .A1(G902), .A2(G237), .ZN(n491) );
  INV_X1 U468 ( .A(n347), .ZN(n445) );
  NAND2_X1 U469 ( .A1(n471), .A2(KEYINPUT89), .ZN(n466) );
  NAND2_X1 U470 ( .A1(KEYINPUT0), .A2(n499), .ZN(n467) );
  INV_X1 U471 ( .A(n468), .ZN(n442) );
  OR2_X1 U472 ( .A1(n345), .A2(n490), .ZN(n393) );
  XNOR2_X1 U473 ( .A(n546), .B(n542), .ZN(n456) );
  XNOR2_X1 U474 ( .A(n401), .B(n399), .ZN(n420) );
  XOR2_X1 U475 ( .A(KEYINPUT100), .B(G122), .Z(n502) );
  XNOR2_X1 U476 ( .A(G113), .B(G143), .ZN(n501) );
  XOR2_X1 U477 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n505) );
  XNOR2_X1 U478 ( .A(n507), .B(n435), .ZN(n434) );
  INV_X1 U479 ( .A(G104), .ZN(n435) );
  XNOR2_X1 U480 ( .A(G131), .B(G140), .ZN(n507) );
  NAND2_X1 U481 ( .A1(n490), .A2(KEYINPUT2), .ZN(n477) );
  XNOR2_X1 U482 ( .A(n446), .B(n447), .ZN(n426) );
  NAND2_X1 U483 ( .A1(n752), .A2(G224), .ZN(n446) );
  XNOR2_X1 U484 ( .A(n485), .B(KEYINPUT17), .ZN(n447) );
  BUF_X1 U485 ( .A(n662), .Z(n672) );
  INV_X1 U486 ( .A(KEYINPUT41), .ZN(n431) );
  INV_X1 U487 ( .A(n591), .ZN(n417) );
  XNOR2_X1 U488 ( .A(n536), .B(n372), .ZN(n371) );
  XNOR2_X1 U489 ( .A(n518), .B(n451), .ZN(n718) );
  XNOR2_X1 U490 ( .A(n453), .B(n517), .ZN(n452) );
  XNOR2_X1 U491 ( .A(n390), .B(n348), .ZN(n437) );
  NAND2_X1 U492 ( .A1(n479), .A2(n749), .ZN(n476) );
  XNOR2_X1 U493 ( .A(n398), .B(n397), .ZN(n760) );
  INV_X1 U494 ( .A(KEYINPUT110), .ZN(n397) );
  NAND2_X1 U495 ( .A1(n622), .A2(n606), .ZN(n590) );
  INV_X1 U496 ( .A(KEYINPUT35), .ZN(n424) );
  INV_X1 U497 ( .A(n601), .ZN(n427) );
  XNOR2_X1 U498 ( .A(n550), .B(KEYINPUT32), .ZN(n551) );
  INV_X1 U499 ( .A(n637), .ZN(n652) );
  INV_X1 U500 ( .A(n592), .ZN(n418) );
  XNOR2_X1 U501 ( .A(n410), .B(n409), .ZN(n408) );
  INV_X1 U502 ( .A(KEYINPUT96), .ZN(n409) );
  NOR2_X1 U503 ( .A1(n716), .A2(n726), .ZN(n717) );
  XNOR2_X1 U504 ( .A(n702), .B(n703), .ZN(n704) );
  XNOR2_X1 U505 ( .A(n464), .B(n463), .ZN(G75) );
  XNOR2_X1 U506 ( .A(KEYINPUT121), .B(KEYINPUT53), .ZN(n463) );
  OR2_X1 U507 ( .A1(n700), .A2(n465), .ZN(n464) );
  OR2_X1 U508 ( .A1(n701), .A2(G953), .ZN(n465) );
  AND2_X1 U509 ( .A1(n404), .A2(n418), .ZN(n344) );
  BUF_X1 U510 ( .A(n677), .Z(n438) );
  AND2_X1 U511 ( .A1(G210), .A2(n492), .ZN(n345) );
  OR2_X1 U512 ( .A1(KEYINPUT47), .A2(n605), .ZN(n346) );
  OR2_X1 U513 ( .A1(n585), .A2(n498), .ZN(n347) );
  XOR2_X1 U514 ( .A(n525), .B(n531), .Z(n348) );
  AND2_X1 U515 ( .A1(G221), .A2(n537), .ZN(n349) );
  AND2_X1 U516 ( .A1(n476), .A2(n478), .ZN(n350) );
  XOR2_X1 U517 ( .A(n608), .B(KEYINPUT82), .Z(n351) );
  NAND2_X1 U518 ( .A1(n628), .A2(n627), .ZN(n624) );
  XOR2_X1 U519 ( .A(G122), .B(KEYINPUT16), .Z(n352) );
  AND2_X1 U520 ( .A1(n375), .A2(n346), .ZN(n353) );
  XOR2_X1 U521 ( .A(n604), .B(KEYINPUT84), .Z(n354) );
  OR2_X1 U522 ( .A1(n347), .A2(n442), .ZN(n355) );
  INV_X1 U523 ( .A(n438), .ZN(n619) );
  XNOR2_X1 U524 ( .A(KEYINPUT46), .B(KEYINPUT87), .ZN(n356) );
  INV_X1 U525 ( .A(KEYINPUT0), .ZN(n471) );
  XNOR2_X1 U526 ( .A(KEYINPUT77), .B(KEYINPUT34), .ZN(n357) );
  XOR2_X1 U527 ( .A(KEYINPUT38), .B(KEYINPUT78), .Z(n358) );
  AND2_X1 U528 ( .A1(n467), .A2(n466), .ZN(n359) );
  XOR2_X1 U529 ( .A(n630), .B(KEYINPUT62), .Z(n360) );
  INV_X1 U530 ( .A(KEYINPUT2), .ZN(n478) );
  XNOR2_X1 U531 ( .A(G902), .B(KEYINPUT15), .ZN(n625) );
  INV_X1 U532 ( .A(G472), .ZN(n405) );
  BUF_X1 U533 ( .A(n752), .Z(n414) );
  NAND2_X1 U534 ( .A1(n364), .A2(n362), .ZN(n705) );
  NOR2_X1 U535 ( .A1(n699), .A2(n367), .ZN(n362) );
  NAND2_X1 U536 ( .A1(n364), .A2(n363), .ZN(n714) );
  NOR2_X1 U537 ( .A1(n699), .A2(n366), .ZN(n363) );
  INV_X1 U538 ( .A(n629), .ZN(n364) );
  NOR2_X1 U539 ( .A1(n699), .A2(n629), .ZN(n722) );
  NAND2_X1 U540 ( .A1(n365), .A2(n364), .ZN(n631) );
  NOR2_X1 U541 ( .A1(n699), .A2(n405), .ZN(n365) );
  NAND2_X1 U542 ( .A1(n577), .A2(KEYINPUT44), .ZN(n575) );
  NAND2_X1 U543 ( .A1(n558), .A2(n756), .ZN(n577) );
  XNOR2_X2 U544 ( .A(n425), .B(n424), .ZN(n756) );
  XNOR2_X1 U545 ( .A(n553), .B(n459), .ZN(n678) );
  XNOR2_X1 U546 ( .A(n742), .B(n371), .ZN(n419) );
  NAND2_X2 U547 ( .A1(n441), .A2(n439), .ZN(n568) );
  NAND2_X1 U548 ( .A1(n370), .A2(n619), .ZN(n384) );
  XNOR2_X1 U549 ( .A(n614), .B(KEYINPUT36), .ZN(n370) );
  XNOR2_X2 U550 ( .A(G146), .B(G125), .ZN(n500) );
  AND2_X1 U551 ( .A1(n376), .A2(n353), .ZN(n377) );
  NAND2_X1 U552 ( .A1(n759), .A2(n380), .ZN(n376) );
  XNOR2_X2 U553 ( .A(n590), .B(KEYINPUT40), .ZN(n759) );
  NAND2_X1 U554 ( .A1(n381), .A2(n377), .ZN(n616) );
  INV_X1 U555 ( .A(n356), .ZN(n378) );
  INV_X1 U556 ( .A(n758), .ZN(n379) );
  AND2_X1 U557 ( .A1(n758), .A2(n356), .ZN(n380) );
  NOR2_X1 U558 ( .A1(n759), .A2(n356), .ZN(n382) );
  NAND2_X1 U559 ( .A1(n354), .A2(n384), .ZN(n383) );
  INV_X1 U560 ( .A(n384), .ZN(n658) );
  NAND2_X1 U561 ( .A1(n568), .A2(n385), .ZN(n410) );
  NAND2_X1 U562 ( .A1(n385), .A2(n416), .ZN(n415) );
  XNOR2_X1 U563 ( .A(n458), .B(n559), .ZN(n385) );
  NAND2_X1 U564 ( .A1(n389), .A2(n480), .ZN(n386) );
  NAND2_X1 U565 ( .A1(n388), .A2(KEYINPUT68), .ZN(n387) );
  INV_X1 U566 ( .A(n389), .ZN(n388) );
  XNOR2_X2 U567 ( .A(KEYINPUT4), .B(KEYINPUT64), .ZN(n389) );
  OR2_X1 U568 ( .A1(n702), .A2(n393), .ZN(n392) );
  NAND2_X1 U569 ( .A1(n702), .A2(n345), .ZN(n396) );
  OR2_X1 U570 ( .A1(n621), .A2(n406), .ZN(n398) );
  NOR2_X1 U571 ( .A1(n567), .A2(n404), .ZN(n686) );
  NAND2_X1 U572 ( .A1(n408), .A2(n404), .ZN(n407) );
  XNOR2_X2 U573 ( .A(n547), .B(n405), .ZN(n684) );
  XNOR2_X1 U574 ( .A(n406), .B(n358), .ZN(n663) );
  NAND2_X1 U575 ( .A1(n602), .A2(n406), .ZN(n648) );
  XNOR2_X1 U576 ( .A(n411), .B(n452), .ZN(n451) );
  XNOR2_X2 U577 ( .A(n530), .B(n529), .ZN(n412) );
  NOR2_X1 U578 ( .A1(n678), .A2(n412), .ZN(n458) );
  NOR2_X2 U579 ( .A1(n413), .A2(n727), .ZN(n699) );
  XNOR2_X1 U580 ( .A(n617), .B(KEYINPUT111), .ZN(n613) );
  XNOR2_X1 U581 ( .A(n419), .B(n349), .ZN(n724) );
  INV_X1 U582 ( .A(n415), .ZN(n600) );
  AND2_X1 U583 ( .A1(n588), .A2(n417), .ZN(n416) );
  NOR2_X1 U584 ( .A1(n706), .A2(n726), .ZN(n707) );
  NOR2_X2 U585 ( .A1(n611), .A2(n637), .ZN(n617) );
  NOR2_X1 U586 ( .A1(n624), .A2(n625), .ZN(n474) );
  XNOR2_X1 U587 ( .A(n545), .B(n420), .ZN(n546) );
  XNOR2_X1 U588 ( .A(n543), .B(n456), .ZN(n630) );
  XNOR2_X1 U589 ( .A(n515), .B(n426), .ZN(n488) );
  XNOR2_X1 U590 ( .A(n557), .B(n357), .ZN(n428) );
  NAND2_X1 U591 ( .A1(n600), .A2(n663), .ZN(n429) );
  NAND2_X1 U592 ( .A1(n474), .A2(n479), .ZN(n433) );
  NAND2_X1 U593 ( .A1(n568), .A2(n523), .ZN(n524) );
  INV_X1 U594 ( .A(n598), .ZN(n440) );
  NAND2_X1 U595 ( .A1(n598), .A2(n468), .ZN(n443) );
  XNOR2_X2 U596 ( .A(G128), .B(KEYINPUT83), .ZN(n455) );
  XNOR2_X2 U597 ( .A(n462), .B(n460), .ZN(n592) );
  INV_X1 U598 ( .A(n479), .ZN(n727) );
  XNOR2_X1 U599 ( .A(n631), .B(n360), .ZN(n633) );
  INV_X1 U600 ( .A(n608), .ZN(n554) );
  XNOR2_X1 U601 ( .A(KEYINPUT48), .B(KEYINPUT71), .ZN(n615) );
  INV_X1 U602 ( .A(KEYINPUT24), .ZN(n534) );
  XNOR2_X1 U603 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U604 ( .A(n528), .B(n527), .ZN(n529) );
  INV_X1 U605 ( .A(n726), .ZN(n632) );
  NAND2_X1 U606 ( .A1(n633), .A2(n632), .ZN(n634) );
  INV_X1 U607 ( .A(KEYINPUT89), .ZN(n499) );
  INV_X1 U608 ( .A(n625), .ZN(n490) );
  INV_X1 U609 ( .A(KEYINPUT68), .ZN(n480) );
  XNOR2_X2 U610 ( .A(n744), .B(G101), .ZN(n545) );
  XOR2_X1 U611 ( .A(G113), .B(KEYINPUT3), .Z(n483) );
  XNOR2_X1 U612 ( .A(G119), .B(G116), .ZN(n482) );
  INV_X1 U613 ( .A(n500), .ZN(n486) );
  XNOR2_X1 U614 ( .A(n486), .B(KEYINPUT18), .ZN(n487) );
  XNOR2_X1 U615 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U616 ( .A(n491), .B(KEYINPUT79), .ZN(n492) );
  NAND2_X1 U617 ( .A1(G214), .A2(n492), .ZN(n664) );
  INV_X1 U618 ( .A(KEYINPUT19), .ZN(n493) );
  NAND2_X1 U619 ( .A1(G234), .A2(G237), .ZN(n494) );
  XNOR2_X1 U620 ( .A(n494), .B(KEYINPUT14), .ZN(n496) );
  NAND2_X1 U621 ( .A1(n496), .A2(G952), .ZN(n495) );
  XOR2_X1 U622 ( .A(n495), .B(KEYINPUT92), .Z(n694) );
  AND2_X1 U623 ( .A1(n414), .A2(n694), .ZN(n585) );
  NAND2_X1 U624 ( .A1(G902), .A2(n496), .ZN(n581) );
  NOR2_X1 U625 ( .A1(G898), .A2(n414), .ZN(n497) );
  XNOR2_X1 U626 ( .A(KEYINPUT93), .B(n497), .ZN(n739) );
  NOR2_X1 U627 ( .A1(n581), .A2(n739), .ZN(n498) );
  XNOR2_X1 U628 ( .A(KEYINPUT13), .B(G475), .ZN(n511) );
  XNOR2_X1 U629 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U630 ( .A(n532), .B(n503), .ZN(n509) );
  NAND2_X1 U631 ( .A1(G214), .A2(n544), .ZN(n504) );
  XNOR2_X1 U632 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U633 ( .A(n509), .B(n508), .ZN(n713) );
  NOR2_X1 U634 ( .A1(G902), .A2(n713), .ZN(n510) );
  XOR2_X1 U635 ( .A(KEYINPUT8), .B(KEYINPUT69), .Z(n513) );
  NAND2_X1 U636 ( .A1(G234), .A2(n752), .ZN(n512) );
  XNOR2_X1 U637 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U638 ( .A(KEYINPUT85), .B(n514), .ZN(n537) );
  NAND2_X1 U639 ( .A1(n537), .A2(G217), .ZN(n518) );
  XOR2_X1 U640 ( .A(G122), .B(KEYINPUT9), .Z(n517) );
  NOR2_X1 U641 ( .A1(G902), .A2(n718), .ZN(n520) );
  XNOR2_X1 U642 ( .A(KEYINPUT102), .B(KEYINPUT103), .ZN(n519) );
  NAND2_X1 U643 ( .A1(G234), .A2(n625), .ZN(n521) );
  XNOR2_X1 U644 ( .A(KEYINPUT20), .B(n521), .ZN(n538) );
  NAND2_X1 U645 ( .A1(n538), .A2(G221), .ZN(n522) );
  XNOR2_X1 U646 ( .A(n522), .B(KEYINPUT21), .ZN(n552) );
  NOR2_X1 U647 ( .A1(n666), .A2(n552), .ZN(n523) );
  NAND2_X1 U648 ( .A1(G227), .A2(n414), .ZN(n525) );
  XNOR2_X1 U649 ( .A(G137), .B(G140), .ZN(n531) );
  XNOR2_X1 U650 ( .A(KEYINPUT72), .B(KEYINPUT73), .ZN(n528) );
  XNOR2_X1 U651 ( .A(G119), .B(KEYINPUT94), .ZN(n533) );
  XNOR2_X1 U652 ( .A(G128), .B(G110), .ZN(n535) );
  XOR2_X1 U653 ( .A(KEYINPUT25), .B(KEYINPUT80), .Z(n540) );
  NAND2_X1 U654 ( .A1(G217), .A2(n538), .ZN(n539) );
  XNOR2_X1 U655 ( .A(n540), .B(n539), .ZN(n541) );
  XOR2_X1 U656 ( .A(n592), .B(KEYINPUT105), .Z(n675) );
  NOR2_X1 U657 ( .A1(n630), .A2(G902), .ZN(n547) );
  NOR2_X1 U658 ( .A1(n548), .A2(n351), .ZN(n549) );
  INV_X1 U659 ( .A(KEYINPUT66), .ZN(n550) );
  NAND2_X1 U660 ( .A1(n560), .A2(n561), .ZN(n601) );
  INV_X1 U661 ( .A(n552), .ZN(n674) );
  NAND2_X1 U662 ( .A1(n674), .A2(n592), .ZN(n553) );
  INV_X1 U663 ( .A(n567), .ZN(n555) );
  NAND2_X1 U664 ( .A1(n662), .A2(n568), .ZN(n557) );
  XNOR2_X1 U665 ( .A(n560), .B(KEYINPUT101), .ZN(n562) );
  NAND2_X1 U666 ( .A1(n561), .A2(n562), .ZN(n639) );
  INV_X1 U667 ( .A(n561), .ZN(n564) );
  INV_X1 U668 ( .A(n562), .ZN(n563) );
  NAND2_X1 U669 ( .A1(n564), .A2(n563), .ZN(n589) );
  NAND2_X1 U670 ( .A1(n639), .A2(n589), .ZN(n599) );
  INV_X1 U671 ( .A(n599), .ZN(n668) );
  NOR2_X1 U672 ( .A1(n640), .A2(n668), .ZN(n573) );
  AND2_X1 U673 ( .A1(n608), .A2(n675), .ZN(n565) );
  NAND2_X1 U674 ( .A1(n566), .A2(n565), .ZN(n635) );
  XOR2_X1 U675 ( .A(KEYINPUT31), .B(KEYINPUT99), .Z(n570) );
  NAND2_X1 U676 ( .A1(n686), .A2(n568), .ZN(n569) );
  XNOR2_X1 U677 ( .A(n570), .B(n569), .ZN(n656) );
  NAND2_X1 U678 ( .A1(n656), .A2(n599), .ZN(n571) );
  NAND2_X1 U679 ( .A1(n635), .A2(n571), .ZN(n572) );
  NOR2_X1 U680 ( .A1(n573), .A2(n572), .ZN(n574) );
  NAND2_X1 U681 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U682 ( .A(n576), .B(KEYINPUT88), .ZN(n579) );
  NOR2_X1 U683 ( .A1(n577), .A2(KEYINPUT44), .ZN(n578) );
  OR2_X1 U684 ( .A1(n414), .A2(n581), .ZN(n582) );
  XNOR2_X1 U685 ( .A(KEYINPUT108), .B(n582), .ZN(n583) );
  NOR2_X1 U686 ( .A1(G900), .A2(n583), .ZN(n584) );
  NOR2_X1 U687 ( .A1(n585), .A2(n584), .ZN(n591) );
  INV_X1 U688 ( .A(KEYINPUT30), .ZN(n587) );
  NAND2_X1 U689 ( .A1(n684), .A2(n664), .ZN(n586) );
  XNOR2_X1 U690 ( .A(n587), .B(n586), .ZN(n588) );
  INV_X1 U691 ( .A(n589), .ZN(n606) );
  NAND2_X1 U692 ( .A1(n664), .A2(n663), .ZN(n667) );
  NOR2_X1 U693 ( .A1(n592), .A2(n591), .ZN(n593) );
  NAND2_X1 U694 ( .A1(n593), .A2(n674), .ZN(n607) );
  NAND2_X1 U695 ( .A1(n689), .A2(n596), .ZN(n595) );
  INV_X1 U696 ( .A(n596), .ZN(n597) );
  NAND2_X1 U697 ( .A1(n650), .A2(n599), .ZN(n605) );
  NAND2_X1 U698 ( .A1(n605), .A2(KEYINPUT47), .ZN(n603) );
  NOR2_X1 U699 ( .A1(n601), .A2(n415), .ZN(n602) );
  NAND2_X1 U700 ( .A1(n603), .A2(n648), .ZN(n604) );
  INV_X1 U701 ( .A(KEYINPUT109), .ZN(n609) );
  XNOR2_X1 U702 ( .A(n610), .B(n609), .ZN(n611) );
  NAND2_X1 U703 ( .A1(n617), .A2(n664), .ZN(n618) );
  NOR2_X1 U704 ( .A1(n619), .A2(n618), .ZN(n620) );
  XNOR2_X1 U705 ( .A(n620), .B(KEYINPUT43), .ZN(n621) );
  INV_X1 U706 ( .A(n639), .ZN(n655) );
  NAND2_X1 U707 ( .A1(n622), .A2(n655), .ZN(n661) );
  INV_X1 U708 ( .A(n661), .ZN(n623) );
  AND2_X2 U709 ( .A1(n628), .A2(n627), .ZN(n749) );
  XNOR2_X1 U710 ( .A(n634), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U711 ( .A(G101), .B(KEYINPUT112), .ZN(n636) );
  XNOR2_X1 U712 ( .A(n636), .B(n635), .ZN(G3) );
  NOR2_X1 U713 ( .A1(n640), .A2(n637), .ZN(n638) );
  XOR2_X1 U714 ( .A(G104), .B(n638), .Z(G6) );
  NOR2_X1 U715 ( .A1(n640), .A2(n639), .ZN(n642) );
  XNOR2_X1 U716 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n641) );
  XNOR2_X1 U717 ( .A(n642), .B(n641), .ZN(n643) );
  XNOR2_X1 U718 ( .A(G107), .B(n643), .ZN(G9) );
  XOR2_X1 U719 ( .A(n644), .B(G110), .Z(G12) );
  XOR2_X1 U720 ( .A(KEYINPUT113), .B(KEYINPUT29), .Z(n646) );
  NAND2_X1 U721 ( .A1(n650), .A2(n655), .ZN(n645) );
  XNOR2_X1 U722 ( .A(n646), .B(n645), .ZN(n647) );
  XOR2_X1 U723 ( .A(G128), .B(n647), .Z(G30) );
  XNOR2_X1 U724 ( .A(G143), .B(KEYINPUT114), .ZN(n649) );
  XNOR2_X1 U725 ( .A(n649), .B(n648), .ZN(G45) );
  NAND2_X1 U726 ( .A1(n650), .A2(n652), .ZN(n651) );
  XNOR2_X1 U727 ( .A(n651), .B(G146), .ZN(G48) );
  XOR2_X1 U728 ( .A(G113), .B(KEYINPUT115), .Z(n654) );
  NAND2_X1 U729 ( .A1(n652), .A2(n656), .ZN(n653) );
  XNOR2_X1 U730 ( .A(n654), .B(n653), .ZN(G15) );
  NAND2_X1 U731 ( .A1(n656), .A2(n655), .ZN(n657) );
  XNOR2_X1 U732 ( .A(n657), .B(G116), .ZN(G18) );
  XNOR2_X1 U733 ( .A(n658), .B(KEYINPUT116), .ZN(n659) );
  XNOR2_X1 U734 ( .A(n659), .B(KEYINPUT37), .ZN(n660) );
  XNOR2_X1 U735 ( .A(G125), .B(n660), .ZN(G27) );
  XNOR2_X1 U736 ( .A(G134), .B(n661), .ZN(G36) );
  NAND2_X1 U737 ( .A1(n689), .A2(n672), .ZN(n697) );
  NOR2_X1 U738 ( .A1(n664), .A2(n663), .ZN(n665) );
  NOR2_X1 U739 ( .A1(n666), .A2(n665), .ZN(n670) );
  NOR2_X1 U740 ( .A1(n668), .A2(n667), .ZN(n669) );
  NOR2_X1 U741 ( .A1(n670), .A2(n669), .ZN(n671) );
  XNOR2_X1 U742 ( .A(n671), .B(KEYINPUT119), .ZN(n673) );
  NAND2_X1 U743 ( .A1(n673), .A2(n672), .ZN(n692) );
  NOR2_X1 U744 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U745 ( .A(KEYINPUT49), .B(n676), .ZN(n682) );
  XOR2_X1 U746 ( .A(KEYINPUT117), .B(KEYINPUT50), .Z(n680) );
  NAND2_X1 U747 ( .A1(n678), .A2(n438), .ZN(n679) );
  XNOR2_X1 U748 ( .A(n680), .B(n679), .ZN(n681) );
  NAND2_X1 U749 ( .A1(n682), .A2(n681), .ZN(n683) );
  NOR2_X1 U750 ( .A1(n684), .A2(n683), .ZN(n685) );
  NOR2_X1 U751 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U752 ( .A(n687), .B(KEYINPUT118), .ZN(n688) );
  XNOR2_X1 U753 ( .A(n688), .B(KEYINPUT51), .ZN(n690) );
  NAND2_X1 U754 ( .A1(n690), .A2(n689), .ZN(n691) );
  NAND2_X1 U755 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U756 ( .A(KEYINPUT52), .B(n693), .ZN(n695) );
  NAND2_X1 U757 ( .A1(n695), .A2(n694), .ZN(n696) );
  NAND2_X1 U758 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U759 ( .A(n698), .B(KEYINPUT120), .ZN(n701) );
  NOR2_X1 U760 ( .A1(n699), .A2(n350), .ZN(n700) );
  XOR2_X1 U761 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n703) );
  XNOR2_X1 U762 ( .A(n705), .B(n704), .ZN(n706) );
  XNOR2_X1 U763 ( .A(KEYINPUT56), .B(n707), .ZN(G51) );
  NAND2_X1 U764 ( .A1(n722), .A2(G469), .ZN(n711) );
  XOR2_X1 U765 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n708) );
  XNOR2_X1 U766 ( .A(n709), .B(n708), .ZN(n710) );
  XNOR2_X1 U767 ( .A(n711), .B(n710), .ZN(n712) );
  NOR2_X1 U768 ( .A1(n726), .A2(n712), .ZN(G54) );
  XOR2_X1 U769 ( .A(n713), .B(KEYINPUT59), .Z(n715) );
  XNOR2_X1 U770 ( .A(n715), .B(n714), .ZN(n716) );
  XNOR2_X1 U771 ( .A(n717), .B(KEYINPUT60), .ZN(G60) );
  XNOR2_X1 U772 ( .A(n718), .B(KEYINPUT122), .ZN(n720) );
  NAND2_X1 U773 ( .A1(G478), .A2(n722), .ZN(n719) );
  XNOR2_X1 U774 ( .A(n720), .B(n719), .ZN(n721) );
  NOR2_X1 U775 ( .A1(n726), .A2(n721), .ZN(G63) );
  NAND2_X1 U776 ( .A1(G217), .A2(n722), .ZN(n723) );
  XNOR2_X1 U777 ( .A(n724), .B(n723), .ZN(n725) );
  NOR2_X1 U778 ( .A1(n726), .A2(n725), .ZN(G66) );
  NOR2_X1 U779 ( .A1(G953), .A2(n727), .ZN(n728) );
  XNOR2_X1 U780 ( .A(n728), .B(KEYINPUT123), .ZN(n732) );
  NAND2_X1 U781 ( .A1(G953), .A2(G224), .ZN(n729) );
  XNOR2_X1 U782 ( .A(KEYINPUT61), .B(n729), .ZN(n730) );
  NAND2_X1 U783 ( .A1(n730), .A2(G898), .ZN(n731) );
  NAND2_X1 U784 ( .A1(n732), .A2(n731), .ZN(n741) );
  XNOR2_X1 U785 ( .A(n733), .B(KEYINPUT124), .ZN(n736) );
  XNOR2_X1 U786 ( .A(n734), .B(G101), .ZN(n735) );
  XNOR2_X1 U787 ( .A(n736), .B(n735), .ZN(n737) );
  XNOR2_X1 U788 ( .A(KEYINPUT125), .B(n737), .ZN(n738) );
  NAND2_X1 U789 ( .A1(n739), .A2(n738), .ZN(n740) );
  XOR2_X1 U790 ( .A(n741), .B(n740), .Z(G69) );
  XNOR2_X1 U791 ( .A(n742), .B(KEYINPUT126), .ZN(n746) );
  XNOR2_X1 U792 ( .A(n744), .B(n743), .ZN(n745) );
  XNOR2_X1 U793 ( .A(n746), .B(n745), .ZN(n750) );
  XNOR2_X1 U794 ( .A(G227), .B(n750), .ZN(n747) );
  NAND2_X1 U795 ( .A1(n747), .A2(G900), .ZN(n748) );
  NAND2_X1 U796 ( .A1(n748), .A2(G953), .ZN(n755) );
  XNOR2_X1 U797 ( .A(n750), .B(n749), .ZN(n751) );
  XNOR2_X1 U798 ( .A(n751), .B(KEYINPUT127), .ZN(n753) );
  NAND2_X1 U799 ( .A1(n753), .A2(n414), .ZN(n754) );
  NAND2_X1 U800 ( .A1(n755), .A2(n754), .ZN(G72) );
  XNOR2_X1 U801 ( .A(n756), .B(G122), .ZN(G24) );
  XOR2_X1 U802 ( .A(n757), .B(G119), .Z(G21) );
  XNOR2_X1 U803 ( .A(G137), .B(n758), .ZN(G39) );
  XNOR2_X1 U804 ( .A(n759), .B(G131), .ZN(G33) );
  XOR2_X1 U805 ( .A(G140), .B(n760), .Z(G42) );
endmodule

