

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U553 ( .A1(G29), .A2(n959), .ZN(n519) );
  INV_X1 U554 ( .A(n758), .ZN(n730) );
  NOR2_X1 U555 ( .A1(G164), .A2(G1384), .ZN(n710) );
  AND2_X1 U556 ( .A1(G2104), .A2(G2105), .ZN(n873) );
  NAND2_X1 U557 ( .A1(n873), .A2(G114), .ZN(n528) );
  INV_X1 U558 ( .A(G2105), .ZN(n523) );
  NOR2_X1 U559 ( .A1(G2104), .A2(n523), .ZN(n875) );
  NAND2_X1 U560 ( .A1(G126), .A2(n875), .ZN(n522) );
  NOR2_X1 U561 ( .A1(G2104), .A2(G2105), .ZN(n520) );
  XOR2_X2 U562 ( .A(KEYINPUT17), .B(n520), .Z(n880) );
  NAND2_X1 U563 ( .A1(G138), .A2(n880), .ZN(n521) );
  NAND2_X1 U564 ( .A1(n522), .A2(n521), .ZN(n526) );
  AND2_X1 U565 ( .A1(n523), .A2(G2104), .ZN(n879) );
  NAND2_X1 U566 ( .A1(G102), .A2(n879), .ZN(n524) );
  XOR2_X1 U567 ( .A(KEYINPUT86), .B(n524), .Z(n525) );
  NOR2_X1 U568 ( .A1(n526), .A2(n525), .ZN(n527) );
  NAND2_X1 U569 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U570 ( .A(n529), .B(KEYINPUT87), .ZN(G164) );
  INV_X1 U571 ( .A(G651), .ZN(n535) );
  NOR2_X1 U572 ( .A1(G543), .A2(n535), .ZN(n530) );
  XOR2_X1 U573 ( .A(KEYINPUT1), .B(n530), .Z(n629) );
  NAND2_X1 U574 ( .A1(G63), .A2(n629), .ZN(n532) );
  XOR2_X1 U575 ( .A(KEYINPUT0), .B(G543), .Z(n626) );
  NOR2_X2 U576 ( .A1(G651), .A2(n626), .ZN(n630) );
  NAND2_X1 U577 ( .A1(G51), .A2(n630), .ZN(n531) );
  NAND2_X1 U578 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U579 ( .A(KEYINPUT6), .B(n533), .ZN(n540) );
  NOR2_X1 U580 ( .A1(G651), .A2(G543), .ZN(n633) );
  NAND2_X1 U581 ( .A1(n633), .A2(G89), .ZN(n534) );
  XNOR2_X1 U582 ( .A(n534), .B(KEYINPUT4), .ZN(n537) );
  NOR2_X1 U583 ( .A1(n626), .A2(n535), .ZN(n635) );
  NAND2_X1 U584 ( .A1(G76), .A2(n635), .ZN(n536) );
  NAND2_X1 U585 ( .A1(n537), .A2(n536), .ZN(n538) );
  XOR2_X1 U586 ( .A(n538), .B(KEYINPUT5), .Z(n539) );
  NOR2_X1 U587 ( .A1(n540), .A2(n539), .ZN(n541) );
  XOR2_X1 U588 ( .A(KEYINPUT74), .B(n541), .Z(n542) );
  XNOR2_X1 U589 ( .A(KEYINPUT7), .B(n542), .ZN(G168) );
  XOR2_X1 U590 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U591 ( .A1(G64), .A2(n629), .ZN(n544) );
  NAND2_X1 U592 ( .A1(G52), .A2(n630), .ZN(n543) );
  NAND2_X1 U593 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U594 ( .A(KEYINPUT66), .B(n545), .ZN(n550) );
  NAND2_X1 U595 ( .A1(G77), .A2(n635), .ZN(n547) );
  NAND2_X1 U596 ( .A1(G90), .A2(n633), .ZN(n546) );
  NAND2_X1 U597 ( .A1(n547), .A2(n546), .ZN(n548) );
  XOR2_X1 U598 ( .A(KEYINPUT9), .B(n548), .Z(n549) );
  NOR2_X1 U599 ( .A1(n550), .A2(n549), .ZN(G171) );
  NAND2_X1 U600 ( .A1(G72), .A2(n635), .ZN(n552) );
  NAND2_X1 U601 ( .A1(G85), .A2(n633), .ZN(n551) );
  NAND2_X1 U602 ( .A1(n552), .A2(n551), .ZN(n556) );
  NAND2_X1 U603 ( .A1(G60), .A2(n629), .ZN(n554) );
  NAND2_X1 U604 ( .A1(G47), .A2(n630), .ZN(n553) );
  NAND2_X1 U605 ( .A1(n554), .A2(n553), .ZN(n555) );
  OR2_X1 U606 ( .A1(n556), .A2(n555), .ZN(G290) );
  AND2_X1 U607 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U608 ( .A1(G65), .A2(n629), .ZN(n558) );
  NAND2_X1 U609 ( .A1(G78), .A2(n635), .ZN(n557) );
  NAND2_X1 U610 ( .A1(n558), .A2(n557), .ZN(n562) );
  NAND2_X1 U611 ( .A1(G91), .A2(n633), .ZN(n560) );
  NAND2_X1 U612 ( .A1(G53), .A2(n630), .ZN(n559) );
  NAND2_X1 U613 ( .A1(n560), .A2(n559), .ZN(n561) );
  NOR2_X1 U614 ( .A1(n562), .A2(n561), .ZN(n717) );
  INV_X1 U615 ( .A(n717), .ZN(G299) );
  INV_X1 U616 ( .A(G57), .ZN(G237) );
  INV_X1 U617 ( .A(G132), .ZN(G219) );
  INV_X1 U618 ( .A(G82), .ZN(G220) );
  NAND2_X1 U619 ( .A1(G7), .A2(G661), .ZN(n563) );
  XNOR2_X1 U620 ( .A(n563), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U621 ( .A(G223), .ZN(n820) );
  NAND2_X1 U622 ( .A1(n820), .A2(G567), .ZN(n564) );
  XNOR2_X1 U623 ( .A(n564), .B(KEYINPUT67), .ZN(n565) );
  XNOR2_X1 U624 ( .A(KEYINPUT11), .B(n565), .ZN(G234) );
  NAND2_X1 U625 ( .A1(G56), .A2(n629), .ZN(n566) );
  XNOR2_X1 U626 ( .A(n566), .B(KEYINPUT68), .ZN(n567) );
  XNOR2_X1 U627 ( .A(KEYINPUT14), .B(n567), .ZN(n575) );
  NAND2_X1 U628 ( .A1(G68), .A2(n635), .ZN(n571) );
  XOR2_X1 U629 ( .A(KEYINPUT69), .B(KEYINPUT12), .Z(n569) );
  NAND2_X1 U630 ( .A1(G81), .A2(n633), .ZN(n568) );
  XNOR2_X1 U631 ( .A(n569), .B(n568), .ZN(n570) );
  NAND2_X1 U632 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U633 ( .A(n572), .B(KEYINPUT13), .ZN(n573) );
  XNOR2_X1 U634 ( .A(KEYINPUT70), .B(n573), .ZN(n574) );
  NAND2_X1 U635 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U636 ( .A(n576), .B(KEYINPUT71), .ZN(n578) );
  NAND2_X1 U637 ( .A1(G43), .A2(n630), .ZN(n577) );
  NAND2_X1 U638 ( .A1(n578), .A2(n577), .ZN(n982) );
  INV_X1 U639 ( .A(G860), .ZN(n826) );
  OR2_X1 U640 ( .A1(n982), .A2(n826), .ZN(G153) );
  NAND2_X1 U641 ( .A1(G868), .A2(G171), .ZN(n588) );
  NAND2_X1 U642 ( .A1(G66), .A2(n629), .ZN(n580) );
  NAND2_X1 U643 ( .A1(G92), .A2(n633), .ZN(n579) );
  NAND2_X1 U644 ( .A1(n580), .A2(n579), .ZN(n585) );
  NAND2_X1 U645 ( .A1(G79), .A2(n635), .ZN(n582) );
  NAND2_X1 U646 ( .A1(G54), .A2(n630), .ZN(n581) );
  NAND2_X1 U647 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U648 ( .A(KEYINPUT72), .B(n583), .ZN(n584) );
  NOR2_X1 U649 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U650 ( .A(n586), .B(KEYINPUT15), .ZN(n969) );
  INV_X1 U651 ( .A(n969), .ZN(n905) );
  INV_X1 U652 ( .A(G868), .ZN(n652) );
  NAND2_X1 U653 ( .A1(n905), .A2(n652), .ZN(n587) );
  NAND2_X1 U654 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U655 ( .A(n589), .B(KEYINPUT73), .ZN(G284) );
  NAND2_X1 U656 ( .A1(G868), .A2(G286), .ZN(n591) );
  NAND2_X1 U657 ( .A1(G299), .A2(n652), .ZN(n590) );
  NAND2_X1 U658 ( .A1(n591), .A2(n590), .ZN(G297) );
  NAND2_X1 U659 ( .A1(n826), .A2(G559), .ZN(n592) );
  NAND2_X1 U660 ( .A1(n592), .A2(n905), .ZN(n593) );
  XNOR2_X1 U661 ( .A(n593), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U662 ( .A1(G868), .A2(n982), .ZN(n596) );
  NAND2_X1 U663 ( .A1(G868), .A2(n905), .ZN(n594) );
  NOR2_X1 U664 ( .A1(G559), .A2(n594), .ZN(n595) );
  NOR2_X1 U665 ( .A1(n596), .A2(n595), .ZN(G282) );
  NAND2_X1 U666 ( .A1(G123), .A2(n875), .ZN(n597) );
  XNOR2_X1 U667 ( .A(n597), .B(KEYINPUT18), .ZN(n600) );
  NAND2_X1 U668 ( .A1(G135), .A2(n880), .ZN(n598) );
  XOR2_X1 U669 ( .A(KEYINPUT75), .B(n598), .Z(n599) );
  NAND2_X1 U670 ( .A1(n600), .A2(n599), .ZN(n604) );
  NAND2_X1 U671 ( .A1(G99), .A2(n879), .ZN(n602) );
  NAND2_X1 U672 ( .A1(G111), .A2(n873), .ZN(n601) );
  NAND2_X1 U673 ( .A1(n602), .A2(n601), .ZN(n603) );
  NOR2_X1 U674 ( .A1(n604), .A2(n603), .ZN(n944) );
  XNOR2_X1 U675 ( .A(n944), .B(G2096), .ZN(n606) );
  INV_X1 U676 ( .A(G2100), .ZN(n605) );
  NAND2_X1 U677 ( .A1(n606), .A2(n605), .ZN(G156) );
  XOR2_X1 U678 ( .A(KEYINPUT79), .B(KEYINPUT2), .Z(n608) );
  NAND2_X1 U679 ( .A1(G73), .A2(n635), .ZN(n607) );
  XNOR2_X1 U680 ( .A(n608), .B(n607), .ZN(n615) );
  NAND2_X1 U681 ( .A1(G61), .A2(n629), .ZN(n610) );
  NAND2_X1 U682 ( .A1(G86), .A2(n633), .ZN(n609) );
  NAND2_X1 U683 ( .A1(n610), .A2(n609), .ZN(n613) );
  NAND2_X1 U684 ( .A1(n630), .A2(G48), .ZN(n611) );
  XOR2_X1 U685 ( .A(KEYINPUT80), .B(n611), .Z(n612) );
  NOR2_X1 U686 ( .A1(n613), .A2(n612), .ZN(n614) );
  NAND2_X1 U687 ( .A1(n615), .A2(n614), .ZN(G305) );
  NAND2_X1 U688 ( .A1(G62), .A2(n629), .ZN(n617) );
  NAND2_X1 U689 ( .A1(G50), .A2(n630), .ZN(n616) );
  NAND2_X1 U690 ( .A1(n617), .A2(n616), .ZN(n618) );
  XNOR2_X1 U691 ( .A(KEYINPUT81), .B(n618), .ZN(n622) );
  NAND2_X1 U692 ( .A1(G75), .A2(n635), .ZN(n620) );
  NAND2_X1 U693 ( .A1(G88), .A2(n633), .ZN(n619) );
  AND2_X1 U694 ( .A1(n620), .A2(n619), .ZN(n621) );
  NAND2_X1 U695 ( .A1(n622), .A2(n621), .ZN(G303) );
  INV_X1 U696 ( .A(G303), .ZN(G166) );
  NAND2_X1 U697 ( .A1(G49), .A2(n630), .ZN(n624) );
  NAND2_X1 U698 ( .A1(G74), .A2(G651), .ZN(n623) );
  NAND2_X1 U699 ( .A1(n624), .A2(n623), .ZN(n625) );
  NOR2_X1 U700 ( .A1(n629), .A2(n625), .ZN(n628) );
  NAND2_X1 U701 ( .A1(n626), .A2(G87), .ZN(n627) );
  NAND2_X1 U702 ( .A1(n628), .A2(n627), .ZN(G288) );
  NAND2_X1 U703 ( .A1(G67), .A2(n629), .ZN(n632) );
  NAND2_X1 U704 ( .A1(G55), .A2(n630), .ZN(n631) );
  NAND2_X1 U705 ( .A1(n632), .A2(n631), .ZN(n640) );
  NAND2_X1 U706 ( .A1(n633), .A2(G93), .ZN(n634) );
  XNOR2_X1 U707 ( .A(n634), .B(KEYINPUT76), .ZN(n637) );
  NAND2_X1 U708 ( .A1(G80), .A2(n635), .ZN(n636) );
  NAND2_X1 U709 ( .A1(n637), .A2(n636), .ZN(n638) );
  XOR2_X1 U710 ( .A(KEYINPUT77), .B(n638), .Z(n639) );
  NOR2_X1 U711 ( .A1(n640), .A2(n639), .ZN(n641) );
  XOR2_X1 U712 ( .A(KEYINPUT78), .B(n641), .Z(n827) );
  XOR2_X1 U713 ( .A(KEYINPUT82), .B(KEYINPUT19), .Z(n642) );
  XNOR2_X1 U714 ( .A(G305), .B(n642), .ZN(n643) );
  XNOR2_X1 U715 ( .A(n827), .B(n643), .ZN(n645) );
  XNOR2_X1 U716 ( .A(G290), .B(G166), .ZN(n644) );
  XNOR2_X1 U717 ( .A(n645), .B(n644), .ZN(n646) );
  XNOR2_X1 U718 ( .A(n717), .B(n646), .ZN(n647) );
  XNOR2_X1 U719 ( .A(n647), .B(G288), .ZN(n903) );
  NAND2_X1 U720 ( .A1(G559), .A2(n905), .ZN(n648) );
  XOR2_X1 U721 ( .A(n982), .B(n648), .Z(n825) );
  XNOR2_X1 U722 ( .A(n903), .B(n825), .ZN(n649) );
  XNOR2_X1 U723 ( .A(n649), .B(KEYINPUT83), .ZN(n650) );
  NAND2_X1 U724 ( .A1(n650), .A2(G868), .ZN(n651) );
  XNOR2_X1 U725 ( .A(n651), .B(KEYINPUT84), .ZN(n654) );
  NAND2_X1 U726 ( .A1(n827), .A2(n652), .ZN(n653) );
  NAND2_X1 U727 ( .A1(n654), .A2(n653), .ZN(G295) );
  NAND2_X1 U728 ( .A1(G2078), .A2(G2084), .ZN(n655) );
  XOR2_X1 U729 ( .A(KEYINPUT20), .B(n655), .Z(n656) );
  NAND2_X1 U730 ( .A1(G2090), .A2(n656), .ZN(n657) );
  XNOR2_X1 U731 ( .A(KEYINPUT21), .B(n657), .ZN(n658) );
  NAND2_X1 U732 ( .A1(n658), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U733 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U734 ( .A1(G220), .A2(G219), .ZN(n659) );
  XOR2_X1 U735 ( .A(KEYINPUT22), .B(n659), .Z(n660) );
  NOR2_X1 U736 ( .A1(G218), .A2(n660), .ZN(n661) );
  NAND2_X1 U737 ( .A1(G96), .A2(n661), .ZN(n829) );
  NAND2_X1 U738 ( .A1(n829), .A2(G2106), .ZN(n665) );
  NAND2_X1 U739 ( .A1(G120), .A2(G69), .ZN(n662) );
  NOR2_X1 U740 ( .A1(G237), .A2(n662), .ZN(n663) );
  NAND2_X1 U741 ( .A1(G108), .A2(n663), .ZN(n830) );
  NAND2_X1 U742 ( .A1(n830), .A2(G567), .ZN(n664) );
  NAND2_X1 U743 ( .A1(n665), .A2(n664), .ZN(n831) );
  NAND2_X1 U744 ( .A1(G661), .A2(G483), .ZN(n666) );
  XOR2_X1 U745 ( .A(KEYINPUT85), .B(n666), .Z(n667) );
  NOR2_X1 U746 ( .A1(n831), .A2(n667), .ZN(n824) );
  NAND2_X1 U747 ( .A1(n824), .A2(G36), .ZN(G176) );
  NAND2_X1 U748 ( .A1(G101), .A2(n879), .ZN(n668) );
  XNOR2_X1 U749 ( .A(n668), .B(KEYINPUT23), .ZN(n669) );
  XNOR2_X1 U750 ( .A(n669), .B(KEYINPUT65), .ZN(n671) );
  NAND2_X1 U751 ( .A1(G137), .A2(n880), .ZN(n670) );
  NAND2_X1 U752 ( .A1(n671), .A2(n670), .ZN(n675) );
  NAND2_X1 U753 ( .A1(G125), .A2(n875), .ZN(n673) );
  NAND2_X1 U754 ( .A1(G113), .A2(n873), .ZN(n672) );
  NAND2_X1 U755 ( .A1(n673), .A2(n672), .ZN(n674) );
  NOR2_X1 U756 ( .A1(n675), .A2(n674), .ZN(G160) );
  XNOR2_X1 U757 ( .A(G1986), .B(G290), .ZN(n966) );
  NAND2_X1 U758 ( .A1(G160), .A2(G40), .ZN(n708) );
  NOR2_X1 U759 ( .A1(n710), .A2(n708), .ZN(n804) );
  NAND2_X1 U760 ( .A1(n966), .A2(n804), .ZN(n793) );
  XNOR2_X1 U761 ( .A(KEYINPUT88), .B(KEYINPUT34), .ZN(n679) );
  NAND2_X1 U762 ( .A1(G104), .A2(n879), .ZN(n677) );
  NAND2_X1 U763 ( .A1(G140), .A2(n880), .ZN(n676) );
  NAND2_X1 U764 ( .A1(n677), .A2(n676), .ZN(n678) );
  XNOR2_X1 U765 ( .A(n679), .B(n678), .ZN(n684) );
  NAND2_X1 U766 ( .A1(G128), .A2(n875), .ZN(n681) );
  NAND2_X1 U767 ( .A1(G116), .A2(n873), .ZN(n680) );
  NAND2_X1 U768 ( .A1(n681), .A2(n680), .ZN(n682) );
  XOR2_X1 U769 ( .A(KEYINPUT35), .B(n682), .Z(n683) );
  NOR2_X1 U770 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U771 ( .A(KEYINPUT36), .B(n685), .ZN(n887) );
  XNOR2_X1 U772 ( .A(KEYINPUT37), .B(G2067), .ZN(n801) );
  NOR2_X1 U773 ( .A1(n887), .A2(n801), .ZN(n935) );
  NAND2_X1 U774 ( .A1(n804), .A2(n935), .ZN(n799) );
  XNOR2_X1 U775 ( .A(n804), .B(KEYINPUT92), .ZN(n704) );
  NAND2_X1 U776 ( .A1(n873), .A2(G117), .ZN(n692) );
  NAND2_X1 U777 ( .A1(G129), .A2(n875), .ZN(n687) );
  NAND2_X1 U778 ( .A1(G141), .A2(n880), .ZN(n686) );
  NAND2_X1 U779 ( .A1(n687), .A2(n686), .ZN(n690) );
  NAND2_X1 U780 ( .A1(n879), .A2(G105), .ZN(n688) );
  XOR2_X1 U781 ( .A(KEYINPUT38), .B(n688), .Z(n689) );
  NOR2_X1 U782 ( .A1(n690), .A2(n689), .ZN(n691) );
  NAND2_X1 U783 ( .A1(n692), .A2(n691), .ZN(n693) );
  XOR2_X1 U784 ( .A(KEYINPUT91), .B(n693), .Z(n886) );
  NAND2_X1 U785 ( .A1(G1996), .A2(n886), .ZN(n703) );
  NAND2_X1 U786 ( .A1(G95), .A2(n879), .ZN(n694) );
  XNOR2_X1 U787 ( .A(n694), .B(KEYINPUT90), .ZN(n701) );
  NAND2_X1 U788 ( .A1(G131), .A2(n880), .ZN(n696) );
  NAND2_X1 U789 ( .A1(G107), .A2(n873), .ZN(n695) );
  NAND2_X1 U790 ( .A1(n696), .A2(n695), .ZN(n699) );
  NAND2_X1 U791 ( .A1(G119), .A2(n875), .ZN(n697) );
  XNOR2_X1 U792 ( .A(KEYINPUT89), .B(n697), .ZN(n698) );
  NOR2_X1 U793 ( .A1(n699), .A2(n698), .ZN(n700) );
  NAND2_X1 U794 ( .A1(n701), .A2(n700), .ZN(n891) );
  NAND2_X1 U795 ( .A1(G1991), .A2(n891), .ZN(n702) );
  NAND2_X1 U796 ( .A1(n703), .A2(n702), .ZN(n945) );
  NAND2_X1 U797 ( .A1(n704), .A2(n945), .ZN(n705) );
  XNOR2_X1 U798 ( .A(n705), .B(KEYINPUT93), .ZN(n796) );
  INV_X1 U799 ( .A(n796), .ZN(n706) );
  NAND2_X1 U800 ( .A1(n799), .A2(n706), .ZN(n707) );
  XNOR2_X1 U801 ( .A(n707), .B(KEYINPUT94), .ZN(n791) );
  INV_X1 U802 ( .A(n708), .ZN(n709) );
  NAND2_X1 U803 ( .A1(n710), .A2(n709), .ZN(n758) );
  NAND2_X1 U804 ( .A1(G8), .A2(n758), .ZN(n787) );
  NOR2_X1 U805 ( .A1(G2084), .A2(n758), .ZN(n743) );
  NAND2_X1 U806 ( .A1(G8), .A2(n743), .ZN(n756) );
  NOR2_X1 U807 ( .A1(G1966), .A2(n787), .ZN(n754) );
  OR2_X1 U808 ( .A1(n730), .A2(G1961), .ZN(n712) );
  XNOR2_X1 U809 ( .A(G2078), .B(KEYINPUT25), .ZN(n922) );
  NAND2_X1 U810 ( .A1(n730), .A2(n922), .ZN(n711) );
  NAND2_X1 U811 ( .A1(n712), .A2(n711), .ZN(n747) );
  NAND2_X1 U812 ( .A1(n747), .A2(G171), .ZN(n742) );
  NAND2_X1 U813 ( .A1(n730), .A2(G2072), .ZN(n713) );
  XNOR2_X1 U814 ( .A(n713), .B(KEYINPUT27), .ZN(n715) );
  INV_X1 U815 ( .A(G1956), .ZN(n996) );
  NOR2_X1 U816 ( .A1(n996), .A2(n730), .ZN(n714) );
  NOR2_X1 U817 ( .A1(n715), .A2(n714), .ZN(n718) );
  OR2_X1 U818 ( .A1(n718), .A2(n717), .ZN(n716) );
  XNOR2_X1 U819 ( .A(n716), .B(KEYINPUT28), .ZN(n739) );
  NAND2_X1 U820 ( .A1(n718), .A2(n717), .ZN(n737) );
  XNOR2_X1 U821 ( .A(KEYINPUT64), .B(KEYINPUT26), .ZN(n723) );
  NOR2_X1 U822 ( .A1(G1996), .A2(n723), .ZN(n722) );
  NAND2_X1 U823 ( .A1(G1348), .A2(n969), .ZN(n976) );
  NAND2_X1 U824 ( .A1(n976), .A2(n723), .ZN(n719) );
  NOR2_X1 U825 ( .A1(n719), .A2(G1341), .ZN(n720) );
  NOR2_X1 U826 ( .A1(n730), .A2(n720), .ZN(n721) );
  NOR2_X1 U827 ( .A1(n722), .A2(n721), .ZN(n728) );
  NAND2_X1 U828 ( .A1(n969), .A2(G2067), .ZN(n725) );
  NAND2_X1 U829 ( .A1(G1996), .A2(n723), .ZN(n724) );
  NAND2_X1 U830 ( .A1(n725), .A2(n724), .ZN(n726) );
  NAND2_X1 U831 ( .A1(n726), .A2(n730), .ZN(n727) );
  NAND2_X1 U832 ( .A1(n728), .A2(n727), .ZN(n729) );
  NOR2_X1 U833 ( .A1(n982), .A2(n729), .ZN(n735) );
  NAND2_X1 U834 ( .A1(G1348), .A2(n758), .ZN(n732) );
  NAND2_X1 U835 ( .A1(G2067), .A2(n730), .ZN(n731) );
  NAND2_X1 U836 ( .A1(n732), .A2(n731), .ZN(n733) );
  NOR2_X1 U837 ( .A1(n733), .A2(n969), .ZN(n734) );
  NOR2_X1 U838 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U839 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U840 ( .A1(n739), .A2(n738), .ZN(n740) );
  XOR2_X1 U841 ( .A(KEYINPUT29), .B(n740), .Z(n741) );
  NAND2_X1 U842 ( .A1(n742), .A2(n741), .ZN(n752) );
  NOR2_X1 U843 ( .A1(n754), .A2(n743), .ZN(n744) );
  NAND2_X1 U844 ( .A1(G8), .A2(n744), .ZN(n745) );
  XNOR2_X1 U845 ( .A(KEYINPUT30), .B(n745), .ZN(n746) );
  NOR2_X1 U846 ( .A1(G168), .A2(n746), .ZN(n749) );
  NOR2_X1 U847 ( .A1(G171), .A2(n747), .ZN(n748) );
  NOR2_X1 U848 ( .A1(n749), .A2(n748), .ZN(n750) );
  XOR2_X1 U849 ( .A(KEYINPUT31), .B(n750), .Z(n751) );
  NAND2_X1 U850 ( .A1(n752), .A2(n751), .ZN(n757) );
  INV_X1 U851 ( .A(n757), .ZN(n753) );
  NOR2_X1 U852 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U853 ( .A1(n756), .A2(n755), .ZN(n768) );
  NAND2_X1 U854 ( .A1(n757), .A2(G286), .ZN(n764) );
  NOR2_X1 U855 ( .A1(G1971), .A2(n787), .ZN(n760) );
  NOR2_X1 U856 ( .A1(G2090), .A2(n758), .ZN(n759) );
  NOR2_X1 U857 ( .A1(n760), .A2(n759), .ZN(n761) );
  XOR2_X1 U858 ( .A(KEYINPUT95), .B(n761), .Z(n762) );
  NAND2_X1 U859 ( .A1(n762), .A2(G303), .ZN(n763) );
  NAND2_X1 U860 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U861 ( .A1(G8), .A2(n765), .ZN(n766) );
  XNOR2_X1 U862 ( .A(KEYINPUT32), .B(n766), .ZN(n767) );
  NAND2_X1 U863 ( .A1(n768), .A2(n767), .ZN(n781) );
  NOR2_X1 U864 ( .A1(G1976), .A2(G288), .ZN(n972) );
  NOR2_X1 U865 ( .A1(G1971), .A2(G303), .ZN(n769) );
  NOR2_X1 U866 ( .A1(n972), .A2(n769), .ZN(n770) );
  NAND2_X1 U867 ( .A1(n781), .A2(n770), .ZN(n772) );
  NAND2_X1 U868 ( .A1(G288), .A2(G1976), .ZN(n771) );
  XNOR2_X1 U869 ( .A(n771), .B(KEYINPUT96), .ZN(n973) );
  NAND2_X1 U870 ( .A1(n772), .A2(n973), .ZN(n773) );
  NOR2_X1 U871 ( .A1(n787), .A2(n773), .ZN(n774) );
  NOR2_X1 U872 ( .A1(KEYINPUT33), .A2(n774), .ZN(n777) );
  NAND2_X1 U873 ( .A1(n972), .A2(KEYINPUT33), .ZN(n775) );
  NOR2_X1 U874 ( .A1(n775), .A2(n787), .ZN(n776) );
  NOR2_X1 U875 ( .A1(n777), .A2(n776), .ZN(n778) );
  XOR2_X1 U876 ( .A(G1981), .B(G305), .Z(n961) );
  NAND2_X1 U877 ( .A1(n778), .A2(n961), .ZN(n784) );
  NOR2_X1 U878 ( .A1(G2090), .A2(G303), .ZN(n779) );
  NAND2_X1 U879 ( .A1(G8), .A2(n779), .ZN(n780) );
  NAND2_X1 U880 ( .A1(n781), .A2(n780), .ZN(n782) );
  NAND2_X1 U881 ( .A1(n782), .A2(n787), .ZN(n783) );
  NAND2_X1 U882 ( .A1(n784), .A2(n783), .ZN(n789) );
  NOR2_X1 U883 ( .A1(G1981), .A2(G305), .ZN(n785) );
  XOR2_X1 U884 ( .A(n785), .B(KEYINPUT24), .Z(n786) );
  NOR2_X1 U885 ( .A1(n787), .A2(n786), .ZN(n788) );
  NOR2_X1 U886 ( .A1(n789), .A2(n788), .ZN(n790) );
  NOR2_X1 U887 ( .A1(n791), .A2(n790), .ZN(n792) );
  NAND2_X1 U888 ( .A1(n793), .A2(n792), .ZN(n807) );
  NOR2_X1 U889 ( .A1(G1996), .A2(n886), .ZN(n950) );
  NOR2_X1 U890 ( .A1(G1986), .A2(G290), .ZN(n794) );
  NOR2_X1 U891 ( .A1(G1991), .A2(n891), .ZN(n946) );
  NOR2_X1 U892 ( .A1(n794), .A2(n946), .ZN(n795) );
  NOR2_X1 U893 ( .A1(n796), .A2(n795), .ZN(n797) );
  NOR2_X1 U894 ( .A1(n950), .A2(n797), .ZN(n798) );
  XNOR2_X1 U895 ( .A(KEYINPUT39), .B(n798), .ZN(n800) );
  NAND2_X1 U896 ( .A1(n800), .A2(n799), .ZN(n802) );
  NAND2_X1 U897 ( .A1(n887), .A2(n801), .ZN(n937) );
  NAND2_X1 U898 ( .A1(n802), .A2(n937), .ZN(n803) );
  XOR2_X1 U899 ( .A(KEYINPUT97), .B(n803), .Z(n805) );
  NAND2_X1 U900 ( .A1(n805), .A2(n804), .ZN(n806) );
  NAND2_X1 U901 ( .A1(n807), .A2(n806), .ZN(n808) );
  XNOR2_X1 U902 ( .A(KEYINPUT40), .B(n808), .ZN(G329) );
  XNOR2_X1 U903 ( .A(KEYINPUT98), .B(G2446), .ZN(n818) );
  XOR2_X1 U904 ( .A(KEYINPUT99), .B(G2427), .Z(n810) );
  XNOR2_X1 U905 ( .A(G2435), .B(G2438), .ZN(n809) );
  XNOR2_X1 U906 ( .A(n810), .B(n809), .ZN(n814) );
  XOR2_X1 U907 ( .A(G2454), .B(G2430), .Z(n812) );
  XNOR2_X1 U908 ( .A(G1348), .B(G1341), .ZN(n811) );
  XNOR2_X1 U909 ( .A(n812), .B(n811), .ZN(n813) );
  XOR2_X1 U910 ( .A(n814), .B(n813), .Z(n816) );
  XNOR2_X1 U911 ( .A(G2451), .B(G2443), .ZN(n815) );
  XNOR2_X1 U912 ( .A(n816), .B(n815), .ZN(n817) );
  XNOR2_X1 U913 ( .A(n818), .B(n817), .ZN(n819) );
  NAND2_X1 U914 ( .A1(n819), .A2(G14), .ZN(n909) );
  XOR2_X1 U915 ( .A(KEYINPUT100), .B(n909), .Z(G401) );
  NAND2_X1 U916 ( .A1(G2106), .A2(n820), .ZN(G217) );
  AND2_X1 U917 ( .A1(G15), .A2(G2), .ZN(n821) );
  NAND2_X1 U918 ( .A1(G661), .A2(n821), .ZN(G259) );
  NAND2_X1 U919 ( .A1(G3), .A2(G1), .ZN(n822) );
  XOR2_X1 U920 ( .A(KEYINPUT101), .B(n822), .Z(n823) );
  NAND2_X1 U921 ( .A1(n824), .A2(n823), .ZN(G188) );
  XOR2_X1 U922 ( .A(G69), .B(KEYINPUT102), .Z(G235) );
  NAND2_X1 U924 ( .A1(n826), .A2(n825), .ZN(n828) );
  XNOR2_X1 U925 ( .A(n828), .B(n827), .ZN(G145) );
  INV_X1 U926 ( .A(G120), .ZN(G236) );
  INV_X1 U927 ( .A(G96), .ZN(G221) );
  NOR2_X1 U928 ( .A1(n830), .A2(n829), .ZN(G325) );
  INV_X1 U929 ( .A(G325), .ZN(G261) );
  INV_X1 U930 ( .A(n831), .ZN(G319) );
  XOR2_X1 U931 ( .A(KEYINPUT107), .B(KEYINPUT106), .Z(n833) );
  XNOR2_X1 U932 ( .A(G2067), .B(KEYINPUT105), .ZN(n832) );
  XNOR2_X1 U933 ( .A(n833), .B(n832), .ZN(n837) );
  XOR2_X1 U934 ( .A(KEYINPUT104), .B(KEYINPUT43), .Z(n835) );
  XNOR2_X1 U935 ( .A(G2678), .B(KEYINPUT103), .ZN(n834) );
  XNOR2_X1 U936 ( .A(n835), .B(n834), .ZN(n836) );
  XNOR2_X1 U937 ( .A(n837), .B(n836), .ZN(n844) );
  XOR2_X1 U938 ( .A(G2100), .B(KEYINPUT42), .Z(n839) );
  XNOR2_X1 U939 ( .A(G2078), .B(G2084), .ZN(n838) );
  XNOR2_X1 U940 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U941 ( .A(n840), .B(G2096), .Z(n842) );
  XNOR2_X1 U942 ( .A(G2072), .B(G2090), .ZN(n841) );
  XNOR2_X1 U943 ( .A(n842), .B(n841), .ZN(n843) );
  XNOR2_X1 U944 ( .A(n844), .B(n843), .ZN(G227) );
  XOR2_X1 U945 ( .A(G1981), .B(G1971), .Z(n846) );
  XNOR2_X1 U946 ( .A(G1966), .B(G1961), .ZN(n845) );
  XNOR2_X1 U947 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U948 ( .A(n847), .B(G2474), .Z(n849) );
  XNOR2_X1 U949 ( .A(G1986), .B(G1976), .ZN(n848) );
  XNOR2_X1 U950 ( .A(n849), .B(n848), .ZN(n853) );
  XOR2_X1 U951 ( .A(KEYINPUT41), .B(G1956), .Z(n851) );
  XNOR2_X1 U952 ( .A(G1996), .B(G1991), .ZN(n850) );
  XNOR2_X1 U953 ( .A(n851), .B(n850), .ZN(n852) );
  XNOR2_X1 U954 ( .A(n853), .B(n852), .ZN(G229) );
  NAND2_X1 U955 ( .A1(n873), .A2(G112), .ZN(n860) );
  NAND2_X1 U956 ( .A1(G100), .A2(n879), .ZN(n855) );
  NAND2_X1 U957 ( .A1(G136), .A2(n880), .ZN(n854) );
  NAND2_X1 U958 ( .A1(n855), .A2(n854), .ZN(n858) );
  NAND2_X1 U959 ( .A1(n875), .A2(G124), .ZN(n856) );
  XOR2_X1 U960 ( .A(KEYINPUT44), .B(n856), .Z(n857) );
  NOR2_X1 U961 ( .A1(n858), .A2(n857), .ZN(n859) );
  NAND2_X1 U962 ( .A1(n860), .A2(n859), .ZN(n861) );
  XOR2_X1 U963 ( .A(KEYINPUT108), .B(n861), .Z(G162) );
  NAND2_X1 U964 ( .A1(n873), .A2(G115), .ZN(n862) );
  XOR2_X1 U965 ( .A(KEYINPUT113), .B(n862), .Z(n864) );
  NAND2_X1 U966 ( .A1(n875), .A2(G127), .ZN(n863) );
  NAND2_X1 U967 ( .A1(n864), .A2(n863), .ZN(n865) );
  XNOR2_X1 U968 ( .A(n865), .B(KEYINPUT47), .ZN(n871) );
  NAND2_X1 U969 ( .A1(n880), .A2(G139), .ZN(n866) );
  XOR2_X1 U970 ( .A(KEYINPUT111), .B(n866), .Z(n868) );
  NAND2_X1 U971 ( .A1(n879), .A2(G103), .ZN(n867) );
  NAND2_X1 U972 ( .A1(n868), .A2(n867), .ZN(n869) );
  XOR2_X1 U973 ( .A(KEYINPUT112), .B(n869), .Z(n870) );
  NAND2_X1 U974 ( .A1(n871), .A2(n870), .ZN(n872) );
  XNOR2_X1 U975 ( .A(n872), .B(KEYINPUT114), .ZN(n938) );
  NAND2_X1 U976 ( .A1(G118), .A2(n873), .ZN(n874) );
  XNOR2_X1 U977 ( .A(n874), .B(KEYINPUT110), .ZN(n878) );
  NAND2_X1 U978 ( .A1(G130), .A2(n875), .ZN(n876) );
  XOR2_X1 U979 ( .A(KEYINPUT109), .B(n876), .Z(n877) );
  NAND2_X1 U980 ( .A1(n878), .A2(n877), .ZN(n885) );
  NAND2_X1 U981 ( .A1(G106), .A2(n879), .ZN(n882) );
  NAND2_X1 U982 ( .A1(G142), .A2(n880), .ZN(n881) );
  NAND2_X1 U983 ( .A1(n882), .A2(n881), .ZN(n883) );
  XOR2_X1 U984 ( .A(KEYINPUT45), .B(n883), .Z(n884) );
  NOR2_X1 U985 ( .A1(n885), .A2(n884), .ZN(n890) );
  XOR2_X1 U986 ( .A(n887), .B(n886), .Z(n888) );
  XNOR2_X1 U987 ( .A(G162), .B(n888), .ZN(n889) );
  XNOR2_X1 U988 ( .A(n890), .B(n889), .ZN(n893) );
  XNOR2_X1 U989 ( .A(n891), .B(n944), .ZN(n892) );
  XNOR2_X1 U990 ( .A(n893), .B(n892), .ZN(n897) );
  XOR2_X1 U991 ( .A(KEYINPUT46), .B(KEYINPUT115), .Z(n895) );
  XNOR2_X1 U992 ( .A(KEYINPUT48), .B(KEYINPUT116), .ZN(n894) );
  XNOR2_X1 U993 ( .A(n895), .B(n894), .ZN(n896) );
  XOR2_X1 U994 ( .A(n897), .B(n896), .Z(n899) );
  XNOR2_X1 U995 ( .A(G164), .B(G160), .ZN(n898) );
  XNOR2_X1 U996 ( .A(n899), .B(n898), .ZN(n900) );
  XOR2_X1 U997 ( .A(n938), .B(n900), .Z(n901) );
  NOR2_X1 U998 ( .A1(G37), .A2(n901), .ZN(G395) );
  XOR2_X1 U999 ( .A(n982), .B(G286), .Z(n902) );
  XNOR2_X1 U1000 ( .A(n903), .B(n902), .ZN(n904) );
  XOR2_X1 U1001 ( .A(n904), .B(KEYINPUT117), .Z(n907) );
  XNOR2_X1 U1002 ( .A(G171), .B(n905), .ZN(n906) );
  XNOR2_X1 U1003 ( .A(n907), .B(n906), .ZN(n908) );
  NOR2_X1 U1004 ( .A1(G37), .A2(n908), .ZN(G397) );
  NAND2_X1 U1005 ( .A1(G319), .A2(n909), .ZN(n912) );
  NOR2_X1 U1006 ( .A1(G227), .A2(G229), .ZN(n910) );
  XNOR2_X1 U1007 ( .A(KEYINPUT49), .B(n910), .ZN(n911) );
  NOR2_X1 U1008 ( .A1(n912), .A2(n911), .ZN(n914) );
  NOR2_X1 U1009 ( .A1(G395), .A2(G397), .ZN(n913) );
  NAND2_X1 U1010 ( .A1(n914), .A2(n913), .ZN(G225) );
  INV_X1 U1011 ( .A(G225), .ZN(G308) );
  INV_X1 U1012 ( .A(G171), .ZN(G301) );
  INV_X1 U1013 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1014 ( .A(KEYINPUT55), .B(KEYINPUT119), .ZN(n934) );
  XOR2_X1 U1015 ( .A(G2090), .B(G35), .Z(n928) );
  XOR2_X1 U1016 ( .A(KEYINPUT53), .B(KEYINPUT120), .Z(n926) );
  XNOR2_X1 U1017 ( .A(G1996), .B(G32), .ZN(n916) );
  XNOR2_X1 U1018 ( .A(G33), .B(G2072), .ZN(n915) );
  NOR2_X1 U1019 ( .A1(n916), .A2(n915), .ZN(n921) );
  XOR2_X1 U1020 ( .A(G2067), .B(G26), .Z(n917) );
  NAND2_X1 U1021 ( .A1(n917), .A2(G28), .ZN(n919) );
  XNOR2_X1 U1022 ( .A(G25), .B(G1991), .ZN(n918) );
  NOR2_X1 U1023 ( .A1(n919), .A2(n918), .ZN(n920) );
  NAND2_X1 U1024 ( .A1(n921), .A2(n920), .ZN(n924) );
  XOR2_X1 U1025 ( .A(G27), .B(n922), .Z(n923) );
  NOR2_X1 U1026 ( .A1(n924), .A2(n923), .ZN(n925) );
  XNOR2_X1 U1027 ( .A(n926), .B(n925), .ZN(n927) );
  NAND2_X1 U1028 ( .A1(n928), .A2(n927), .ZN(n931) );
  XNOR2_X1 U1029 ( .A(G34), .B(G2084), .ZN(n929) );
  XNOR2_X1 U1030 ( .A(KEYINPUT54), .B(n929), .ZN(n930) );
  NOR2_X1 U1031 ( .A1(n931), .A2(n930), .ZN(n932) );
  OR2_X1 U1032 ( .A1(G29), .A2(n932), .ZN(n933) );
  XNOR2_X1 U1033 ( .A(n934), .B(n933), .ZN(n960) );
  INV_X1 U1034 ( .A(n935), .ZN(n936) );
  NAND2_X1 U1035 ( .A1(n937), .A2(n936), .ZN(n957) );
  XOR2_X1 U1036 ( .A(G164), .B(G2078), .Z(n940) );
  XNOR2_X1 U1037 ( .A(G2072), .B(n938), .ZN(n939) );
  NOR2_X1 U1038 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1039 ( .A(KEYINPUT50), .B(n941), .ZN(n955) );
  XOR2_X1 U1040 ( .A(G2084), .B(G160), .Z(n942) );
  XNOR2_X1 U1041 ( .A(KEYINPUT118), .B(n942), .ZN(n943) );
  NOR2_X1 U1042 ( .A1(n944), .A2(n943), .ZN(n948) );
  NOR2_X1 U1043 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1044 ( .A1(n948), .A2(n947), .ZN(n953) );
  XOR2_X1 U1045 ( .A(G2090), .B(G162), .Z(n949) );
  NOR2_X1 U1046 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1047 ( .A(n951), .B(KEYINPUT51), .ZN(n952) );
  NOR2_X1 U1048 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1049 ( .A1(n955), .A2(n954), .ZN(n956) );
  NOR2_X1 U1050 ( .A1(n957), .A2(n956), .ZN(n958) );
  XOR2_X1 U1051 ( .A(n958), .B(KEYINPUT52), .Z(n959) );
  NAND2_X1 U1052 ( .A1(n960), .A2(n519), .ZN(n1019) );
  XNOR2_X1 U1053 ( .A(G16), .B(KEYINPUT56), .ZN(n988) );
  XNOR2_X1 U1054 ( .A(G1966), .B(G168), .ZN(n962) );
  NAND2_X1 U1055 ( .A1(n962), .A2(n961), .ZN(n964) );
  XOR2_X1 U1056 ( .A(KEYINPUT57), .B(KEYINPUT121), .Z(n963) );
  XNOR2_X1 U1057 ( .A(n964), .B(n963), .ZN(n986) );
  XNOR2_X1 U1058 ( .A(G171), .B(G1961), .ZN(n968) );
  XNOR2_X1 U1059 ( .A(G1956), .B(G299), .ZN(n965) );
  NOR2_X1 U1060 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1061 ( .A1(n968), .A2(n967), .ZN(n971) );
  NOR2_X1 U1062 ( .A1(G1348), .A2(n969), .ZN(n970) );
  NOR2_X1 U1063 ( .A1(n971), .A2(n970), .ZN(n981) );
  XOR2_X1 U1064 ( .A(n972), .B(KEYINPUT122), .Z(n974) );
  NAND2_X1 U1065 ( .A1(n974), .A2(n973), .ZN(n975) );
  XNOR2_X1 U1066 ( .A(n975), .B(KEYINPUT123), .ZN(n977) );
  NAND2_X1 U1067 ( .A1(n977), .A2(n976), .ZN(n979) );
  XNOR2_X1 U1068 ( .A(G1971), .B(G303), .ZN(n978) );
  NOR2_X1 U1069 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1070 ( .A1(n981), .A2(n980), .ZN(n984) );
  XNOR2_X1 U1071 ( .A(G1341), .B(n982), .ZN(n983) );
  NOR2_X1 U1072 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1073 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1074 ( .A1(n988), .A2(n987), .ZN(n1016) );
  INV_X1 U1075 ( .A(G16), .ZN(n1014) );
  XNOR2_X1 U1076 ( .A(KEYINPUT125), .B(G1966), .ZN(n989) );
  XNOR2_X1 U1077 ( .A(n989), .B(G21), .ZN(n1009) );
  XOR2_X1 U1078 ( .A(G1976), .B(KEYINPUT126), .Z(n990) );
  XNOR2_X1 U1079 ( .A(G23), .B(n990), .ZN(n994) );
  XNOR2_X1 U1080 ( .A(G1986), .B(G24), .ZN(n992) );
  XNOR2_X1 U1081 ( .A(G1971), .B(G22), .ZN(n991) );
  NOR2_X1 U1082 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1083 ( .A1(n994), .A2(n993), .ZN(n995) );
  XNOR2_X1 U1084 ( .A(n995), .B(KEYINPUT58), .ZN(n1007) );
  XNOR2_X1 U1085 ( .A(G20), .B(n996), .ZN(n1000) );
  XNOR2_X1 U1086 ( .A(G1341), .B(G19), .ZN(n998) );
  XNOR2_X1 U1087 ( .A(G6), .B(G1981), .ZN(n997) );
  NOR2_X1 U1088 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1089 ( .A1(n1000), .A2(n999), .ZN(n1003) );
  XOR2_X1 U1090 ( .A(KEYINPUT59), .B(G1348), .Z(n1001) );
  XNOR2_X1 U1091 ( .A(G4), .B(n1001), .ZN(n1002) );
  NOR2_X1 U1092 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XOR2_X1 U1093 ( .A(n1004), .B(KEYINPUT60), .Z(n1005) );
  XNOR2_X1 U1094 ( .A(KEYINPUT124), .B(n1005), .ZN(n1006) );
  NOR2_X1 U1095 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1096 ( .A1(n1009), .A2(n1008), .ZN(n1011) );
  XNOR2_X1 U1097 ( .A(G5), .B(G1961), .ZN(n1010) );
  NOR2_X1 U1098 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1099 ( .A(KEYINPUT61), .B(n1012), .ZN(n1013) );
  NAND2_X1 U1100 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1101 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XOR2_X1 U1102 ( .A(KEYINPUT127), .B(n1017), .Z(n1018) );
  NOR2_X1 U1103 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1104 ( .A1(n1020), .A2(G11), .ZN(n1021) );
  XOR2_X1 U1105 ( .A(KEYINPUT62), .B(n1021), .Z(G311) );
  INV_X1 U1106 ( .A(G311), .ZN(G150) );
endmodule

