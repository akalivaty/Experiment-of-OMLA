//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 0 0 0 0 0 1 1 1 1 0 1 1 0 1 1 0 0 0 1 0 0 0 0 0 1 0 0 1 0 1 0 0 0 1 1 1 1 1 0 1 0 1 0 0 0 0 1 0 1 1 0 0 1 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:12 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1229, new_n1230, new_n1231,
    new_n1232, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1280, new_n1281,
    new_n1282, new_n1283, new_n1284;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  AOI22_X1  g0003(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n204));
  INV_X1    g0004(.A(G68), .ZN(new_n205));
  INV_X1    g0005(.A(G238), .ZN(new_n206));
  INV_X1    g0006(.A(G77), .ZN(new_n207));
  INV_X1    g0007(.A(G244), .ZN(new_n208));
  OAI221_X1 g0008(.A(new_n204), .B1(new_n205), .B2(new_n206), .C1(new_n207), .C2(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n209), .A2(KEYINPUT66), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n212));
  NAND3_X1  g0012(.A1(new_n210), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n209), .A2(KEYINPUT66), .ZN(new_n214));
  OAI21_X1  g0014(.A(new_n203), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT67), .ZN(new_n216));
  INV_X1    g0016(.A(KEYINPUT1), .ZN(new_n217));
  OR2_X1    g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n216), .A2(new_n217), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n203), .A2(G13), .ZN(new_n220));
  OAI211_X1 g0020(.A(new_n220), .B(G250), .C1(G257), .C2(G264), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT64), .Z(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT0), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G13), .ZN(new_n224));
  INV_X1    g0024(.A(G20), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NOR2_X1   g0026(.A1(G58), .A2(G68), .ZN(new_n227));
  INV_X1    g0027(.A(KEYINPUT65), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(KEYINPUT65), .B1(G58), .B2(G68), .ZN(new_n230));
  NAND3_X1  g0030(.A1(new_n229), .A2(G50), .A3(new_n230), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n223), .B1(new_n226), .B2(new_n232), .ZN(new_n233));
  AND3_X1   g0033(.A1(new_n218), .A2(new_n219), .A3(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT68), .ZN(new_n236));
  XOR2_X1   g0036(.A(G264), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  INV_X1    g0039(.A(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(KEYINPUT2), .B(G226), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n238), .B(new_n243), .ZN(G358));
  XOR2_X1   g0044(.A(G68), .B(G77), .Z(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G58), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G107), .B(G116), .Z(new_n248));
  XNOR2_X1  g0048(.A(G87), .B(G97), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  INV_X1    g0051(.A(G41), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(KEYINPUT69), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT69), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(G41), .ZN(new_n255));
  INV_X1    g0055(.A(G45), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n253), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  AND2_X1   g0057(.A1(G33), .A2(G41), .ZN(new_n258));
  OAI21_X1  g0058(.A(KEYINPUT70), .B1(new_n258), .B2(new_n224), .ZN(new_n259));
  NAND2_X1  g0059(.A1(G33), .A2(G41), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT70), .ZN(new_n261));
  NAND4_X1  g0061(.A1(new_n260), .A2(new_n261), .A3(G1), .A4(G13), .ZN(new_n262));
  INV_X1    g0062(.A(G1), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G274), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  NAND4_X1  g0065(.A1(new_n257), .A2(new_n259), .A3(new_n262), .A4(new_n265), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n263), .B1(G41), .B2(G45), .ZN(new_n267));
  NAND4_X1  g0067(.A1(new_n259), .A2(G232), .A3(new_n262), .A4(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G190), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n258), .A2(new_n224), .ZN(new_n272));
  AND2_X1   g0072(.A1(KEYINPUT3), .A2(G33), .ZN(new_n273));
  NOR2_X1   g0073(.A1(KEYINPUT3), .A2(G33), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G1698), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(KEYINPUT72), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT72), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G1698), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n277), .A2(new_n279), .A3(G223), .ZN(new_n280));
  NAND2_X1  g0080(.A1(G226), .A2(G1698), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n275), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G33), .ZN(new_n283));
  INV_X1    g0083(.A(G87), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n272), .B1(new_n282), .B2(new_n285), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n270), .A2(new_n271), .A3(new_n286), .ZN(new_n287));
  XNOR2_X1  g0087(.A(KEYINPUT72), .B(G1698), .ZN(new_n288));
  AOI22_X1  g0088(.A1(new_n288), .A2(G223), .B1(G226), .B2(G1698), .ZN(new_n289));
  OAI22_X1  g0089(.A1(new_n289), .A2(new_n275), .B1(new_n283), .B2(new_n284), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n269), .B1(new_n290), .B2(new_n272), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n287), .B1(new_n291), .B2(G200), .ZN(new_n292));
  NAND3_X1  g0092(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT74), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND4_X1  g0095(.A1(KEYINPUT74), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n295), .A2(new_n224), .A3(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G13), .ZN(new_n298));
  NOR3_X1   g0098(.A1(new_n298), .A2(new_n225), .A3(G1), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  XNOR2_X1  g0100(.A(KEYINPUT8), .B(G58), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n301), .B1(new_n263), .B2(G20), .ZN(new_n302));
  AOI22_X1  g0102(.A1(new_n300), .A2(new_n302), .B1(new_n299), .B2(new_n301), .ZN(new_n303));
  INV_X1    g0103(.A(G58), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n304), .A2(new_n205), .ZN(new_n305));
  OAI21_X1  g0105(.A(G20), .B1(new_n305), .B2(new_n227), .ZN(new_n306));
  NOR2_X1   g0106(.A1(G20), .A2(G33), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(G159), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  AOI21_X1  g0109(.A(KEYINPUT7), .B1(new_n275), .B2(new_n225), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT7), .ZN(new_n311));
  NOR4_X1   g0111(.A1(new_n273), .A2(new_n274), .A3(new_n311), .A4(G20), .ZN(new_n312));
  OAI21_X1  g0112(.A(G68), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT82), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n309), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  OR2_X1    g0115(.A1(KEYINPUT3), .A2(G33), .ZN(new_n316));
  NAND2_X1  g0116(.A1(KEYINPUT3), .A2(G33), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n316), .A2(new_n225), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(new_n311), .ZN(new_n319));
  NAND4_X1  g0119(.A1(new_n316), .A2(KEYINPUT7), .A3(new_n225), .A4(new_n317), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n205), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(KEYINPUT82), .ZN(new_n322));
  AOI21_X1  g0122(.A(KEYINPUT16), .B1(new_n315), .B2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n309), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n313), .A2(KEYINPUT16), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(new_n297), .ZN(new_n326));
  OAI211_X1 g0126(.A(new_n292), .B(new_n303), .C1(new_n323), .C2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT17), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n303), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT16), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n324), .B1(new_n321), .B2(KEYINPUT82), .ZN(new_n332));
  AOI211_X1 g0132(.A(new_n314), .B(new_n205), .C1(new_n319), .C2(new_n320), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n331), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(new_n297), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n321), .A2(new_n309), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n335), .B1(new_n336), .B2(KEYINPUT16), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n330), .B1(new_n334), .B2(new_n337), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n270), .A2(G179), .A3(new_n286), .ZN(new_n339));
  INV_X1    g0139(.A(G169), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n339), .B1(new_n291), .B2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  OAI21_X1  g0142(.A(KEYINPUT18), .B1(new_n338), .B2(new_n342), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n303), .B1(new_n323), .B2(new_n326), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT18), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n344), .A2(new_n345), .A3(new_n341), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n338), .A2(KEYINPUT17), .A3(new_n292), .ZN(new_n347));
  NAND4_X1  g0147(.A1(new_n329), .A2(new_n343), .A3(new_n346), .A4(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n316), .A2(new_n317), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n350), .B1(new_n206), .B2(new_n276), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n351), .B1(G232), .B2(new_n288), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n272), .B1(new_n350), .B2(G107), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n266), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n259), .A2(new_n262), .A3(new_n267), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(KEYINPUT71), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT71), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n259), .A2(new_n357), .A3(new_n262), .A4(new_n267), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n208), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n354), .A2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(new_n340), .ZN(new_n362));
  INV_X1    g0162(.A(G179), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n360), .A2(new_n363), .ZN(new_n364));
  XNOR2_X1  g0164(.A(KEYINPUT15), .B(G87), .ZN(new_n365));
  INV_X1    g0165(.A(new_n365), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n283), .A2(G20), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT77), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n369), .B1(new_n225), .B2(new_n207), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  XNOR2_X1  g0171(.A(new_n301), .B(KEYINPUT76), .ZN(new_n372));
  INV_X1    g0172(.A(new_n307), .ZN(new_n373));
  OAI221_X1 g0173(.A(new_n371), .B1(KEYINPUT77), .B2(new_n368), .C1(new_n372), .C2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(new_n297), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n263), .A2(G20), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n300), .A2(G77), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n299), .A2(new_n207), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n375), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  AND3_X1   g0179(.A1(new_n362), .A2(new_n364), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n361), .A2(G200), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n379), .B1(G190), .B2(new_n360), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n380), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  AND2_X1   g0183(.A1(new_n349), .A2(new_n383), .ZN(new_n384));
  OAI211_X1 g0184(.A(new_n277), .B(new_n279), .C1(new_n273), .C2(new_n274), .ZN(new_n385));
  INV_X1    g0185(.A(G222), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  XNOR2_X1  g0187(.A(new_n387), .B(KEYINPUT73), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n350), .A2(G223), .A3(G1698), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n389), .B1(new_n207), .B2(new_n350), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n272), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n356), .A2(new_n358), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(G226), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n391), .A2(new_n266), .A3(new_n393), .ZN(new_n394));
  OR2_X1    g0194(.A1(new_n394), .A2(G179), .ZN(new_n395));
  NOR2_X1   g0195(.A1(G50), .A2(G58), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n225), .B1(new_n396), .B2(new_n205), .ZN(new_n397));
  XOR2_X1   g0197(.A(new_n397), .B(KEYINPUT75), .Z(new_n398));
  INV_X1    g0198(.A(new_n301), .ZN(new_n399));
  AOI22_X1  g0199(.A1(new_n399), .A2(new_n367), .B1(G150), .B2(new_n307), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(G50), .ZN(new_n402));
  AOI22_X1  g0202(.A1(new_n401), .A2(new_n297), .B1(new_n402), .B2(new_n299), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n300), .A2(G50), .A3(new_n376), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n394), .A2(new_n340), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n395), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT9), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n405), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n403), .A2(KEYINPUT9), .A3(new_n404), .ZN(new_n411));
  AND2_X1   g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT10), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n394), .A2(G200), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n391), .A2(G190), .A3(new_n266), .A4(new_n393), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n412), .A2(new_n413), .A3(new_n414), .A4(new_n415), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n414), .A2(new_n410), .A3(new_n415), .A4(new_n411), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(KEYINPUT10), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n408), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  AND3_X1   g0219(.A1(KEYINPUT78), .A2(G33), .A3(G97), .ZN(new_n420));
  AOI21_X1  g0220(.A(KEYINPUT78), .B1(G33), .B2(G97), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n277), .A2(new_n279), .ZN(new_n424));
  INV_X1    g0224(.A(G226), .ZN(new_n425));
  OAI22_X1  g0225(.A1(new_n424), .A2(new_n425), .B1(new_n240), .B2(new_n276), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n423), .B1(new_n426), .B2(new_n350), .ZN(new_n427));
  INV_X1    g0227(.A(new_n272), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n266), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n206), .B1(new_n356), .B2(new_n358), .ZN(new_n430));
  OAI21_X1  g0230(.A(KEYINPUT13), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  AOI22_X1  g0231(.A1(new_n288), .A2(G226), .B1(G232), .B2(G1698), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n422), .B1(new_n432), .B2(new_n275), .ZN(new_n433));
  AND2_X1   g0233(.A1(new_n259), .A2(new_n262), .ZN(new_n434));
  XNOR2_X1  g0234(.A(KEYINPUT69), .B(G41), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n264), .B1(new_n435), .B2(new_n256), .ZN(new_n436));
  AOI22_X1  g0236(.A1(new_n433), .A2(new_n272), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n392), .A2(G238), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT13), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n437), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n340), .B1(new_n431), .B2(new_n440), .ZN(new_n441));
  OR2_X1    g0241(.A1(new_n441), .A2(KEYINPUT14), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(KEYINPUT14), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  OAI21_X1  g0244(.A(KEYINPUT80), .B1(new_n429), .B2(new_n430), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT80), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n437), .A2(new_n438), .A3(new_n446), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n445), .A2(new_n447), .A3(KEYINPUT13), .ZN(new_n448));
  AND2_X1   g0248(.A1(new_n448), .A2(new_n440), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(G179), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n444), .A2(new_n450), .ZN(new_n451));
  AOI22_X1  g0251(.A1(new_n367), .A2(G77), .B1(G20), .B2(new_n205), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n452), .B1(new_n402), .B2(new_n373), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(new_n297), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT81), .ZN(new_n455));
  XNOR2_X1  g0255(.A(new_n454), .B(new_n455), .ZN(new_n456));
  OR2_X1    g0256(.A1(new_n456), .A2(KEYINPUT11), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(KEYINPUT11), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n299), .A2(new_n205), .ZN(new_n459));
  XNOR2_X1  g0259(.A(new_n459), .B(KEYINPUT12), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n300), .A2(G68), .A3(new_n376), .ZN(new_n461));
  AND2_X1   g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n457), .A2(new_n458), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n451), .A2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(new_n463), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n448), .A2(G190), .A3(new_n440), .ZN(new_n466));
  INV_X1    g0266(.A(G200), .ZN(new_n467));
  AOI211_X1 g0267(.A(KEYINPUT79), .B(new_n467), .C1(new_n431), .C2(new_n440), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT79), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n431), .A2(new_n440), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n469), .B1(new_n470), .B2(G200), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n465), .B(new_n466), .C1(new_n468), .C2(new_n471), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n384), .A2(new_n419), .A3(new_n464), .A4(new_n472), .ZN(new_n473));
  OAI211_X1 g0273(.A(G250), .B(G1698), .C1(new_n273), .C2(new_n274), .ZN(new_n474));
  NAND2_X1  g0274(.A1(G33), .A2(G283), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n385), .A2(new_n208), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n476), .B1(new_n477), .B2(KEYINPUT4), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n350), .A2(new_n288), .A3(G244), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT4), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n479), .A2(KEYINPUT83), .A3(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  AOI21_X1  g0282(.A(KEYINPUT83), .B1(new_n479), .B2(new_n480), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n478), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(new_n272), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n252), .A2(KEYINPUT5), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n259), .A2(G274), .A3(new_n262), .A4(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT84), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT5), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n254), .A2(G41), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n252), .A2(KEYINPUT69), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n490), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n256), .A2(G1), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n489), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  AOI21_X1  g0295(.A(KEYINPUT5), .B1(new_n253), .B2(new_n255), .ZN(new_n496));
  INV_X1    g0296(.A(new_n494), .ZN(new_n497));
  NOR3_X1   g0297(.A1(new_n496), .A2(KEYINPUT84), .A3(new_n497), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n488), .B1(new_n495), .B2(new_n498), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n486), .B(new_n494), .C1(new_n435), .C2(KEYINPUT5), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n434), .A2(new_n500), .A3(G257), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n485), .A2(new_n503), .A3(G190), .ZN(new_n504));
  INV_X1    g0304(.A(G107), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n505), .A2(KEYINPUT6), .A3(G97), .ZN(new_n506));
  INV_X1    g0306(.A(G97), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n507), .A2(new_n505), .ZN(new_n508));
  NOR2_X1   g0308(.A1(G97), .A2(G107), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n506), .B1(new_n510), .B2(KEYINPUT6), .ZN(new_n511));
  AOI22_X1  g0311(.A1(new_n511), .A2(G20), .B1(G77), .B2(new_n307), .ZN(new_n512));
  OAI21_X1  g0312(.A(G107), .B1(new_n310), .B2(new_n312), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n335), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n299), .A2(new_n507), .ZN(new_n515));
  AOI22_X1  g0315(.A1(new_n293), .A2(new_n294), .B1(G1), .B2(G13), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n298), .A2(G1), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(G20), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n263), .A2(G33), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n516), .A2(new_n518), .A3(new_n296), .A4(new_n519), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n515), .B1(new_n520), .B2(new_n507), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n514), .A2(new_n521), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n480), .B1(new_n385), .B2(new_n208), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT83), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n481), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n428), .B1(new_n526), .B2(new_n478), .ZN(new_n527));
  INV_X1    g0327(.A(new_n501), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n493), .A2(new_n489), .A3(new_n494), .ZN(new_n529));
  OAI21_X1  g0329(.A(KEYINPUT84), .B1(new_n496), .B2(new_n497), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n487), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  OAI21_X1  g0331(.A(KEYINPUT85), .B1(new_n528), .B2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT85), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n499), .A2(new_n533), .A3(new_n501), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n527), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n504), .B(new_n522), .C1(new_n535), .C2(new_n467), .ZN(new_n536));
  NOR3_X1   g0336(.A1(new_n528), .A2(new_n531), .A3(KEYINPUT85), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n533), .B1(new_n499), .B2(new_n501), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n485), .B(new_n363), .C1(new_n537), .C2(new_n538), .ZN(new_n539));
  OR2_X1    g0339(.A1(new_n514), .A2(new_n521), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n340), .B1(new_n527), .B2(new_n502), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n536), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(KEYINPUT86), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n434), .A2(new_n500), .A3(G264), .ZN(new_n545));
  OAI211_X1 g0345(.A(G257), .B(G1698), .C1(new_n273), .C2(new_n274), .ZN(new_n546));
  NAND2_X1  g0346(.A1(G33), .A2(G294), .ZN(new_n547));
  INV_X1    g0347(.A(G250), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n546), .B(new_n547), .C1(new_n385), .C2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n272), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n499), .A2(new_n545), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(new_n340), .ZN(new_n552));
  AND2_X1   g0352(.A1(new_n550), .A2(new_n545), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n553), .A2(new_n363), .A3(new_n499), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n299), .A2(new_n505), .ZN(new_n556));
  XNOR2_X1  g0356(.A(new_n556), .B(KEYINPUT25), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n520), .A2(new_n505), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(new_n559), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n225), .B(G87), .C1(new_n273), .C2(new_n274), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(KEYINPUT22), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT22), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n350), .A2(new_n563), .A3(new_n225), .A4(G87), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(G33), .A2(G116), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n566), .A2(G20), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT23), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n568), .B1(new_n225), .B2(G107), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n505), .A2(KEYINPUT23), .A3(G20), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n567), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n565), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(KEYINPUT24), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT24), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n565), .A2(new_n574), .A3(new_n571), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n560), .B1(new_n576), .B2(new_n297), .ZN(new_n577));
  OAI21_X1  g0377(.A(KEYINPUT91), .B1(new_n555), .B2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(new_n575), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n574), .B1(new_n565), .B2(new_n571), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n297), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(new_n559), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT91), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n582), .A2(new_n583), .A3(new_n554), .A4(new_n552), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n366), .A2(new_n518), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n520), .A2(new_n284), .ZN(new_n586));
  XNOR2_X1  g0386(.A(KEYINPUT87), .B(G87), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n509), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT19), .ZN(new_n589));
  NAND2_X1  g0389(.A1(G33), .A2(G97), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT78), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(KEYINPUT78), .A2(G33), .A3(G97), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n589), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n588), .B1(new_n594), .B2(G20), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(KEYINPUT88), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT88), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n588), .B(new_n597), .C1(new_n594), .C2(G20), .ZN(new_n598));
  AOI21_X1  g0398(.A(KEYINPUT19), .B1(new_n367), .B2(G97), .ZN(new_n599));
  AOI21_X1  g0399(.A(G20), .B1(new_n316), .B2(new_n317), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n599), .B1(G68), .B2(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n596), .A2(new_n598), .A3(new_n601), .ZN(new_n602));
  AOI211_X1 g0402(.A(new_n585), .B(new_n586), .C1(new_n602), .C2(new_n297), .ZN(new_n603));
  OAI211_X1 g0403(.A(G244), .B(G1698), .C1(new_n273), .C2(new_n274), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n566), .B(new_n604), .C1(new_n385), .C2(new_n206), .ZN(new_n605));
  OAI22_X1  g0405(.A1(new_n494), .A2(new_n548), .B1(new_n264), .B2(new_n256), .ZN(new_n606));
  AOI22_X1  g0406(.A1(new_n605), .A2(new_n272), .B1(new_n434), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n271), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n608), .B1(G200), .B2(new_n607), .ZN(new_n609));
  OAI21_X1  g0409(.A(KEYINPUT19), .B1(new_n420), .B2(new_n421), .ZN(new_n610));
  AOI22_X1  g0410(.A1(new_n610), .A2(new_n225), .B1(new_n509), .B2(new_n587), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n601), .B1(new_n611), .B2(new_n597), .ZN(new_n612));
  INV_X1    g0412(.A(new_n598), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n297), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(new_n585), .ZN(new_n615));
  XNOR2_X1  g0415(.A(new_n365), .B(KEYINPUT89), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n616), .A2(new_n300), .A3(new_n519), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n614), .A2(new_n615), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n607), .A2(G179), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n619), .B1(new_n340), .B2(new_n607), .ZN(new_n620));
  AOI22_X1  g0420(.A1(new_n603), .A2(new_n609), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n553), .A2(G190), .A3(new_n499), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n551), .A2(G200), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n577), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  AND4_X1   g0424(.A1(new_n578), .A2(new_n584), .A3(new_n621), .A4(new_n624), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n434), .A2(new_n500), .A3(G270), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n350), .A2(new_n288), .A3(G257), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n350), .A2(G264), .A3(G1698), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n275), .A2(G303), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n627), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(new_n272), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n499), .A2(new_n626), .A3(new_n631), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n632), .A2(KEYINPUT21), .A3(G169), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n529), .A2(new_n530), .ZN(new_n634));
  AOI22_X1  g0434(.A1(new_n634), .A2(new_n488), .B1(new_n630), .B2(new_n272), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n635), .A2(G179), .A3(new_n626), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n633), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n520), .A2(G116), .ZN(new_n638));
  INV_X1    g0438(.A(G116), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n518), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(G20), .B1(G33), .B2(G283), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n283), .A2(G97), .ZN(new_n643));
  AOI22_X1  g0443(.A1(new_n642), .A2(new_n643), .B1(G20), .B2(new_n639), .ZN(new_n644));
  AOI21_X1  g0444(.A(KEYINPUT20), .B1(new_n297), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n297), .A2(new_n644), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT20), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n641), .B1(new_n645), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n637), .A2(new_n649), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n649), .B1(new_n632), .B2(G200), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n651), .B1(new_n271), .B2(new_n632), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n632), .A2(new_n649), .A3(G169), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT21), .ZN(new_n654));
  AND3_X1   g0454(.A1(new_n653), .A2(KEYINPUT90), .A3(new_n654), .ZN(new_n655));
  AOI21_X1  g0455(.A(KEYINPUT90), .B1(new_n653), .B2(new_n654), .ZN(new_n656));
  OAI211_X1 g0456(.A(new_n650), .B(new_n652), .C1(new_n655), .C2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT86), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n536), .A2(new_n542), .A3(new_n659), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n544), .A2(new_n625), .A3(new_n658), .A4(new_n660), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n473), .A2(new_n661), .ZN(G372));
  NAND2_X1  g0462(.A1(new_n416), .A2(new_n418), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n329), .A2(new_n347), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n472), .A2(new_n380), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n664), .B1(new_n464), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n343), .A2(new_n346), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n663), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n668), .A2(new_n407), .ZN(new_n669));
  INV_X1    g0469(.A(new_n473), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT92), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n582), .A2(new_n554), .A3(new_n552), .ZN(new_n672));
  OAI211_X1 g0472(.A(new_n650), .B(new_n672), .C1(new_n655), .C2(new_n656), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n536), .A2(new_n542), .A3(new_n624), .A4(new_n621), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n671), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n527), .A2(new_n502), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n540), .B1(new_n677), .B2(G190), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n485), .B1(new_n537), .B2(new_n538), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(G200), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n485), .A2(new_n503), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n522), .B1(new_n681), .B2(new_n340), .ZN(new_n682));
  AOI22_X1  g0482(.A1(new_n678), .A2(new_n680), .B1(new_n682), .B2(new_n539), .ZN(new_n683));
  AND2_X1   g0483(.A1(new_n621), .A2(new_n624), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n683), .A2(new_n684), .A3(new_n673), .A4(KEYINPUT92), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT26), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n603), .A2(new_n609), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n618), .A2(new_n620), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n686), .B1(new_n689), .B2(new_n542), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n621), .A2(new_n682), .A3(KEYINPUT26), .A4(new_n539), .ZN(new_n691));
  AOI22_X1  g0491(.A1(new_n690), .A2(new_n691), .B1(new_n618), .B2(new_n620), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n676), .A2(new_n685), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n670), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n669), .A2(new_n694), .ZN(G369));
  OAI21_X1  g0495(.A(new_n650), .B1(new_n655), .B2(new_n656), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n517), .A2(new_n225), .ZN(new_n698));
  OR2_X1    g0498(.A1(new_n698), .A2(KEYINPUT27), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(KEYINPUT27), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n699), .A2(new_n700), .A3(G213), .ZN(new_n701));
  INV_X1    g0501(.A(G343), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n649), .A2(new_n703), .ZN(new_n704));
  MUX2_X1   g0504(.A(new_n697), .B(new_n657), .S(new_n704), .Z(new_n705));
  XNOR2_X1  g0505(.A(new_n705), .B(KEYINPUT93), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(G330), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  AND3_X1   g0508(.A1(new_n578), .A2(new_n584), .A3(new_n624), .ZN(new_n709));
  INV_X1    g0509(.A(new_n703), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n709), .B1(new_n577), .B2(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n711), .B1(new_n672), .B2(new_n710), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n708), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n672), .A2(new_n703), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n697), .A2(new_n703), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n714), .B1(new_n715), .B2(new_n709), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n713), .A2(new_n716), .ZN(G399));
  INV_X1    g0517(.A(new_n435), .ZN(new_n718));
  INV_X1    g0518(.A(new_n220), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n588), .A2(G116), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n721), .A2(new_n722), .A3(G1), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n723), .B1(new_n231), .B2(new_n721), .ZN(new_n724));
  XNOR2_X1  g0524(.A(new_n724), .B(KEYINPUT28), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n693), .A2(new_n710), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT29), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n578), .A2(new_n584), .ZN(new_n729));
  OAI211_X1 g0529(.A(new_n683), .B(new_n684), .C1(new_n729), .C2(new_n696), .ZN(new_n730));
  AOI211_X1 g0530(.A(new_n727), .B(new_n703), .C1(new_n692), .C2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n728), .A2(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n607), .A2(G179), .ZN(new_n734));
  AND2_X1   g0534(.A1(new_n551), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n679), .A2(new_n632), .A3(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT30), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n605), .A2(new_n272), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n434), .A2(new_n606), .ZN(new_n739));
  AND3_X1   g0539(.A1(new_n738), .A2(G179), .A3(new_n739), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n740), .A2(new_n553), .A3(new_n635), .A4(new_n626), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n737), .B1(new_n681), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n550), .A2(new_n545), .ZN(new_n743));
  NOR3_X1   g0543(.A1(new_n632), .A2(new_n619), .A3(new_n743), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n744), .A2(new_n677), .A3(KEYINPUT30), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n736), .A2(new_n742), .A3(new_n745), .ZN(new_n746));
  AND3_X1   g0546(.A1(new_n746), .A2(KEYINPUT31), .A3(new_n703), .ZN(new_n747));
  AOI21_X1  g0547(.A(KEYINPUT31), .B1(new_n746), .B2(new_n703), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n749), .B1(new_n661), .B2(new_n703), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(G330), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n733), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n725), .B1(new_n753), .B2(G1), .ZN(G364));
  AOI21_X1  g0554(.A(new_n224), .B1(G20), .B2(new_n340), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n225), .A2(new_n363), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(G200), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(G190), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT32), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n225), .A2(G179), .ZN(new_n762));
  NOR2_X1   g0562(.A1(G190), .A2(G200), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(G159), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  OAI22_X1  g0566(.A1(new_n760), .A2(new_n205), .B1(new_n761), .B2(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(new_n761), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n762), .A2(G190), .A3(G200), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n768), .B1(new_n587), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n757), .A2(new_n763), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n757), .A2(G190), .A3(new_n467), .ZN(new_n772));
  OAI221_X1 g0572(.A(new_n350), .B1(new_n771), .B2(new_n207), .C1(new_n304), .C2(new_n772), .ZN(new_n773));
  NOR3_X1   g0573(.A1(new_n767), .A2(new_n770), .A3(new_n773), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n762), .A2(new_n271), .A3(G200), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(new_n505), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n758), .A2(new_n271), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n776), .B1(G50), .B2(new_n777), .ZN(new_n778));
  NOR3_X1   g0578(.A1(new_n271), .A2(G179), .A3(G200), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(new_n225), .ZN(new_n780));
  OAI211_X1 g0580(.A(new_n774), .B(new_n778), .C1(new_n507), .C2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n772), .ZN(new_n782));
  INV_X1    g0582(.A(new_n764), .ZN(new_n783));
  AOI22_X1  g0583(.A1(new_n782), .A2(G322), .B1(new_n783), .B2(G329), .ZN(new_n784));
  INV_X1    g0584(.A(new_n771), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n350), .B1(new_n785), .B2(G311), .ZN(new_n786));
  AND2_X1   g0586(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n775), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(G283), .ZN(new_n789));
  INV_X1    g0589(.A(new_n780), .ZN(new_n790));
  XNOR2_X1  g0590(.A(KEYINPUT33), .B(G317), .ZN(new_n791));
  AOI22_X1  g0591(.A1(G294), .A2(new_n790), .B1(new_n759), .B2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n769), .ZN(new_n793));
  AOI22_X1  g0593(.A1(new_n777), .A2(G326), .B1(new_n793), .B2(G303), .ZN(new_n794));
  NAND4_X1  g0594(.A1(new_n787), .A2(new_n789), .A3(new_n792), .A4(new_n794), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n756), .B1(new_n781), .B2(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n298), .A2(G20), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n263), .B1(new_n797), .B2(G45), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n721), .A2(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(G13), .A2(G33), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(G20), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n802), .A2(new_n755), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n719), .A2(new_n350), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n806), .B1(new_n232), .B2(new_n256), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n807), .B1(new_n256), .B2(new_n247), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n350), .A2(new_n220), .ZN(new_n809));
  INV_X1    g0609(.A(G355), .ZN(new_n810));
  OAI22_X1  g0610(.A1(new_n809), .A2(new_n810), .B1(G116), .B2(new_n220), .ZN(new_n811));
  XNOR2_X1  g0611(.A(new_n811), .B(KEYINPUT94), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n804), .B1(new_n808), .B2(new_n812), .ZN(new_n813));
  NOR3_X1   g0613(.A1(new_n796), .A2(new_n799), .A3(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n802), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n814), .B1(new_n706), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n707), .A2(new_n799), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n706), .A2(G330), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n816), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  XNOR2_X1  g0619(.A(KEYINPUT95), .B(KEYINPUT96), .ZN(new_n820));
  XNOR2_X1  g0620(.A(new_n819), .B(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(G396));
  INV_X1    g0622(.A(new_n799), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n380), .A2(new_n710), .ZN(new_n824));
  AOI22_X1  g0624(.A1(new_n382), .A2(new_n381), .B1(new_n379), .B2(new_n703), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n824), .B1(new_n825), .B2(new_n380), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n726), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n693), .A2(new_n383), .A3(new_n710), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n823), .B1(new_n829), .B2(new_n751), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n830), .B1(new_n751), .B2(new_n829), .ZN(new_n831));
  AOI22_X1  g0631(.A1(new_n782), .A2(G143), .B1(new_n785), .B2(G159), .ZN(new_n832));
  INV_X1    g0632(.A(new_n777), .ZN(new_n833));
  INV_X1    g0633(.A(G137), .ZN(new_n834));
  INV_X1    g0634(.A(G150), .ZN(new_n835));
  OAI221_X1 g0635(.A(new_n832), .B1(new_n833), .B2(new_n834), .C1(new_n835), .C2(new_n760), .ZN(new_n836));
  XOR2_X1   g0636(.A(new_n836), .B(KEYINPUT34), .Z(new_n837));
  NAND2_X1  g0637(.A1(new_n788), .A2(G68), .ZN(new_n838));
  INV_X1    g0638(.A(G132), .ZN(new_n839));
  OAI211_X1 g0639(.A(new_n838), .B(new_n350), .C1(new_n839), .C2(new_n764), .ZN(new_n840));
  OAI22_X1  g0640(.A1(new_n780), .A2(new_n304), .B1(new_n769), .B2(new_n402), .ZN(new_n841));
  NOR3_X1   g0641(.A1(new_n837), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n775), .A2(new_n284), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n843), .B1(G303), .B2(new_n777), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n844), .B1(new_n505), .B2(new_n769), .ZN(new_n845));
  AOI22_X1  g0645(.A1(G116), .A2(new_n785), .B1(new_n783), .B2(G311), .ZN(new_n846));
  INV_X1    g0646(.A(G294), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n846), .B(new_n275), .C1(new_n847), .C2(new_n772), .ZN(new_n848));
  INV_X1    g0648(.A(G283), .ZN(new_n849));
  OAI22_X1  g0649(.A1(new_n760), .A2(new_n849), .B1(new_n507), .B2(new_n780), .ZN(new_n850));
  NOR3_X1   g0650(.A1(new_n845), .A2(new_n848), .A3(new_n850), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n755), .B1(new_n842), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n756), .A2(new_n801), .ZN(new_n853));
  OAI211_X1 g0653(.A(new_n852), .B(new_n823), .C1(G77), .C2(new_n853), .ZN(new_n854));
  XOR2_X1   g0654(.A(new_n854), .B(KEYINPUT97), .Z(new_n855));
  INV_X1    g0655(.A(new_n826), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n855), .B1(new_n801), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n831), .A2(new_n857), .ZN(G384));
  OR2_X1    g0658(.A1(new_n511), .A2(KEYINPUT35), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n511), .A2(KEYINPUT35), .ZN(new_n860));
  NAND4_X1  g0660(.A1(new_n859), .A2(G116), .A3(new_n226), .A4(new_n860), .ZN(new_n861));
  XOR2_X1   g0661(.A(new_n861), .B(KEYINPUT36), .Z(new_n862));
  NOR3_X1   g0662(.A1(new_n231), .A2(new_n207), .A3(new_n305), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(new_n864));
  OR2_X1    g0664(.A1(new_n864), .A2(KEYINPUT98), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n402), .A2(G68), .ZN(new_n866));
  XNOR2_X1  g0666(.A(new_n866), .B(KEYINPUT99), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n867), .B1(new_n864), .B2(KEYINPUT98), .ZN(new_n868));
  AOI211_X1 g0668(.A(new_n263), .B(G13), .C1(new_n865), .C2(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n862), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT39), .ZN(new_n871));
  XOR2_X1   g0671(.A(KEYINPUT101), .B(KEYINPUT38), .Z(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n344), .A2(new_n341), .ZN(new_n874));
  INV_X1    g0674(.A(new_n701), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n344), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n874), .A2(new_n876), .A3(new_n327), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(KEYINPUT37), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT37), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n874), .A2(new_n876), .A3(new_n879), .A4(new_n327), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n348), .A2(new_n344), .A3(new_n875), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n873), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n331), .B1(new_n321), .B2(new_n309), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n884), .A2(new_n325), .A3(new_n297), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n701), .B1(new_n885), .B2(new_n303), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n348), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n885), .A2(new_n303), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n888), .B1(new_n341), .B2(new_n875), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(new_n327), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(KEYINPUT37), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n880), .A2(new_n891), .ZN(new_n892));
  AND3_X1   g0692(.A1(new_n887), .A2(KEYINPUT38), .A3(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n871), .B1(new_n883), .B2(new_n893), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n887), .A2(KEYINPUT38), .A3(new_n892), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(KEYINPUT100), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT100), .ZN(new_n897));
  NAND4_X1  g0697(.A1(new_n887), .A2(new_n897), .A3(new_n892), .A4(KEYINPUT38), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n887), .A2(new_n892), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT38), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n896), .A2(new_n898), .A3(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n894), .B1(new_n902), .B2(new_n871), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n451), .A2(new_n463), .A3(new_n710), .ZN(new_n904));
  OR2_X1    g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n463), .A2(new_n703), .ZN(new_n906));
  AOI22_X1  g0706(.A1(new_n442), .A2(new_n443), .B1(new_n449), .B2(G179), .ZN(new_n907));
  OAI211_X1 g0707(.A(new_n472), .B(new_n906), .C1(new_n907), .C2(new_n465), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n451), .A2(new_n463), .A3(new_n703), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n911), .B1(new_n828), .B2(new_n824), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n902), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n667), .A2(new_n701), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n905), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n728), .A2(new_n670), .A3(new_n732), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(new_n669), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n915), .B(new_n917), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n826), .B1(new_n908), .B2(new_n909), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n902), .A2(new_n750), .A3(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT40), .ZN(new_n921));
  AND2_X1   g0721(.A1(new_n919), .A2(new_n750), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n881), .A2(new_n882), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n872), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n921), .B1(new_n924), .B2(new_n895), .ZN(new_n925));
  AOI22_X1  g0725(.A1(new_n920), .A2(new_n921), .B1(new_n922), .B2(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n926), .A2(new_n670), .A3(new_n750), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(G330), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n926), .B1(new_n670), .B2(new_n750), .ZN(new_n929));
  OR2_X1    g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n918), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n931), .B1(new_n263), .B2(new_n797), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n918), .A2(new_n930), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n870), .B1(new_n932), .B2(new_n933), .ZN(G367));
  OAI21_X1  g0734(.A(new_n683), .B1(new_n522), .B2(new_n710), .ZN(new_n935));
  INV_X1    g0735(.A(new_n542), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(new_n703), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n938), .A2(new_n715), .A3(new_n709), .ZN(new_n939));
  OR2_X1    g0739(.A1(new_n939), .A2(KEYINPUT42), .ZN(new_n940));
  AND2_X1   g0740(.A1(new_n729), .A2(new_n536), .ZN(new_n941));
  OR2_X1    g0741(.A1(new_n941), .A2(new_n936), .ZN(new_n942));
  AOI22_X1  g0742(.A1(new_n939), .A2(KEYINPUT42), .B1(new_n710), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n940), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(KEYINPUT103), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n944), .A2(KEYINPUT103), .ZN(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n603), .A2(new_n710), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n948), .A2(new_n618), .A3(new_n620), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n949), .B1(new_n689), .B2(new_n948), .ZN(new_n950));
  OR2_X1    g0750(.A1(new_n950), .A2(KEYINPUT102), .ZN(new_n951));
  AOI21_X1  g0751(.A(KEYINPUT43), .B1(new_n950), .B2(KEYINPUT102), .ZN(new_n952));
  NAND4_X1  g0752(.A1(new_n945), .A2(new_n947), .A3(new_n951), .A4(new_n952), .ZN(new_n953));
  AOI22_X1  g0753(.A1(new_n951), .A2(new_n952), .B1(KEYINPUT43), .B2(new_n950), .ZN(new_n954));
  INV_X1    g0754(.A(new_n945), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n954), .B1(new_n946), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n953), .A2(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(new_n713), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n958), .A2(new_n938), .ZN(new_n959));
  XOR2_X1   g0759(.A(new_n957), .B(new_n959), .Z(new_n960));
  XOR2_X1   g0760(.A(new_n720), .B(KEYINPUT41), .Z(new_n961));
  NOR2_X1   g0761(.A1(new_n716), .A2(new_n938), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n962), .B(KEYINPUT44), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n716), .A2(new_n938), .ZN(new_n964));
  XOR2_X1   g0764(.A(KEYINPUT104), .B(KEYINPUT45), .Z(new_n965));
  XNOR2_X1  g0765(.A(new_n964), .B(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n963), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n958), .A2(new_n967), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n713), .A2(new_n963), .A3(new_n966), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n715), .A2(new_n709), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n972), .B1(new_n712), .B2(new_n715), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n707), .B(new_n973), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n974), .A2(new_n752), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n971), .A2(new_n975), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n961), .B1(new_n976), .B2(new_n753), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n798), .B(KEYINPUT105), .ZN(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n960), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  AND2_X1   g0780(.A1(new_n238), .A2(new_n805), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n803), .B1(new_n220), .B2(new_n365), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n823), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n793), .A2(G116), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT46), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  XOR2_X1   g0786(.A(new_n986), .B(KEYINPUT107), .Z(new_n987));
  INV_X1    g0787(.A(G311), .ZN(new_n988));
  INV_X1    g0788(.A(G303), .ZN(new_n989));
  OAI22_X1  g0789(.A1(new_n833), .A2(new_n988), .B1(new_n989), .B2(new_n772), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT106), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n775), .A2(new_n507), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n780), .A2(new_n505), .ZN(new_n993));
  AOI211_X1 g0793(.A(new_n992), .B(new_n993), .C1(G294), .C2(new_n759), .ZN(new_n994));
  INV_X1    g0794(.A(G317), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n275), .B1(new_n764), .B2(new_n995), .C1(new_n849), .C2(new_n771), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n996), .B1(new_n985), .B2(new_n984), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n987), .A2(new_n991), .A3(new_n994), .A4(new_n997), .ZN(new_n998));
  OAI22_X1  g0798(.A1(new_n780), .A2(new_n205), .B1(new_n772), .B2(new_n835), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT108), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n999), .A2(new_n1000), .B1(G143), .B2(new_n777), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1001), .B1(new_n1000), .B2(new_n999), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1002), .B(KEYINPUT109), .ZN(new_n1003));
  OAI221_X1 g0803(.A(new_n350), .B1(new_n402), .B2(new_n771), .C1(new_n760), .C2(new_n765), .ZN(new_n1004));
  OAI22_X1  g0804(.A1(new_n769), .A2(new_n304), .B1(new_n764), .B2(new_n834), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT110), .ZN(new_n1006));
  AND2_X1   g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n775), .A2(new_n207), .ZN(new_n1008));
  NOR3_X1   g0808(.A1(new_n1004), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1009), .B1(new_n1006), .B2(new_n1005), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n998), .B1(new_n1003), .B2(new_n1010), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1011), .B(KEYINPUT47), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n983), .B1(new_n1012), .B2(new_n755), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(new_n815), .B2(new_n950), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n980), .A2(new_n1014), .ZN(G387));
  INV_X1    g0815(.A(new_n975), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n974), .A2(new_n752), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1016), .A2(new_n720), .A3(new_n1017), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n712), .A2(new_n815), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n722), .A2(new_n809), .B1(G107), .B2(new_n220), .ZN(new_n1020));
  XOR2_X1   g0820(.A(new_n1020), .B(KEYINPUT111), .Z(new_n1021));
  NOR2_X1   g0821(.A1(new_n372), .A2(G50), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT50), .ZN(new_n1023));
  AOI21_X1  g0823(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1023), .A2(new_n722), .A3(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n806), .B1(new_n243), .B2(G45), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1021), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n782), .A2(G317), .B1(new_n785), .B2(G303), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(KEYINPUT113), .B(G322), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n1028), .B1(new_n833), .B2(new_n1029), .C1(new_n988), .C2(new_n760), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT48), .ZN(new_n1031));
  OR2_X1    g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n790), .A2(G283), .B1(new_n793), .B2(G294), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1032), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT49), .ZN(new_n1036));
  OR2_X1    g0836(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n775), .A2(new_n639), .ZN(new_n1039));
  AOI211_X1 g0839(.A(new_n350), .B(new_n1039), .C1(G326), .C2(new_n783), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1037), .A2(new_n1038), .A3(new_n1040), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(KEYINPUT112), .B(G150), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n771), .A2(new_n205), .B1(new_n764), .B2(new_n1042), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n275), .B(new_n1043), .C1(G50), .C2(new_n782), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n992), .B1(G159), .B2(new_n777), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n759), .A2(new_n399), .B1(new_n793), .B2(G77), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n616), .A2(new_n790), .ZN(new_n1047));
  NAND4_X1  g0847(.A1(new_n1044), .A2(new_n1045), .A3(new_n1046), .A4(new_n1047), .ZN(new_n1048));
  AND2_X1   g0848(.A1(new_n1041), .A2(new_n1048), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n823), .B1(new_n804), .B2(new_n1027), .C1(new_n1049), .C2(new_n756), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n1018), .B1(new_n974), .B2(new_n978), .C1(new_n1019), .C2(new_n1050), .ZN(G393));
  NAND2_X1  g0851(.A1(new_n1016), .A2(new_n970), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n976), .A2(new_n720), .A3(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n971), .A2(new_n979), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n803), .B1(new_n507), .B2(new_n220), .C1(new_n250), .C2(new_n806), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1055), .A2(new_n823), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n790), .A2(G116), .B1(new_n785), .B2(G294), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1057), .B1(new_n989), .B2(new_n760), .ZN(new_n1058));
  XOR2_X1   g0858(.A(new_n1058), .B(KEYINPUT115), .Z(new_n1059));
  OAI22_X1  g0859(.A1(new_n833), .A2(new_n995), .B1(new_n988), .B2(new_n772), .ZN(new_n1060));
  XOR2_X1   g0860(.A(KEYINPUT114), .B(KEYINPUT52), .Z(new_n1061));
  OR2_X1    g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n793), .A2(G283), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n275), .B1(new_n764), .B2(new_n1029), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n1065), .A2(new_n776), .ZN(new_n1066));
  NAND4_X1  g0866(.A1(new_n1062), .A2(new_n1063), .A3(new_n1064), .A4(new_n1066), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(G150), .A2(new_n777), .B1(new_n782), .B2(G159), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1068), .B(KEYINPUT51), .ZN(new_n1069));
  AOI211_X1 g0869(.A(new_n275), .B(new_n843), .C1(G143), .C2(new_n783), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n790), .A2(G77), .ZN(new_n1071));
  OR2_X1    g0871(.A1(new_n372), .A2(new_n771), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n759), .A2(G50), .B1(new_n793), .B2(G68), .ZN(new_n1073));
  NAND4_X1  g0873(.A1(new_n1070), .A2(new_n1071), .A3(new_n1072), .A4(new_n1073), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n1059), .A2(new_n1067), .B1(new_n1069), .B2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1056), .B1(new_n1075), .B2(new_n755), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1076), .B1(new_n938), .B2(new_n815), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1053), .A2(new_n1054), .A3(new_n1077), .ZN(G390));
  INV_X1    g0878(.A(new_n904), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n903), .B1(new_n912), .B2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n703), .B1(new_n692), .B2(new_n730), .ZN(new_n1081));
  OR2_X1    g0881(.A1(new_n825), .A2(new_n380), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n1081), .A2(new_n1082), .B1(new_n380), .B2(new_n710), .ZN(new_n1083));
  OAI221_X1 g0883(.A(new_n904), .B1(new_n893), .B2(new_n883), .C1(new_n1083), .C2(new_n911), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1080), .A2(new_n1084), .ZN(new_n1085));
  NAND4_X1  g0885(.A1(new_n750), .A2(G330), .A3(new_n856), .A4(new_n910), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1080), .A2(new_n1086), .A3(new_n1084), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n670), .A2(G330), .A3(new_n750), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n916), .A2(new_n669), .A3(new_n1090), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n750), .A2(G330), .A3(new_n856), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(new_n911), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1093), .A2(new_n1086), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n828), .A2(new_n824), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1093), .A2(new_n1086), .A3(new_n1083), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1091), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g0898(.A(KEYINPUT116), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n1088), .B(new_n1089), .C1(new_n1098), .C2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(KEYINPUT29), .B1(new_n693), .B2(new_n710), .ZN(new_n1101));
  NOR3_X1   g0901(.A1(new_n1101), .A2(new_n473), .A3(new_n731), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n751), .A2(new_n473), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n668), .A2(new_n407), .ZN(new_n1104));
  NOR3_X1   g0904(.A1(new_n1102), .A2(new_n1103), .A3(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1097), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n1093), .A2(new_n1086), .B1(new_n824), .B2(new_n828), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1105), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  AND3_X1   g0908(.A1(new_n1080), .A2(new_n1086), .A3(new_n1084), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1086), .B1(new_n1080), .B2(new_n1084), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n1108), .B(KEYINPUT116), .C1(new_n1109), .C2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1100), .A2(new_n1111), .A3(new_n720), .ZN(new_n1112));
  OAI22_X1  g0912(.A1(new_n505), .A2(new_n760), .B1(new_n833), .B2(new_n849), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1113), .B1(G87), .B2(new_n793), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n772), .A2(new_n639), .B1(new_n771), .B2(new_n507), .ZN(new_n1115));
  AOI211_X1 g0915(.A(new_n350), .B(new_n1115), .C1(G294), .C2(new_n783), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n1114), .A2(new_n838), .A3(new_n1071), .A4(new_n1116), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(KEYINPUT54), .B(G143), .ZN(new_n1118));
  INV_X1    g0918(.A(G125), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n771), .A2(new_n1118), .B1(new_n764), .B2(new_n1119), .ZN(new_n1120));
  AOI211_X1 g0920(.A(new_n275), .B(new_n1120), .C1(G132), .C2(new_n782), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n769), .A2(new_n1042), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(new_n1122), .B(KEYINPUT53), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n777), .A2(G128), .B1(new_n788), .B2(G50), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(G159), .A2(new_n790), .B1(new_n759), .B2(G137), .ZN(new_n1125));
  NAND4_X1  g0925(.A1(new_n1121), .A2(new_n1123), .A3(new_n1124), .A4(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n756), .B1(new_n1117), .B2(new_n1126), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n823), .B1(new_n399), .B2(new_n853), .ZN(new_n1128));
  AOI211_X1 g0928(.A(new_n1127), .B(new_n1128), .C1(new_n903), .C2(new_n800), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1129), .B1(new_n1130), .B2(new_n979), .ZN(new_n1131));
  AND2_X1   g0931(.A1(new_n1131), .A2(KEYINPUT117), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n1131), .A2(KEYINPUT117), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1112), .B1(new_n1132), .B2(new_n1133), .ZN(G378));
  AND3_X1   g0934(.A1(new_n896), .A2(new_n898), .A3(new_n901), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n919), .A2(new_n750), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n921), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(KEYINPUT120), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n925), .A2(new_n750), .A3(new_n919), .ZN(new_n1139));
  NAND4_X1  g0939(.A1(new_n1137), .A2(new_n1138), .A3(G330), .A4(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n405), .A2(new_n875), .ZN(new_n1141));
  XOR2_X1   g0941(.A(new_n419), .B(new_n1141), .Z(new_n1142));
  XNOR2_X1  g0942(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(new_n1142), .B(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1140), .A2(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1138), .B1(new_n926), .B2(G330), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  XNOR2_X1  g0948(.A(new_n1142), .B(new_n1143), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1137), .A2(G330), .A3(new_n1139), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1149), .A2(new_n1150), .A3(KEYINPUT120), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n915), .B1(new_n1148), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1150), .A2(KEYINPUT120), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1154), .A2(new_n1140), .A3(new_n1145), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n915), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1155), .A2(new_n1156), .A3(new_n1151), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1153), .A2(new_n979), .A3(new_n1157), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n823), .B1(G50), .B2(new_n853), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(G33), .A2(G41), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(new_n1160), .B(KEYINPUT118), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1161), .A2(new_n402), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1162), .B1(new_n435), .B2(new_n275), .ZN(new_n1163));
  AOI211_X1 g0963(.A(new_n718), .B(new_n350), .C1(new_n782), .C2(G107), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1164), .B1(new_n849), .B2(new_n764), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1165), .B1(new_n616), .B2(new_n785), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n775), .A2(new_n304), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(new_n1167), .B(KEYINPUT119), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n790), .A2(G68), .B1(new_n793), .B2(G77), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(G97), .A2(new_n759), .B1(new_n777), .B2(G116), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n1166), .A2(new_n1168), .A3(new_n1169), .A4(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT58), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1163), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1161), .B1(G124), .B2(new_n783), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n1119), .A2(new_n833), .B1(new_n760), .B2(new_n839), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(new_n782), .A2(G128), .B1(new_n785), .B2(G137), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1176), .B1(new_n769), .B2(new_n1118), .ZN(new_n1177));
  AOI211_X1 g0977(.A(new_n1175), .B(new_n1177), .C1(G150), .C2(new_n790), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT59), .ZN(new_n1179));
  OAI221_X1 g0979(.A(new_n1174), .B1(new_n765), .B2(new_n775), .C1(new_n1178), .C2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1178), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n1181), .A2(KEYINPUT59), .ZN(new_n1182));
  OAI221_X1 g0982(.A(new_n1173), .B1(new_n1172), .B2(new_n1171), .C1(new_n1180), .C2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1159), .B1(new_n1183), .B2(new_n755), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1184), .B1(new_n1149), .B2(new_n801), .ZN(new_n1185));
  AND2_X1   g0985(.A1(new_n1158), .A2(new_n1185), .ZN(new_n1186));
  AND2_X1   g0986(.A1(new_n1153), .A2(new_n1157), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1088), .A2(new_n1089), .A3(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1189), .A2(new_n1105), .ZN(new_n1190));
  AOI21_X1  g0990(.A(KEYINPUT57), .B1(new_n1187), .B2(new_n1190), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1153), .A2(new_n1190), .A3(KEYINPUT57), .A4(new_n1157), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1192), .A2(new_n720), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1186), .B1(new_n1191), .B2(new_n1193), .ZN(G375));
  NAND3_X1  g0994(.A1(new_n1096), .A2(new_n1091), .A3(new_n1097), .ZN(new_n1195));
  AND2_X1   g0995(.A1(new_n1108), .A2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n961), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  XNOR2_X1  g0998(.A(new_n1198), .B(KEYINPUT121), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n910), .A2(new_n801), .ZN(new_n1200));
  XNOR2_X1  g1000(.A(new_n1200), .B(KEYINPUT122), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n823), .B1(G68), .B2(new_n853), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n772), .A2(new_n834), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n350), .B1(new_n771), .B2(new_n835), .ZN(new_n1204));
  AOI211_X1 g1004(.A(new_n1203), .B(new_n1204), .C1(G128), .C2(new_n783), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1118), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(new_n759), .A2(new_n1206), .B1(new_n793), .B2(G159), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(G50), .A2(new_n790), .B1(new_n777), .B2(G132), .ZN(new_n1208));
  NAND4_X1  g1008(.A1(new_n1205), .A2(new_n1168), .A3(new_n1207), .A4(new_n1208), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n759), .A2(G116), .B1(new_n785), .B2(G107), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1210), .B1(new_n847), .B2(new_n833), .ZN(new_n1211));
  XNOR2_X1  g1011(.A(new_n1211), .B(KEYINPUT123), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n275), .B1(new_n764), .B2(new_n989), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(G283), .B2(new_n782), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1008), .B1(G97), .B2(new_n793), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1047), .A2(new_n1214), .A3(new_n1215), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1209), .B1(new_n1212), .B2(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1202), .B1(new_n1217), .B2(new_n755), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n1188), .A2(new_n979), .B1(new_n1201), .B2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1199), .A2(new_n1219), .ZN(G381));
  OR4_X1    g1020(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT124), .ZN(new_n1222));
  AND3_X1   g1022(.A1(new_n1112), .A2(new_n1222), .A3(new_n1131), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1222), .B1(new_n1112), .B2(new_n1131), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  NOR4_X1   g1025(.A1(new_n1221), .A2(G387), .A3(G381), .A4(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(G375), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1226), .A2(new_n1227), .ZN(G407));
  NAND2_X1  g1028(.A1(new_n702), .A2(G213), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1225), .A2(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(KEYINPUT125), .B1(new_n1227), .B2(new_n1230), .ZN(new_n1231));
  AND3_X1   g1031(.A1(new_n1227), .A2(KEYINPUT125), .A3(new_n1230), .ZN(new_n1232));
  OAI211_X1 g1032(.A(G407), .B(G213), .C1(new_n1231), .C2(new_n1232), .ZN(G409));
  NAND4_X1  g1033(.A1(new_n1153), .A2(new_n1190), .A3(new_n1197), .A4(new_n1157), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1234), .A2(new_n1158), .A3(new_n1185), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1235), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(KEYINPUT126), .ZN(new_n1237));
  OAI211_X1 g1037(.A(G378), .B(new_n1186), .C1(new_n1191), .C2(new_n1193), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT126), .ZN(new_n1239));
  OAI211_X1 g1039(.A(new_n1235), .B(new_n1239), .C1(new_n1223), .C2(new_n1224), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1237), .A2(new_n1238), .A3(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT60), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n1196), .A2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1195), .A2(new_n1242), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1244), .A2(new_n720), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1219), .B1(new_n1243), .B2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(G384), .ZN(new_n1247));
  OR2_X1    g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1241), .A2(new_n1229), .A3(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(KEYINPUT62), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1241), .A2(new_n1229), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n702), .A2(G213), .A3(G2897), .ZN(new_n1255));
  XNOR2_X1  g1055(.A(new_n1250), .B(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1254), .A2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT61), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT62), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1241), .A2(new_n1259), .A3(new_n1229), .A4(new_n1251), .ZN(new_n1260));
  NAND4_X1  g1060(.A1(new_n1253), .A2(new_n1257), .A3(new_n1258), .A4(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(G390), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(G387), .A2(new_n1262), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n980), .A2(new_n1014), .A3(G390), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  XNOR2_X1  g1065(.A(G393), .B(new_n821), .ZN(new_n1266));
  AOI21_X1  g1066(.A(G390), .B1(new_n980), .B2(new_n1014), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1266), .B1(new_n1267), .B2(KEYINPUT127), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1265), .A2(new_n1268), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1263), .A2(KEYINPUT127), .A3(new_n1264), .A4(new_n1266), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1261), .A2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1271), .ZN(new_n1273));
  AOI21_X1  g1073(.A(KEYINPUT61), .B1(new_n1254), .B2(new_n1256), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT63), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1252), .A2(new_n1275), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1241), .A2(KEYINPUT63), .A3(new_n1229), .A4(new_n1251), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1273), .A2(new_n1274), .A3(new_n1276), .A4(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1272), .A2(new_n1278), .ZN(G405));
  NOR2_X1   g1079(.A1(new_n1227), .A2(new_n1225), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1238), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1251), .B1(new_n1280), .B2(new_n1281), .ZN(new_n1282));
  OAI211_X1 g1082(.A(new_n1250), .B(new_n1238), .C1(new_n1227), .C2(new_n1225), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  XNOR2_X1  g1084(.A(new_n1284), .B(new_n1271), .ZN(G402));
endmodule


