//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 1 1 0 0 0 0 1 0 1 0 0 1 0 1 0 0 1 1 1 0 1 1 1 0 0 1 0 0 1 1 1 1 0 1 0 0 1 0 1 1 0 0 0 1 0 1 1 0 1 1 0 1 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:34:58 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n241, new_n242, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n257, new_n258, new_n259, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1251, new_n1252, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338, new_n1339;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XOR2_X1   g0003(.A(new_n203), .B(KEYINPUT64), .Z(new_n204));
  INV_X1    g0004(.A(G77), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n204), .A2(new_n205), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  XOR2_X1   g0008(.A(KEYINPUT67), .B(G77), .Z(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n210), .A2(G244), .ZN(new_n211));
  INV_X1    g0011(.A(G226), .ZN(new_n212));
  INV_X1    g0012(.A(G68), .ZN(new_n213));
  INV_X1    g0013(.A(G238), .ZN(new_n214));
  OAI22_X1  g0014(.A1(new_n202), .A2(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  AOI21_X1  g0015(.A(new_n215), .B1(G116), .B2(G270), .ZN(new_n216));
  NAND3_X1  g0016(.A1(new_n211), .A2(KEYINPUT68), .A3(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n219));
  NAND3_X1  g0019(.A1(new_n217), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  AOI21_X1  g0020(.A(KEYINPUT68), .B1(new_n211), .B2(new_n216), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n208), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT1), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n208), .A2(G13), .ZN(new_n224));
  INV_X1    g0024(.A(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(G250), .B1(G257), .B2(G264), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OR2_X1    g0027(.A1(new_n227), .A2(KEYINPUT0), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n229), .A2(KEYINPUT65), .ZN(new_n230));
  INV_X1    g0030(.A(KEYINPUT65), .ZN(new_n231));
  NAND3_X1  g0031(.A1(new_n231), .A2(G1), .A3(G13), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  INV_X1    g0033(.A(G20), .ZN(new_n234));
  NOR2_X1   g0034(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  INV_X1    g0035(.A(new_n201), .ZN(new_n236));
  NAND2_X1  g0036(.A1(new_n236), .A2(G50), .ZN(new_n237));
  INV_X1    g0037(.A(new_n237), .ZN(new_n238));
  NAND2_X1  g0038(.A1(new_n235), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g0039(.A1(new_n227), .A2(KEYINPUT0), .ZN(new_n240));
  NAND3_X1  g0040(.A1(new_n228), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT66), .ZN(new_n242));
  NOR2_X1   g0042(.A1(new_n223), .A2(new_n242), .ZN(G361));
  XNOR2_X1  g0043(.A(G238), .B(G244), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(G232), .ZN(new_n245));
  XOR2_X1   g0045(.A(KEYINPUT2), .B(G226), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G250), .B(G257), .Z(new_n248));
  XNOR2_X1  g0048(.A(G264), .B(G270), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(new_n247), .B(new_n250), .Z(G358));
  XOR2_X1   g0051(.A(G87), .B(G97), .Z(new_n252));
  XNOR2_X1  g0052(.A(G107), .B(G116), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n202), .A2(G68), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n213), .A2(G50), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  XNOR2_X1  g0057(.A(G58), .B(G77), .ZN(new_n258));
  XNOR2_X1  g0058(.A(new_n257), .B(new_n258), .ZN(new_n259));
  XNOR2_X1  g0059(.A(new_n254), .B(new_n259), .ZN(G351));
  INV_X1    g0060(.A(G33), .ZN(new_n261));
  INV_X1    g0061(.A(G41), .ZN(new_n262));
  OAI211_X1 g0062(.A(G1), .B(G13), .C1(new_n261), .C2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G1), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n264), .B1(G41), .B2(G45), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G232), .ZN(new_n267));
  INV_X1    g0067(.A(G274), .ZN(new_n268));
  OAI22_X1  g0068(.A1(new_n266), .A2(new_n267), .B1(new_n268), .B2(new_n265), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n261), .A2(KEYINPUT3), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT3), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G33), .ZN(new_n272));
  NAND4_X1  g0072(.A1(new_n270), .A2(new_n272), .A3(G226), .A4(G1698), .ZN(new_n273));
  INV_X1    g0073(.A(G1698), .ZN(new_n274));
  NAND4_X1  g0074(.A1(new_n270), .A2(new_n272), .A3(G223), .A4(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G87), .ZN(new_n276));
  OAI211_X1 g0076(.A(new_n273), .B(new_n275), .C1(new_n261), .C2(new_n276), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n261), .A2(new_n262), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n233), .A2(new_n278), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n269), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G169), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n282), .B1(G179), .B2(new_n280), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n208), .A2(new_n261), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n285), .B1(new_n230), .B2(new_n232), .ZN(new_n286));
  AND2_X1   g0086(.A1(G58), .A2(G68), .ZN(new_n287));
  OAI21_X1  g0087(.A(G20), .B1(new_n287), .B2(new_n201), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(KEYINPUT76), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT76), .ZN(new_n290));
  OAI211_X1 g0090(.A(new_n290), .B(G20), .C1(new_n287), .C2(new_n201), .ZN(new_n291));
  NOR2_X1   g0091(.A1(G20), .A2(G33), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(G159), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n289), .A2(new_n291), .A3(new_n293), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n271), .A2(G33), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n261), .A2(KEYINPUT3), .ZN(new_n296));
  OAI211_X1 g0096(.A(KEYINPUT7), .B(new_n234), .C1(new_n295), .C2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT75), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT7), .ZN(new_n300));
  XNOR2_X1  g0100(.A(KEYINPUT3), .B(G33), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n300), .B1(new_n301), .B2(G20), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n270), .A2(new_n272), .ZN(new_n303));
  NAND4_X1  g0103(.A1(new_n303), .A2(KEYINPUT75), .A3(KEYINPUT7), .A4(new_n234), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n299), .A2(new_n302), .A3(new_n304), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n294), .B1(new_n305), .B2(G68), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n286), .B1(new_n306), .B2(KEYINPUT16), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n302), .A2(KEYINPUT77), .A3(new_n297), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT77), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n303), .A2(new_n309), .A3(KEYINPUT7), .A4(new_n234), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n308), .A2(G68), .A3(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n294), .ZN(new_n312));
  AOI21_X1  g0112(.A(KEYINPUT16), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n307), .A2(new_n314), .ZN(new_n315));
  XOR2_X1   g0115(.A(KEYINPUT8), .B(G58), .Z(new_n316));
  NAND3_X1  g0116(.A1(new_n264), .A2(G13), .A3(G20), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n285), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n233), .A2(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n321), .B1(new_n264), .B2(G20), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n319), .B1(new_n323), .B2(new_n316), .ZN(new_n324));
  INV_X1    g0124(.A(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(KEYINPUT78), .B1(new_n315), .B2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT78), .ZN(new_n327));
  AOI211_X1 g0127(.A(new_n327), .B(new_n324), .C1(new_n307), .C2(new_n314), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n284), .B1(new_n326), .B2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT79), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n277), .A2(new_n279), .ZN(new_n331));
  INV_X1    g0131(.A(G190), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n265), .A2(new_n268), .ZN(new_n333));
  AND2_X1   g0133(.A1(new_n263), .A2(new_n265), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n333), .B1(new_n334), .B2(G232), .ZN(new_n335));
  AND3_X1   g0135(.A1(new_n331), .A2(new_n332), .A3(new_n335), .ZN(new_n336));
  AOI21_X1  g0136(.A(G200), .B1(new_n331), .B2(new_n335), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n330), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n331), .A2(new_n332), .A3(new_n335), .ZN(new_n339));
  OAI211_X1 g0139(.A(new_n339), .B(KEYINPUT79), .C1(new_n280), .C2(G200), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n341), .A2(new_n315), .A3(new_n325), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(KEYINPUT17), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT17), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n341), .A2(new_n315), .A3(new_n344), .A4(new_n325), .ZN(new_n345));
  AOI22_X1  g0145(.A1(new_n329), .A2(KEYINPUT18), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT16), .ZN(new_n347));
  AOI211_X1 g0147(.A(new_n347), .B(new_n294), .C1(new_n305), .C2(G68), .ZN(new_n348));
  NOR3_X1   g0148(.A1(new_n348), .A2(new_n313), .A3(new_n286), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n327), .B1(new_n349), .B2(new_n324), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n315), .A2(KEYINPUT78), .A3(new_n325), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n283), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT18), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n346), .A2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT80), .ZN(new_n356));
  XNOR2_X1  g0156(.A(new_n355), .B(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT81), .ZN(new_n358));
  NAND2_X1  g0158(.A1(G33), .A2(G97), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n301), .A2(G1698), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n301), .A2(new_n274), .ZN(new_n361));
  OAI221_X1 g0161(.A(new_n359), .B1(new_n360), .B2(new_n267), .C1(new_n212), .C2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(new_n279), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT13), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n333), .B1(new_n334), .B2(G238), .ZN(new_n365));
  AND3_X1   g0165(.A1(new_n363), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n364), .B1(new_n363), .B2(new_n365), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  OAI21_X1  g0168(.A(KEYINPUT14), .B1(new_n368), .B2(new_n281), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT14), .ZN(new_n370));
  OAI211_X1 g0170(.A(new_n370), .B(G169), .C1(new_n366), .C2(new_n367), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n368), .A2(G179), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n369), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n234), .A2(G33), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT71), .ZN(new_n375));
  XNOR2_X1  g0175(.A(new_n374), .B(new_n375), .ZN(new_n376));
  OR2_X1    g0176(.A1(new_n376), .A2(new_n205), .ZN(new_n377));
  AOI22_X1  g0177(.A1(new_n292), .A2(G50), .B1(G20), .B2(new_n213), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n286), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  XOR2_X1   g0179(.A(KEYINPUT74), .B(KEYINPUT11), .Z(new_n380));
  OR2_X1    g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n379), .A2(new_n380), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n322), .A2(G68), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n318), .A2(new_n213), .ZN(new_n384));
  XNOR2_X1  g0184(.A(new_n384), .B(KEYINPUT12), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n381), .A2(new_n382), .A3(new_n383), .A4(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n373), .A2(new_n386), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n204), .A2(new_n234), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n292), .A2(G150), .ZN(new_n389));
  INV_X1    g0189(.A(new_n316), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n389), .B1(new_n376), .B2(new_n390), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n321), .B1(new_n388), .B2(new_n391), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n317), .A2(G50), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n393), .B1(new_n322), .B2(G50), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  XNOR2_X1  g0196(.A(KEYINPUT69), .B(G226), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n333), .B1(new_n334), .B2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT70), .ZN(new_n399));
  OR2_X1    g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n301), .A2(G222), .A3(new_n274), .ZN(new_n401));
  INV_X1    g0201(.A(G223), .ZN(new_n402));
  OAI221_X1 g0202(.A(new_n401), .B1(new_n209), .B2(new_n301), .C1(new_n360), .C2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(new_n279), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n398), .A2(new_n399), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n400), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n406), .A2(G179), .ZN(new_n407));
  AOI211_X1 g0207(.A(new_n396), .B(new_n407), .C1(new_n281), .C2(new_n406), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n406), .A2(new_n332), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n409), .B1(KEYINPUT9), .B2(new_n396), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT9), .ZN(new_n411));
  AOI22_X1  g0211(.A1(new_n395), .A2(new_n411), .B1(new_n406), .B2(G200), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(KEYINPUT10), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT10), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n410), .A2(new_n415), .A3(new_n412), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n408), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n386), .B1(new_n368), .B2(G190), .ZN(new_n418));
  INV_X1    g0218(.A(G200), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n418), .B1(new_n419), .B2(new_n368), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n303), .A2(G107), .ZN(new_n421));
  OAI221_X1 g0221(.A(new_n421), .B1(new_n360), .B2(new_n214), .C1(new_n267), .C2(new_n361), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(new_n279), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n333), .B1(new_n334), .B2(G244), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n423), .A2(G190), .A3(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT72), .ZN(new_n426));
  XNOR2_X1  g0226(.A(new_n425), .B(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT73), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n316), .A2(new_n292), .ZN(new_n429));
  XOR2_X1   g0229(.A(KEYINPUT15), .B(G87), .Z(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  OAI221_X1 g0231(.A(new_n429), .B1(new_n234), .B2(new_n209), .C1(new_n431), .C2(new_n374), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(new_n321), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n322), .A2(G77), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n209), .A2(new_n318), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n428), .B1(new_n434), .B2(new_n437), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n433), .A2(KEYINPUT73), .A3(new_n435), .A4(new_n436), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n423), .A2(new_n424), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(G200), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n427), .A2(new_n438), .A3(new_n439), .A4(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n440), .A2(G179), .ZN(new_n444));
  AOI21_X1  g0244(.A(G169), .B1(new_n423), .B2(new_n424), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n438), .A2(new_n439), .ZN(new_n447));
  AND2_X1   g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n443), .A2(new_n448), .ZN(new_n449));
  AND4_X1   g0249(.A1(new_n387), .A2(new_n417), .A3(new_n420), .A4(new_n449), .ZN(new_n450));
  AND3_X1   g0250(.A1(new_n357), .A2(new_n358), .A3(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n358), .B1(new_n357), .B2(new_n450), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  OAI21_X1  g0253(.A(KEYINPUT83), .B1(new_n261), .B2(G1), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT83), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n455), .A2(new_n264), .A3(G33), .ZN(new_n456));
  AND3_X1   g0256(.A1(new_n454), .A2(new_n456), .A3(new_n317), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n286), .A2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(G107), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n318), .A2(new_n459), .ZN(new_n461));
  XNOR2_X1  g0261(.A(new_n461), .B(KEYINPUT25), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n270), .A2(new_n272), .A3(new_n234), .A4(G87), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(KEYINPUT22), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT22), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n301), .A2(new_n466), .A3(new_n234), .A4(G87), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  XOR2_X1   g0268(.A(KEYINPUT87), .B(KEYINPUT24), .Z(new_n469));
  NAND2_X1  g0269(.A1(G33), .A2(G116), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n470), .A2(G20), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT23), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n472), .B1(new_n234), .B2(G107), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n459), .A2(KEYINPUT23), .A3(G20), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n471), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n468), .A2(new_n469), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(KEYINPUT88), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n468), .A2(new_n475), .ZN(new_n478));
  INV_X1    g0278(.A(new_n469), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT88), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n468), .A2(new_n481), .A3(new_n469), .A4(new_n475), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n477), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT89), .ZN(new_n484));
  AND3_X1   g0284(.A1(new_n483), .A2(new_n484), .A3(new_n321), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n484), .B1(new_n483), .B2(new_n321), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n463), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n301), .A2(G257), .A3(G1698), .ZN(new_n488));
  INV_X1    g0288(.A(G294), .ZN(new_n489));
  INV_X1    g0289(.A(G250), .ZN(new_n490));
  OAI221_X1 g0290(.A(new_n488), .B1(new_n261), .B2(new_n489), .C1(new_n361), .C2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(new_n279), .ZN(new_n492));
  NAND2_X1  g0292(.A1(KEYINPUT5), .A2(G41), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  NOR2_X1   g0294(.A1(KEYINPUT5), .A2(G41), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(G45), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n497), .A2(G1), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(G274), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n496), .A2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(new_n500), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n229), .B1(G33), .B2(G41), .ZN(new_n502));
  INV_X1    g0302(.A(new_n495), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(new_n493), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n502), .B1(new_n504), .B2(new_n498), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(G264), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n492), .A2(new_n501), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(new_n281), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n506), .A2(new_n501), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n509), .B1(new_n491), .B2(new_n279), .ZN(new_n510));
  INV_X1    g0310(.A(G179), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n508), .A2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n487), .A2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT20), .ZN(new_n516));
  AOI21_X1  g0316(.A(G20), .B1(G33), .B2(G283), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n261), .A2(G97), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(G116), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(G20), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n516), .B1(new_n286), .B2(new_n522), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n517), .A2(new_n518), .B1(G20), .B2(new_n520), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n321), .A2(KEYINPUT20), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n286), .A2(new_n457), .A3(G116), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n318), .A2(new_n520), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n500), .B1(new_n505), .B2(G270), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n270), .A2(new_n272), .A3(G257), .A4(new_n274), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n270), .A2(new_n272), .A3(G264), .A4(G1698), .ZN(new_n532));
  INV_X1    g0332(.A(G303), .ZN(new_n533));
  OAI211_X1 g0333(.A(new_n531), .B(new_n532), .C1(new_n533), .C2(new_n301), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(new_n279), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n281), .B1(new_n530), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n529), .A2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT21), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AND3_X1   g0339(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n530), .A2(new_n535), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(G200), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n530), .A2(new_n535), .A3(G190), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n540), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n529), .A2(new_n536), .A3(KEYINPUT21), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n541), .A2(new_n511), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(new_n529), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n539), .A2(new_n544), .A3(new_n545), .A4(new_n547), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n270), .A2(new_n272), .A3(G238), .A4(new_n274), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n270), .A2(new_n272), .A3(G244), .A4(G1698), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n549), .A2(new_n550), .A3(new_n470), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(new_n279), .ZN(new_n552));
  OAI21_X1  g0352(.A(G250), .B1(new_n497), .B2(G1), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n499), .B1(new_n502), .B2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(new_n281), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n286), .A2(new_n457), .A3(new_n430), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT85), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n430), .A2(new_n317), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT19), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n234), .B1(new_n359), .B2(new_n562), .ZN(new_n563));
  NOR2_X1   g0363(.A1(G97), .A2(G107), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n276), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n270), .A2(new_n272), .A3(new_n234), .A4(G68), .ZN(new_n567));
  INV_X1    g0367(.A(G97), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n562), .B1(new_n374), .B2(new_n568), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n566), .A2(new_n567), .A3(new_n569), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n561), .B1(new_n570), .B2(new_n321), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n286), .A2(new_n457), .A3(KEYINPUT85), .A4(new_n430), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n560), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n554), .B1(new_n551), .B2(new_n279), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n511), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n557), .A2(new_n573), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n556), .A2(G200), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n570), .A2(new_n321), .ZN(new_n578));
  INV_X1    g0378(.A(new_n561), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n286), .A2(new_n457), .A3(G87), .ZN(new_n580));
  AND3_X1   g0380(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n574), .A2(G190), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n577), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT86), .ZN(new_n584));
  AND3_X1   g0384(.A1(new_n576), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n584), .B1(new_n576), .B2(new_n583), .ZN(new_n586));
  NOR3_X1   g0386(.A1(new_n548), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n510), .A2(new_n332), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n588), .B1(G200), .B2(new_n510), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n589), .B(new_n463), .C1(new_n485), .C2(new_n486), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n270), .A2(new_n272), .A3(G244), .A4(new_n274), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT4), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n301), .A2(KEYINPUT4), .A3(G244), .A4(new_n274), .ZN(new_n594));
  NAND2_X1  g0394(.A1(G33), .A2(G283), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n301), .A2(G250), .A3(G1698), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n593), .A2(new_n594), .A3(new_n595), .A4(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n279), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n498), .B1(new_n494), .B2(new_n495), .ZN(new_n599));
  AND3_X1   g0399(.A1(new_n599), .A2(G257), .A3(new_n263), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n598), .A2(G190), .A3(new_n501), .A4(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(KEYINPUT84), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n318), .A2(new_n568), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n604), .B1(new_n458), .B2(new_n568), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n308), .A2(G107), .A3(new_n310), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT6), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n568), .A2(new_n459), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n607), .B1(new_n608), .B2(new_n564), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n459), .A2(KEYINPUT82), .A3(KEYINPUT6), .A4(G97), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT82), .ZN(new_n611));
  NAND2_X1  g0411(.A1(KEYINPUT6), .A2(G97), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n611), .B1(new_n612), .B2(G107), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n609), .A2(new_n610), .A3(new_n613), .ZN(new_n614));
  AOI22_X1  g0414(.A1(new_n614), .A2(G20), .B1(G77), .B2(new_n292), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n606), .A2(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n605), .B1(new_n616), .B2(new_n321), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n598), .A2(new_n501), .A3(new_n601), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(G200), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n600), .B1(new_n597), .B2(new_n279), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT84), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n620), .A2(new_n621), .A3(G190), .A4(new_n501), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n603), .A2(new_n617), .A3(new_n619), .A4(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n618), .A2(new_n281), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n620), .A2(new_n511), .A3(new_n501), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n286), .B1(new_n606), .B2(new_n615), .ZN(new_n626));
  OAI211_X1 g0426(.A(new_n624), .B(new_n625), .C1(new_n626), .C2(new_n605), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n623), .A2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n628), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n515), .A2(new_n587), .A3(new_n590), .A4(new_n629), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n453), .A2(new_n630), .ZN(G372));
  NAND2_X1  g0431(.A1(new_n420), .A2(new_n448), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(new_n387), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n343), .A2(new_n345), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n283), .B1(new_n315), .B2(new_n325), .ZN(new_n636));
  XNOR2_X1  g0436(.A(new_n636), .B(KEYINPUT18), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n414), .A2(new_n416), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n408), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  XOR2_X1   g0440(.A(new_n576), .B(KEYINPUT90), .Z(new_n641));
  AND2_X1   g0441(.A1(new_n576), .A2(new_n583), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n623), .A2(new_n627), .A3(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n463), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n473), .A2(new_n474), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n645), .B1(G20), .B2(new_n470), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n646), .B1(new_n465), .B2(new_n467), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n482), .B1(new_n469), .B2(new_n647), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n481), .B1(new_n647), .B2(new_n469), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n321), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(KEYINPUT89), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n483), .A2(new_n484), .A3(new_n321), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n644), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n643), .B1(new_n653), .B2(new_n589), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n539), .A2(new_n545), .A3(new_n547), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n656), .B1(new_n653), .B2(new_n513), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n641), .B1(new_n654), .B2(new_n657), .ZN(new_n658));
  AOI211_X1 g0458(.A(new_n500), .B(new_n600), .C1(new_n597), .C2(new_n279), .ZN(new_n659));
  OAI22_X1  g0459(.A1(G169), .A2(new_n659), .B1(new_n626), .B2(new_n605), .ZN(new_n660));
  INV_X1    g0460(.A(new_n625), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n576), .A2(new_n583), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(KEYINPUT86), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n576), .A2(new_n583), .A3(new_n584), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n662), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(KEYINPUT26), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n663), .B1(new_n627), .B2(KEYINPUT91), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT26), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n616), .A2(new_n321), .ZN(new_n670));
  INV_X1    g0470(.A(new_n605), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT91), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n672), .A2(new_n673), .A3(new_n625), .A4(new_n624), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n668), .A2(new_n669), .A3(new_n674), .ZN(new_n675));
  AND2_X1   g0475(.A1(new_n667), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n658), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n640), .B1(new_n453), .B2(new_n678), .ZN(G369));
  NOR2_X1   g0479(.A1(new_n653), .A2(new_n513), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n264), .A2(new_n234), .A3(G13), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(KEYINPUT27), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT27), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n683), .A2(new_n264), .A3(new_n234), .A4(G13), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n682), .A2(G213), .A3(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT92), .ZN(new_n686));
  XNOR2_X1  g0486(.A(new_n685), .B(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(G343), .ZN(new_n688));
  NOR3_X1   g0488(.A1(new_n687), .A2(KEYINPUT93), .A3(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT93), .ZN(new_n690));
  XNOR2_X1  g0490(.A(new_n685), .B(KEYINPUT92), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n690), .B1(new_n691), .B2(G343), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n680), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n656), .A2(new_n694), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n515), .A2(new_n590), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n653), .A2(new_n693), .ZN(new_n699));
  OAI211_X1 g0499(.A(new_n695), .B(new_n697), .C1(new_n698), .C2(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n693), .A2(new_n540), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n655), .A2(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n702), .B1(new_n548), .B2(new_n701), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(G330), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n700), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT94), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n707), .B1(new_n689), .B2(new_n692), .ZN(new_n708));
  OAI21_X1  g0508(.A(KEYINPUT93), .B1(new_n687), .B2(new_n688), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n691), .A2(new_n690), .A3(G343), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n709), .A2(KEYINPUT94), .A3(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n708), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n680), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n515), .A2(new_n696), .A3(new_n590), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n706), .A2(new_n713), .A3(new_n714), .ZN(G399));
  INV_X1    g0515(.A(KEYINPUT95), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n716), .B1(new_n225), .B2(G41), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n224), .A2(KEYINPUT95), .A3(new_n262), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n565), .A2(G116), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n719), .A2(G1), .A3(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n721), .B1(new_n237), .B2(new_n719), .ZN(new_n722));
  XNOR2_X1  g0522(.A(new_n722), .B(KEYINPUT28), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n507), .A2(new_n556), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n724), .A2(KEYINPUT30), .A3(new_n620), .A4(new_n546), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n510), .A2(G179), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n726), .A2(new_n618), .A3(new_n541), .A4(new_n556), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n546), .A2(new_n510), .A3(new_n620), .A4(new_n574), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT30), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n725), .A2(new_n727), .A3(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n712), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n731), .A2(new_n732), .A3(KEYINPUT31), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n731), .A2(new_n694), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT31), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  OAI211_X1 g0536(.A(new_n733), .B(new_n736), .C1(new_n630), .C2(new_n732), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(G330), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT29), .ZN(new_n739));
  INV_X1    g0539(.A(new_n641), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n629), .A2(new_n590), .A3(new_n642), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n655), .B1(new_n487), .B2(new_n514), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n740), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n667), .A2(new_n675), .ZN(new_n744));
  OAI211_X1 g0544(.A(new_n739), .B(new_n712), .C1(new_n743), .C2(new_n744), .ZN(new_n745));
  OAI21_X1  g0545(.A(KEYINPUT91), .B1(new_n660), .B2(new_n661), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n746), .A2(KEYINPUT26), .A3(new_n642), .A4(new_n674), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(KEYINPUT96), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT96), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n668), .A2(new_n749), .A3(KEYINPUT26), .A4(new_n674), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n666), .A2(new_n669), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n748), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n694), .B1(new_n658), .B2(new_n752), .ZN(new_n753));
  OAI211_X1 g0553(.A(new_n738), .B(new_n745), .C1(new_n739), .C2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n723), .B1(new_n755), .B2(G1), .ZN(G364));
  INV_X1    g0556(.A(new_n719), .ZN(new_n757));
  AND2_X1   g0557(.A1(new_n234), .A2(G13), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n264), .B1(new_n758), .B2(G45), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n757), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n705), .A2(new_n761), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n762), .B1(G330), .B2(new_n703), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n233), .B1(G20), .B2(new_n281), .ZN(new_n764));
  OR2_X1    g0564(.A1(new_n764), .A2(KEYINPUT99), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(KEYINPUT99), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n332), .A2(G20), .ZN(new_n769));
  NOR3_X1   g0569(.A1(new_n769), .A2(G179), .A3(G200), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(G159), .ZN(new_n772));
  NOR3_X1   g0572(.A1(new_n771), .A2(KEYINPUT32), .A3(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n769), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n419), .A2(G179), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(new_n459), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n511), .A2(new_n419), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n234), .A2(new_n332), .ZN(new_n779));
  AND2_X1   g0579(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n777), .B1(G50), .B2(new_n780), .ZN(new_n781));
  NOR3_X1   g0581(.A1(new_n769), .A2(new_n511), .A3(G200), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n781), .B1(new_n209), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n774), .A2(new_n778), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n779), .A2(new_n775), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  AOI22_X1  g0588(.A1(new_n786), .A2(G68), .B1(new_n788), .B2(G87), .ZN(new_n789));
  INV_X1    g0589(.A(G58), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n779), .A2(G179), .A3(new_n419), .ZN(new_n791));
  OAI211_X1 g0591(.A(new_n789), .B(new_n301), .C1(new_n790), .C2(new_n791), .ZN(new_n792));
  OAI21_X1  g0592(.A(KEYINPUT32), .B1(new_n771), .B2(new_n772), .ZN(new_n793));
  NOR3_X1   g0593(.A1(new_n332), .A2(G179), .A3(G200), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(new_n234), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n793), .B1(new_n568), .B2(new_n795), .ZN(new_n796));
  OR4_X1    g0596(.A1(new_n773), .A2(new_n784), .A3(new_n792), .A4(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n776), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n301), .B1(new_n798), .B2(G283), .ZN(new_n799));
  XOR2_X1   g0599(.A(KEYINPUT33), .B(G317), .Z(new_n800));
  OAI221_X1 g0600(.A(new_n799), .B1(new_n533), .B2(new_n787), .C1(new_n785), .C2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n795), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n801), .B1(G294), .B2(new_n802), .ZN(new_n803));
  AOI22_X1  g0603(.A1(new_n780), .A2(G326), .B1(new_n770), .B2(G329), .ZN(new_n804));
  INV_X1    g0604(.A(new_n791), .ZN(new_n805));
  AOI22_X1  g0605(.A1(new_n805), .A2(G322), .B1(G311), .B2(new_n782), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n803), .A2(new_n804), .A3(new_n806), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n768), .B1(new_n797), .B2(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(G13), .A2(G33), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n810), .A2(G20), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n767), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n238), .A2(new_n497), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n225), .A2(new_n301), .ZN(new_n814));
  OAI211_X1 g0614(.A(new_n813), .B(new_n814), .C1(new_n259), .C2(new_n497), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n301), .A2(G355), .A3(new_n224), .ZN(new_n816));
  OAI211_X1 g0616(.A(new_n815), .B(new_n816), .C1(G116), .C2(new_n224), .ZN(new_n817));
  INV_X1    g0617(.A(KEYINPUT98), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n812), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n819), .B1(new_n818), .B2(new_n817), .ZN(new_n820));
  XOR2_X1   g0620(.A(new_n761), .B(KEYINPUT97), .Z(new_n821));
  NOR3_X1   g0621(.A1(new_n808), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n811), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n822), .B1(new_n703), .B2(new_n823), .ZN(new_n824));
  AND2_X1   g0624(.A1(new_n763), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(G396));
  NAND2_X1  g0626(.A1(new_n448), .A2(new_n694), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n447), .A2(new_n694), .ZN(new_n828));
  INV_X1    g0628(.A(KEYINPUT100), .ZN(new_n829));
  AND3_X1   g0629(.A1(new_n446), .A2(new_n829), .A3(new_n447), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n829), .B1(new_n446), .B2(new_n447), .ZN(new_n831));
  OAI211_X1 g0631(.A(new_n442), .B(new_n828), .C1(new_n830), .C2(new_n831), .ZN(new_n832));
  OAI211_X1 g0632(.A(new_n827), .B(new_n832), .C1(new_n678), .C2(new_n732), .ZN(new_n833));
  AND2_X1   g0633(.A1(new_n737), .A2(G330), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n832), .A2(new_n827), .ZN(new_n835));
  OAI211_X1 g0635(.A(new_n835), .B(new_n712), .C1(new_n743), .C2(new_n744), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n833), .A2(new_n834), .A3(new_n836), .ZN(new_n837));
  AND2_X1   g0637(.A1(new_n837), .A2(KEYINPUT101), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n834), .B1(new_n833), .B2(new_n836), .ZN(new_n839));
  NOR3_X1   g0639(.A1(new_n838), .A2(new_n761), .A3(new_n839), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n840), .B1(KEYINPUT101), .B2(new_n837), .ZN(new_n841));
  INV_X1    g0641(.A(new_n821), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n768), .A2(new_n810), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n842), .B1(new_n843), .B2(G77), .ZN(new_n844));
  INV_X1    g0644(.A(new_n780), .ZN(new_n845));
  INV_X1    g0645(.A(G311), .ZN(new_n846));
  OAI22_X1  g0646(.A1(new_n845), .A2(new_n533), .B1(new_n771), .B2(new_n846), .ZN(new_n847));
  AOI211_X1 g0647(.A(new_n301), .B(new_n847), .C1(G294), .C2(new_n805), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n802), .A2(G97), .ZN(new_n849));
  AOI22_X1  g0649(.A1(new_n798), .A2(G87), .B1(new_n788), .B2(G107), .ZN(new_n850));
  AOI22_X1  g0650(.A1(new_n786), .A2(G283), .B1(G116), .B2(new_n782), .ZN(new_n851));
  NAND4_X1  g0651(.A1(new_n848), .A2(new_n849), .A3(new_n850), .A4(new_n851), .ZN(new_n852));
  AOI22_X1  g0652(.A1(new_n780), .A2(G137), .B1(new_n782), .B2(G159), .ZN(new_n853));
  INV_X1    g0653(.A(G143), .ZN(new_n854));
  INV_X1    g0654(.A(G150), .ZN(new_n855));
  OAI221_X1 g0655(.A(new_n853), .B1(new_n854), .B2(new_n791), .C1(new_n855), .C2(new_n785), .ZN(new_n856));
  XOR2_X1   g0656(.A(new_n856), .B(KEYINPUT34), .Z(new_n857));
  AOI22_X1  g0657(.A1(new_n798), .A2(G68), .B1(G132), .B2(new_n770), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n303), .B1(new_n788), .B2(G50), .ZN(new_n859));
  OAI211_X1 g0659(.A(new_n858), .B(new_n859), .C1(new_n790), .C2(new_n795), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n852), .B1(new_n857), .B2(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n844), .B1(new_n861), .B2(new_n767), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n862), .B1(new_n835), .B2(new_n810), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n841), .A2(new_n863), .ZN(G384));
  OAI211_X1 g0664(.A(G116), .B(new_n235), .C1(new_n614), .C2(KEYINPUT35), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n865), .B1(KEYINPUT35), .B2(new_n614), .ZN(new_n866));
  XNOR2_X1  g0666(.A(new_n866), .B(KEYINPUT36), .ZN(new_n867));
  OR3_X1    g0667(.A1(new_n209), .A2(new_n237), .A3(new_n287), .ZN(new_n868));
  AOI211_X1 g0668(.A(new_n264), .B(G13), .C1(new_n868), .C2(new_n255), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n731), .A2(KEYINPUT31), .A3(new_n694), .ZN(new_n871));
  OAI211_X1 g0671(.A(new_n736), .B(new_n871), .C1(new_n630), .C2(new_n732), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT104), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NOR4_X1   g0674(.A1(new_n628), .A2(new_n548), .A3(new_n585), .A4(new_n586), .ZN(new_n875));
  NAND4_X1  g0675(.A1(new_n875), .A2(new_n515), .A3(new_n590), .A4(new_n712), .ZN(new_n876));
  NAND4_X1  g0676(.A1(new_n876), .A2(KEYINPUT104), .A3(new_n736), .A4(new_n871), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n386), .A2(new_n694), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n387), .A2(new_n420), .A3(new_n879), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n373), .A2(new_n386), .A3(new_n694), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND4_X1  g0682(.A1(new_n878), .A2(KEYINPUT40), .A3(new_n835), .A4(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n687), .B1(new_n350), .B2(new_n351), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n349), .A2(new_n324), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n342), .B1(new_n885), .B2(new_n283), .ZN(new_n886));
  OAI21_X1  g0686(.A(KEYINPUT37), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT102), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n691), .B1(new_n326), .B2(new_n328), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT37), .ZN(new_n891));
  NAND4_X1  g0691(.A1(new_n329), .A2(new_n890), .A3(new_n891), .A4(new_n342), .ZN(new_n892));
  OAI211_X1 g0692(.A(KEYINPUT102), .B(KEYINPUT37), .C1(new_n884), .C2(new_n886), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n889), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n890), .B1(new_n637), .B2(new_n634), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(KEYINPUT38), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n307), .B1(KEYINPUT16), .B2(new_n306), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(new_n325), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(new_n691), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n900), .B1(new_n346), .B2(new_n354), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n342), .A2(new_n891), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n352), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n899), .A2(new_n284), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n900), .A2(new_n904), .A3(new_n342), .ZN(new_n905));
  AOI22_X1  g0705(.A1(new_n903), .A2(new_n890), .B1(new_n905), .B2(KEYINPUT37), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT38), .ZN(new_n907));
  NOR3_X1   g0707(.A1(new_n901), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(KEYINPUT105), .B1(new_n897), .B2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT105), .ZN(new_n910));
  INV_X1    g0710(.A(new_n900), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n634), .B1(new_n352), .B2(new_n353), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n329), .A2(KEYINPUT18), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n911), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n905), .A2(KEYINPUT37), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n892), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n914), .A2(KEYINPUT38), .A3(new_n916), .ZN(new_n917));
  AOI22_X1  g0717(.A1(new_n887), .A2(new_n888), .B1(new_n903), .B2(new_n890), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n895), .B1(new_n918), .B2(new_n893), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n910), .B(new_n917), .C1(new_n919), .C2(KEYINPUT38), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n883), .B1(new_n909), .B2(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(KEYINPUT38), .B1(new_n914), .B2(new_n916), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n917), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n882), .A2(new_n835), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n925), .B1(new_n874), .B2(new_n877), .ZN(new_n926));
  AOI21_X1  g0726(.A(KEYINPUT40), .B1(new_n924), .B2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(new_n878), .ZN(new_n928));
  OR4_X1    g0728(.A1(new_n453), .A2(new_n921), .A3(new_n927), .A4(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(G330), .ZN(new_n930));
  NOR3_X1   g0730(.A1(new_n921), .A2(new_n927), .A3(new_n930), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n928), .A2(new_n930), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(new_n451), .B2(new_n452), .ZN(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n929), .B1(new_n931), .B2(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT39), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n936), .B(new_n917), .C1(new_n919), .C2(KEYINPUT38), .ZN(new_n937));
  OAI21_X1  g0737(.A(KEYINPUT39), .B1(new_n908), .B2(new_n922), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n387), .A2(new_n694), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n830), .A2(new_n831), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(new_n693), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n836), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(new_n882), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(new_n637), .ZN(new_n947));
  AOI22_X1  g0747(.A1(new_n946), .A2(new_n924), .B1(new_n947), .B2(new_n687), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT103), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n941), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(new_n940), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n951), .B1(new_n937), .B2(new_n938), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n947), .A2(new_n687), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n908), .A2(new_n922), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n953), .B1(new_n954), .B2(new_n945), .ZN(new_n955));
  OAI21_X1  g0755(.A(KEYINPUT103), .B1(new_n952), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n950), .A2(new_n956), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n935), .B(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n658), .A2(new_n752), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n739), .B1(new_n959), .B2(new_n693), .ZN(new_n960));
  AOI211_X1 g0760(.A(KEYINPUT29), .B(new_n732), .C1(new_n658), .C2(new_n676), .ZN(new_n961));
  OAI22_X1  g0761(.A1(new_n451), .A2(new_n452), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  AND2_X1   g0762(.A1(new_n962), .A2(new_n640), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n958), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n964), .B1(new_n264), .B2(new_n758), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n958), .A2(new_n963), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n870), .B1(new_n965), .B2(new_n966), .ZN(G367));
  OR2_X1    g0767(.A1(new_n693), .A2(new_n581), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n968), .A2(new_n642), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n969), .B1(new_n740), .B2(new_n968), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n970), .A2(KEYINPUT43), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n732), .A2(new_n662), .ZN(new_n972));
  OAI211_X1 g0772(.A(new_n627), .B(new_n623), .C1(new_n712), .C2(new_n617), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n974), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n975), .A2(new_n714), .ZN(new_n976));
  XOR2_X1   g0776(.A(new_n976), .B(KEYINPUT42), .Z(new_n977));
  INV_X1    g0777(.A(KEYINPUT106), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n974), .B(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(new_n680), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n732), .B1(new_n980), .B2(new_n627), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n971), .B1(new_n977), .B2(new_n981), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n970), .A2(KEYINPUT43), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(new_n983), .ZN(new_n985));
  OAI211_X1 g0785(.A(new_n985), .B(new_n971), .C1(new_n977), .C2(new_n981), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n984), .A2(new_n986), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n979), .A2(new_n705), .A3(new_n700), .ZN(new_n988));
  INV_X1    g0788(.A(new_n988), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n987), .B(new_n989), .ZN(new_n990));
  XOR2_X1   g0790(.A(new_n719), .B(KEYINPUT41), .Z(new_n991));
  INV_X1    g0791(.A(new_n991), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n960), .A2(new_n961), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT107), .ZN(new_n994));
  OAI211_X1 g0794(.A(new_n515), .B(new_n590), .C1(new_n653), .C2(new_n693), .ZN(new_n995));
  NAND4_X1  g0795(.A1(new_n995), .A2(new_n704), .A3(new_n697), .A4(new_n695), .ZN(new_n996));
  AND3_X1   g0796(.A1(new_n706), .A2(new_n714), .A3(new_n996), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n993), .A2(new_n994), .A3(new_n738), .A4(new_n997), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n706), .A2(new_n714), .A3(new_n996), .ZN(new_n999));
  OAI21_X1  g0799(.A(KEYINPUT107), .B1(new_n754), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1001), .A2(KEYINPUT108), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT108), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n998), .A2(new_n1000), .A3(new_n1003), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n714), .A2(new_n713), .A3(new_n974), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT45), .ZN(new_n1006));
  AND2_X1   g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n714), .A2(new_n713), .ZN(new_n1009));
  AOI21_X1  g0809(.A(KEYINPUT44), .B1(new_n1009), .B2(new_n975), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT44), .ZN(new_n1011));
  AOI211_X1 g0811(.A(new_n1011), .B(new_n974), .C1(new_n714), .C2(new_n713), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n1007), .A2(new_n1008), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1013), .A2(new_n705), .A3(new_n700), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n706), .B1(new_n1010), .B2(new_n1012), .C1(new_n1008), .C2(new_n1007), .ZN(new_n1015));
  AND2_X1   g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1002), .A2(new_n1004), .A3(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n992), .B1(new_n1017), .B2(new_n755), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n990), .B1(new_n1018), .B2(new_n760), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n814), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n812), .B1(new_n224), .B2(new_n431), .C1(new_n250), .C2(new_n1020), .ZN(new_n1021));
  AND2_X1   g0821(.A1(new_n1021), .A2(KEYINPUT109), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n1021), .A2(KEYINPUT109), .ZN(new_n1023));
  NOR3_X1   g0823(.A1(new_n1022), .A2(new_n1023), .A3(new_n821), .ZN(new_n1024));
  INV_X1    g0824(.A(G137), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n771), .A2(new_n1025), .B1(new_n790), .B2(new_n787), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT111), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n783), .A2(new_n202), .B1(new_n772), .B2(new_n785), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT110), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n802), .A2(G68), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n845), .A2(new_n854), .B1(new_n776), .B2(new_n209), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n301), .B1(new_n791), .B2(new_n855), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND4_X1  g0833(.A1(new_n1027), .A2(new_n1029), .A3(new_n1030), .A4(new_n1033), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT112), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n788), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1036));
  INV_X1    g0836(.A(KEYINPUT46), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1037), .B1(new_n787), .B2(new_n520), .ZN(new_n1038));
  OAI211_X1 g0838(.A(new_n1036), .B(new_n1038), .C1(new_n459), .C2(new_n795), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n798), .A2(G97), .B1(G317), .B2(new_n770), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1040), .B1(new_n846), .B2(new_n845), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n303), .B1(new_n791), .B2(new_n533), .ZN(new_n1042));
  INV_X1    g0842(.A(G283), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n783), .A2(new_n1043), .B1(new_n489), .B2(new_n785), .ZN(new_n1044));
  OR3_X1    g0844(.A1(new_n1041), .A2(new_n1042), .A3(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1035), .B1(new_n1039), .B2(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n1046), .ZN(new_n1047));
  AND2_X1   g0847(.A1(new_n1047), .A2(KEYINPUT47), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n767), .B1(new_n1047), .B2(KEYINPUT47), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n1024), .B1(new_n823), .B2(new_n970), .C1(new_n1048), .C2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1019), .A2(new_n1050), .ZN(G387));
  AOI22_X1  g0851(.A1(new_n780), .A2(G322), .B1(new_n782), .B2(G303), .ZN(new_n1052));
  INV_X1    g0852(.A(G317), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n1052), .B1(new_n846), .B2(new_n785), .C1(new_n1053), .C2(new_n791), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT48), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n1055), .B1(new_n1043), .B2(new_n795), .C1(new_n489), .C2(new_n787), .ZN(new_n1056));
  INV_X1    g0856(.A(KEYINPUT49), .ZN(new_n1057));
  OR2_X1    g0857(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n776), .A2(new_n520), .ZN(new_n1060));
  AOI211_X1 g0860(.A(new_n301), .B(new_n1060), .C1(G326), .C2(new_n770), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1058), .A2(new_n1059), .A3(new_n1061), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n845), .A2(new_n772), .B1(new_n771), .B2(new_n855), .ZN(new_n1063));
  AOI211_X1 g0863(.A(new_n303), .B(new_n1063), .C1(G97), .C2(new_n798), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n316), .A2(new_n786), .B1(new_n805), .B2(G50), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n209), .A2(new_n787), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(G68), .B2(new_n782), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n802), .A2(new_n430), .ZN(new_n1068));
  NAND4_X1  g0868(.A1(new_n1064), .A2(new_n1065), .A3(new_n1067), .A4(new_n1068), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n768), .B1(new_n1062), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n812), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n247), .A2(G45), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(KEYINPUT113), .B(KEYINPUT50), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1073), .B1(new_n316), .B2(new_n202), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n316), .A2(new_n202), .A3(new_n1073), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n1075), .B(new_n497), .C1(new_n213), .C2(new_n205), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n1072), .B(new_n814), .C1(new_n1074), .C2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1077), .A2(new_n720), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n1078), .B(new_n224), .C1(new_n301), .C2(new_n1072), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n225), .A2(new_n459), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1071), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  NOR3_X1   g0881(.A1(new_n1070), .A2(new_n821), .A3(new_n1081), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n995), .A2(new_n695), .A3(new_n811), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  XOR2_X1   g0884(.A(new_n1084), .B(KEYINPUT114), .Z(new_n1085));
  AOI21_X1  g0885(.A(new_n1085), .B1(new_n760), .B2(new_n997), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n1001), .B(new_n757), .C1(new_n755), .C2(new_n997), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1086), .A2(new_n1087), .ZN(G393));
  NAND2_X1  g0888(.A1(new_n1016), .A2(new_n760), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n254), .A2(new_n1020), .B1(new_n568), .B2(new_n224), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n842), .B1(new_n1071), .B2(new_n1090), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n845), .A2(new_n1053), .B1(new_n791), .B2(new_n846), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(new_n1092), .B(KEYINPUT52), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(G294), .A2(new_n782), .B1(new_n770), .B2(G322), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n786), .A2(G303), .B1(new_n788), .B2(G283), .ZN(new_n1095));
  AOI211_X1 g0895(.A(new_n301), .B(new_n777), .C1(G116), .C2(new_n802), .ZN(new_n1096));
  NAND4_X1  g0896(.A1(new_n1093), .A2(new_n1094), .A3(new_n1095), .A4(new_n1096), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n845), .A2(new_n855), .B1(new_n791), .B2(new_n772), .ZN(new_n1098));
  XNOR2_X1  g0898(.A(new_n1098), .B(KEYINPUT51), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n802), .A2(G77), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(new_n786), .A2(G50), .B1(new_n782), .B2(new_n316), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1099), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n788), .A2(G68), .B1(new_n770), .B2(G143), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n1103), .B(new_n301), .C1(new_n276), .C2(new_n776), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(new_n1104), .B(KEYINPUT115), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1097), .B1(new_n1102), .B2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1091), .B1(new_n1106), .B2(new_n767), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1107), .B1(new_n979), .B2(new_n823), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1089), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n719), .B1(new_n1001), .B2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1109), .B1(new_n1017), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1112), .ZN(G390));
  OAI211_X1 g0913(.A(new_n753), .B(new_n442), .C1(new_n831), .C2(new_n830), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(new_n943), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n940), .B1(new_n1115), .B2(new_n882), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n909), .A2(new_n920), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n938), .B(new_n937), .C1(new_n946), .C2(new_n940), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NAND4_X1  g0920(.A1(new_n878), .A2(G330), .A3(new_n835), .A4(new_n882), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n925), .A2(new_n738), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1118), .A2(new_n1119), .A3(new_n1125), .ZN(new_n1126));
  AND2_X1   g0926(.A1(new_n1123), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1127), .A2(new_n760), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n771), .A2(new_n489), .B1(new_n213), .B2(new_n776), .ZN(new_n1129));
  AOI211_X1 g0929(.A(new_n301), .B(new_n1129), .C1(G87), .C2(new_n788), .ZN(new_n1130));
  AOI22_X1  g0930(.A1(new_n805), .A2(G116), .B1(new_n780), .B2(G283), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n786), .A2(G107), .B1(G97), .B2(new_n782), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n1130), .A2(new_n1100), .A3(new_n1131), .A4(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n770), .A2(G125), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1134), .B1(new_n202), .B2(new_n776), .ZN(new_n1135));
  AOI211_X1 g0935(.A(new_n303), .B(new_n1135), .C1(G128), .C2(new_n780), .ZN(new_n1136));
  OAI21_X1  g0936(.A(KEYINPUT53), .B1(new_n787), .B2(new_n855), .ZN(new_n1137));
  NOR3_X1   g0937(.A1(new_n787), .A2(KEYINPUT53), .A3(new_n855), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(G159), .B2(new_n802), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(KEYINPUT54), .B(G143), .ZN(new_n1140));
  INV_X1    g0940(.A(G132), .ZN(new_n1141));
  OAI22_X1  g0941(.A1(new_n783), .A2(new_n1140), .B1(new_n1141), .B2(new_n791), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1142), .B1(G137), .B2(new_n786), .ZN(new_n1143));
  NAND4_X1  g0943(.A1(new_n1136), .A2(new_n1137), .A3(new_n1139), .A4(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n768), .B1(new_n1133), .B2(new_n1144), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n843), .A2(new_n316), .ZN(new_n1146));
  NOR3_X1   g0946(.A1(new_n1145), .A2(new_n821), .A3(new_n1146), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1147), .B1(new_n939), .B2(new_n810), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1128), .A2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n878), .A2(G330), .A3(new_n835), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n882), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1115), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1152), .A2(new_n1153), .A3(new_n1125), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n835), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1151), .B1(new_n738), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1121), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1157), .A2(new_n944), .ZN(new_n1158));
  AND2_X1   g0958(.A1(new_n1154), .A2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n962), .A2(new_n933), .A3(new_n640), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  OR2_X1    g0961(.A1(new_n1127), .A2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n719), .B1(new_n1127), .B2(new_n1161), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1149), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(G378));
  OAI211_X1 g0965(.A(new_n950), .B(new_n956), .C1(new_n931), .C2(KEYINPUT119), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n883), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1117), .A2(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n927), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1168), .A2(new_n1169), .A3(G330), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT119), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n949), .B1(new_n941), .B2(new_n948), .ZN(new_n1172));
  NOR3_X1   g0972(.A1(new_n952), .A2(new_n955), .A3(KEYINPUT103), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n1170), .B(new_n1171), .C1(new_n1172), .C2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1166), .A2(new_n1174), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(new_n417), .B(KEYINPUT118), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n396), .A2(new_n687), .ZN(new_n1177));
  OR2_X1    g0977(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1180));
  AND3_X1   g0980(.A1(new_n1178), .A2(new_n1179), .A3(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1179), .B1(new_n1178), .B2(new_n1180), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(new_n931), .B2(KEYINPUT119), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1175), .A2(new_n1185), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1166), .A2(new_n1174), .A3(new_n1184), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n809), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n761), .B1(new_n843), .B2(G50), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(new_n1190), .B(KEYINPUT117), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n202), .B1(G33), .B2(G41), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1192), .B1(new_n303), .B2(new_n262), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n790), .A2(new_n776), .B1(new_n791), .B2(new_n459), .ZN(new_n1194));
  NOR4_X1   g0994(.A1(new_n1194), .A2(new_n1066), .A3(G41), .A4(new_n301), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n780), .A2(G116), .B1(new_n770), .B2(G283), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(new_n786), .A2(G97), .B1(new_n782), .B2(new_n430), .ZN(new_n1197));
  NAND4_X1  g0997(.A1(new_n1195), .A2(new_n1030), .A3(new_n1196), .A4(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(KEYINPUT58), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1193), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(G128), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n791), .A2(new_n1201), .B1(new_n787), .B2(new_n1140), .ZN(new_n1202));
  XNOR2_X1  g1002(.A(new_n1202), .B(KEYINPUT116), .ZN(new_n1203));
  OAI22_X1  g1003(.A1(new_n783), .A2(new_n1025), .B1(new_n1141), .B2(new_n785), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1204), .B1(G125), .B2(new_n780), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n1203), .B(new_n1205), .C1(new_n855), .C2(new_n795), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1206), .A2(KEYINPUT59), .ZN(new_n1207));
  AOI211_X1 g1007(.A(G33), .B(G41), .C1(new_n770), .C2(G124), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n1207), .B(new_n1208), .C1(new_n772), .C2(new_n776), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n1206), .A2(KEYINPUT59), .ZN(new_n1210));
  OAI221_X1 g1010(.A(new_n1200), .B1(new_n1199), .B2(new_n1198), .C1(new_n1209), .C2(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1191), .B1(new_n1211), .B2(new_n767), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n1188), .A2(new_n760), .B1(new_n1189), .B2(new_n1212), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1161), .A2(new_n1126), .A3(new_n1123), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1160), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  AND3_X1   g1016(.A1(new_n1166), .A2(new_n1174), .A3(new_n1184), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1184), .B1(new_n1166), .B2(new_n1174), .ZN(new_n1218));
  OAI211_X1 g1018(.A(new_n1216), .B(KEYINPUT57), .C1(new_n1217), .C2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1219), .A2(new_n757), .ZN(new_n1220));
  AOI21_X1  g1020(.A(KEYINPUT57), .B1(new_n1188), .B2(new_n1216), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1213), .B1(new_n1220), .B2(new_n1221), .ZN(G375));
  INV_X1    g1022(.A(new_n1161), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1223), .A2(new_n1224), .A3(new_n991), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1151), .A2(KEYINPUT120), .A3(new_n809), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT120), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1227), .B1(new_n882), .B2(new_n810), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n842), .B1(new_n843), .B2(G68), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n788), .A2(G97), .B1(new_n780), .B2(G294), .ZN(new_n1230));
  OAI221_X1 g1030(.A(new_n1230), .B1(new_n459), .B2(new_n783), .C1(new_n520), .C2(new_n785), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(new_n805), .A2(G283), .B1(G303), .B2(new_n770), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n301), .B1(new_n798), .B2(G77), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1232), .A2(new_n1233), .A3(new_n1068), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(new_n805), .A2(G137), .B1(G128), .B2(new_n770), .ZN(new_n1235));
  OAI221_X1 g1035(.A(new_n1235), .B1(new_n772), .B2(new_n787), .C1(new_n785), .C2(new_n1140), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n303), .B1(new_n798), .B2(G58), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n780), .A2(G132), .B1(new_n782), .B2(G150), .ZN(new_n1238));
  OAI211_X1 g1038(.A(new_n1237), .B(new_n1238), .C1(new_n202), .C2(new_n795), .ZN(new_n1239));
  OAI22_X1  g1039(.A1(new_n1231), .A2(new_n1234), .B1(new_n1236), .B2(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1229), .B1(new_n767), .B2(new_n1240), .ZN(new_n1241));
  AND3_X1   g1041(.A1(new_n1226), .A2(new_n1228), .A3(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1159), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1242), .B1(new_n1243), .B2(new_n760), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1225), .A2(new_n1244), .ZN(G381));
  OAI211_X1 g1045(.A(new_n1164), .B(new_n1213), .C1(new_n1220), .C2(new_n1221), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1086), .A2(new_n825), .A3(new_n1087), .ZN(new_n1248));
  NOR4_X1   g1048(.A1(G381), .A2(G390), .A3(G384), .A4(new_n1248), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1247), .A2(new_n1019), .A3(new_n1050), .A4(new_n1249), .ZN(G407));
  NAND2_X1  g1050(.A1(new_n688), .A2(G213), .ZN(new_n1251));
  XNOR2_X1  g1051(.A(new_n1251), .B(KEYINPUT121), .ZN(new_n1252));
  OAI211_X1 g1052(.A(G407), .B(G213), .C1(new_n1246), .C2(new_n1252), .ZN(G409));
  XNOR2_X1  g1053(.A(new_n987), .B(new_n988), .ZN(new_n1254));
  AND3_X1   g1054(.A1(new_n998), .A2(new_n1000), .A3(new_n1003), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1003), .B1(new_n998), .B2(new_n1000), .ZN(new_n1256));
  NOR3_X1   g1056(.A1(new_n1255), .A2(new_n1256), .A3(new_n1110), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n991), .B1(new_n1257), .B2(new_n754), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1254), .B1(new_n1258), .B2(new_n759), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1050), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1112), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1019), .A2(new_n1050), .A3(G390), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(G393), .A2(G396), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1263), .A2(new_n1248), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1261), .A2(new_n1262), .A3(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT126), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1261), .A2(KEYINPUT126), .A3(new_n1262), .A4(new_n1264), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT125), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1261), .A2(new_n1269), .A3(new_n1262), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1110), .B1(new_n1001), .B2(KEYINPUT108), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n754), .B1(new_n1271), .B2(new_n1004), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n759), .B1(new_n1272), .B2(new_n992), .ZN(new_n1273));
  AOI211_X1 g1073(.A(new_n1260), .B(new_n1112), .C1(new_n1273), .C2(new_n990), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1264), .B1(new_n1274), .B2(KEYINPUT125), .ZN(new_n1275));
  AOI22_X1  g1075(.A1(new_n1267), .A2(new_n1268), .B1(new_n1270), .B2(new_n1275), .ZN(new_n1276));
  AOI21_X1  g1076(.A(KEYINPUT60), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT122), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1278), .A2(new_n1279), .A3(new_n1223), .ZN(new_n1280));
  OAI21_X1  g1080(.A(KEYINPUT122), .B1(new_n1277), .B2(new_n1161), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1224), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n719), .B1(new_n1282), .B2(KEYINPUT60), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1280), .A2(new_n1281), .A3(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1284), .A2(new_n1244), .ZN(new_n1285));
  INV_X1    g1085(.A(G384), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1284), .A2(G384), .A3(new_n1244), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(KEYINPUT61), .B1(new_n1289), .B2(KEYINPUT62), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT123), .ZN(new_n1291));
  INV_X1    g1091(.A(G2897), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1251), .B1(new_n1291), .B2(new_n1292), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1293), .B1(new_n1291), .B2(new_n1292), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1287), .A2(new_n1288), .A3(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT124), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  NAND4_X1  g1097(.A1(new_n1287), .A2(KEYINPUT124), .A3(new_n1288), .A4(new_n1294), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  NOR2_X1   g1099(.A1(new_n1252), .A2(new_n1292), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1289), .A2(new_n1300), .ZN(new_n1301));
  AOI21_X1  g1101(.A(KEYINPUT62), .B1(new_n1299), .B2(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(G375), .A2(G378), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1216), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1304));
  OAI211_X1 g1104(.A(new_n1213), .B(new_n1164), .C1(new_n992), .C2(new_n1304), .ZN(new_n1305));
  AND3_X1   g1105(.A1(new_n1303), .A2(new_n1252), .A3(new_n1305), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1290), .B1(new_n1302), .B2(new_n1306), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1303), .A2(new_n1251), .A3(new_n1305), .ZN(new_n1308));
  NOR3_X1   g1108(.A1(new_n1308), .A2(KEYINPUT62), .A3(new_n1289), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1276), .B1(new_n1307), .B2(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1289), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1306), .A2(KEYINPUT63), .A3(new_n1311), .ZN(new_n1312));
  NOR2_X1   g1112(.A1(new_n1276), .A2(KEYINPUT61), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT63), .ZN(new_n1314));
  AOI22_X1  g1114(.A1(new_n1297), .A2(new_n1298), .B1(new_n1289), .B2(new_n1300), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1314), .B1(new_n1315), .B2(new_n1308), .ZN(new_n1316));
  NOR2_X1   g1116(.A1(new_n1308), .A2(new_n1289), .ZN(new_n1317));
  OAI211_X1 g1117(.A(new_n1312), .B(new_n1313), .C1(new_n1316), .C2(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1310), .A2(new_n1318), .ZN(G405));
  NAND2_X1  g1119(.A1(new_n1275), .A2(new_n1270), .ZN(new_n1320));
  AOI21_X1  g1120(.A(G390), .B1(new_n1019), .B2(new_n1050), .ZN(new_n1321));
  NOR2_X1   g1121(.A1(new_n1274), .A2(new_n1321), .ZN(new_n1322));
  AOI21_X1  g1122(.A(KEYINPUT126), .B1(new_n1322), .B2(new_n1264), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1268), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n1320), .B1(new_n1323), .B2(new_n1324), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1325), .A2(new_n1246), .A3(new_n1303), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT57), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1304), .A2(new_n1327), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1328), .A2(new_n757), .A3(new_n1219), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1164), .B1(new_n1329), .B2(new_n1213), .ZN(new_n1330));
  OAI21_X1  g1130(.A(new_n1276), .B1(new_n1247), .B2(new_n1330), .ZN(new_n1331));
  INV_X1    g1131(.A(KEYINPUT127), .ZN(new_n1332));
  AND3_X1   g1132(.A1(new_n1326), .A2(new_n1331), .A3(new_n1332), .ZN(new_n1333));
  AOI21_X1  g1133(.A(new_n1332), .B1(new_n1326), .B2(new_n1331), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1289), .B1(new_n1333), .B2(new_n1334), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1326), .A2(new_n1331), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1336), .A2(KEYINPUT127), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n1326), .A2(new_n1331), .A3(new_n1332), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1337), .A2(new_n1311), .A3(new_n1338), .ZN(new_n1339));
  AND2_X1   g1139(.A1(new_n1335), .A2(new_n1339), .ZN(G402));
endmodule


