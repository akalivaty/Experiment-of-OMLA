//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 0 0 1 1 1 1 1 0 1 1 0 1 0 0 0 1 0 1 0 0 1 0 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 0 1 0 1 1 0 0 0 1 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:05 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1238, new_n1239, new_n1240, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311,
    new_n1312;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  NOR2_X1   g0003(.A1(G97), .A2(G107), .ZN(new_n204));
  INV_X1    g0004(.A(new_n204), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n205), .A2(G87), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(new_n208), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n202), .A2(G50), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(new_n213), .A2(KEYINPUT0), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n218), .B1(KEYINPUT0), .B2(new_n213), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT64), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n221));
  INV_X1    g0021(.A(G77), .ZN(new_n222));
  INV_X1    g0022(.A(G244), .ZN(new_n223));
  INV_X1    g0023(.A(G107), .ZN(new_n224));
  INV_X1    g0024(.A(G264), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n221), .B1(new_n222), .B2(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n210), .B1(new_n226), .B2(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT1), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n220), .A2(new_n231), .ZN(G361));
  XOR2_X1   g0032(.A(G238), .B(G244), .Z(new_n233));
  XNOR2_X1  g0033(.A(G226), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n237), .B(new_n240), .Z(G358));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT66), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G68), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G58), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n245), .B(new_n248), .Z(G351));
  NAND2_X1  g0049(.A1(G33), .A2(G41), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n250), .A2(G1), .A3(G13), .ZN(new_n251));
  OR2_X1    g0051(.A1(KEYINPUT3), .A2(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(KEYINPUT3), .A2(G33), .ZN(new_n253));
  AOI21_X1  g0053(.A(G1698), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  AND2_X1   g0054(.A1(KEYINPUT3), .A2(G33), .ZN(new_n255));
  NOR2_X1   g0055(.A1(KEYINPUT3), .A2(G33), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  AOI22_X1  g0057(.A1(new_n254), .A2(G222), .B1(new_n257), .B2(G77), .ZN(new_n258));
  XNOR2_X1  g0058(.A(KEYINPUT3), .B(G33), .ZN(new_n259));
  XNOR2_X1  g0059(.A(KEYINPUT68), .B(G223), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n259), .A2(new_n260), .A3(G1698), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n258), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(KEYINPUT69), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT69), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n258), .A2(new_n264), .A3(new_n261), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n251), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT70), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n251), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  XNOR2_X1  g0070(.A(KEYINPUT67), .B(G226), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G41), .ZN(new_n273));
  INV_X1    g0073(.A(G45), .ZN(new_n274));
  AOI21_X1  g0074(.A(G1), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n275), .A2(new_n251), .A3(G274), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n272), .A2(new_n276), .ZN(new_n277));
  NOR3_X1   g0077(.A1(new_n266), .A2(new_n267), .A3(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n267), .B1(new_n266), .B2(new_n277), .ZN(new_n280));
  INV_X1    g0080(.A(G169), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n279), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(new_n214), .ZN(new_n284));
  XNOR2_X1  g0084(.A(KEYINPUT8), .B(G58), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n208), .A2(G33), .ZN(new_n286));
  INV_X1    g0086(.A(G150), .ZN(new_n287));
  NOR2_X1   g0087(.A1(G20), .A2(G33), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  OAI22_X1  g0089(.A1(new_n285), .A2(new_n286), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G50), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n208), .B1(new_n201), .B2(new_n291), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n284), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n207), .A2(G13), .A3(G20), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n295), .A2(new_n284), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n291), .B1(new_n207), .B2(G20), .ZN(new_n297));
  AOI22_X1  g0097(.A1(new_n296), .A2(new_n297), .B1(new_n291), .B2(new_n295), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n293), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n282), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(KEYINPUT71), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT71), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n282), .A2(new_n302), .A3(new_n299), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT72), .ZN(new_n304));
  INV_X1    g0104(.A(G179), .ZN(new_n305));
  INV_X1    g0105(.A(new_n280), .ZN(new_n306));
  OAI211_X1 g0106(.A(new_n304), .B(new_n305), .C1(new_n306), .C2(new_n278), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n305), .B1(new_n306), .B2(new_n278), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(KEYINPUT72), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n301), .A2(new_n303), .A3(new_n307), .A4(new_n309), .ZN(new_n310));
  OAI21_X1  g0110(.A(G190), .B1(new_n306), .B2(new_n278), .ZN(new_n311));
  XOR2_X1   g0111(.A(KEYINPUT74), .B(G200), .Z(new_n312));
  NAND3_X1  g0112(.A1(new_n279), .A2(new_n280), .A3(new_n312), .ZN(new_n313));
  XNOR2_X1  g0113(.A(new_n299), .B(KEYINPUT9), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n311), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(KEYINPUT10), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT10), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n311), .A2(new_n313), .A3(new_n317), .A4(new_n314), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n310), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT16), .ZN(new_n321));
  INV_X1    g0121(.A(G68), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT7), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n323), .B1(new_n259), .B2(G20), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n257), .A2(KEYINPUT7), .A3(new_n208), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n322), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(G58), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n327), .A2(new_n322), .ZN(new_n328));
  OAI21_X1  g0128(.A(G20), .B1(new_n328), .B2(new_n201), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n288), .A2(G159), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n321), .B1(new_n326), .B2(new_n331), .ZN(new_n332));
  AOI21_X1  g0132(.A(KEYINPUT7), .B1(new_n257), .B2(new_n208), .ZN(new_n333));
  NOR4_X1   g0133(.A1(new_n255), .A2(new_n256), .A3(new_n323), .A4(G20), .ZN(new_n334));
  OAI21_X1  g0134(.A(G68), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n331), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n335), .A2(KEYINPUT16), .A3(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n332), .A2(new_n337), .A3(new_n284), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n285), .B1(new_n207), .B2(G20), .ZN(new_n339));
  AOI22_X1  g0139(.A1(new_n339), .A2(new_n296), .B1(new_n295), .B2(new_n285), .ZN(new_n340));
  AND2_X1   g0140(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  OAI211_X1 g0141(.A(G226), .B(G1698), .C1(new_n255), .C2(new_n256), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(KEYINPUT75), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT75), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n259), .A2(new_n344), .A3(G226), .A4(G1698), .ZN(new_n345));
  NAND2_X1  g0145(.A1(G33), .A2(G87), .ZN(new_n346));
  INV_X1    g0146(.A(G1698), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n259), .A2(G223), .A3(new_n347), .ZN(new_n348));
  NAND4_X1  g0148(.A1(new_n343), .A2(new_n345), .A3(new_n346), .A4(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n251), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(G232), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n276), .B1(new_n269), .B2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n351), .A2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(G200), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n353), .B1(new_n349), .B2(new_n350), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT76), .ZN(new_n359));
  INV_X1    g0159(.A(G190), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n358), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n357), .A2(new_n361), .ZN(new_n362));
  AOI211_X1 g0162(.A(G190), .B(new_n353), .C1(new_n349), .C2(new_n350), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n363), .A2(new_n359), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n341), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT17), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  OAI211_X1 g0167(.A(new_n341), .B(KEYINPUT17), .C1(new_n362), .C2(new_n364), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n351), .A2(new_n305), .A3(new_n354), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n370), .B1(G169), .B2(new_n358), .ZN(new_n371));
  OAI21_X1  g0171(.A(KEYINPUT18), .B1(new_n341), .B2(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(G169), .B1(new_n351), .B2(new_n354), .ZN(new_n373));
  AOI211_X1 g0173(.A(G179), .B(new_n353), .C1(new_n349), .C2(new_n350), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n338), .A2(new_n340), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT18), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n375), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n372), .A2(new_n378), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n369), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n295), .A2(new_n322), .ZN(new_n381));
  XNOR2_X1  g0181(.A(new_n381), .B(KEYINPUT12), .ZN(new_n382));
  AOI22_X1  g0182(.A1(new_n288), .A2(G50), .B1(G20), .B2(new_n322), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n383), .B1(new_n222), .B2(new_n286), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n384), .A2(KEYINPUT11), .A3(new_n284), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n207), .A2(G20), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n296), .A2(G68), .A3(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n382), .A2(new_n385), .A3(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(KEYINPUT11), .B1(new_n384), .B2(new_n284), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT14), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n254), .A2(G226), .ZN(new_n393));
  NAND2_X1  g0193(.A1(G33), .A2(G97), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n259), .A2(G232), .A3(G1698), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n393), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(new_n350), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT13), .ZN(new_n398));
  INV_X1    g0198(.A(new_n276), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n399), .B1(G238), .B2(new_n270), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n397), .A2(new_n398), .A3(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n398), .B1(new_n397), .B2(new_n400), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n392), .B(G169), .C1(new_n402), .C2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n403), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n405), .A2(G179), .A3(new_n401), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n405), .A2(new_n401), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n392), .B1(new_n408), .B2(G169), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n391), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n402), .A2(new_n403), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(G190), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n408), .A2(G200), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n412), .A2(new_n413), .A3(new_n390), .ZN(new_n414));
  NAND2_X1  g0214(.A1(G20), .A2(G77), .ZN(new_n415));
  XNOR2_X1  g0215(.A(KEYINPUT15), .B(G87), .ZN(new_n416));
  OAI221_X1 g0216(.A(new_n415), .B1(new_n416), .B2(new_n286), .C1(new_n289), .C2(new_n285), .ZN(new_n417));
  AOI22_X1  g0217(.A1(new_n417), .A2(new_n284), .B1(new_n222), .B2(new_n295), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n296), .A2(G77), .A3(new_n386), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT73), .ZN(new_n420));
  AND2_X1   g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n419), .A2(new_n420), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n418), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n276), .B1(new_n269), .B2(new_n223), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n259), .A2(G232), .A3(new_n347), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n259), .A2(G238), .A3(G1698), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n425), .B(new_n426), .C1(new_n224), .C2(new_n259), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n424), .B1(new_n427), .B2(new_n350), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n423), .B1(new_n312), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n428), .A2(G190), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n429), .A2(new_n281), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n428), .A2(new_n305), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n433), .A2(new_n434), .A3(new_n423), .ZN(new_n435));
  AND2_X1   g0235(.A1(new_n432), .A2(new_n435), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n380), .A2(new_n410), .A3(new_n414), .A4(new_n436), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n320), .A2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT6), .ZN(new_n439));
  AND2_X1   g0239(.A1(G97), .A2(G107), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n439), .B1(new_n440), .B2(new_n204), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n224), .A2(KEYINPUT6), .A3(G97), .ZN(new_n442));
  AND2_X1   g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  OAI22_X1  g0243(.A1(new_n443), .A2(new_n208), .B1(new_n222), .B2(new_n289), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n224), .B1(new_n324), .B2(new_n325), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n284), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n294), .A2(G97), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n207), .A2(G33), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n294), .A2(new_n448), .A3(new_n214), .A4(new_n283), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n447), .B1(new_n450), .B2(G97), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n446), .A2(new_n451), .ZN(new_n452));
  OAI211_X1 g0252(.A(G250), .B(G1698), .C1(new_n255), .C2(new_n256), .ZN(new_n453));
  NAND2_X1  g0253(.A1(G33), .A2(G283), .ZN(new_n454));
  OAI211_X1 g0254(.A(G244), .B(new_n347), .C1(new_n255), .C2(new_n256), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT4), .ZN(new_n456));
  OAI211_X1 g0256(.A(new_n453), .B(new_n454), .C1(new_n455), .C2(new_n456), .ZN(new_n457));
  AOI21_X1  g0257(.A(KEYINPUT4), .B1(new_n254), .B2(G244), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n350), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n207), .A2(G45), .ZN(new_n460));
  NOR2_X1   g0260(.A1(KEYINPUT5), .A2(G41), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(KEYINPUT5), .A2(G41), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n460), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(G274), .ZN(new_n465));
  INV_X1    g0265(.A(new_n214), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n465), .B1(new_n466), .B2(new_n250), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n274), .A2(G1), .ZN(new_n469));
  INV_X1    g0269(.A(new_n463), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n469), .B1(new_n470), .B2(new_n461), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n471), .A2(G257), .A3(new_n251), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n468), .A2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n459), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(new_n281), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n455), .A2(new_n456), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n259), .A2(KEYINPUT4), .A3(G244), .A4(new_n347), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n477), .A2(new_n478), .A3(new_n453), .A4(new_n454), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n473), .B1(new_n479), .B2(new_n350), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(new_n305), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n452), .A2(new_n476), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n475), .A2(G200), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n480), .A2(G190), .ZN(new_n484));
  INV_X1    g0284(.A(new_n451), .ZN(new_n485));
  OAI21_X1  g0285(.A(G107), .B1(new_n333), .B2(new_n334), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n441), .A2(new_n442), .ZN(new_n487));
  AOI22_X1  g0287(.A1(new_n487), .A2(G20), .B1(G77), .B2(new_n288), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n485), .B1(new_n489), .B2(new_n284), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n483), .A2(new_n484), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n254), .A2(G238), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n259), .A2(G244), .A3(G1698), .ZN(new_n493));
  NAND2_X1  g0293(.A1(G33), .A2(G116), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n492), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(new_n350), .ZN(new_n496));
  AND2_X1   g0296(.A1(new_n460), .A2(G250), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(new_n251), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n251), .A2(G274), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n498), .B1(new_n460), .B2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n496), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(new_n312), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n259), .A2(new_n208), .A3(G68), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT19), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n208), .B1(new_n394), .B2(new_n505), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n506), .B1(G87), .B2(new_n205), .ZN(new_n507));
  INV_X1    g0307(.A(G97), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n505), .B1(new_n286), .B2(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n504), .A2(new_n507), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(new_n284), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n416), .A2(new_n295), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n450), .A2(G87), .ZN(new_n513));
  AND3_X1   g0313(.A1(new_n511), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n500), .B1(new_n350), .B2(new_n495), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(G190), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n503), .A2(new_n514), .A3(new_n516), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n511), .B(new_n512), .C1(new_n449), .C2(new_n416), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n496), .A2(new_n305), .A3(new_n501), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n518), .B(new_n519), .C1(new_n515), .C2(G169), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n482), .A2(new_n491), .A3(new_n517), .A4(new_n520), .ZN(new_n521));
  AOI21_X1  g0321(.A(KEYINPUT25), .B1(new_n295), .B2(new_n224), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n295), .A2(KEYINPUT25), .A3(new_n224), .ZN(new_n524));
  AOI22_X1  g0324(.A1(new_n523), .A2(new_n524), .B1(G107), .B2(new_n450), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  OAI21_X1  g0326(.A(KEYINPUT23), .B1(new_n208), .B2(G107), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT23), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n528), .A2(new_n224), .A3(G20), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n208), .A2(G33), .A3(G116), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n527), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT78), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n527), .A2(new_n529), .A3(new_n530), .A4(KEYINPUT78), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n208), .B(G87), .C1(new_n255), .C2(new_n256), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(KEYINPUT22), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT22), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n259), .A2(new_n538), .A3(new_n208), .A4(G87), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n535), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(KEYINPUT79), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT79), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n535), .A2(new_n540), .A3(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n542), .A2(KEYINPUT24), .A3(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(new_n284), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n543), .B1(new_n535), .B2(new_n540), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT24), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n526), .B1(new_n545), .B2(new_n549), .ZN(new_n550));
  NOR3_X1   g0350(.A1(new_n464), .A2(new_n225), .A3(new_n350), .ZN(new_n551));
  OAI211_X1 g0351(.A(G257), .B(G1698), .C1(new_n255), .C2(new_n256), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT80), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n259), .A2(KEYINPUT80), .A3(G257), .A4(G1698), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n259), .A2(G250), .A3(new_n347), .ZN(new_n556));
  NAND2_X1  g0356(.A1(G33), .A2(G294), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n554), .A2(new_n555), .A3(new_n556), .A4(new_n557), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n551), .B1(new_n558), .B2(new_n350), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n559), .A2(new_n360), .A3(new_n468), .ZN(new_n560));
  INV_X1    g0360(.A(new_n468), .ZN(new_n561));
  AOI211_X1 g0361(.A(new_n551), .B(new_n561), .C1(new_n558), .C2(new_n350), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n560), .B1(new_n562), .B2(G200), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n550), .A2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT82), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n550), .A2(KEYINPUT82), .A3(new_n563), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n521), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT81), .ZN(new_n569));
  AND3_X1   g0369(.A1(new_n559), .A2(G179), .A3(new_n468), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n281), .B1(new_n559), .B2(new_n468), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n569), .B1(new_n572), .B2(new_n550), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n454), .B(new_n208), .C1(G33), .C2(new_n508), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT77), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT20), .ZN(new_n576));
  INV_X1    g0376(.A(G116), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n575), .A2(new_n576), .B1(new_n577), .B2(G20), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n574), .A2(new_n578), .A3(new_n284), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n575), .A2(new_n576), .ZN(new_n580));
  OR2_X1    g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n294), .A2(new_n577), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n582), .B1(new_n450), .B2(new_n577), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n579), .A2(new_n580), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n581), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  XNOR2_X1  g0385(.A(KEYINPUT5), .B(G41), .ZN(new_n586));
  AOI22_X1  g0386(.A1(new_n586), .A2(new_n469), .B1(new_n466), .B2(new_n250), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n587), .A2(G270), .B1(new_n464), .B2(new_n467), .ZN(new_n588));
  OAI211_X1 g0388(.A(G264), .B(G1698), .C1(new_n255), .C2(new_n256), .ZN(new_n589));
  OAI211_X1 g0389(.A(G257), .B(new_n347), .C1(new_n255), .C2(new_n256), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n252), .A2(G303), .A3(new_n253), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n350), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n588), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n585), .A2(new_n594), .A3(G169), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT21), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n594), .A2(G200), .ZN(new_n598));
  INV_X1    g0398(.A(new_n585), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n598), .B(new_n599), .C1(new_n360), .C2(new_n594), .ZN(new_n600));
  AND3_X1   g0400(.A1(new_n588), .A2(G179), .A3(new_n593), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n585), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n585), .A2(new_n594), .A3(KEYINPUT21), .A4(G169), .ZN(new_n603));
  AND4_X1   g0403(.A1(new_n597), .A2(new_n600), .A3(new_n602), .A4(new_n603), .ZN(new_n604));
  AND3_X1   g0404(.A1(new_n535), .A2(new_n540), .A3(new_n543), .ZN(new_n605));
  NOR3_X1   g0405(.A1(new_n605), .A2(new_n547), .A3(new_n548), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n541), .A2(KEYINPUT79), .A3(new_n548), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n284), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n525), .B1(new_n606), .B2(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n559), .A2(G179), .A3(new_n468), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n610), .B1(new_n562), .B2(new_n281), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n609), .A2(KEYINPUT81), .A3(new_n611), .ZN(new_n612));
  AND3_X1   g0412(.A1(new_n573), .A2(new_n604), .A3(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n438), .A2(new_n568), .A3(new_n613), .ZN(new_n614));
  XOR2_X1   g0414(.A(new_n614), .B(KEYINPUT83), .Z(G372));
  INV_X1    g0415(.A(new_n319), .ZN(new_n616));
  AND3_X1   g0416(.A1(new_n412), .A2(new_n413), .A3(new_n390), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n435), .A2(KEYINPUT84), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT84), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n433), .A2(new_n619), .A3(new_n423), .A4(new_n434), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n410), .B1(new_n617), .B2(new_n621), .ZN(new_n622));
  AND2_X1   g0422(.A1(new_n367), .A2(new_n368), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n379), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n310), .B1(new_n616), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(KEYINPUT85), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT85), .ZN(new_n627));
  OAI211_X1 g0427(.A(new_n627), .B(new_n310), .C1(new_n616), .C2(new_n624), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n609), .A2(new_n611), .ZN(new_n630));
  AND3_X1   g0430(.A1(new_n597), .A2(new_n602), .A3(new_n603), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  AND4_X1   g0432(.A1(new_n482), .A2(new_n491), .A3(new_n517), .A4(new_n520), .ZN(new_n633));
  AOI21_X1  g0433(.A(KEYINPUT82), .B1(new_n550), .B2(new_n563), .ZN(new_n634));
  AND3_X1   g0434(.A1(new_n550), .A2(KEYINPUT82), .A3(new_n563), .ZN(new_n635));
  OAI211_X1 g0435(.A(new_n632), .B(new_n633), .C1(new_n634), .C2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n520), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT26), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n517), .A2(new_n520), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n638), .B1(new_n639), .B2(new_n482), .ZN(new_n640));
  INV_X1    g0440(.A(new_n482), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n641), .A2(KEYINPUT26), .A3(new_n520), .A4(new_n517), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n637), .B1(new_n640), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n636), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n438), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n629), .A2(new_n645), .ZN(G369));
  NAND3_X1  g0446(.A1(new_n207), .A2(new_n208), .A3(G13), .ZN(new_n647));
  OR2_X1    g0447(.A1(new_n647), .A2(KEYINPUT27), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(KEYINPUT27), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n648), .A2(new_n649), .A3(G213), .ZN(new_n650));
  INV_X1    g0450(.A(G343), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  OAI22_X1  g0453(.A1(new_n635), .A2(new_n634), .B1(new_n550), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n573), .A2(new_n612), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT87), .ZN(new_n656));
  NOR3_X1   g0456(.A1(new_n630), .A2(new_n656), .A3(new_n653), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n572), .A2(new_n550), .ZN(new_n658));
  AOI21_X1  g0458(.A(KEYINPUT87), .B1(new_n658), .B2(new_n652), .ZN(new_n659));
  OAI22_X1  g0459(.A1(new_n654), .A2(new_n655), .B1(new_n657), .B2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n599), .A2(new_n653), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n631), .A2(new_n600), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT86), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n662), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n604), .A2(KEYINPUT86), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n631), .A2(new_n662), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n667), .A2(G330), .A3(new_n668), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n661), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n630), .A2(new_n652), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n631), .A2(new_n652), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n672), .B1(new_n660), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n671), .A2(new_n674), .ZN(G399));
  INV_X1    g0475(.A(new_n211), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n676), .A2(G41), .ZN(new_n677));
  INV_X1    g0477(.A(G87), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n204), .A2(new_n678), .A3(new_n577), .ZN(new_n679));
  XOR2_X1   g0479(.A(new_n679), .B(KEYINPUT88), .Z(new_n680));
  NOR3_X1   g0480(.A1(new_n677), .A2(new_n680), .A3(new_n207), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n681), .B1(new_n217), .B2(new_n677), .ZN(new_n682));
  XNOR2_X1  g0482(.A(KEYINPUT89), .B(KEYINPUT28), .ZN(new_n683));
  XNOR2_X1  g0483(.A(new_n682), .B(new_n683), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n601), .A2(new_n559), .A3(new_n480), .A4(new_n515), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT30), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  AND3_X1   g0487(.A1(new_n459), .A2(new_n474), .A3(KEYINPUT30), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n688), .A2(new_n559), .A3(new_n515), .A4(new_n601), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n559), .A2(new_n468), .ZN(new_n690));
  AOI21_X1  g0490(.A(G179), .B1(new_n496), .B2(new_n501), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n690), .A2(new_n691), .A3(new_n475), .A4(new_n594), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n687), .A2(new_n689), .A3(new_n692), .ZN(new_n693));
  AND3_X1   g0493(.A1(new_n693), .A2(KEYINPUT31), .A3(new_n652), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT90), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n687), .A2(KEYINPUT90), .A3(new_n692), .A4(new_n689), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n696), .A2(new_n652), .A3(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT31), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n694), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(KEYINPUT91), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT91), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n653), .B1(new_n693), .B2(new_n695), .ZN(new_n703));
  AOI21_X1  g0503(.A(KEYINPUT31), .B1(new_n703), .B2(new_n697), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n702), .B1(new_n704), .B2(new_n694), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n613), .A2(new_n568), .A3(new_n653), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n701), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(G330), .ZN(new_n708));
  AOI211_X1 g0508(.A(KEYINPUT29), .B(new_n652), .C1(new_n636), .C2(new_n643), .ZN(new_n709));
  AND3_X1   g0509(.A1(new_n573), .A2(new_n612), .A3(new_n631), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n633), .B1(new_n635), .B2(new_n634), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n643), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(new_n653), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n709), .B1(KEYINPUT29), .B2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n708), .A2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n684), .B1(new_n716), .B2(G1), .ZN(G364));
  AND2_X1   g0517(.A1(new_n208), .A2(G13), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n207), .B1(new_n718), .B2(G45), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n677), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(G13), .A2(G33), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n723), .A2(G20), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n214), .B1(G20), .B2(new_n281), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n676), .A2(new_n257), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(G355), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n729), .B1(G116), .B2(new_n211), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n676), .A2(new_n259), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n732), .B1(new_n274), .B2(new_n217), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n248), .A2(G45), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n730), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n208), .A2(G179), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n312), .A2(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(G190), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(G107), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n737), .A2(new_n360), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n739), .B1(new_n741), .B2(new_n678), .ZN(new_n742));
  NOR2_X1   g0542(.A1(G190), .A2(G200), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n736), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(G159), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT32), .ZN(new_n747));
  NAND2_X1  g0547(.A1(G20), .A2(G179), .ZN(new_n748));
  NOR3_X1   g0548(.A1(new_n748), .A2(new_n360), .A3(new_n356), .ZN(new_n749));
  AOI22_X1  g0549(.A1(new_n746), .A2(new_n747), .B1(G50), .B2(new_n749), .ZN(new_n750));
  NOR3_X1   g0550(.A1(new_n360), .A2(G179), .A3(G200), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(new_n208), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n750), .B1(new_n508), .B2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n748), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(new_n743), .ZN(new_n755));
  NOR3_X1   g0555(.A1(new_n748), .A2(new_n360), .A3(G200), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  OAI221_X1 g0557(.A(new_n259), .B1(new_n755), .B2(new_n222), .C1(new_n757), .C2(new_n327), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n754), .A2(new_n360), .A3(G200), .ZN(new_n759));
  OAI22_X1  g0559(.A1(new_n746), .A2(new_n747), .B1(new_n322), .B2(new_n759), .ZN(new_n760));
  NOR4_X1   g0560(.A1(new_n742), .A2(new_n753), .A3(new_n758), .A4(new_n760), .ZN(new_n761));
  OR2_X1    g0561(.A1(new_n741), .A2(KEYINPUT92), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n741), .A2(KEYINPUT92), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(G303), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g0566(.A(KEYINPUT33), .B(G317), .ZN(new_n767));
  AND2_X1   g0567(.A1(new_n767), .A2(KEYINPUT94), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n767), .A2(KEYINPUT94), .ZN(new_n769));
  NOR3_X1   g0569(.A1(new_n768), .A2(new_n769), .A3(new_n759), .ZN(new_n770));
  INV_X1    g0570(.A(G311), .ZN(new_n771));
  INV_X1    g0571(.A(G322), .ZN(new_n772));
  OAI221_X1 g0572(.A(new_n257), .B1(new_n755), .B2(new_n771), .C1(new_n757), .C2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(G326), .ZN(new_n774));
  INV_X1    g0574(.A(new_n749), .ZN(new_n775));
  INV_X1    g0575(.A(G294), .ZN(new_n776));
  OAI22_X1  g0576(.A1(new_n774), .A2(new_n775), .B1(new_n752), .B2(new_n776), .ZN(new_n777));
  NOR4_X1   g0577(.A1(new_n766), .A2(new_n770), .A3(new_n773), .A4(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n744), .ZN(new_n779));
  AOI22_X1  g0579(.A1(new_n738), .A2(G283), .B1(G329), .B2(new_n779), .ZN(new_n780));
  XOR2_X1   g0580(.A(new_n780), .B(KEYINPUT93), .Z(new_n781));
  AOI21_X1  g0581(.A(new_n761), .B1(new_n778), .B2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n725), .ZN(new_n783));
  OAI221_X1 g0583(.A(new_n721), .B1(new_n727), .B2(new_n735), .C1(new_n782), .C2(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n667), .A2(new_n668), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n784), .B1(new_n785), .B2(new_n724), .ZN(new_n786));
  XNOR2_X1  g0586(.A(new_n786), .B(KEYINPUT95), .ZN(new_n787));
  INV_X1    g0587(.A(new_n721), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n669), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(G330), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n789), .B1(new_n790), .B2(new_n785), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n787), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(G396));
  AOI21_X1  g0593(.A(new_n652), .B1(new_n636), .B2(new_n643), .ZN(new_n794));
  NAND4_X1  g0594(.A1(new_n618), .A2(new_n423), .A3(new_n620), .A4(new_n652), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n423), .A2(new_n652), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n432), .A2(new_n435), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  XNOR2_X1  g0598(.A(new_n794), .B(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n721), .B1(new_n708), .B2(new_n799), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n800), .B1(new_n708), .B2(new_n799), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n783), .A2(new_n723), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n721), .B1(G77), .B2(new_n802), .ZN(new_n803));
  XOR2_X1   g0603(.A(new_n803), .B(KEYINPUT96), .Z(new_n804));
  INV_X1    g0604(.A(new_n764), .ZN(new_n805));
  INV_X1    g0605(.A(new_n755), .ZN(new_n806));
  AOI22_X1  g0606(.A1(new_n806), .A2(G159), .B1(G143), .B2(new_n756), .ZN(new_n807));
  INV_X1    g0607(.A(G137), .ZN(new_n808));
  OAI221_X1 g0608(.A(new_n807), .B1(new_n808), .B2(new_n775), .C1(new_n287), .C2(new_n759), .ZN(new_n809));
  INV_X1    g0609(.A(KEYINPUT34), .ZN(new_n810));
  AOI22_X1  g0610(.A1(new_n805), .A2(G50), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(G132), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n259), .B1(new_n744), .B2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n738), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n814), .A2(new_n322), .ZN(new_n815));
  INV_X1    g0615(.A(new_n752), .ZN(new_n816));
  AOI211_X1 g0616(.A(new_n813), .B(new_n815), .C1(G58), .C2(new_n816), .ZN(new_n817));
  OAI211_X1 g0617(.A(new_n811), .B(new_n817), .C1(new_n810), .C2(new_n809), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n257), .B1(new_n764), .B2(new_n224), .ZN(new_n819));
  XOR2_X1   g0619(.A(new_n819), .B(KEYINPUT98), .Z(new_n820));
  AOI22_X1  g0620(.A1(new_n816), .A2(G97), .B1(new_n756), .B2(G294), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n821), .B(KEYINPUT99), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n738), .A2(G87), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n749), .A2(G303), .ZN(new_n824));
  XOR2_X1   g0624(.A(KEYINPUT97), .B(G283), .Z(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n759), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  AOI22_X1  g0628(.A1(G311), .A2(new_n779), .B1(new_n806), .B2(G116), .ZN(new_n829));
  NAND4_X1  g0629(.A1(new_n823), .A2(new_n824), .A3(new_n828), .A4(new_n829), .ZN(new_n830));
  OR2_X1    g0630(.A1(new_n822), .A2(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n818), .B1(new_n820), .B2(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n804), .B1(new_n832), .B2(new_n725), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n833), .B1(new_n723), .B2(new_n798), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n801), .A2(new_n834), .ZN(G384));
  OR2_X1    g0635(.A1(new_n487), .A2(KEYINPUT35), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n487), .A2(KEYINPUT35), .ZN(new_n837));
  NAND4_X1  g0637(.A1(new_n836), .A2(G116), .A3(new_n215), .A4(new_n837), .ZN(new_n838));
  XOR2_X1   g0638(.A(new_n838), .B(KEYINPUT36), .Z(new_n839));
  OR3_X1    g0639(.A1(new_n216), .A2(new_n222), .A3(new_n328), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n291), .A2(G68), .ZN(new_n841));
  AOI211_X1 g0641(.A(new_n207), .B(G13), .C1(new_n840), .C2(new_n841), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT39), .ZN(new_n844));
  INV_X1    g0644(.A(new_n650), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n376), .A2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n847), .B1(new_n369), .B2(new_n379), .ZN(new_n848));
  AOI22_X1  g0648(.A1(new_n363), .A2(new_n359), .B1(new_n355), .B2(new_n356), .ZN(new_n849));
  OAI21_X1  g0649(.A(KEYINPUT76), .B1(new_n355), .B2(G190), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n376), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  AOI22_X1  g0651(.A1(new_n371), .A2(new_n650), .B1(new_n338), .B2(new_n340), .ZN(new_n852));
  OAI21_X1  g0652(.A(KEYINPUT37), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n376), .B1(new_n375), .B2(new_n845), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT37), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n365), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n853), .A2(KEYINPUT100), .A3(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT100), .ZN(new_n858));
  OAI211_X1 g0658(.A(new_n858), .B(KEYINPUT37), .C1(new_n851), .C2(new_n852), .ZN(new_n859));
  AND4_X1   g0659(.A1(KEYINPUT38), .A2(new_n848), .A3(new_n857), .A4(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n853), .A2(KEYINPUT101), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n856), .A2(KEYINPUT102), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT102), .ZN(new_n863));
  NAND4_X1  g0663(.A1(new_n365), .A2(new_n854), .A3(new_n863), .A4(new_n855), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT101), .ZN(new_n865));
  OAI211_X1 g0665(.A(new_n865), .B(KEYINPUT37), .C1(new_n851), .C2(new_n852), .ZN(new_n866));
  NAND4_X1  g0666(.A1(new_n861), .A2(new_n862), .A3(new_n864), .A4(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(KEYINPUT38), .B1(new_n867), .B2(new_n848), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n844), .B1(new_n860), .B2(new_n868), .ZN(new_n869));
  OAI21_X1  g0669(.A(KEYINPUT14), .B1(new_n411), .B2(new_n281), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n870), .A2(new_n406), .A3(new_n404), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n871), .A2(new_n391), .A3(new_n653), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT38), .ZN(new_n874));
  INV_X1    g0674(.A(new_n379), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n846), .B1(new_n623), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n857), .A2(new_n859), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n874), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND4_X1  g0678(.A1(new_n848), .A2(KEYINPUT38), .A3(new_n857), .A4(new_n859), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n878), .A2(KEYINPUT39), .A3(new_n879), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n869), .A2(new_n873), .A3(new_n880), .ZN(new_n881));
  OAI211_X1 g0681(.A(new_n410), .B(new_n414), .C1(new_n390), .C2(new_n653), .ZN(new_n882));
  OAI211_X1 g0682(.A(new_n391), .B(new_n652), .C1(new_n617), .C2(new_n871), .ZN(new_n883));
  AND2_X1   g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n794), .A2(new_n798), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n435), .A2(new_n652), .ZN(new_n886));
  INV_X1    g0686(.A(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n884), .B1(new_n885), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n878), .A2(new_n879), .ZN(new_n889));
  AOI22_X1  g0689(.A1(new_n888), .A2(new_n889), .B1(new_n379), .B2(new_n650), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n881), .A2(new_n890), .ZN(new_n891));
  AND2_X1   g0691(.A1(new_n713), .A2(KEYINPUT29), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n438), .B1(new_n892), .B2(new_n709), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n629), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g0694(.A(new_n891), .B(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n860), .A2(new_n868), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n698), .A2(new_n699), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n703), .A2(KEYINPUT31), .A3(new_n697), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n706), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(new_n798), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n901), .B1(new_n882), .B2(new_n883), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  OAI21_X1  g0703(.A(KEYINPUT40), .B1(new_n897), .B2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT103), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  OAI211_X1 g0706(.A(new_n900), .B(new_n902), .C1(KEYINPUT103), .C2(KEYINPUT40), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n906), .A2(new_n889), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n904), .A2(new_n908), .ZN(new_n909));
  AND2_X1   g0709(.A1(new_n438), .A2(new_n900), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n909), .A2(new_n910), .ZN(new_n913));
  NOR3_X1   g0713(.A1(new_n912), .A2(new_n913), .A3(new_n790), .ZN(new_n914));
  OAI22_X1  g0714(.A1(new_n896), .A2(new_n914), .B1(new_n207), .B2(new_n718), .ZN(new_n915));
  AND2_X1   g0715(.A1(new_n896), .A2(new_n914), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n843), .B1(new_n915), .B2(new_n916), .ZN(G367));
  INV_X1    g0717(.A(new_n673), .ZN(new_n918));
  AOI22_X1  g0718(.A1(new_n566), .A2(new_n567), .B1(new_n609), .B2(new_n652), .ZN(new_n919));
  INV_X1    g0719(.A(new_n655), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n656), .B1(new_n630), .B2(new_n653), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n658), .A2(KEYINPUT87), .A3(new_n652), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n918), .B1(new_n921), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n641), .A2(new_n652), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n482), .B(new_n491), .C1(new_n490), .C2(new_n653), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n925), .A2(new_n928), .ZN(new_n929));
  OR2_X1    g0729(.A1(new_n929), .A2(KEYINPUT42), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n482), .B1(new_n920), .B2(new_n927), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n653), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n929), .A2(KEYINPUT42), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n930), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n514), .A2(new_n653), .ZN(new_n935));
  OR2_X1    g0735(.A1(new_n639), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n637), .A2(new_n935), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT43), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n938), .A2(KEYINPUT43), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n934), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(new_n928), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n671), .A2(new_n944), .ZN(new_n945));
  AND2_X1   g0745(.A1(new_n933), .A2(new_n932), .ZN(new_n946));
  NAND4_X1  g0746(.A1(new_n946), .A2(new_n940), .A3(new_n939), .A4(new_n930), .ZN(new_n947));
  AND3_X1   g0747(.A1(new_n943), .A2(new_n945), .A3(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n945), .B1(new_n943), .B2(new_n947), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  XOR2_X1   g0750(.A(new_n677), .B(KEYINPUT41), .Z(new_n951));
  INV_X1    g0751(.A(KEYINPUT44), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n952), .B1(new_n674), .B2(new_n928), .ZN(new_n953));
  OAI211_X1 g0753(.A(KEYINPUT44), .B(new_n944), .C1(new_n925), .C2(new_n672), .ZN(new_n954));
  AND2_X1   g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n660), .A2(new_n673), .ZN(new_n956));
  INV_X1    g0756(.A(new_n672), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n956), .A2(new_n957), .A3(new_n928), .ZN(new_n958));
  XOR2_X1   g0758(.A(KEYINPUT104), .B(KEYINPUT45), .Z(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n674), .A2(new_n928), .A3(new_n959), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  OAI211_X1 g0763(.A(KEYINPUT105), .B(new_n670), .C1(new_n955), .C2(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(new_n962), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n959), .B1(new_n674), .B2(new_n928), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n953), .A2(new_n954), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n967), .A2(new_n671), .A3(new_n968), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n921), .A2(new_n924), .A3(new_n918), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n669), .B1(new_n970), .B2(KEYINPUT106), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n970), .A2(new_n669), .A3(KEYINPUT106), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n972), .A2(new_n925), .A3(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n973), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n956), .B1(new_n975), .B2(new_n971), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n715), .B1(new_n974), .B2(new_n976), .ZN(new_n977));
  OR2_X1    g0777(.A1(new_n670), .A2(KEYINPUT105), .ZN(new_n978));
  NAND4_X1  g0778(.A1(new_n964), .A2(new_n969), .A3(new_n977), .A4(new_n978), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n951), .B1(new_n979), .B2(new_n716), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n950), .B1(new_n980), .B2(new_n720), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n731), .A2(new_n240), .ZN(new_n982));
  INV_X1    g0782(.A(new_n416), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n727), .B1(new_n676), .B2(new_n983), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n788), .B1(new_n982), .B2(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(new_n724), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n805), .A2(KEYINPUT46), .A3(G116), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT46), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n988), .B1(new_n741), .B2(new_n577), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n257), .B1(new_n825), .B2(new_n755), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n990), .B1(G317), .B2(new_n779), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n738), .A2(G97), .ZN(new_n992));
  AOI22_X1  g0792(.A1(new_n816), .A2(G107), .B1(new_n827), .B2(G294), .ZN(new_n993));
  AND3_X1   g0793(.A1(new_n991), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  AOI22_X1  g0794(.A1(G311), .A2(new_n749), .B1(new_n756), .B2(G303), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT107), .ZN(new_n996));
  NAND4_X1  g0796(.A1(new_n987), .A2(new_n989), .A3(new_n994), .A4(new_n996), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n752), .A2(new_n322), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n998), .B1(G143), .B2(new_n749), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n999), .B1(new_n745), .B2(new_n759), .ZN(new_n1000));
  OAI22_X1  g0800(.A1(new_n757), .A2(new_n287), .B1(new_n755), .B2(new_n291), .ZN(new_n1001));
  XOR2_X1   g0801(.A(KEYINPUT108), .B(G137), .Z(new_n1002));
  INV_X1    g0802(.A(new_n1002), .ZN(new_n1003));
  AOI211_X1 g0803(.A(new_n257), .B(new_n1001), .C1(new_n779), .C2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n738), .A2(G77), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n740), .A2(G58), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n1004), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n997), .B1(new_n1000), .B2(new_n1007), .ZN(new_n1008));
  XOR2_X1   g0808(.A(new_n1008), .B(KEYINPUT47), .Z(new_n1009));
  OAI221_X1 g0809(.A(new_n985), .B1(new_n986), .B2(new_n938), .C1(new_n1009), .C2(new_n783), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n981), .A2(new_n1010), .ZN(G387));
  INV_X1    g0811(.A(new_n977), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n974), .A2(new_n976), .A3(new_n715), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1012), .A2(new_n677), .A3(new_n1013), .ZN(new_n1014));
  OR2_X1    g0814(.A1(new_n237), .A2(new_n274), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n1015), .A2(new_n731), .B1(new_n680), .B2(new_n728), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n285), .A2(G50), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT50), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n274), .B1(new_n322), .B2(new_n222), .C1(new_n1017), .C2(new_n1018), .ZN(new_n1019));
  AOI211_X1 g0819(.A(new_n680), .B(new_n1019), .C1(new_n1018), .C2(new_n1017), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n1016), .A2(new_n1020), .B1(G107), .B2(new_n211), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n788), .B1(new_n1021), .B2(new_n726), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n740), .A2(G77), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n257), .B1(new_n806), .B2(G68), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n779), .A2(G150), .B1(G50), .B2(new_n756), .ZN(new_n1025));
  NAND4_X1  g0825(.A1(new_n992), .A2(new_n1023), .A3(new_n1024), .A4(new_n1025), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n752), .A2(new_n416), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n775), .A2(new_n745), .B1(new_n285), .B2(new_n759), .ZN(new_n1028));
  NOR3_X1   g0828(.A1(new_n1026), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(new_n806), .A2(G303), .B1(G317), .B2(new_n756), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n1030), .B1(new_n771), .B2(new_n759), .C1(new_n772), .C2(new_n775), .ZN(new_n1031));
  XOR2_X1   g0831(.A(new_n1031), .B(KEYINPUT109), .Z(new_n1032));
  INV_X1    g0832(.A(new_n1032), .ZN(new_n1033));
  OR2_X1    g0833(.A1(new_n1033), .A2(KEYINPUT48), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1033), .A2(KEYINPUT48), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n740), .A2(G294), .B1(new_n816), .B2(new_n826), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1034), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n1037), .ZN(new_n1038));
  OR2_X1    g0838(.A1(new_n1038), .A2(KEYINPUT49), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n257), .B1(new_n774), .B2(new_n744), .C1(new_n814), .C2(new_n577), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1040), .B1(new_n1038), .B2(KEYINPUT49), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1029), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1022), .B1(new_n1042), .B2(new_n783), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1043), .B1(new_n661), .B2(new_n724), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n719), .B1(new_n974), .B2(new_n976), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1014), .A2(new_n1046), .ZN(G393));
  NAND3_X1  g0847(.A1(new_n968), .A2(new_n962), .A3(new_n961), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n1048), .A2(new_n670), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n671), .B1(new_n967), .B2(new_n968), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1012), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1051), .A2(new_n979), .A3(new_n677), .ZN(new_n1052));
  OAI21_X1  g0852(.A(KEYINPUT110), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1048), .A2(new_n670), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT110), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1054), .A2(new_n1055), .A3(new_n969), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1053), .A2(new_n720), .A3(new_n1056), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n245), .A2(new_n732), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n726), .B1(new_n508), .B2(new_n211), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n721), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  INV_X1    g0860(.A(G143), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n259), .B1(new_n744), .B2(new_n1061), .C1(new_n285), .C2(new_n755), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n740), .A2(G68), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n816), .A2(G77), .B1(new_n827), .B2(G50), .ZN(new_n1065));
  NAND4_X1  g0865(.A1(new_n823), .A2(new_n1063), .A3(new_n1064), .A4(new_n1065), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(G150), .A2(new_n749), .B1(new_n756), .B2(G159), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1067), .B(KEYINPUT51), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n740), .A2(new_n826), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n257), .B1(new_n755), .B2(new_n776), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(G322), .B2(new_n779), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n816), .A2(G116), .B1(new_n827), .B2(G303), .ZN(new_n1072));
  NAND4_X1  g0872(.A1(new_n739), .A2(new_n1069), .A3(new_n1071), .A4(new_n1072), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(G317), .A2(new_n749), .B1(new_n756), .B2(G311), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(KEYINPUT111), .B(KEYINPUT52), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n1074), .B(new_n1075), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n1066), .A2(new_n1068), .B1(new_n1073), .B2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1060), .B1(new_n725), .B2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1078), .B1(new_n928), .B2(new_n986), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1052), .A2(new_n1057), .A3(new_n1079), .ZN(G390));
  NAND2_X1  g0880(.A1(new_n869), .A2(new_n880), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n886), .B1(new_n794), .B2(new_n798), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n872), .B1(new_n1082), .B2(new_n884), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n884), .ZN(new_n1085));
  NAND4_X1  g0885(.A1(new_n707), .A2(G330), .A3(new_n798), .A4(new_n1085), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT113), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(new_n872), .B(KEYINPUT112), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n867), .A2(new_n848), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(new_n874), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1088), .B1(new_n1090), .B2(new_n879), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n712), .A2(new_n653), .A3(new_n798), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n884), .B1(new_n1092), .B2(new_n887), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1087), .B1(new_n1091), .B2(new_n1094), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1088), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1096), .B1(new_n860), .B2(new_n868), .ZN(new_n1097));
  NOR3_X1   g0897(.A1(new_n1097), .A2(KEYINPUT113), .A3(new_n1093), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n1084), .B(new_n1086), .C1(new_n1095), .C2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1091), .A2(new_n1094), .A3(new_n1087), .ZN(new_n1100));
  OAI21_X1  g0900(.A(KEYINPUT113), .B1(new_n1097), .B2(new_n1093), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n1100), .A2(new_n1101), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n900), .A2(G330), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(new_n902), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1099), .B1(new_n1102), .B2(new_n1105), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n884), .B1(new_n1103), .B2(new_n901), .ZN(new_n1107));
  NAND4_X1  g0907(.A1(new_n1086), .A2(new_n1107), .A3(new_n887), .A4(new_n1092), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n707), .A2(G330), .A3(new_n798), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n1109), .A2(new_n884), .B1(new_n902), .B2(new_n1104), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1108), .B1(new_n1110), .B2(new_n1082), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1104), .A2(new_n438), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n629), .A2(new_n893), .A3(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1111), .A2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n677), .B1(new_n1106), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(KEYINPUT114), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1106), .A2(new_n1115), .ZN(new_n1119));
  OAI211_X1 g0919(.A(KEYINPUT114), .B(new_n677), .C1(new_n1106), .C2(new_n1115), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1118), .A2(new_n1119), .A3(new_n1120), .ZN(new_n1121));
  OR2_X1    g0921(.A1(new_n1106), .A2(new_n719), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1081), .A2(new_n722), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n740), .A2(G150), .ZN(new_n1124));
  XOR2_X1   g0924(.A(KEYINPUT115), .B(KEYINPUT53), .Z(new_n1125));
  XNOR2_X1  g0925(.A(new_n1124), .B(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(G128), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n1127), .A2(new_n775), .B1(new_n752), .B2(new_n745), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1128), .B1(new_n827), .B2(new_n1003), .ZN(new_n1129));
  INV_X1    g0929(.A(G125), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n259), .B1(new_n744), .B2(new_n1130), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(KEYINPUT54), .B(G143), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n757), .A2(new_n812), .B1(new_n755), .B2(new_n1132), .ZN(new_n1133));
  AOI211_X1 g0933(.A(new_n1131), .B(new_n1133), .C1(G50), .C2(new_n738), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1126), .A2(new_n1129), .A3(new_n1134), .ZN(new_n1135));
  OAI221_X1 g0935(.A(new_n257), .B1(new_n744), .B2(new_n776), .C1(new_n757), .C2(new_n577), .ZN(new_n1136));
  AOI211_X1 g0936(.A(new_n1136), .B(new_n815), .C1(G77), .C2(new_n816), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1137), .B1(new_n678), .B2(new_n764), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n806), .A2(G97), .B1(new_n749), .B2(G283), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1139), .B1(new_n224), .B2(new_n759), .ZN(new_n1140));
  XNOR2_X1  g0940(.A(new_n1140), .B(KEYINPUT116), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1135), .B1(new_n1138), .B2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n783), .B1(new_n1142), .B2(KEYINPUT117), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1143), .B1(KEYINPUT117), .B2(new_n1142), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n783), .A2(new_n285), .A3(new_n723), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n1123), .A2(new_n721), .A3(new_n1144), .A4(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1122), .A2(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1121), .A2(new_n1148), .ZN(G378));
  NAND2_X1  g0949(.A1(new_n299), .A2(new_n845), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(new_n320), .B(new_n1150), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n1151), .B(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1154), .A2(KEYINPUT120), .ZN(new_n1155));
  AND3_X1   g0955(.A1(new_n891), .A2(new_n909), .A3(G330), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n790), .B1(new_n904), .B2(new_n908), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n1157), .A2(new_n891), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1155), .B1(new_n1156), .B2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n909), .A2(G330), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n891), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  XOR2_X1   g0962(.A(new_n320), .B(new_n1150), .Z(new_n1163));
  NAND2_X1  g0963(.A1(new_n1163), .A2(new_n1153), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1165));
  AND3_X1   g0965(.A1(new_n1164), .A2(KEYINPUT120), .A3(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1157), .A2(new_n891), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1162), .A2(new_n1166), .A3(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1159), .A2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1154), .A2(new_n722), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n721), .B1(G50), .B2(new_n802), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n259), .A2(G41), .ZN(new_n1172));
  INV_X1    g0972(.A(G283), .ZN(new_n1173));
  OAI221_X1 g0973(.A(new_n1172), .B1(new_n1173), .B2(new_n744), .C1(new_n224), .C2(new_n757), .ZN(new_n1174));
  AOI211_X1 g0974(.A(new_n998), .B(new_n1174), .C1(G116), .C2(new_n749), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n759), .A2(new_n508), .B1(new_n755), .B2(new_n416), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(new_n1176), .B(KEYINPUT118), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n738), .A2(G58), .ZN(new_n1178));
  NAND4_X1  g0978(.A1(new_n1175), .A2(new_n1023), .A3(new_n1177), .A4(new_n1178), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(new_n1179), .B(KEYINPUT119), .ZN(new_n1180));
  OR2_X1    g0980(.A1(new_n1180), .A2(KEYINPUT58), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1180), .A2(KEYINPUT58), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(G33), .A2(G41), .ZN(new_n1183));
  NOR3_X1   g0983(.A1(new_n1172), .A2(G50), .A3(new_n1183), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n757), .A2(new_n1127), .B1(new_n755), .B2(new_n808), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(G132), .B2(new_n827), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n816), .A2(G150), .B1(G125), .B2(new_n749), .ZN(new_n1187));
  OAI211_X1 g0987(.A(new_n1186), .B(new_n1187), .C1(new_n741), .C2(new_n1132), .ZN(new_n1188));
  OR2_X1    g0988(.A1(new_n1188), .A2(KEYINPUT59), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n779), .A2(G124), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n1183), .B(new_n1190), .C1(new_n814), .C2(new_n745), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1191), .B1(new_n1188), .B2(KEYINPUT59), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1184), .B1(new_n1189), .B2(new_n1192), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1181), .A2(new_n1182), .A3(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1171), .B1(new_n1194), .B2(new_n725), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n1169), .A2(new_n720), .B1(new_n1170), .B2(new_n1195), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1114), .B1(new_n1106), .B2(new_n1115), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1169), .A2(new_n1197), .A3(KEYINPUT57), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1198), .A2(new_n677), .ZN(new_n1199));
  AOI21_X1  g0999(.A(KEYINPUT57), .B1(new_n1169), .B2(new_n1197), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1196), .B1(new_n1199), .B2(new_n1200), .ZN(G375));
  OAI211_X1 g1001(.A(new_n1113), .B(new_n1108), .C1(new_n1082), .C2(new_n1110), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n951), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1115), .A2(new_n1202), .A3(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n884), .A2(new_n722), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n721), .B1(G68), .B2(new_n802), .ZN(new_n1206));
  OAI221_X1 g1006(.A(new_n259), .B1(new_n755), .B2(new_n287), .C1(new_n1127), .C2(new_n744), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1207), .B1(G50), .B2(new_n816), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n1208), .B(new_n1178), .C1(new_n764), .C2(new_n745), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT123), .ZN(new_n1210));
  OR2_X1    g1010(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n757), .A2(new_n1002), .B1(new_n759), .B2(new_n1132), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(G132), .B2(new_n749), .ZN(new_n1214));
  XNOR2_X1  g1014(.A(new_n1214), .B(KEYINPUT122), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1211), .A2(new_n1212), .A3(new_n1215), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n759), .A2(new_n577), .ZN(new_n1217));
  AOI211_X1 g1017(.A(new_n1217), .B(new_n1027), .C1(G294), .C2(new_n749), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n257), .B1(new_n755), .B2(new_n224), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n757), .A2(new_n1173), .B1(new_n744), .B2(new_n765), .ZN(new_n1220));
  AOI211_X1 g1020(.A(new_n1219), .B(new_n1220), .C1(G77), .C2(new_n738), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n1218), .B(new_n1221), .C1(new_n764), .C2(new_n508), .ZN(new_n1222));
  XNOR2_X1  g1022(.A(new_n1222), .B(KEYINPUT121), .ZN(new_n1223));
  AOI21_X1  g1023(.A(KEYINPUT124), .B1(new_n1216), .B2(new_n1223), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n1224), .A2(new_n783), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1216), .A2(KEYINPUT124), .A3(new_n1223), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1206), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n1111), .A2(new_n720), .B1(new_n1205), .B2(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1204), .A2(new_n1228), .ZN(G381));
  INV_X1    g1029(.A(G375), .ZN(new_n1230));
  AND2_X1   g1030(.A1(new_n1120), .A2(new_n1119), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1147), .B1(new_n1231), .B2(new_n1118), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(G393), .A2(G396), .ZN(new_n1233));
  INV_X1    g1033(.A(G384), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  NOR4_X1   g1035(.A1(G387), .A2(new_n1235), .A3(G390), .A4(G381), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1230), .A2(new_n1232), .A3(new_n1236), .ZN(G407));
  NAND2_X1  g1037(.A1(new_n651), .A2(G213), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1230), .A2(new_n1232), .A3(new_n1239), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(G407), .A2(new_n1240), .A3(G213), .ZN(G409));
  NAND3_X1  g1041(.A1(new_n1169), .A2(new_n1197), .A3(new_n1203), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1196), .A2(new_n1242), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1243), .A2(new_n1121), .A3(new_n1148), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1244), .B1(G375), .B2(new_n1232), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1115), .A2(KEYINPUT60), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(new_n1202), .ZN(new_n1247));
  OR2_X1    g1047(.A1(new_n1110), .A2(new_n1082), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1248), .A2(KEYINPUT60), .A3(new_n1113), .A4(new_n1108), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1247), .A2(new_n677), .A3(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(G384), .B1(new_n1250), .B2(new_n1228), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1202), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT60), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1253), .B1(new_n1111), .B2(new_n1114), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1252), .A2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1249), .A2(new_n677), .ZN(new_n1256));
  OAI211_X1 g1056(.A(G384), .B(new_n1228), .C1(new_n1255), .C2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1251), .A2(new_n1258), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1245), .A2(new_n1238), .A3(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(KEYINPUT62), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1245), .A2(new_n1238), .ZN(new_n1262));
  INV_X1    g1062(.A(G2897), .ZN(new_n1263));
  OAI22_X1  g1063(.A1(new_n1251), .A2(new_n1258), .B1(new_n1263), .B2(new_n1238), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1228), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(new_n1234), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1238), .A2(new_n1263), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1266), .A2(new_n1257), .A3(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1264), .A2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1262), .A2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT61), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT62), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1245), .A2(new_n1272), .A3(new_n1238), .A4(new_n1259), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1261), .A2(new_n1270), .A3(new_n1271), .A4(new_n1273), .ZN(new_n1274));
  AND3_X1   g1074(.A1(new_n981), .A2(G390), .A3(new_n1010), .ZN(new_n1275));
  AOI21_X1  g1075(.A(G390), .B1(new_n981), .B2(new_n1010), .ZN(new_n1276));
  OAI21_X1  g1076(.A(KEYINPUT127), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n792), .B1(new_n1014), .B2(new_n1046), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1233), .A2(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1277), .A2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1279), .ZN(new_n1281));
  OAI211_X1 g1081(.A(KEYINPUT127), .B(new_n1281), .C1(new_n1275), .C2(new_n1276), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1280), .A2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1274), .A2(new_n1283), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1280), .A2(new_n1271), .A3(new_n1282), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT63), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1285), .B1(new_n1286), .B2(new_n1260), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1169), .A2(new_n1197), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT57), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1290), .A2(new_n677), .A3(new_n1198), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1291), .A2(G378), .A3(new_n1196), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1239), .B1(new_n1292), .B2(new_n1244), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1293), .A2(KEYINPUT63), .A3(new_n1259), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(new_n1262), .A2(KEYINPUT125), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT126), .ZN(new_n1296));
  AND3_X1   g1096(.A1(new_n1266), .A2(new_n1257), .A3(new_n1267), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1267), .B1(new_n1266), .B2(new_n1257), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1296), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1264), .A2(KEYINPUT126), .A3(new_n1268), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT125), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1301), .B1(new_n1302), .B2(new_n1293), .ZN(new_n1303));
  OAI211_X1 g1103(.A(new_n1287), .B(new_n1294), .C1(new_n1295), .C2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1284), .A2(new_n1304), .ZN(G405));
  NAND2_X1  g1105(.A1(G375), .A2(new_n1232), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1283), .A2(new_n1292), .A3(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1306), .A2(new_n1292), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1308), .A2(new_n1280), .A3(new_n1282), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1307), .A2(new_n1309), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1310), .B1(new_n1251), .B2(new_n1258), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1307), .A2(new_n1259), .A3(new_n1309), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1311), .A2(new_n1312), .ZN(G402));
endmodule


