//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 1 0 0 0 1 0 0 0 1 1 1 1 1 0 0 0 0 1 1 0 1 1 1 0 0 0 0 1 0 1 0 1 0 1 1 0 0 1 0 1 0 0 1 1 0 0 0 1 0 1 0 0 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:39 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n590, new_n591, new_n592, new_n593, new_n594, new_n595,
    new_n596, new_n597, new_n598, new_n599, new_n601, new_n602, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n632, new_n633,
    new_n634, new_n636, new_n637, new_n638, new_n639, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n663, new_n664, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n691,
    new_n692, new_n693, new_n694, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n748, new_n749, new_n750,
    new_n752, new_n753, new_n754, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n827, new_n828, new_n830, new_n831, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n841, new_n842,
    new_n844, new_n845, new_n846, new_n847, new_n849, new_n850, new_n851,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n898, new_n899;
  XOR2_X1   g000(.A(G211gat), .B(G218gat), .Z(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  OR2_X1    g002(.A1(new_n203), .A2(KEYINPUT70), .ZN(new_n204));
  XOR2_X1   g003(.A(G197gat), .B(G204gat), .Z(new_n205));
  AOI21_X1  g004(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(new_n204), .B(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  XOR2_X1   g009(.A(KEYINPUT72), .B(G155gat), .Z(new_n211));
  INV_X1    g010(.A(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G162gat), .ZN(new_n213));
  OAI21_X1  g012(.A(KEYINPUT2), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(G155gat), .B(G162gat), .ZN(new_n215));
  XOR2_X1   g014(.A(G141gat), .B(G148gat), .Z(new_n216));
  NAND3_X1  g015(.A1(new_n214), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  XNOR2_X1  g016(.A(KEYINPUT71), .B(KEYINPUT2), .ZN(new_n218));
  AND2_X1   g017(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  OR2_X1    g018(.A1(new_n219), .A2(new_n215), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n217), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT3), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT29), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n210), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  AOI21_X1  g025(.A(KEYINPUT29), .B1(new_n208), .B2(new_n203), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n227), .B1(new_n203), .B2(new_n208), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n222), .B1(new_n223), .B2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(G228gat), .ZN(new_n230));
  INV_X1    g029(.A(G233gat), .ZN(new_n231));
  OAI22_X1  g030(.A1(new_n226), .A2(new_n229), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n232), .B(KEYINPUT77), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n223), .B1(new_n209), .B2(KEYINPUT29), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(new_n221), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT78), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n226), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n230), .A2(new_n231), .ZN(new_n238));
  OAI211_X1 g037(.A(new_n237), .B(new_n238), .C1(new_n236), .C2(new_n235), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n233), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(G22gat), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(G78gat), .B(G106gat), .ZN(new_n243));
  XNOR2_X1  g042(.A(KEYINPUT31), .B(G50gat), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n243), .B(new_n244), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n241), .B1(new_n233), .B2(new_n239), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n245), .B1(new_n246), .B2(KEYINPUT79), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n242), .B(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT25), .ZN(new_n250));
  NOR2_X1   g049(.A1(G169gat), .A2(G176gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(KEYINPUT23), .ZN(new_n252));
  NAND2_X1  g051(.A1(G169gat), .A2(G176gat), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT23), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n254), .B1(G169gat), .B2(G176gat), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n252), .A2(new_n253), .A3(new_n255), .ZN(new_n256));
  AOI21_X1  g055(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n257), .A2(KEYINPUT66), .ZN(new_n258));
  NAND3_X1  g057(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n259), .B1(G183gat), .B2(G190gat), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n257), .A2(KEYINPUT66), .ZN(new_n262));
  AOI211_X1 g061(.A(new_n250), .B(new_n256), .C1(new_n261), .C2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT64), .ZN(new_n264));
  OAI22_X1  g063(.A1(new_n256), .A2(new_n264), .B1(new_n260), .B2(new_n257), .ZN(new_n265));
  AND2_X1   g064(.A1(new_n256), .A2(new_n264), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n250), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT65), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n263), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n269), .B1(new_n268), .B2(new_n267), .ZN(new_n270));
  XNOR2_X1  g069(.A(KEYINPUT27), .B(G183gat), .ZN(new_n271));
  INV_X1    g070(.A(G190gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  XOR2_X1   g072(.A(new_n273), .B(KEYINPUT28), .Z(new_n274));
  AOI22_X1  g073(.A1(new_n251), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n275));
  INV_X1    g074(.A(new_n253), .ZN(new_n276));
  OR2_X1    g075(.A1(new_n251), .A2(KEYINPUT26), .ZN(new_n277));
  OAI211_X1 g076(.A(new_n274), .B(new_n275), .C1(new_n276), .C2(new_n277), .ZN(new_n278));
  AND2_X1   g077(.A1(new_n270), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(G226gat), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n279), .B1(new_n280), .B2(new_n231), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n280), .A2(new_n231), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n282), .A2(KEYINPUT29), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n281), .B1(new_n279), .B2(new_n283), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n284), .B(new_n210), .ZN(new_n285));
  XNOR2_X1  g084(.A(G8gat), .B(G36gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(G64gat), .B(G92gat), .ZN(new_n287));
  XOR2_X1   g086(.A(new_n286), .B(new_n287), .Z(new_n288));
  NAND2_X1  g087(.A1(new_n285), .A2(new_n288), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n284), .B(new_n209), .ZN(new_n290));
  INV_X1    g089(.A(new_n288), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n289), .A2(new_n292), .A3(KEYINPUT30), .ZN(new_n293));
  OR3_X1    g092(.A1(new_n290), .A2(KEYINPUT30), .A3(new_n291), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  XNOR2_X1  g095(.A(G1gat), .B(G29gat), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n297), .B(KEYINPUT0), .ZN(new_n298));
  XOR2_X1   g097(.A(G57gat), .B(G85gat), .Z(new_n299));
  XNOR2_X1  g098(.A(new_n298), .B(new_n299), .ZN(new_n300));
  XNOR2_X1  g099(.A(G113gat), .B(G120gat), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n301), .A2(KEYINPUT1), .ZN(new_n302));
  XNOR2_X1  g101(.A(G127gat), .B(G134gat), .ZN(new_n303));
  XNOR2_X1  g102(.A(new_n302), .B(new_n303), .ZN(new_n304));
  OR3_X1    g103(.A1(new_n221), .A2(KEYINPUT4), .A3(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT74), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  OAI21_X1  g106(.A(KEYINPUT4), .B1(new_n221), .B2(new_n304), .ZN(new_n308));
  XNOR2_X1  g107(.A(new_n307), .B(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n221), .A2(KEYINPUT3), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n224), .A2(new_n304), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(G225gat), .A2(G233gat), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n300), .B1(new_n315), .B2(KEYINPUT39), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n221), .B(new_n304), .ZN(new_n317));
  OR2_X1    g116(.A1(new_n317), .A2(new_n314), .ZN(new_n318));
  AND2_X1   g117(.A1(new_n318), .A2(KEYINPUT39), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n316), .B1(new_n315), .B2(new_n319), .ZN(new_n320));
  OR2_X1    g119(.A1(new_n320), .A2(KEYINPUT40), .ZN(new_n321));
  AND2_X1   g120(.A1(new_n311), .A2(new_n313), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n305), .A2(KEYINPUT73), .A3(new_n308), .ZN(new_n323));
  OAI211_X1 g122(.A(new_n322), .B(new_n323), .C1(KEYINPUT73), .C2(new_n308), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT5), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n325), .B1(new_n317), .B2(new_n314), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n309), .A2(new_n325), .A3(new_n322), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n300), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n329), .B1(new_n320), .B2(KEYINPUT40), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n296), .A2(new_n321), .A3(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT38), .ZN(new_n332));
  OR2_X1    g131(.A1(new_n290), .A2(KEYINPUT37), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n288), .B1(new_n290), .B2(KEYINPUT37), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n332), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n329), .ZN(new_n336));
  XNOR2_X1  g135(.A(KEYINPUT75), .B(KEYINPUT6), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n327), .A2(new_n328), .A3(new_n300), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(new_n337), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n338), .B1(new_n336), .B2(new_n341), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n333), .A2(new_n332), .A3(new_n334), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n342), .A2(new_n289), .A3(new_n343), .ZN(new_n344));
  OAI211_X1 g143(.A(new_n249), .B(new_n331), .C1(new_n335), .C2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n341), .A2(KEYINPUT76), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT76), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n329), .B1(new_n340), .B2(new_n347), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n338), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n248), .B1(new_n296), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n345), .A2(new_n350), .ZN(new_n351));
  XNOR2_X1  g150(.A(G15gat), .B(G43gat), .ZN(new_n352));
  XNOR2_X1  g151(.A(G71gat), .B(G99gat), .ZN(new_n353));
  XNOR2_X1  g152(.A(new_n352), .B(new_n353), .ZN(new_n354));
  XNOR2_X1  g153(.A(new_n279), .B(new_n304), .ZN(new_n355));
  NAND2_X1  g154(.A1(G227gat), .A2(G233gat), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n354), .B1(new_n358), .B2(KEYINPUT32), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT67), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT33), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n360), .B1(new_n358), .B2(new_n361), .ZN(new_n362));
  NOR3_X1   g161(.A1(new_n357), .A2(KEYINPUT67), .A3(KEYINPUT33), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n359), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  OAI211_X1 g163(.A(new_n358), .B(KEYINPUT32), .C1(new_n361), .C2(new_n354), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT68), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n355), .A2(new_n356), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT34), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT69), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n369), .B1(new_n356), .B2(new_n370), .ZN(new_n371));
  XNOR2_X1  g170(.A(new_n368), .B(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n366), .B1(new_n367), .B2(new_n373), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n364), .A2(KEYINPUT68), .A3(new_n372), .A4(new_n365), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n374), .A2(KEYINPUT36), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n366), .A2(new_n372), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT36), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n364), .A2(new_n373), .A3(new_n365), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n377), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n376), .A2(new_n380), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n351), .A2(new_n381), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n248), .B1(new_n374), .B2(new_n375), .ZN(new_n383));
  INV_X1    g182(.A(new_n349), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n383), .A2(new_n384), .A3(new_n295), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n377), .A2(new_n379), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n386), .A2(new_n248), .ZN(new_n387));
  NOR3_X1   g186(.A1(new_n296), .A2(KEYINPUT35), .A3(new_n342), .ZN(new_n388));
  AOI22_X1  g187(.A1(new_n385), .A2(KEYINPUT35), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n382), .A2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT14), .ZN(new_n391));
  INV_X1    g190(.A(G29gat), .ZN(new_n392));
  INV_X1    g191(.A(G36gat), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n391), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT81), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NOR3_X1   g195(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(KEYINPUT81), .ZN(new_n398));
  OAI21_X1  g197(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n396), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  XNOR2_X1  g199(.A(G43gat), .B(G50gat), .ZN(new_n401));
  AOI22_X1  g200(.A1(new_n401), .A2(KEYINPUT15), .B1(G29gat), .B2(G36gat), .ZN(new_n402));
  AOI21_X1  g201(.A(KEYINPUT15), .B1(G43gat), .B2(G50gat), .ZN(new_n403));
  XNOR2_X1  g202(.A(KEYINPUT80), .B(G43gat), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n403), .B1(new_n404), .B2(G50gat), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n400), .A2(new_n402), .A3(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n399), .ZN(new_n407));
  OAI22_X1  g206(.A1(new_n407), .A2(new_n397), .B1(new_n392), .B2(new_n393), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n408), .A2(KEYINPUT15), .A3(new_n401), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n406), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n241), .A2(G15gat), .ZN(new_n411));
  INV_X1    g210(.A(G15gat), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(G22gat), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT16), .ZN(new_n414));
  OAI211_X1 g213(.A(new_n411), .B(new_n413), .C1(new_n414), .C2(G1gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(G15gat), .B(G22gat), .ZN(new_n416));
  OAI221_X1 g215(.A(new_n415), .B1(KEYINPUT82), .B2(G8gat), .C1(G1gat), .C2(new_n416), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n415), .B1(G1gat), .B2(new_n416), .ZN(new_n418));
  INV_X1    g217(.A(G8gat), .ZN(new_n419));
  OAI21_X1  g218(.A(KEYINPUT82), .B1(new_n416), .B2(G1gat), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n418), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n410), .A2(new_n417), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(G229gat), .A2(G233gat), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n410), .A2(KEYINPUT17), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT17), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n406), .A2(new_n427), .A3(new_n409), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n421), .A2(new_n417), .ZN(new_n430));
  AOI21_X1  g229(.A(KEYINPUT83), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  AND3_X1   g230(.A1(new_n406), .A2(new_n427), .A3(new_n409), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n427), .B1(new_n406), .B2(new_n409), .ZN(new_n433));
  OAI211_X1 g232(.A(KEYINPUT83), .B(new_n430), .C1(new_n432), .C2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  OAI211_X1 g234(.A(KEYINPUT18), .B(new_n425), .C1(new_n431), .C2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT85), .ZN(new_n437));
  XNOR2_X1  g236(.A(new_n430), .B(new_n410), .ZN(new_n438));
  XOR2_X1   g237(.A(new_n423), .B(KEYINPUT13), .Z(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n437), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(new_n422), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n410), .B1(new_n417), .B2(new_n421), .ZN(new_n443));
  OAI211_X1 g242(.A(KEYINPUT85), .B(new_n439), .C1(new_n442), .C2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n441), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n436), .A2(new_n445), .A3(KEYINPUT84), .ZN(new_n446));
  XNOR2_X1  g245(.A(G113gat), .B(G141gat), .ZN(new_n447));
  XNOR2_X1  g246(.A(new_n447), .B(G197gat), .ZN(new_n448));
  XOR2_X1   g247(.A(KEYINPUT11), .B(G169gat), .Z(new_n449));
  XNOR2_X1  g248(.A(new_n448), .B(new_n449), .ZN(new_n450));
  XOR2_X1   g249(.A(new_n450), .B(KEYINPUT12), .Z(new_n451));
  NAND2_X1  g250(.A1(new_n436), .A2(new_n445), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n430), .B1(new_n432), .B2(new_n433), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT83), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n424), .B1(new_n455), .B2(new_n434), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n456), .A2(KEYINPUT18), .ZN(new_n457));
  OAI211_X1 g256(.A(new_n446), .B(new_n451), .C1(new_n452), .C2(new_n457), .ZN(new_n458));
  OR2_X1    g257(.A1(new_n456), .A2(KEYINPUT18), .ZN(new_n459));
  AOI22_X1  g258(.A1(new_n456), .A2(KEYINPUT18), .B1(new_n441), .B2(new_n444), .ZN(new_n460));
  INV_X1    g259(.A(new_n451), .ZN(new_n461));
  OAI211_X1 g260(.A(new_n459), .B(new_n460), .C1(KEYINPUT84), .C2(new_n461), .ZN(new_n462));
  AND2_X1   g261(.A1(new_n458), .A2(new_n462), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n390), .A2(new_n463), .ZN(new_n464));
  XNOR2_X1  g263(.A(G190gat), .B(G218gat), .ZN(new_n465));
  XNOR2_X1  g264(.A(new_n465), .B(KEYINPUT90), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(G85gat), .ZN(new_n468));
  INV_X1    g267(.A(G92gat), .ZN(new_n469));
  OAI21_X1  g268(.A(KEYINPUT7), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT7), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n471), .A2(G85gat), .A3(G92gat), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  XOR2_X1   g272(.A(G99gat), .B(G106gat), .Z(new_n474));
  NAND2_X1  g273(.A1(G99gat), .A2(G106gat), .ZN(new_n475));
  AOI22_X1  g274(.A1(KEYINPUT8), .A2(new_n475), .B1(new_n468), .B2(new_n469), .ZN(new_n476));
  AND3_X1   g275(.A1(new_n473), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n474), .B1(new_n473), .B2(new_n476), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n429), .A2(new_n479), .ZN(new_n480));
  OR2_X1    g279(.A1(new_n477), .A2(new_n478), .ZN(new_n481));
  AND2_X1   g280(.A1(G232gat), .A2(G233gat), .ZN(new_n482));
  AOI22_X1  g281(.A1(new_n481), .A2(new_n410), .B1(KEYINPUT41), .B2(new_n482), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n467), .B1(new_n480), .B2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(new_n484), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n482), .A2(KEYINPUT41), .ZN(new_n486));
  XNOR2_X1  g285(.A(G134gat), .B(G162gat), .ZN(new_n487));
  XOR2_X1   g286(.A(new_n486), .B(new_n487), .Z(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n480), .A2(new_n467), .A3(new_n483), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n485), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT91), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n490), .B1(new_n484), .B2(new_n493), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n480), .A2(KEYINPUT91), .A3(new_n467), .A4(new_n483), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(new_n488), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT92), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n496), .A2(KEYINPUT92), .A3(new_n488), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n492), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(G71gat), .A2(G78gat), .ZN(new_n502));
  OR2_X1    g301(.A1(G71gat), .A2(G78gat), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT9), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT86), .ZN(new_n506));
  INV_X1    g305(.A(G57gat), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(KEYINPUT86), .A2(G57gat), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n508), .A2(KEYINPUT87), .A3(G64gat), .A4(new_n509), .ZN(new_n510));
  OAI21_X1  g309(.A(KEYINPUT88), .B1(new_n507), .B2(G64gat), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT88), .ZN(new_n512));
  INV_X1    g311(.A(G64gat), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n512), .A2(new_n513), .A3(G57gat), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n510), .A2(new_n511), .A3(new_n514), .ZN(new_n515));
  AND2_X1   g314(.A1(KEYINPUT86), .A2(G57gat), .ZN(new_n516));
  NOR2_X1   g315(.A1(KEYINPUT86), .A2(G57gat), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(KEYINPUT87), .B1(new_n518), .B2(G64gat), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n505), .B1(new_n515), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n503), .A2(new_n502), .ZN(new_n521));
  XOR2_X1   g320(.A(G57gat), .B(G64gat), .Z(new_n522));
  AOI21_X1  g321(.A(new_n521), .B1(new_n522), .B2(KEYINPUT9), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n520), .A2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT21), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n430), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  XOR2_X1   g326(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n528));
  XNOR2_X1  g327(.A(new_n527), .B(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n525), .A2(new_n526), .ZN(new_n531));
  NAND2_X1  g330(.A1(G231gat), .A2(G233gat), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n531), .B(new_n532), .ZN(new_n533));
  XNOR2_X1  g332(.A(G127gat), .B(G155gat), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n534), .B(KEYINPUT89), .ZN(new_n535));
  AND2_X1   g334(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n533), .A2(new_n535), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  XOR2_X1   g337(.A(G183gat), .B(G211gat), .Z(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n533), .B(new_n535), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n542), .A2(new_n539), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n530), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n538), .A2(new_n540), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n542), .A2(new_n539), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n545), .A2(new_n529), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n501), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(G230gat), .A2(G233gat), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n473), .A2(new_n476), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(KEYINPUT93), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n520), .A2(new_n524), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n553), .A2(new_n481), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n508), .A2(G64gat), .A3(new_n509), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT87), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  AND2_X1   g356(.A1(new_n511), .A2(new_n514), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n557), .A2(new_n510), .A3(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n523), .B1(new_n559), .B2(new_n505), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n560), .A2(new_n479), .A3(new_n552), .ZN(new_n561));
  AOI21_X1  g360(.A(KEYINPUT10), .B1(new_n554), .B2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT10), .ZN(new_n563));
  NOR3_X1   g362(.A1(new_n525), .A2(new_n563), .A3(new_n479), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n550), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n550), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n554), .A2(new_n566), .A3(new_n561), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(G120gat), .B(G148gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n569), .B(KEYINPUT94), .ZN(new_n570));
  XNOR2_X1  g369(.A(G176gat), .B(G204gat), .ZN(new_n571));
  XOR2_X1   g370(.A(new_n570), .B(new_n571), .Z(new_n572));
  OR2_X1    g371(.A1(new_n568), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n568), .A2(new_n572), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n549), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n464), .A2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n578), .A2(new_n349), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n579), .B(G1gat), .ZN(G1324gat));
  OAI21_X1  g379(.A(G8gat), .B1(new_n577), .B2(new_n295), .ZN(new_n581));
  OR2_X1    g380(.A1(new_n581), .A2(KEYINPUT95), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(KEYINPUT95), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n577), .A2(new_n295), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT42), .ZN(new_n585));
  XOR2_X1   g384(.A(KEYINPUT16), .B(G8gat), .Z(new_n586));
  AND3_X1   g385(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n585), .B1(new_n584), .B2(new_n586), .ZN(new_n588));
  OAI211_X1 g387(.A(new_n582), .B(new_n583), .C1(new_n587), .C2(new_n588), .ZN(G1325gat));
  OR3_X1    g388(.A1(new_n577), .A2(G15gat), .A3(new_n386), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n381), .A2(KEYINPUT96), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT96), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n376), .A2(new_n380), .A3(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g395(.A(G15gat), .B1(new_n577), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n590), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT97), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(G1326gat));
  NOR2_X1   g399(.A1(new_n577), .A2(new_n249), .ZN(new_n601));
  XOR2_X1   g400(.A(KEYINPUT43), .B(G22gat), .Z(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(G1327gat));
  INV_X1    g402(.A(KEYINPUT100), .ZN(new_n604));
  AOI21_X1  g403(.A(KEYINPUT92), .B1(new_n496), .B2(new_n488), .ZN(new_n605));
  AOI211_X1 g404(.A(new_n498), .B(new_n489), .C1(new_n494), .C2(new_n495), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n491), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n607), .B1(new_n382), .B2(new_n389), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n604), .B1(new_n608), .B2(KEYINPUT44), .ZN(new_n609));
  INV_X1    g408(.A(new_n389), .ZN(new_n610));
  NAND4_X1  g409(.A1(new_n591), .A2(new_n350), .A3(new_n345), .A4(new_n594), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT44), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n612), .A2(new_n613), .A3(new_n607), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n609), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n608), .A2(new_n604), .A3(KEYINPUT44), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n548), .B(KEYINPUT99), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  AND2_X1   g417(.A1(new_n463), .A2(KEYINPUT98), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n463), .A2(KEYINPUT98), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NOR3_X1   g421(.A1(new_n618), .A2(new_n622), .A3(new_n575), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n615), .A2(new_n616), .A3(new_n623), .ZN(new_n624));
  OAI21_X1  g423(.A(G29gat), .B1(new_n624), .B2(new_n384), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n458), .A2(new_n462), .ZN(new_n626));
  NOR3_X1   g425(.A1(new_n501), .A2(new_n548), .A3(new_n575), .ZN(new_n627));
  OAI211_X1 g426(.A(new_n626), .B(new_n627), .C1(new_n382), .C2(new_n389), .ZN(new_n628));
  NOR3_X1   g427(.A1(new_n628), .A2(G29gat), .A3(new_n384), .ZN(new_n629));
  XOR2_X1   g428(.A(new_n629), .B(KEYINPUT45), .Z(new_n630));
  NAND2_X1  g429(.A1(new_n625), .A2(new_n630), .ZN(G1328gat));
  OAI21_X1  g430(.A(G36gat), .B1(new_n624), .B2(new_n295), .ZN(new_n632));
  NOR3_X1   g431(.A1(new_n628), .A2(G36gat), .A3(new_n295), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(KEYINPUT46), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n632), .A2(new_n634), .ZN(G1329gat));
  INV_X1    g434(.A(new_n596), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n636), .A2(new_n404), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n628), .A2(new_n386), .ZN(new_n638));
  OAI22_X1  g437(.A1(new_n624), .A2(new_n637), .B1(new_n404), .B2(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g439(.A(KEYINPUT101), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n249), .B1(new_n628), .B2(new_n641), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n642), .B1(new_n641), .B2(new_n628), .ZN(new_n643));
  INV_X1    g442(.A(G50gat), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n248), .A2(G50gat), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n645), .B1(new_n624), .B2(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(KEYINPUT48), .ZN(G1331gat));
  NOR2_X1   g447(.A1(new_n621), .A2(new_n549), .ZN(new_n649));
  AND3_X1   g448(.A1(new_n612), .A2(new_n575), .A3(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(new_n349), .ZN(new_n651));
  XOR2_X1   g450(.A(new_n651), .B(new_n518), .Z(G1332gat));
  AOI21_X1  g451(.A(new_n295), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(KEYINPUT102), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n650), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(KEYINPUT103), .ZN(new_n656));
  OR2_X1    g455(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n656), .B(new_n657), .ZN(G1333gat));
  NAND2_X1  g457(.A1(new_n650), .A2(new_n636), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n386), .A2(G71gat), .ZN(new_n660));
  AOI22_X1  g459(.A1(new_n659), .A2(G71gat), .B1(new_n650), .B2(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g461(.A1(new_n650), .A2(new_n248), .ZN(new_n663));
  XOR2_X1   g462(.A(KEYINPUT104), .B(G78gat), .Z(new_n664));
  XNOR2_X1  g463(.A(new_n663), .B(new_n664), .ZN(G1335gat));
  INV_X1    g464(.A(new_n575), .ZN(new_n666));
  NOR3_X1   g465(.A1(new_n384), .A2(G85gat), .A3(new_n666), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n621), .A2(new_n548), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n612), .A2(new_n607), .A3(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT51), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND4_X1  g470(.A1(new_n612), .A2(KEYINPUT51), .A3(new_n607), .A4(new_n668), .ZN(new_n672));
  AND3_X1   g471(.A1(new_n671), .A2(KEYINPUT105), .A3(new_n672), .ZN(new_n673));
  AOI21_X1  g472(.A(KEYINPUT105), .B1(new_n671), .B2(new_n672), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n667), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n668), .A2(new_n575), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n615), .A2(new_n616), .A3(new_n677), .ZN(new_n678));
  OAI21_X1  g477(.A(G85gat), .B1(new_n678), .B2(new_n384), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n675), .A2(new_n679), .ZN(G1336gat));
  NAND4_X1  g479(.A1(new_n615), .A2(new_n296), .A3(new_n616), .A4(new_n677), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n681), .A2(G92gat), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n671), .A2(new_n672), .ZN(new_n683));
  NOR3_X1   g482(.A1(new_n295), .A2(G92gat), .A3(new_n666), .ZN(new_n684));
  AOI21_X1  g483(.A(KEYINPUT52), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n684), .B(KEYINPUT106), .ZN(new_n687));
  AOI22_X1  g486(.A1(new_n681), .A2(G92gat), .B1(new_n683), .B2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT52), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n686), .B1(new_n688), .B2(new_n689), .ZN(G1337gat));
  XOR2_X1   g489(.A(KEYINPUT107), .B(G99gat), .Z(new_n691));
  NOR3_X1   g490(.A1(new_n386), .A2(new_n666), .A3(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n692), .B1(new_n673), .B2(new_n674), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n691), .B1(new_n678), .B2(new_n596), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(G1338gat));
  NAND4_X1  g494(.A1(new_n615), .A2(new_n248), .A3(new_n616), .A4(new_n677), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(G106gat), .ZN(new_n697));
  NOR3_X1   g496(.A1(new_n249), .A2(G106gat), .A3(new_n666), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n683), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g498(.A(KEYINPUT108), .B(KEYINPUT53), .ZN(new_n700));
  AND3_X1   g499(.A1(new_n697), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n700), .B1(new_n697), .B2(new_n699), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n701), .A2(new_n702), .ZN(G1339gat));
  NOR2_X1   g502(.A1(new_n553), .A2(new_n481), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n479), .B1(new_n560), .B2(new_n552), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n563), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(new_n564), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n706), .A2(new_n566), .A3(new_n707), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n708), .A2(new_n565), .A3(KEYINPUT54), .ZN(new_n709));
  XNOR2_X1  g508(.A(KEYINPUT109), .B(KEYINPUT54), .ZN(new_n710));
  OAI211_X1 g509(.A(new_n550), .B(new_n710), .C1(new_n562), .C2(new_n564), .ZN(new_n711));
  NAND4_X1  g510(.A1(new_n709), .A2(KEYINPUT55), .A3(new_n572), .A4(new_n711), .ZN(new_n712));
  AND2_X1   g511(.A1(new_n712), .A2(new_n573), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT55), .ZN(new_n714));
  AND3_X1   g513(.A1(new_n708), .A2(new_n565), .A3(KEYINPUT54), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n711), .A2(new_n572), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n714), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  AND2_X1   g516(.A1(new_n713), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n621), .A2(new_n718), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n442), .B1(new_n455), .B2(new_n434), .ZN(new_n720));
  OAI21_X1  g519(.A(KEYINPUT110), .B1(new_n720), .B2(new_n423), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n438), .A2(new_n440), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NOR3_X1   g522(.A1(new_n720), .A2(KEYINPUT110), .A3(new_n423), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n450), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n460), .A2(new_n459), .A3(new_n461), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n725), .A2(new_n575), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n719), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(new_n501), .ZN(new_n729));
  AND2_X1   g528(.A1(new_n725), .A2(new_n726), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n718), .A2(new_n730), .A3(new_n607), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(KEYINPUT111), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n618), .B1(new_n729), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n649), .A2(new_n666), .ZN(new_n734));
  INV_X1    g533(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  NOR3_X1   g535(.A1(new_n736), .A2(new_n386), .A3(new_n248), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n384), .A2(new_n296), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g538(.A(G113gat), .B1(new_n739), .B2(new_n463), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(KEYINPUT112), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n736), .A2(new_n384), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n742), .A2(new_n295), .A3(new_n383), .ZN(new_n743));
  OR3_X1    g542(.A1(new_n743), .A2(G113gat), .A3(new_n622), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n741), .A2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT113), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n745), .B(new_n746), .ZN(G1340gat));
  INV_X1    g546(.A(G120gat), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n748), .B1(new_n743), .B2(new_n666), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n737), .A2(G120gat), .A3(new_n575), .A4(new_n738), .ZN(new_n750));
  AND2_X1   g549(.A1(new_n749), .A2(new_n750), .ZN(G1341gat));
  OAI21_X1  g550(.A(G127gat), .B1(new_n739), .B2(new_n617), .ZN(new_n752));
  INV_X1    g551(.A(new_n548), .ZN(new_n753));
  OR2_X1    g552(.A1(new_n753), .A2(G127gat), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n752), .B1(new_n743), .B2(new_n754), .ZN(G1342gat));
  NOR3_X1   g554(.A1(new_n743), .A2(G134gat), .A3(new_n501), .ZN(new_n756));
  INV_X1    g555(.A(new_n756), .ZN(new_n757));
  OR2_X1    g556(.A1(new_n757), .A2(KEYINPUT56), .ZN(new_n758));
  OAI21_X1  g557(.A(G134gat), .B1(new_n739), .B2(new_n501), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n757), .A2(KEYINPUT56), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n758), .A2(new_n759), .A3(new_n760), .ZN(G1343gat));
  INV_X1    g560(.A(new_n742), .ZN(new_n762));
  OR2_X1    g561(.A1(new_n762), .A2(KEYINPUT116), .ZN(new_n763));
  NOR3_X1   g562(.A1(new_n636), .A2(new_n249), .A3(new_n296), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n762), .A2(KEYINPUT116), .ZN(new_n765));
  AND3_X1   g564(.A1(new_n763), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n463), .A2(G141gat), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n596), .A2(new_n738), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT57), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n770), .B1(new_n736), .B2(new_n249), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n248), .A2(KEYINPUT57), .ZN(new_n772));
  INV_X1    g571(.A(new_n772), .ZN(new_n773));
  OAI21_X1  g572(.A(KEYINPUT114), .B1(new_n715), .B2(new_n716), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT114), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n709), .A2(new_n775), .A3(new_n572), .A4(new_n711), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n774), .A2(new_n714), .A3(new_n776), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n626), .A2(new_n777), .A3(new_n713), .ZN(new_n778));
  AND3_X1   g577(.A1(new_n778), .A2(KEYINPUT115), .A3(new_n727), .ZN(new_n779));
  AOI21_X1  g578(.A(KEYINPUT115), .B1(new_n778), .B2(new_n727), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n501), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n548), .B1(new_n732), .B2(new_n781), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n773), .B1(new_n782), .B2(new_n735), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n769), .B1(new_n771), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(new_n626), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(G141gat), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT58), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n768), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n784), .A2(new_n621), .ZN(new_n789));
  AOI22_X1  g588(.A1(new_n766), .A2(new_n767), .B1(new_n789), .B2(G141gat), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n788), .B1(new_n790), .B2(new_n787), .ZN(G1344gat));
  INV_X1    g590(.A(G148gat), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n766), .A2(new_n792), .A3(new_n575), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT59), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n736), .A2(new_n772), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n778), .A2(new_n727), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT115), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n778), .A2(KEYINPUT115), .A3(new_n727), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n607), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n713), .A2(new_n717), .ZN(new_n801));
  OAI21_X1  g600(.A(KEYINPUT118), .B1(new_n501), .B2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT118), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n718), .A2(new_n803), .A3(new_n607), .ZN(new_n804));
  AND3_X1   g603(.A1(new_n802), .A2(new_n804), .A3(new_n730), .ZN(new_n805));
  OAI21_X1  g604(.A(KEYINPUT119), .B1(new_n800), .B2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT119), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n802), .A2(new_n804), .A3(new_n730), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n781), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n806), .A2(new_n753), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n576), .A2(new_n463), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT117), .ZN(new_n812));
  XNOR2_X1  g611(.A(new_n811), .B(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n810), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(KEYINPUT120), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT120), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n810), .A2(new_n816), .A3(new_n813), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n815), .A2(new_n248), .A3(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n795), .B1(new_n818), .B2(new_n770), .ZN(new_n819));
  NOR3_X1   g618(.A1(new_n819), .A2(new_n666), .A3(new_n769), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT121), .ZN(new_n821));
  OR2_X1    g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n792), .B1(new_n820), .B2(new_n821), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n794), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  AOI211_X1 g623(.A(KEYINPUT59), .B(new_n792), .C1(new_n784), .C2(new_n575), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n793), .B1(new_n824), .B2(new_n825), .ZN(G1345gat));
  NAND3_X1  g625(.A1(new_n766), .A2(new_n212), .A3(new_n548), .ZN(new_n827));
  AND2_X1   g626(.A1(new_n784), .A2(new_n618), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n827), .B1(new_n212), .B2(new_n828), .ZN(G1346gat));
  AOI21_X1  g628(.A(G162gat), .B1(new_n766), .B2(new_n607), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n501), .A2(new_n213), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n830), .B1(new_n784), .B2(new_n831), .ZN(G1347gat));
  NOR2_X1   g631(.A1(new_n349), .A2(new_n295), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n737), .A2(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(G169gat), .B1(new_n834), .B2(new_n463), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n736), .A2(new_n349), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n836), .A2(new_n296), .A3(new_n383), .ZN(new_n837));
  OR2_X1    g636(.A1(new_n622), .A2(G169gat), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n835), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  XOR2_X1   g638(.A(new_n839), .B(KEYINPUT122), .Z(G1348gat));
  OAI21_X1  g639(.A(G176gat), .B1(new_n834), .B2(new_n666), .ZN(new_n841));
  OR2_X1    g640(.A1(new_n666), .A2(G176gat), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n841), .B1(new_n837), .B2(new_n842), .ZN(G1349gat));
  INV_X1    g642(.A(new_n837), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n844), .A2(new_n271), .A3(new_n548), .ZN(new_n845));
  OAI21_X1  g644(.A(G183gat), .B1(new_n834), .B2(new_n617), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g646(.A(new_n847), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g647(.A(G190gat), .B1(new_n834), .B2(new_n501), .ZN(new_n849));
  XNOR2_X1  g648(.A(new_n849), .B(KEYINPUT61), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n844), .A2(new_n272), .A3(new_n607), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(G1351gat));
  NAND4_X1  g651(.A1(new_n591), .A2(new_n248), .A3(new_n296), .A4(new_n594), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT123), .ZN(new_n854));
  OR2_X1    g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n853), .A2(new_n854), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n855), .A2(new_n836), .A3(new_n856), .ZN(new_n857));
  NOR3_X1   g656(.A1(new_n857), .A2(G197gat), .A3(new_n622), .ZN(new_n858));
  OR2_X1    g657(.A1(new_n819), .A2(KEYINPUT124), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n819), .A2(KEYINPUT124), .ZN(new_n860));
  AND2_X1   g659(.A1(new_n596), .A2(new_n833), .ZN(new_n861));
  NAND4_X1  g660(.A1(new_n859), .A2(new_n626), .A3(new_n860), .A4(new_n861), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n858), .B1(new_n862), .B2(G197gat), .ZN(new_n863));
  XNOR2_X1  g662(.A(new_n863), .B(KEYINPUT125), .ZN(G1352gat));
  AND3_X1   g663(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(new_n575), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(G204gat), .ZN(new_n867));
  NOR3_X1   g666(.A1(new_n857), .A2(G204gat), .A3(new_n666), .ZN(new_n868));
  XNOR2_X1  g667(.A(new_n868), .B(KEYINPUT62), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n867), .A2(new_n869), .ZN(G1353gat));
  INV_X1    g669(.A(new_n857), .ZN(new_n871));
  INV_X1    g670(.A(G211gat), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n871), .A2(new_n872), .A3(new_n548), .ZN(new_n873));
  NAND4_X1  g672(.A1(new_n591), .A2(new_n548), .A3(new_n594), .A4(new_n833), .ZN(new_n874));
  XNOR2_X1  g673(.A(new_n811), .B(KEYINPUT117), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n781), .A2(new_n808), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n548), .B1(new_n876), .B2(KEYINPUT119), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n875), .B1(new_n877), .B2(new_n809), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n248), .B1(new_n878), .B2(new_n816), .ZN(new_n879));
  INV_X1    g678(.A(new_n817), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n770), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(new_n795), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n874), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n872), .B1(new_n883), .B2(KEYINPUT126), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT126), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n885), .B1(new_n819), .B2(new_n874), .ZN(new_n886));
  AOI21_X1  g685(.A(KEYINPUT63), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(new_n874), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n249), .B1(new_n814), .B2(KEYINPUT120), .ZN(new_n889));
  AOI21_X1  g688(.A(KEYINPUT57), .B1(new_n889), .B2(new_n817), .ZN(new_n890));
  OAI211_X1 g689(.A(new_n888), .B(KEYINPUT126), .C1(new_n890), .C2(new_n795), .ZN(new_n891));
  AND4_X1   g690(.A1(KEYINPUT63), .A2(new_n886), .A3(G211gat), .A4(new_n891), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n873), .B1(new_n887), .B2(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT127), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  OAI211_X1 g694(.A(KEYINPUT127), .B(new_n873), .C1(new_n887), .C2(new_n892), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(G1354gat));
  AOI21_X1  g696(.A(G218gat), .B1(new_n871), .B2(new_n607), .ZN(new_n898));
  AND2_X1   g697(.A1(new_n607), .A2(G218gat), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n898), .B1(new_n865), .B2(new_n899), .ZN(G1355gat));
endmodule


