

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759;

  AND2_X1 U361 ( .A1(n354), .A2(n355), .ZN(n352) );
  AND2_X1 U362 ( .A1(n641), .A2(n640), .ZN(n355) );
  XNOR2_X1 U363 ( .A(n627), .B(n339), .ZN(n672) );
  XNOR2_X1 U364 ( .A(n628), .B(KEYINPUT96), .ZN(n339) );
  AND2_X1 U365 ( .A1(n403), .A2(n460), .ZN(n697) );
  XNOR2_X1 U366 ( .A(n612), .B(n611), .ZN(n757) );
  XNOR2_X1 U367 ( .A(n623), .B(KEYINPUT73), .ZN(n403) );
  XNOR2_X1 U368 ( .A(n548), .B(n547), .ZN(n586) );
  XNOR2_X1 U369 ( .A(n423), .B(KEYINPUT90), .ZN(n422) );
  XNOR2_X2 U370 ( .A(n742), .B(n556), .ZN(n651) );
  XNOR2_X1 U371 ( .A(n405), .B(n404), .ZN(n390) );
  NAND2_X1 U372 ( .A1(n389), .A2(n373), .ZN(n405) );
  INV_X2 U373 ( .A(KEYINPUT3), .ZN(n423) );
  NOR2_X2 U374 ( .A1(n576), .A2(n630), .ZN(n577) );
  XOR2_X2 U375 ( .A(n493), .B(n492), .Z(n372) );
  XOR2_X2 U376 ( .A(n645), .B(n647), .Z(n341) );
  XOR2_X2 U377 ( .A(n711), .B(n710), .Z(n370) );
  XNOR2_X2 U378 ( .A(n715), .B(n714), .ZN(n716) );
  XNOR2_X2 U379 ( .A(n462), .B(n461), .ZN(n724) );
  NAND2_X2 U380 ( .A1(n418), .A2(n472), .ZN(n470) );
  NOR2_X2 U381 ( .A1(n682), .A2(n679), .ZN(n429) );
  NOR2_X1 U382 ( .A1(n671), .A2(n669), .ZN(n681) );
  XNOR2_X1 U383 ( .A(KEYINPUT86), .B(KEYINPUT63), .ZN(n340) );
  XNOR2_X1 U384 ( .A(n350), .B(KEYINPUT45), .ZN(n728) );
  NOR2_X2 U385 ( .A1(n596), .A2(n559), .ZN(n560) );
  XNOR2_X2 U386 ( .A(n594), .B(n427), .ZN(n395) );
  NAND2_X1 U387 ( .A1(n363), .A2(n362), .ZN(n361) );
  INV_X1 U388 ( .A(n704), .ZN(n360) );
  INV_X1 U389 ( .A(n583), .ZN(n630) );
  XNOR2_X1 U390 ( .A(n443), .B(G125), .ZN(n518) );
  NOR2_X1 U391 ( .A1(n457), .A2(G953), .ZN(n456) );
  XNOR2_X1 U392 ( .A(G140), .B(G137), .ZN(n549) );
  INV_X1 U393 ( .A(KEYINPUT60), .ZN(n344) );
  INV_X1 U394 ( .A(KEYINPUT56), .ZN(n347) );
  XNOR2_X1 U395 ( .A(KEYINPUT8), .B(KEYINPUT68), .ZN(n458) );
  INV_X1 U396 ( .A(G146), .ZN(n443) );
  NOR2_X1 U397 ( .A1(n708), .A2(G953), .ZN(n343) );
  NAND2_X1 U398 ( .A1(n361), .A2(n360), .ZN(n705) );
  XNOR2_X1 U399 ( .A(n700), .B(n364), .ZN(n363) );
  AND2_X1 U400 ( .A1(n400), .A2(n398), .ZN(n397) );
  NOR2_X1 U401 ( .A1(n757), .A2(n755), .ZN(n430) );
  XNOR2_X1 U402 ( .A(n597), .B(KEYINPUT112), .ZN(n758) );
  XNOR2_X1 U403 ( .A(n359), .B(n357), .ZN(n356) );
  NOR2_X1 U404 ( .A1(n592), .A2(n591), .ZN(n604) );
  XNOR2_X1 U405 ( .A(n437), .B(KEYINPUT103), .ZN(n671) );
  XNOR2_X1 U406 ( .A(n564), .B(n421), .ZN(n669) );
  XNOR2_X1 U407 ( .A(n583), .B(KEYINPUT6), .ZN(n636) );
  XNOR2_X1 U408 ( .A(n407), .B(n549), .ZN(n742) );
  INV_X1 U409 ( .A(n701), .ZN(n362) );
  XNOR2_X1 U410 ( .A(n486), .B(n487), .ZN(n531) );
  XNOR2_X1 U411 ( .A(n456), .B(n458), .ZN(n534) );
  XNOR2_X1 U412 ( .A(n422), .B(n484), .ZN(n487) );
  XNOR2_X1 U413 ( .A(n518), .B(n442), .ZN(n740) );
  XNOR2_X1 U414 ( .A(n358), .B(KEYINPUT118), .ZN(n357) );
  INV_X1 U415 ( .A(n727), .ZN(n342) );
  XNOR2_X1 U416 ( .A(n485), .B(G116), .ZN(n486) );
  INV_X1 U417 ( .A(G953), .ZN(n749) );
  XOR2_X1 U418 ( .A(G101), .B(G113), .Z(n485) );
  NOR2_X1 U419 ( .A1(G953), .A2(G237), .ZN(n529) );
  XNOR2_X1 U420 ( .A(KEYINPUT120), .B(KEYINPUT52), .ZN(n364) );
  NAND2_X1 U421 ( .A1(n713), .A2(n342), .ZN(n348) );
  XNOR2_X1 U422 ( .A(n343), .B(KEYINPUT53), .ZN(G75) );
  OR2_X2 U423 ( .A1(n705), .A2(n706), .ZN(n707) );
  XNOR2_X1 U424 ( .A(n345), .B(n344), .ZN(G60) );
  NAND2_X1 U425 ( .A1(n718), .A2(n342), .ZN(n345) );
  XNOR2_X1 U426 ( .A(n346), .B(n340), .ZN(G57) );
  NAND2_X1 U427 ( .A1(n349), .A2(n342), .ZN(n346) );
  BUF_X2 U428 ( .A(n365), .Z(n385) );
  XNOR2_X2 U429 ( .A(n644), .B(KEYINPUT65), .ZN(n365) );
  XNOR2_X2 U430 ( .A(n451), .B(n419), .ZN(n406) );
  XNOR2_X2 U431 ( .A(n644), .B(KEYINPUT65), .ZN(n723) );
  XNOR2_X1 U432 ( .A(n348), .B(n347), .ZN(G51) );
  NAND2_X2 U433 ( .A1(n706), .A2(n643), .ZN(n644) );
  XNOR2_X2 U434 ( .A(n382), .B(KEYINPUT2), .ZN(n706) );
  XNOR2_X1 U435 ( .A(n648), .B(n341), .ZN(n349) );
  NAND2_X1 U436 ( .A1(n352), .A2(n351), .ZN(n350) );
  NAND2_X1 U437 ( .A1(n353), .A2(n386), .ZN(n351) );
  NAND2_X1 U438 ( .A1(n479), .A2(n621), .ZN(n353) );
  NAND2_X1 U439 ( .A1(n478), .A2(KEYINPUT44), .ZN(n354) );
  NAND2_X1 U440 ( .A1(n356), .A2(n703), .ZN(n698) );
  INV_X1 U441 ( .A(KEYINPUT51), .ZN(n358) );
  OR2_X1 U442 ( .A1(n696), .A2(n697), .ZN(n359) );
  XNOR2_X1 U443 ( .A(n481), .B(KEYINPUT19), .ZN(n366) );
  NAND2_X2 U444 ( .A1(n603), .A2(n677), .ZN(n481) );
  BUF_X1 U445 ( .A(n754), .Z(n367) );
  XNOR2_X1 U446 ( .A(n405), .B(n404), .ZN(n368) );
  XNOR2_X1 U447 ( .A(n528), .B(n527), .ZN(n407) );
  XNOR2_X2 U448 ( .A(n494), .B(n372), .ZN(n603) );
  OR2_X1 U449 ( .A1(G237), .A2(G902), .ZN(n491) );
  NAND2_X1 U450 ( .A1(n473), .A2(KEYINPUT48), .ZN(n472) );
  XNOR2_X1 U451 ( .A(n441), .B(G104), .ZN(n516) );
  INV_X1 U452 ( .A(G122), .ZN(n441) );
  XNOR2_X1 U453 ( .A(G134), .B(G131), .ZN(n527) );
  NAND2_X1 U454 ( .A1(n469), .A2(n474), .ZN(n468) );
  INV_X1 U455 ( .A(KEYINPUT82), .ZN(n416) );
  NOR2_X1 U456 ( .A1(n470), .A2(n675), .ZN(n392) );
  INV_X1 U457 ( .A(KEYINPUT38), .ZN(n427) );
  AND2_X1 U458 ( .A1(G953), .A2(G902), .ZN(n496) );
  NAND2_X1 U459 ( .A1(G214), .A2(n491), .ZN(n677) );
  INV_X1 U460 ( .A(G234), .ZN(n457) );
  XOR2_X1 U461 ( .A(n376), .B(n518), .Z(n369) );
  NAND2_X1 U462 ( .A1(n586), .A2(n569), .ZN(n576) );
  XNOR2_X1 U463 ( .A(n531), .B(n476), .ZN(n475) );
  XNOR2_X1 U464 ( .A(n477), .B(n532), .ZN(n476) );
  XOR2_X1 U465 ( .A(KEYINPUT5), .B(G137), .Z(n532) );
  XNOR2_X1 U466 ( .A(G107), .B(G110), .ZN(n734) );
  XNOR2_X1 U467 ( .A(n531), .B(n483), .ZN(n733) );
  XNOR2_X1 U468 ( .A(n516), .B(KEYINPUT16), .ZN(n483) );
  XNOR2_X1 U469 ( .A(G116), .B(G122), .ZN(n503) );
  XOR2_X1 U470 ( .A(KEYINPUT7), .B(G107), .Z(n504) );
  XOR2_X1 U471 ( .A(KEYINPUT98), .B(KEYINPUT11), .Z(n511) );
  XNOR2_X1 U472 ( .A(G131), .B(G113), .ZN(n510) );
  INV_X1 U473 ( .A(KEYINPUT10), .ZN(n442) );
  XNOR2_X1 U474 ( .A(n516), .B(n440), .ZN(n439) );
  XNOR2_X1 U475 ( .A(n517), .B(G140), .ZN(n440) );
  XOR2_X1 U476 ( .A(G143), .B(KEYINPUT99), .Z(n513) );
  XNOR2_X1 U477 ( .A(n734), .B(KEYINPUT71), .ZN(n555) );
  XNOR2_X1 U478 ( .A(G104), .B(G101), .ZN(n551) );
  NAND2_X1 U479 ( .A1(n384), .A2(n383), .ZN(n746) );
  NAND2_X1 U480 ( .A1(n391), .A2(n615), .ZN(n384) );
  NOR2_X1 U481 ( .A1(n468), .A2(n416), .ZN(n413) );
  XNOR2_X1 U482 ( .A(n622), .B(n453), .ZN(n596) );
  INV_X1 U483 ( .A(KEYINPUT88), .ZN(n453) );
  INV_X1 U484 ( .A(KEYINPUT0), .ZN(n404) );
  XNOR2_X1 U485 ( .A(n509), .B(G478), .ZN(n581) );
  NAND2_X1 U486 ( .A1(n557), .A2(G902), .ZN(n449) );
  INV_X1 U487 ( .A(KEYINPUT35), .ZN(n387) );
  NAND2_X1 U488 ( .A1(n397), .A2(n377), .ZN(n402) );
  INV_X1 U489 ( .A(KEYINPUT85), .ZN(n419) );
  XNOR2_X1 U490 ( .A(n430), .B(n424), .ZN(n393) );
  INV_X1 U491 ( .A(KEYINPUT46), .ZN(n424) );
  INV_X1 U492 ( .A(n394), .ZN(n678) );
  XNOR2_X1 U493 ( .A(n530), .B(G146), .ZN(n477) );
  XNOR2_X1 U494 ( .A(KEYINPUT15), .B(G902), .ZN(n642) );
  NAND2_X1 U495 ( .A1(n415), .A2(n414), .ZN(n391) );
  NAND2_X1 U496 ( .A1(G234), .A2(G237), .ZN(n495) );
  NOR2_X1 U497 ( .A1(n576), .A2(n636), .ZN(n570) );
  AND2_X1 U498 ( .A1(n634), .A2(n455), .ZN(n399) );
  NAND2_X1 U499 ( .A1(G469), .A2(n447), .ZN(n446) );
  XNOR2_X1 U500 ( .A(n381), .B(n380), .ZN(n482) );
  XNOR2_X1 U501 ( .A(n490), .B(n555), .ZN(n380) );
  XNOR2_X1 U502 ( .A(n528), .B(n369), .ZN(n381) );
  NAND2_X1 U503 ( .A1(n403), .A2(n459), .ZN(n624) );
  INV_X1 U504 ( .A(n636), .ZN(n459) );
  INV_X1 U505 ( .A(n690), .ZN(n454) );
  INV_X1 U506 ( .A(KEYINPUT41), .ZN(n428) );
  XNOR2_X1 U507 ( .A(KEYINPUT83), .B(KEYINPUT39), .ZN(n605) );
  OR2_X1 U508 ( .A1(n634), .A2(n455), .ZN(n396) );
  INV_X1 U509 ( .A(n465), .ZN(n662) );
  INV_X1 U510 ( .A(n630), .ZN(n460) );
  AND2_X1 U511 ( .A1(n686), .A2(n687), .ZN(n689) );
  INV_X1 U512 ( .A(KEYINPUT22), .ZN(n425) );
  XNOR2_X1 U513 ( .A(n543), .B(n540), .ZN(n461) );
  XNOR2_X1 U514 ( .A(G119), .B(G110), .ZN(n540) );
  XNOR2_X1 U515 ( .A(n420), .B(n502), .ZN(n508) );
  XOR2_X1 U516 ( .A(G134), .B(KEYINPUT9), .Z(n502) );
  XNOR2_X1 U517 ( .A(n740), .B(n439), .ZN(n519) );
  XNOR2_X1 U518 ( .A(KEYINPUT74), .B(G146), .ZN(n552) );
  AND2_X1 U519 ( .A1(n435), .A2(n434), .ZN(n597) );
  INV_X1 U520 ( .A(n596), .ZN(n434) );
  NAND2_X1 U521 ( .A1(n408), .A2(n626), .ZN(n666) );
  XNOR2_X1 U522 ( .A(n410), .B(n409), .ZN(n408) );
  INV_X1 U523 ( .A(KEYINPUT108), .ZN(n409) );
  INV_X1 U524 ( .A(n581), .ZN(n438) );
  INV_X1 U525 ( .A(KEYINPUT102), .ZN(n421) );
  NAND2_X1 U526 ( .A1(n575), .A2(n581), .ZN(n564) );
  INV_X1 U527 ( .A(n386), .ZN(n753) );
  XNOR2_X1 U528 ( .A(n626), .B(KEYINPUT76), .ZN(n371) );
  XNOR2_X1 U529 ( .A(n524), .B(n523), .ZN(n575) );
  OR2_X1 U530 ( .A1(n568), .A2(n499), .ZN(n373) );
  NOR2_X1 U531 ( .A1(n571), .A2(n433), .ZN(n374) );
  XOR2_X1 U532 ( .A(n681), .B(KEYINPUT80), .Z(n375) );
  NAND2_X1 U533 ( .A1(G224), .A2(n749), .ZN(n376) );
  AND2_X1 U534 ( .A1(n396), .A2(n371), .ZN(n377) );
  INV_X1 U535 ( .A(G902), .ZN(n447) );
  XNOR2_X1 U536 ( .A(KEYINPUT111), .B(KEYINPUT36), .ZN(n378) );
  AND2_X1 U537 ( .A1(n464), .A2(KEYINPUT80), .ZN(n379) );
  XNOR2_X1 U538 ( .A(n482), .B(n733), .ZN(n709) );
  AND2_X1 U539 ( .A1(n649), .A2(G953), .ZN(n727) );
  XNOR2_X2 U540 ( .A(n505), .B(KEYINPUT4), .ZN(n528) );
  XNOR2_X2 U541 ( .A(n444), .B(G143), .ZN(n505) );
  NAND2_X1 U542 ( .A1(n728), .A2(n746), .ZN(n382) );
  NAND2_X1 U543 ( .A1(n392), .A2(n413), .ZN(n383) );
  XNOR2_X2 U544 ( .A(n402), .B(n387), .ZN(n386) );
  XNOR2_X1 U545 ( .A(n481), .B(KEYINPUT19), .ZN(n389) );
  NAND2_X1 U546 ( .A1(n432), .A2(n431), .ZN(n601) );
  BUF_X2 U547 ( .A(n603), .Z(n594) );
  BUF_X1 U548 ( .A(n728), .Z(n388) );
  NAND2_X1 U549 ( .A1(n610), .A2(n366), .ZN(n465) );
  NAND2_X1 U550 ( .A1(n390), .A2(n526), .ZN(n426) );
  NAND2_X1 U551 ( .A1(n697), .A2(n368), .ZN(n627) );
  XNOR2_X1 U552 ( .A(n368), .B(KEYINPUT94), .ZN(n634) );
  NOR2_X1 U553 ( .A1(n393), .A2(KEYINPUT48), .ZN(n471) );
  NAND2_X1 U554 ( .A1(n393), .A2(KEYINPUT48), .ZN(n469) );
  NAND2_X1 U555 ( .A1(n395), .A2(n677), .ZN(n682) );
  OR2_X1 U556 ( .A1(n395), .A2(n677), .ZN(n394) );
  NAND2_X1 U557 ( .A1(n604), .A2(n395), .ZN(n606) );
  NAND2_X1 U558 ( .A1(n399), .A2(n702), .ZN(n398) );
  NAND2_X1 U559 ( .A1(n401), .A2(n625), .ZN(n400) );
  INV_X1 U560 ( .A(n702), .ZN(n401) );
  NAND2_X1 U561 ( .A1(n406), .A2(n386), .ZN(n478) );
  OR2_X2 U562 ( .A1(n406), .A2(KEYINPUT84), .ZN(n479) );
  NAND2_X1 U563 ( .A1(n406), .A2(n620), .ZN(n621) );
  XNOR2_X1 U564 ( .A(n407), .B(n475), .ZN(n645) );
  NAND2_X1 U565 ( .A1(n411), .A2(n666), .ZN(n593) );
  NAND2_X1 U566 ( .A1(n604), .A2(n594), .ZN(n410) );
  NAND2_X1 U567 ( .A1(n412), .A2(n580), .ZN(n411) );
  NAND2_X1 U568 ( .A1(n662), .A2(n579), .ZN(n412) );
  NAND2_X1 U569 ( .A1(n468), .A2(n416), .ZN(n414) );
  NAND2_X1 U570 ( .A1(n470), .A2(n416), .ZN(n415) );
  NAND2_X1 U571 ( .A1(n534), .A2(G221), .ZN(n536) );
  NAND2_X1 U572 ( .A1(n417), .A2(n463), .ZN(n462) );
  NAND2_X1 U573 ( .A1(n539), .A2(n740), .ZN(n417) );
  NOR2_X2 U574 ( .A1(n724), .A2(G902), .ZN(n548) );
  BUF_X1 U575 ( .A(n622), .Z(n690) );
  XNOR2_X2 U576 ( .A(n618), .B(KEYINPUT105), .ZN(n754) );
  NAND2_X1 U577 ( .A1(n450), .A2(n449), .ZN(n448) );
  NAND2_X1 U578 ( .A1(n471), .A2(n467), .ZN(n418) );
  OR2_X2 U579 ( .A1(n448), .A2(n445), .ZN(n631) );
  XNOR2_X1 U580 ( .A(n429), .B(n428), .ZN(n703) );
  NAND2_X1 U581 ( .A1(n602), .A2(n601), .ZN(n473) );
  NAND2_X1 U582 ( .A1(n534), .A2(G217), .ZN(n420) );
  XNOR2_X1 U583 ( .A(n436), .B(n378), .ZN(n435) );
  OR2_X2 U584 ( .A1(n598), .A2(n758), .ZN(n600) );
  XNOR2_X2 U585 ( .A(n426), .B(n425), .ZN(n639) );
  NOR2_X1 U586 ( .A1(n758), .A2(n599), .ZN(n431) );
  INV_X1 U587 ( .A(n598), .ZN(n432) );
  NOR2_X1 U588 ( .A1(n607), .A2(n571), .ZN(n595) );
  NAND2_X1 U589 ( .A1(n669), .A2(n374), .ZN(n436) );
  INV_X1 U590 ( .A(n594), .ZN(n433) );
  XNOR2_X1 U591 ( .A(n681), .B(n379), .ZN(n579) );
  NAND2_X1 U592 ( .A1(n582), .A2(n438), .ZN(n437) );
  XNOR2_X2 U593 ( .A(G128), .B(KEYINPUT64), .ZN(n444) );
  XNOR2_X2 U594 ( .A(n631), .B(n558), .ZN(n622) );
  NOR2_X1 U595 ( .A1(n651), .A2(n446), .ZN(n445) );
  NAND2_X1 U596 ( .A1(n651), .A2(n557), .ZN(n450) );
  NOR2_X2 U597 ( .A1(n619), .A2(n754), .ZN(n451) );
  XNOR2_X2 U598 ( .A(n452), .B(n563), .ZN(n619) );
  NAND2_X1 U599 ( .A1(n639), .A2(n561), .ZN(n452) );
  NAND2_X1 U600 ( .A1(n595), .A2(n454), .ZN(n572) );
  INV_X1 U601 ( .A(n625), .ZN(n455) );
  NAND2_X1 U602 ( .A1(n538), .A2(n537), .ZN(n463) );
  XNOR2_X2 U603 ( .A(n466), .B(KEYINPUT109), .ZN(n610) );
  NAND2_X1 U604 ( .A1(n465), .A2(n464), .ZN(n580) );
  INV_X1 U605 ( .A(KEYINPUT47), .ZN(n464) );
  NAND2_X1 U606 ( .A1(n578), .A2(n590), .ZN(n466) );
  INV_X1 U607 ( .A(n473), .ZN(n467) );
  INV_X1 U608 ( .A(n676), .ZN(n474) );
  INV_X1 U609 ( .A(KEYINPUT84), .ZN(n480) );
  INV_X1 U610 ( .A(KEYINPUT12), .ZN(n517) );
  XNOR2_X1 U611 ( .A(n546), .B(n545), .ZN(n547) );
  INV_X1 U612 ( .A(n575), .ZN(n582) );
  XNOR2_X1 U613 ( .A(n719), .B(KEYINPUT122), .ZN(n720) );
  XNOR2_X1 U614 ( .A(n606), .B(n605), .ZN(n614) );
  XNOR2_X1 U615 ( .A(n721), .B(n720), .ZN(n722) );
  XNOR2_X1 U616 ( .A(G119), .B(KEYINPUT70), .ZN(n484) );
  XOR2_X1 U617 ( .A(KEYINPUT75), .B(KEYINPUT91), .Z(n489) );
  XNOR2_X1 U618 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n488) );
  XNOR2_X1 U619 ( .A(n489), .B(n488), .ZN(n490) );
  NAND2_X1 U620 ( .A1(n709), .A2(n642), .ZN(n494) );
  XOR2_X1 U621 ( .A(KEYINPUT79), .B(KEYINPUT92), .Z(n493) );
  NAND2_X1 U622 ( .A1(G210), .A2(n491), .ZN(n492) );
  XNOR2_X1 U623 ( .A(n495), .B(KEYINPUT14), .ZN(n497) );
  NAND2_X1 U624 ( .A1(G952), .A2(n497), .ZN(n701) );
  NOR2_X1 U625 ( .A1(G953), .A2(n701), .ZN(n568) );
  NAND2_X1 U626 ( .A1(n497), .A2(n496), .ZN(n565) );
  NOR2_X1 U627 ( .A1(G898), .A2(n565), .ZN(n498) );
  XOR2_X1 U628 ( .A(KEYINPUT93), .B(n498), .Z(n499) );
  NAND2_X1 U629 ( .A1(G234), .A2(n642), .ZN(n500) );
  XNOR2_X1 U630 ( .A(KEYINPUT20), .B(n500), .ZN(n544) );
  NAND2_X1 U631 ( .A1(n544), .A2(G221), .ZN(n501) );
  XNOR2_X1 U632 ( .A(KEYINPUT21), .B(n501), .ZN(n585) );
  XNOR2_X1 U633 ( .A(n504), .B(n503), .ZN(n506) );
  XNOR2_X1 U634 ( .A(n505), .B(n506), .ZN(n507) );
  XNOR2_X1 U635 ( .A(n508), .B(n507), .ZN(n719) );
  NOR2_X1 U636 ( .A1(n719), .A2(G902), .ZN(n509) );
  XNOR2_X1 U637 ( .A(n511), .B(n510), .ZN(n515) );
  NAND2_X1 U638 ( .A1(G214), .A2(n529), .ZN(n512) );
  XNOR2_X1 U639 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U640 ( .A(n515), .B(n514), .ZN(n520) );
  XNOR2_X1 U641 ( .A(n520), .B(n519), .ZN(n715) );
  NOR2_X1 U642 ( .A1(n715), .A2(G902), .ZN(n524) );
  XOR2_X1 U643 ( .A(KEYINPUT101), .B(KEYINPUT13), .Z(n522) );
  XNOR2_X1 U644 ( .A(KEYINPUT100), .B(G475), .ZN(n521) );
  XNOR2_X1 U645 ( .A(n522), .B(n521), .ZN(n523) );
  NAND2_X1 U646 ( .A1(n581), .A2(n582), .ZN(n525) );
  XNOR2_X1 U647 ( .A(n525), .B(KEYINPUT104), .ZN(n679) );
  NOR2_X1 U648 ( .A1(n585), .A2(n679), .ZN(n526) );
  NAND2_X1 U649 ( .A1(G210), .A2(n529), .ZN(n530) );
  NAND2_X1 U650 ( .A1(n645), .A2(n447), .ZN(n533) );
  XNOR2_X2 U651 ( .A(n533), .B(G472), .ZN(n583) );
  XNOR2_X1 U652 ( .A(n549), .B(KEYINPUT95), .ZN(n535) );
  XNOR2_X1 U653 ( .A(n536), .B(n535), .ZN(n538) );
  INV_X1 U654 ( .A(n740), .ZN(n537) );
  INV_X1 U655 ( .A(n538), .ZN(n539) );
  XOR2_X1 U656 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n542) );
  XNOR2_X1 U657 ( .A(G128), .B(KEYINPUT81), .ZN(n541) );
  XNOR2_X1 U658 ( .A(n542), .B(n541), .ZN(n543) );
  NAND2_X1 U659 ( .A1(n544), .A2(G217), .ZN(n546) );
  INV_X1 U660 ( .A(KEYINPUT25), .ZN(n545) );
  NAND2_X1 U661 ( .A1(n636), .A2(n586), .ZN(n559) );
  NAND2_X1 U662 ( .A1(n749), .A2(G227), .ZN(n550) );
  XNOR2_X1 U663 ( .A(n551), .B(n550), .ZN(n553) );
  XNOR2_X1 U664 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X1 U665 ( .A(n555), .B(n554), .ZN(n556) );
  INV_X1 U666 ( .A(G469), .ZN(n557) );
  XNOR2_X1 U667 ( .A(KEYINPUT67), .B(KEYINPUT1), .ZN(n558) );
  XNOR2_X1 U668 ( .A(n560), .B(KEYINPUT78), .ZN(n561) );
  INV_X1 U669 ( .A(KEYINPUT66), .ZN(n562) );
  XNOR2_X1 U670 ( .A(n562), .B(KEYINPUT32), .ZN(n563) );
  XOR2_X1 U671 ( .A(n619), .B(G119), .Z(G21) );
  INV_X1 U672 ( .A(n669), .ZN(n607) );
  XNOR2_X1 U673 ( .A(KEYINPUT106), .B(n565), .ZN(n566) );
  NOR2_X1 U674 ( .A1(G900), .A2(n566), .ZN(n567) );
  NOR2_X1 U675 ( .A1(n568), .A2(n567), .ZN(n588) );
  NOR2_X1 U676 ( .A1(n588), .A2(n585), .ZN(n569) );
  NAND2_X1 U677 ( .A1(n570), .A2(n677), .ZN(n571) );
  XNOR2_X1 U678 ( .A(n572), .B(KEYINPUT107), .ZN(n573) );
  XNOR2_X1 U679 ( .A(n573), .B(KEYINPUT43), .ZN(n574) );
  NOR2_X1 U680 ( .A1(n594), .A2(n574), .ZN(n676) );
  XNOR2_X1 U681 ( .A(n577), .B(KEYINPUT28), .ZN(n578) );
  INV_X1 U682 ( .A(n631), .ZN(n590) );
  NOR2_X1 U683 ( .A1(n582), .A2(n581), .ZN(n626) );
  NAND2_X1 U684 ( .A1(n583), .A2(n677), .ZN(n584) );
  XOR2_X1 U685 ( .A(KEYINPUT30), .B(n584), .Z(n587) );
  INV_X1 U686 ( .A(n585), .ZN(n686) );
  INV_X1 U687 ( .A(n586), .ZN(n687) );
  NAND2_X1 U688 ( .A1(n587), .A2(n689), .ZN(n592) );
  INV_X1 U689 ( .A(n588), .ZN(n589) );
  NAND2_X1 U690 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U691 ( .A(n593), .B(KEYINPUT72), .ZN(n598) );
  INV_X1 U692 ( .A(KEYINPUT69), .ZN(n599) );
  NAND2_X1 U693 ( .A1(n600), .A2(n599), .ZN(n602) );
  XNOR2_X1 U694 ( .A(KEYINPUT110), .B(KEYINPUT40), .ZN(n609) );
  NOR2_X1 U695 ( .A1(n614), .A2(n607), .ZN(n608) );
  XNOR2_X1 U696 ( .A(n609), .B(n608), .ZN(n755) );
  INV_X1 U697 ( .A(KEYINPUT42), .ZN(n612) );
  NAND2_X1 U698 ( .A1(n703), .A2(n610), .ZN(n611) );
  INV_X1 U699 ( .A(n671), .ZN(n613) );
  NOR2_X1 U700 ( .A1(n614), .A2(n613), .ZN(n675) );
  INV_X1 U701 ( .A(n675), .ZN(n615) );
  OR2_X1 U702 ( .A1(n460), .A2(n687), .ZN(n616) );
  NOR2_X1 U703 ( .A1(n690), .A2(n616), .ZN(n617) );
  NAND2_X1 U704 ( .A1(n639), .A2(n617), .ZN(n618) );
  NOR2_X1 U705 ( .A1(n480), .A2(KEYINPUT44), .ZN(n620) );
  XOR2_X1 U706 ( .A(KEYINPUT77), .B(KEYINPUT34), .Z(n625) );
  NAND2_X1 U707 ( .A1(n622), .A2(n689), .ZN(n623) );
  XNOR2_X2 U708 ( .A(n624), .B(KEYINPUT33), .ZN(n702) );
  XOR2_X1 U709 ( .A(KEYINPUT97), .B(KEYINPUT31), .Z(n628) );
  NAND2_X1 U710 ( .A1(n630), .A2(n689), .ZN(n632) );
  NOR2_X1 U711 ( .A1(n632), .A2(n631), .ZN(n633) );
  AND2_X1 U712 ( .A1(n634), .A2(n633), .ZN(n657) );
  OR2_X1 U713 ( .A1(n672), .A2(n657), .ZN(n635) );
  NAND2_X1 U714 ( .A1(n635), .A2(n375), .ZN(n641) );
  NAND2_X1 U715 ( .A1(n636), .A2(n687), .ZN(n637) );
  NOR2_X1 U716 ( .A1(n637), .A2(n690), .ZN(n638) );
  AND2_X1 U717 ( .A1(n639), .A2(n638), .ZN(n655) );
  INV_X1 U718 ( .A(n655), .ZN(n640) );
  INV_X1 U719 ( .A(n642), .ZN(n643) );
  NAND2_X1 U720 ( .A1(n723), .A2(G472), .ZN(n648) );
  XOR2_X1 U721 ( .A(KEYINPUT87), .B(KEYINPUT113), .Z(n646) );
  XNOR2_X1 U722 ( .A(n646), .B(KEYINPUT62), .ZN(n647) );
  INV_X1 U723 ( .A(G952), .ZN(n649) );
  NAND2_X1 U724 ( .A1(n385), .A2(G469), .ZN(n653) );
  XOR2_X1 U725 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n650) );
  XNOR2_X1 U726 ( .A(n651), .B(n650), .ZN(n652) );
  XNOR2_X1 U727 ( .A(n653), .B(n652), .ZN(n654) );
  NOR2_X1 U728 ( .A1(n654), .A2(n727), .ZN(G54) );
  XOR2_X1 U729 ( .A(G101), .B(n655), .Z(G3) );
  NAND2_X1 U730 ( .A1(n657), .A2(n669), .ZN(n656) );
  XNOR2_X1 U731 ( .A(G104), .B(n656), .ZN(G6) );
  XNOR2_X1 U732 ( .A(KEYINPUT26), .B(KEYINPUT114), .ZN(n661) );
  XOR2_X1 U733 ( .A(G107), .B(KEYINPUT27), .Z(n659) );
  NAND2_X1 U734 ( .A1(n657), .A2(n671), .ZN(n658) );
  XNOR2_X1 U735 ( .A(n659), .B(n658), .ZN(n660) );
  XNOR2_X1 U736 ( .A(n661), .B(n660), .ZN(G9) );
  XOR2_X1 U737 ( .A(KEYINPUT115), .B(KEYINPUT29), .Z(n664) );
  BUF_X1 U738 ( .A(n662), .Z(n667) );
  NAND2_X1 U739 ( .A1(n667), .A2(n671), .ZN(n663) );
  XNOR2_X1 U740 ( .A(n664), .B(n663), .ZN(n665) );
  XOR2_X1 U741 ( .A(G128), .B(n665), .Z(G30) );
  XNOR2_X1 U742 ( .A(G143), .B(n666), .ZN(G45) );
  NAND2_X1 U743 ( .A1(n669), .A2(n667), .ZN(n668) );
  XNOR2_X1 U744 ( .A(n668), .B(G146), .ZN(G48) );
  NAND2_X1 U745 ( .A1(n672), .A2(n669), .ZN(n670) );
  XNOR2_X1 U746 ( .A(n670), .B(G113), .ZN(G15) );
  NAND2_X1 U747 ( .A1(n672), .A2(n671), .ZN(n673) );
  XNOR2_X1 U748 ( .A(n673), .B(KEYINPUT116), .ZN(n674) );
  XNOR2_X1 U749 ( .A(G116), .B(n674), .ZN(G18) );
  XOR2_X1 U750 ( .A(G134), .B(n675), .Z(G36) );
  XOR2_X1 U751 ( .A(G140), .B(n676), .Z(G42) );
  NOR2_X1 U752 ( .A1(n679), .A2(n678), .ZN(n680) );
  XNOR2_X1 U753 ( .A(n680), .B(KEYINPUT119), .ZN(n684) );
  OR2_X1 U754 ( .A1(n682), .A2(n681), .ZN(n683) );
  NAND2_X1 U755 ( .A1(n684), .A2(n683), .ZN(n685) );
  NAND2_X1 U756 ( .A1(n685), .A2(n702), .ZN(n699) );
  NOR2_X1 U757 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U758 ( .A(KEYINPUT49), .B(n688), .ZN(n694) );
  XOR2_X1 U759 ( .A(KEYINPUT117), .B(KEYINPUT50), .Z(n692) );
  NOR2_X1 U760 ( .A1(n690), .A2(n689), .ZN(n691) );
  XOR2_X1 U761 ( .A(n692), .B(n691), .Z(n693) );
  NAND2_X1 U762 ( .A1(n694), .A2(n693), .ZN(n695) );
  NOR2_X1 U763 ( .A1(n460), .A2(n695), .ZN(n696) );
  NAND2_X1 U764 ( .A1(n699), .A2(n698), .ZN(n700) );
  AND2_X1 U765 ( .A1(n703), .A2(n702), .ZN(n704) );
  XOR2_X1 U766 ( .A(KEYINPUT121), .B(n707), .Z(n708) );
  NAND2_X1 U767 ( .A1(n723), .A2(G210), .ZN(n712) );
  INV_X1 U768 ( .A(n709), .ZN(n711) );
  XOR2_X1 U769 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n710) );
  XNOR2_X1 U770 ( .A(n712), .B(n370), .ZN(n713) );
  NAND2_X1 U771 ( .A1(n365), .A2(G475), .ZN(n717) );
  XOR2_X1 U772 ( .A(KEYINPUT59), .B(KEYINPUT89), .Z(n714) );
  XNOR2_X1 U773 ( .A(n717), .B(n716), .ZN(n718) );
  NAND2_X1 U774 ( .A1(n385), .A2(G478), .ZN(n721) );
  NOR2_X1 U775 ( .A1(n727), .A2(n722), .ZN(G63) );
  NAND2_X1 U776 ( .A1(n385), .A2(G217), .ZN(n725) );
  XNOR2_X1 U777 ( .A(n725), .B(n724), .ZN(n726) );
  NOR2_X1 U778 ( .A1(n727), .A2(n726), .ZN(G66) );
  NAND2_X1 U779 ( .A1(n388), .A2(n749), .ZN(n732) );
  NAND2_X1 U780 ( .A1(G953), .A2(G224), .ZN(n729) );
  XNOR2_X1 U781 ( .A(KEYINPUT61), .B(n729), .ZN(n730) );
  NAND2_X1 U782 ( .A1(n730), .A2(G898), .ZN(n731) );
  NAND2_X1 U783 ( .A1(n732), .A2(n731), .ZN(n739) );
  XNOR2_X1 U784 ( .A(n733), .B(KEYINPUT123), .ZN(n735) );
  XNOR2_X1 U785 ( .A(n735), .B(n734), .ZN(n737) );
  NOR2_X1 U786 ( .A1(G898), .A2(n749), .ZN(n736) );
  NOR2_X1 U787 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U788 ( .A(n739), .B(n738), .ZN(G69) );
  XNOR2_X1 U789 ( .A(n740), .B(KEYINPUT124), .ZN(n741) );
  XNOR2_X1 U790 ( .A(n742), .B(n741), .ZN(n748) );
  XNOR2_X1 U791 ( .A(KEYINPUT125), .B(n748), .ZN(n743) );
  XNOR2_X1 U792 ( .A(G227), .B(n743), .ZN(n744) );
  NAND2_X1 U793 ( .A1(n744), .A2(G900), .ZN(n745) );
  NAND2_X1 U794 ( .A1(n745), .A2(G953), .ZN(n752) );
  BUF_X1 U795 ( .A(n746), .Z(n747) );
  XNOR2_X1 U796 ( .A(n748), .B(n747), .ZN(n750) );
  NAND2_X1 U797 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U798 ( .A1(n752), .A2(n751), .ZN(G72) );
  XOR2_X1 U799 ( .A(n753), .B(G122), .Z(G24) );
  XOR2_X1 U800 ( .A(n367), .B(G110), .Z(G12) );
  XOR2_X1 U801 ( .A(G131), .B(n755), .Z(n756) );
  XNOR2_X1 U802 ( .A(KEYINPUT126), .B(n756), .ZN(G33) );
  XOR2_X1 U803 ( .A(G137), .B(n757), .Z(G39) );
  XNOR2_X1 U804 ( .A(G125), .B(KEYINPUT37), .ZN(n759) );
  XNOR2_X1 U805 ( .A(n759), .B(n758), .ZN(G27) );
endmodule

