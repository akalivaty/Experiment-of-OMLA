

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XOR2_X1 U551 ( .A(n701), .B(n700), .Z(n517) );
  NOR2_X2 U552 ( .A1(n760), .A2(n759), .ZN(n761) );
  XOR2_X1 U553 ( .A(KEYINPUT15), .B(n593), .Z(n991) );
  XNOR2_X1 U554 ( .A(KEYINPUT69), .B(KEYINPUT17), .ZN(n527) );
  NOR2_X1 U555 ( .A1(n702), .A2(n793), .ZN(n717) );
  OR2_X2 U556 ( .A1(n702), .A2(n793), .ZN(n741) );
  XNOR2_X1 U557 ( .A(G2104), .B(KEYINPUT66), .ZN(n524) );
  INV_X1 U558 ( .A(KEYINPUT33), .ZN(n773) );
  NOR2_X1 U559 ( .A1(n790), .A2(n789), .ZN(n792) );
  XNOR2_X1 U560 ( .A(n534), .B(n533), .ZN(n536) );
  AND2_X1 U561 ( .A1(n995), .A2(n519), .ZN(n518) );
  OR2_X1 U562 ( .A1(n775), .A2(n788), .ZN(n519) );
  INV_X1 U563 ( .A(KEYINPUT26), .ZN(n714) );
  XNOR2_X1 U564 ( .A(n714), .B(KEYINPUT65), .ZN(n715) );
  XNOR2_X1 U565 ( .A(n716), .B(n715), .ZN(n721) );
  INV_X1 U566 ( .A(KEYINPUT96), .ZN(n733) );
  XNOR2_X1 U567 ( .A(n734), .B(n733), .ZN(n735) );
  NOR2_X1 U568 ( .A1(G2084), .A2(n741), .ZN(n696) );
  INV_X1 U569 ( .A(KEYINPUT23), .ZN(n533) );
  INV_X1 U570 ( .A(KEYINPUT103), .ZN(n791) );
  INV_X1 U571 ( .A(G2105), .ZN(n523) );
  AND2_X1 U572 ( .A1(n524), .A2(n523), .ZN(n613) );
  AND2_X1 U573 ( .A1(n539), .A2(n538), .ZN(n695) );
  NOR2_X1 U574 ( .A1(n532), .A2(n531), .ZN(G164) );
  AND2_X1 U575 ( .A1(G2104), .A2(G2105), .ZN(n893) );
  NAND2_X1 U576 ( .A1(G114), .A2(n893), .ZN(n522) );
  XOR2_X1 U577 ( .A(G2104), .B(KEYINPUT66), .Z(n520) );
  AND2_X1 U578 ( .A1(n520), .A2(G2105), .ZN(n617) );
  NAND2_X1 U579 ( .A1(G126), .A2(n617), .ZN(n521) );
  NAND2_X1 U580 ( .A1(n522), .A2(n521), .ZN(n532) );
  NAND2_X1 U581 ( .A1(G102), .A2(n613), .ZN(n525) );
  XNOR2_X1 U582 ( .A(n525), .B(KEYINPUT86), .ZN(n530) );
  NOR2_X1 U583 ( .A1(G2104), .A2(G2105), .ZN(n526) );
  XNOR2_X1 U584 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U585 ( .A(KEYINPUT68), .B(n528), .ZN(n621) );
  NAND2_X1 U586 ( .A1(G138), .A2(n621), .ZN(n529) );
  NAND2_X1 U587 ( .A1(n530), .A2(n529), .ZN(n531) );
  NAND2_X1 U588 ( .A1(n613), .A2(G101), .ZN(n534) );
  NAND2_X1 U589 ( .A1(n617), .A2(G125), .ZN(n535) );
  NAND2_X1 U590 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U591 ( .A(n537), .B(KEYINPUT67), .ZN(n539) );
  NAND2_X1 U592 ( .A1(G113), .A2(n893), .ZN(n538) );
  NAND2_X1 U593 ( .A1(n621), .A2(G137), .ZN(n540) );
  XNOR2_X1 U594 ( .A(KEYINPUT70), .B(n540), .ZN(n693) );
  AND2_X1 U595 ( .A1(n695), .A2(n693), .ZN(G160) );
  XNOR2_X1 U596 ( .A(G2451), .B(G2443), .ZN(n550) );
  XOR2_X1 U597 ( .A(G2446), .B(G2454), .Z(n542) );
  XNOR2_X1 U598 ( .A(KEYINPUT107), .B(G2435), .ZN(n541) );
  XNOR2_X1 U599 ( .A(n542), .B(n541), .ZN(n546) );
  XOR2_X1 U600 ( .A(KEYINPUT106), .B(G2438), .Z(n544) );
  XNOR2_X1 U601 ( .A(G1348), .B(G1341), .ZN(n543) );
  XNOR2_X1 U602 ( .A(n544), .B(n543), .ZN(n545) );
  XOR2_X1 U603 ( .A(n546), .B(n545), .Z(n548) );
  XNOR2_X1 U604 ( .A(G2430), .B(G2427), .ZN(n547) );
  XNOR2_X1 U605 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U606 ( .A(n550), .B(n549), .ZN(n551) );
  AND2_X1 U607 ( .A1(n551), .A2(G14), .ZN(G401) );
  AND2_X1 U608 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U609 ( .A(G57), .ZN(G237) );
  INV_X1 U610 ( .A(G132), .ZN(G219) );
  INV_X1 U611 ( .A(G82), .ZN(G220) );
  INV_X1 U612 ( .A(G651), .ZN(n554) );
  NOR2_X1 U613 ( .A1(G543), .A2(n554), .ZN(n552) );
  XOR2_X1 U614 ( .A(KEYINPUT1), .B(n552), .Z(n663) );
  NAND2_X1 U615 ( .A1(n663), .A2(G64), .ZN(n553) );
  XNOR2_X1 U616 ( .A(KEYINPUT73), .B(n553), .ZN(n562) );
  NOR2_X1 U617 ( .A1(G651), .A2(G543), .ZN(n649) );
  NAND2_X1 U618 ( .A1(G90), .A2(n649), .ZN(n556) );
  XOR2_X1 U619 ( .A(KEYINPUT0), .B(G543), .Z(n664) );
  NOR2_X2 U620 ( .A1(n664), .A2(n554), .ZN(n652) );
  NAND2_X1 U621 ( .A1(G77), .A2(n652), .ZN(n555) );
  NAND2_X1 U622 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U623 ( .A(n557), .B(KEYINPUT9), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n558), .B(KEYINPUT74), .ZN(n560) );
  NOR2_X2 U625 ( .A1(G651), .A2(n664), .ZN(n659) );
  NAND2_X1 U626 ( .A1(n659), .A2(G52), .ZN(n559) );
  NAND2_X1 U627 ( .A1(n560), .A2(n559), .ZN(n561) );
  NOR2_X1 U628 ( .A1(n562), .A2(n561), .ZN(G171) );
  NAND2_X1 U629 ( .A1(G89), .A2(n649), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n563), .B(KEYINPUT78), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n564), .B(KEYINPUT4), .ZN(n566) );
  NAND2_X1 U632 ( .A1(G76), .A2(n652), .ZN(n565) );
  NAND2_X1 U633 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n567), .B(KEYINPUT5), .ZN(n572) );
  NAND2_X1 U635 ( .A1(G63), .A2(n663), .ZN(n569) );
  NAND2_X1 U636 ( .A1(G51), .A2(n659), .ZN(n568) );
  NAND2_X1 U637 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U638 ( .A(KEYINPUT6), .B(n570), .Z(n571) );
  NAND2_X1 U639 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n573), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U641 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U642 ( .A1(G7), .A2(G661), .ZN(n574) );
  XOR2_X1 U643 ( .A(n574), .B(KEYINPUT10), .Z(n846) );
  NAND2_X1 U644 ( .A1(n846), .A2(G567), .ZN(n575) );
  XOR2_X1 U645 ( .A(KEYINPUT11), .B(n575), .Z(G234) );
  XOR2_X1 U646 ( .A(KEYINPUT14), .B(KEYINPUT76), .Z(n577) );
  NAND2_X1 U647 ( .A1(G56), .A2(n663), .ZN(n576) );
  XNOR2_X1 U648 ( .A(n577), .B(n576), .ZN(n585) );
  NAND2_X1 U649 ( .A1(n649), .A2(G81), .ZN(n578) );
  XNOR2_X1 U650 ( .A(n578), .B(KEYINPUT12), .ZN(n580) );
  NAND2_X1 U651 ( .A1(G68), .A2(n652), .ZN(n579) );
  NAND2_X1 U652 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U653 ( .A(n581), .B(KEYINPUT13), .ZN(n583) );
  NAND2_X1 U654 ( .A1(G43), .A2(n659), .ZN(n582) );
  NAND2_X1 U655 ( .A1(n583), .A2(n582), .ZN(n584) );
  NOR2_X1 U656 ( .A1(n585), .A2(n584), .ZN(n974) );
  NAND2_X1 U657 ( .A1(n974), .A2(G860), .ZN(G153) );
  INV_X1 U658 ( .A(G171), .ZN(G301) );
  NAND2_X1 U659 ( .A1(G868), .A2(G301), .ZN(n595) );
  NAND2_X1 U660 ( .A1(G92), .A2(n649), .ZN(n587) );
  NAND2_X1 U661 ( .A1(G66), .A2(n663), .ZN(n586) );
  NAND2_X1 U662 ( .A1(n587), .A2(n586), .ZN(n592) );
  NAND2_X1 U663 ( .A1(G79), .A2(n652), .ZN(n589) );
  NAND2_X1 U664 ( .A1(G54), .A2(n659), .ZN(n588) );
  NAND2_X1 U665 ( .A1(n589), .A2(n588), .ZN(n590) );
  XOR2_X1 U666 ( .A(KEYINPUT77), .B(n590), .Z(n591) );
  NOR2_X1 U667 ( .A1(n592), .A2(n591), .ZN(n593) );
  INV_X1 U668 ( .A(n991), .ZN(n727) );
  INV_X1 U669 ( .A(G868), .ZN(n610) );
  NAND2_X1 U670 ( .A1(n727), .A2(n610), .ZN(n594) );
  NAND2_X1 U671 ( .A1(n595), .A2(n594), .ZN(G284) );
  NAND2_X1 U672 ( .A1(G78), .A2(n652), .ZN(n597) );
  NAND2_X1 U673 ( .A1(G65), .A2(n663), .ZN(n596) );
  NAND2_X1 U674 ( .A1(n597), .A2(n596), .ZN(n600) );
  NAND2_X1 U675 ( .A1(G91), .A2(n649), .ZN(n598) );
  XNOR2_X1 U676 ( .A(KEYINPUT75), .B(n598), .ZN(n599) );
  NOR2_X1 U677 ( .A1(n600), .A2(n599), .ZN(n602) );
  NAND2_X1 U678 ( .A1(n659), .A2(G53), .ZN(n601) );
  NAND2_X1 U679 ( .A1(n602), .A2(n601), .ZN(G299) );
  NOR2_X1 U680 ( .A1(G286), .A2(n610), .ZN(n604) );
  NOR2_X1 U681 ( .A1(G868), .A2(G299), .ZN(n603) );
  NOR2_X1 U682 ( .A1(n604), .A2(n603), .ZN(G297) );
  INV_X1 U683 ( .A(G860), .ZN(n605) );
  NAND2_X1 U684 ( .A1(n605), .A2(G559), .ZN(n606) );
  NAND2_X1 U685 ( .A1(n606), .A2(n991), .ZN(n607) );
  XNOR2_X1 U686 ( .A(n607), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U687 ( .A1(n727), .A2(n610), .ZN(n608) );
  XNOR2_X1 U688 ( .A(n608), .B(KEYINPUT79), .ZN(n609) );
  NOR2_X1 U689 ( .A1(G559), .A2(n609), .ZN(n612) );
  AND2_X1 U690 ( .A1(n610), .A2(n974), .ZN(n611) );
  NOR2_X1 U691 ( .A1(n612), .A2(n611), .ZN(G282) );
  NAND2_X1 U692 ( .A1(G111), .A2(n893), .ZN(n615) );
  BUF_X1 U693 ( .A(n613), .Z(n896) );
  NAND2_X1 U694 ( .A1(G99), .A2(n896), .ZN(n614) );
  NAND2_X1 U695 ( .A1(n615), .A2(n614), .ZN(n616) );
  XNOR2_X1 U696 ( .A(KEYINPUT80), .B(n616), .ZN(n620) );
  NAND2_X1 U697 ( .A1(n617), .A2(G123), .ZN(n618) );
  XOR2_X1 U698 ( .A(KEYINPUT18), .B(n618), .Z(n619) );
  NOR2_X1 U699 ( .A1(n620), .A2(n619), .ZN(n623) );
  BUF_X1 U700 ( .A(n621), .Z(n897) );
  NAND2_X1 U701 ( .A1(G135), .A2(n897), .ZN(n622) );
  NAND2_X1 U702 ( .A1(n623), .A2(n622), .ZN(n933) );
  XNOR2_X1 U703 ( .A(G2096), .B(n933), .ZN(n624) );
  NOR2_X1 U704 ( .A1(n624), .A2(G2100), .ZN(n625) );
  XNOR2_X1 U705 ( .A(n625), .B(KEYINPUT81), .ZN(G156) );
  NAND2_X1 U706 ( .A1(n991), .A2(G559), .ZN(n673) );
  XOR2_X1 U707 ( .A(n673), .B(n974), .Z(n626) );
  NOR2_X1 U708 ( .A1(G860), .A2(n626), .ZN(n627) );
  XOR2_X1 U709 ( .A(KEYINPUT82), .B(n627), .Z(n634) );
  NAND2_X1 U710 ( .A1(G67), .A2(n663), .ZN(n629) );
  NAND2_X1 U711 ( .A1(G55), .A2(n659), .ZN(n628) );
  NAND2_X1 U712 ( .A1(n629), .A2(n628), .ZN(n633) );
  NAND2_X1 U713 ( .A1(G93), .A2(n649), .ZN(n631) );
  NAND2_X1 U714 ( .A1(G80), .A2(n652), .ZN(n630) );
  NAND2_X1 U715 ( .A1(n631), .A2(n630), .ZN(n632) );
  NOR2_X1 U716 ( .A1(n633), .A2(n632), .ZN(n676) );
  XOR2_X1 U717 ( .A(n634), .B(n676), .Z(G145) );
  NAND2_X1 U718 ( .A1(G60), .A2(n663), .ZN(n636) );
  NAND2_X1 U719 ( .A1(G47), .A2(n659), .ZN(n635) );
  NAND2_X1 U720 ( .A1(n636), .A2(n635), .ZN(n641) );
  NAND2_X1 U721 ( .A1(G85), .A2(n649), .ZN(n638) );
  NAND2_X1 U722 ( .A1(G72), .A2(n652), .ZN(n637) );
  NAND2_X1 U723 ( .A1(n638), .A2(n637), .ZN(n639) );
  XOR2_X1 U724 ( .A(KEYINPUT71), .B(n639), .Z(n640) );
  NOR2_X1 U725 ( .A1(n641), .A2(n640), .ZN(n642) );
  XOR2_X1 U726 ( .A(KEYINPUT72), .B(n642), .Z(G290) );
  NAND2_X1 U727 ( .A1(G88), .A2(n649), .ZN(n644) );
  NAND2_X1 U728 ( .A1(G75), .A2(n652), .ZN(n643) );
  NAND2_X1 U729 ( .A1(n644), .A2(n643), .ZN(n648) );
  NAND2_X1 U730 ( .A1(G62), .A2(n663), .ZN(n646) );
  NAND2_X1 U731 ( .A1(G50), .A2(n659), .ZN(n645) );
  NAND2_X1 U732 ( .A1(n646), .A2(n645), .ZN(n647) );
  NOR2_X1 U733 ( .A1(n648), .A2(n647), .ZN(G166) );
  INV_X1 U734 ( .A(G166), .ZN(G303) );
  NAND2_X1 U735 ( .A1(G86), .A2(n649), .ZN(n651) );
  NAND2_X1 U736 ( .A1(G61), .A2(n663), .ZN(n650) );
  NAND2_X1 U737 ( .A1(n651), .A2(n650), .ZN(n655) );
  NAND2_X1 U738 ( .A1(n652), .A2(G73), .ZN(n653) );
  XOR2_X1 U739 ( .A(KEYINPUT2), .B(n653), .Z(n654) );
  NOR2_X1 U740 ( .A1(n655), .A2(n654), .ZN(n656) );
  XOR2_X1 U741 ( .A(KEYINPUT83), .B(n656), .Z(n658) );
  NAND2_X1 U742 ( .A1(n659), .A2(G48), .ZN(n657) );
  NAND2_X1 U743 ( .A1(n658), .A2(n657), .ZN(G305) );
  NAND2_X1 U744 ( .A1(G49), .A2(n659), .ZN(n661) );
  NAND2_X1 U745 ( .A1(G74), .A2(G651), .ZN(n660) );
  NAND2_X1 U746 ( .A1(n661), .A2(n660), .ZN(n662) );
  NOR2_X1 U747 ( .A1(n663), .A2(n662), .ZN(n666) );
  NAND2_X1 U748 ( .A1(n664), .A2(G87), .ZN(n665) );
  NAND2_X1 U749 ( .A1(n666), .A2(n665), .ZN(G288) );
  XOR2_X1 U750 ( .A(G303), .B(n676), .Z(n667) );
  XNOR2_X1 U751 ( .A(n667), .B(KEYINPUT19), .ZN(n668) );
  XNOR2_X1 U752 ( .A(n668), .B(G305), .ZN(n671) );
  XOR2_X1 U753 ( .A(n974), .B(G299), .Z(n669) );
  XNOR2_X1 U754 ( .A(G288), .B(n669), .ZN(n670) );
  XNOR2_X1 U755 ( .A(n671), .B(n670), .ZN(n672) );
  XNOR2_X1 U756 ( .A(G290), .B(n672), .ZN(n853) );
  XOR2_X1 U757 ( .A(n853), .B(n673), .Z(n674) );
  NAND2_X1 U758 ( .A1(G868), .A2(n674), .ZN(n675) );
  XNOR2_X1 U759 ( .A(n675), .B(KEYINPUT84), .ZN(n678) );
  OR2_X1 U760 ( .A1(n676), .A2(G868), .ZN(n677) );
  NAND2_X1 U761 ( .A1(n678), .A2(n677), .ZN(G295) );
  NAND2_X1 U762 ( .A1(G2084), .A2(G2078), .ZN(n679) );
  XOR2_X1 U763 ( .A(KEYINPUT20), .B(n679), .Z(n680) );
  NAND2_X1 U764 ( .A1(G2090), .A2(n680), .ZN(n681) );
  XNOR2_X1 U765 ( .A(KEYINPUT21), .B(n681), .ZN(n682) );
  NAND2_X1 U766 ( .A1(n682), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U767 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U768 ( .A1(G220), .A2(G219), .ZN(n683) );
  XOR2_X1 U769 ( .A(KEYINPUT22), .B(n683), .Z(n684) );
  NOR2_X1 U770 ( .A1(G218), .A2(n684), .ZN(n685) );
  NAND2_X1 U771 ( .A1(G96), .A2(n685), .ZN(n850) );
  NAND2_X1 U772 ( .A1(G2106), .A2(n850), .ZN(n689) );
  NAND2_X1 U773 ( .A1(G108), .A2(G120), .ZN(n686) );
  NOR2_X1 U774 ( .A1(G237), .A2(n686), .ZN(n687) );
  NAND2_X1 U775 ( .A1(G69), .A2(n687), .ZN(n851) );
  NAND2_X1 U776 ( .A1(G567), .A2(n851), .ZN(n688) );
  NAND2_X1 U777 ( .A1(n689), .A2(n688), .ZN(n690) );
  XOR2_X1 U778 ( .A(KEYINPUT85), .B(n690), .Z(n924) );
  NAND2_X1 U779 ( .A1(G661), .A2(G483), .ZN(n691) );
  NOR2_X1 U780 ( .A1(n924), .A2(n691), .ZN(n849) );
  NAND2_X1 U781 ( .A1(n849), .A2(G36), .ZN(G176) );
  INV_X1 U782 ( .A(KEYINPUT31), .ZN(n709) );
  XNOR2_X1 U783 ( .A(KEYINPUT98), .B(KEYINPUT99), .ZN(n692) );
  XNOR2_X1 U784 ( .A(n692), .B(KEYINPUT30), .ZN(n701) );
  NOR2_X1 U785 ( .A1(G164), .A2(G1384), .ZN(n794) );
  INV_X1 U786 ( .A(n794), .ZN(n702) );
  AND2_X1 U787 ( .A1(G40), .A2(n693), .ZN(n694) );
  NAND2_X1 U788 ( .A1(n695), .A2(n694), .ZN(n793) );
  XOR2_X1 U789 ( .A(KEYINPUT93), .B(n696), .Z(n762) );
  NAND2_X1 U790 ( .A1(G8), .A2(n741), .ZN(n788) );
  NOR2_X1 U791 ( .A1(G1966), .A2(n788), .ZN(n759) );
  NOR2_X1 U792 ( .A1(n762), .A2(n759), .ZN(n698) );
  INV_X1 U793 ( .A(KEYINPUT97), .ZN(n697) );
  XNOR2_X1 U794 ( .A(n698), .B(n697), .ZN(n699) );
  NAND2_X1 U795 ( .A1(n699), .A2(G8), .ZN(n700) );
  NOR2_X1 U796 ( .A1(G168), .A2(n517), .ZN(n707) );
  XNOR2_X1 U797 ( .A(G2078), .B(KEYINPUT25), .ZN(n957) );
  NAND2_X1 U798 ( .A1(n717), .A2(n957), .ZN(n703) );
  XNOR2_X1 U799 ( .A(n703), .B(KEYINPUT94), .ZN(n705) );
  INV_X1 U800 ( .A(G1961), .ZN(n864) );
  NAND2_X1 U801 ( .A1(n864), .A2(n741), .ZN(n704) );
  NAND2_X1 U802 ( .A1(n705), .A2(n704), .ZN(n738) );
  NOR2_X1 U803 ( .A1(G171), .A2(n738), .ZN(n706) );
  NOR2_X1 U804 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U805 ( .A(n709), .B(n708), .ZN(n757) );
  NAND2_X1 U806 ( .A1(n717), .A2(G2072), .ZN(n710) );
  XOR2_X1 U807 ( .A(KEYINPUT27), .B(n710), .Z(n712) );
  NAND2_X1 U808 ( .A1(G1956), .A2(n741), .ZN(n711) );
  NAND2_X1 U809 ( .A1(n712), .A2(n711), .ZN(n728) );
  NAND2_X1 U810 ( .A1(G299), .A2(n728), .ZN(n713) );
  XOR2_X1 U811 ( .A(KEYINPUT28), .B(n713), .Z(n736) );
  NAND2_X1 U812 ( .A1(n717), .A2(G1996), .ZN(n716) );
  NAND2_X1 U813 ( .A1(G1348), .A2(n741), .ZN(n719) );
  NAND2_X1 U814 ( .A1(G2067), .A2(n717), .ZN(n718) );
  NAND2_X1 U815 ( .A1(n719), .A2(n718), .ZN(n726) );
  NAND2_X1 U816 ( .A1(n726), .A2(n727), .ZN(n720) );
  NAND2_X1 U817 ( .A1(n721), .A2(n720), .ZN(n724) );
  NAND2_X1 U818 ( .A1(G1341), .A2(n741), .ZN(n722) );
  XNOR2_X1 U819 ( .A(KEYINPUT95), .B(n722), .ZN(n723) );
  NOR2_X1 U820 ( .A1(n724), .A2(n723), .ZN(n725) );
  NAND2_X1 U821 ( .A1(n725), .A2(n974), .ZN(n732) );
  NOR2_X1 U822 ( .A1(n727), .A2(n726), .ZN(n730) );
  NOR2_X1 U823 ( .A1(n728), .A2(G299), .ZN(n729) );
  NOR2_X1 U824 ( .A1(n730), .A2(n729), .ZN(n731) );
  NAND2_X1 U825 ( .A1(n732), .A2(n731), .ZN(n734) );
  NOR2_X1 U826 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U827 ( .A(n737), .B(KEYINPUT29), .ZN(n740) );
  NAND2_X1 U828 ( .A1(G171), .A2(n738), .ZN(n739) );
  NAND2_X1 U829 ( .A1(n740), .A2(n739), .ZN(n758) );
  INV_X1 U830 ( .A(G8), .ZN(n747) );
  NOR2_X1 U831 ( .A1(G2090), .A2(n741), .ZN(n742) );
  XNOR2_X1 U832 ( .A(KEYINPUT101), .B(n742), .ZN(n745) );
  NOR2_X1 U833 ( .A1(G1971), .A2(n788), .ZN(n743) );
  NOR2_X1 U834 ( .A1(G166), .A2(n743), .ZN(n744) );
  NAND2_X1 U835 ( .A1(n745), .A2(n744), .ZN(n746) );
  OR2_X1 U836 ( .A1(n747), .A2(n746), .ZN(n749) );
  AND2_X1 U837 ( .A1(n758), .A2(n749), .ZN(n748) );
  NAND2_X1 U838 ( .A1(n757), .A2(n748), .ZN(n753) );
  INV_X1 U839 ( .A(n749), .ZN(n751) );
  AND2_X1 U840 ( .A1(G286), .A2(G8), .ZN(n750) );
  OR2_X1 U841 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U842 ( .A1(n753), .A2(n752), .ZN(n754) );
  XNOR2_X1 U843 ( .A(n754), .B(KEYINPUT32), .ZN(n779) );
  NAND2_X1 U844 ( .A1(G1976), .A2(G288), .ZN(n980) );
  INV_X1 U845 ( .A(n788), .ZN(n755) );
  NAND2_X1 U846 ( .A1(n980), .A2(n755), .ZN(n768) );
  INV_X1 U847 ( .A(n768), .ZN(n756) );
  AND2_X1 U848 ( .A1(n779), .A2(n756), .ZN(n765) );
  AND2_X1 U849 ( .A1(n758), .A2(n757), .ZN(n760) );
  XNOR2_X1 U850 ( .A(n761), .B(KEYINPUT100), .ZN(n764) );
  NAND2_X1 U851 ( .A1(n762), .A2(G8), .ZN(n763) );
  NAND2_X1 U852 ( .A1(n764), .A2(n763), .ZN(n780) );
  NAND2_X1 U853 ( .A1(n765), .A2(n780), .ZN(n770) );
  NOR2_X1 U854 ( .A1(G1976), .A2(G288), .ZN(n978) );
  NOR2_X1 U855 ( .A1(G1971), .A2(G303), .ZN(n766) );
  NOR2_X1 U856 ( .A1(n978), .A2(n766), .ZN(n767) );
  OR2_X1 U857 ( .A1(n768), .A2(n767), .ZN(n769) );
  NAND2_X1 U858 ( .A1(n770), .A2(n769), .ZN(n771) );
  XNOR2_X1 U859 ( .A(n771), .B(KEYINPUT64), .ZN(n772) );
  INV_X1 U860 ( .A(n772), .ZN(n774) );
  NAND2_X1 U861 ( .A1(n774), .A2(n773), .ZN(n776) );
  XOR2_X1 U862 ( .A(G1981), .B(G305), .Z(n995) );
  NAND2_X1 U863 ( .A1(n978), .A2(KEYINPUT33), .ZN(n775) );
  NAND2_X1 U864 ( .A1(n776), .A2(n518), .ZN(n785) );
  NOR2_X1 U865 ( .A1(G2090), .A2(G303), .ZN(n777) );
  NAND2_X1 U866 ( .A1(G8), .A2(n777), .ZN(n778) );
  XNOR2_X1 U867 ( .A(n778), .B(KEYINPUT102), .ZN(n782) );
  NAND2_X1 U868 ( .A1(n780), .A2(n779), .ZN(n781) );
  NAND2_X1 U869 ( .A1(n782), .A2(n781), .ZN(n783) );
  NAND2_X1 U870 ( .A1(n783), .A2(n788), .ZN(n784) );
  NAND2_X1 U871 ( .A1(n785), .A2(n784), .ZN(n790) );
  NOR2_X1 U872 ( .A1(G1981), .A2(G305), .ZN(n786) );
  XOR2_X1 U873 ( .A(n786), .B(KEYINPUT24), .Z(n787) );
  NOR2_X1 U874 ( .A1(n788), .A2(n787), .ZN(n789) );
  XNOR2_X1 U875 ( .A(n792), .B(n791), .ZN(n825) );
  NOR2_X1 U876 ( .A1(n794), .A2(n793), .ZN(n841) );
  NAND2_X1 U877 ( .A1(n896), .A2(G104), .ZN(n796) );
  NAND2_X1 U878 ( .A1(G140), .A2(n897), .ZN(n795) );
  NAND2_X1 U879 ( .A1(n796), .A2(n795), .ZN(n797) );
  XNOR2_X1 U880 ( .A(KEYINPUT34), .B(n797), .ZN(n802) );
  NAND2_X1 U881 ( .A1(G116), .A2(n893), .ZN(n799) );
  NAND2_X1 U882 ( .A1(G128), .A2(n617), .ZN(n798) );
  NAND2_X1 U883 ( .A1(n799), .A2(n798), .ZN(n800) );
  XOR2_X1 U884 ( .A(n800), .B(KEYINPUT35), .Z(n801) );
  NOR2_X1 U885 ( .A1(n802), .A2(n801), .ZN(n803) );
  XOR2_X1 U886 ( .A(KEYINPUT36), .B(n803), .Z(n804) );
  XOR2_X1 U887 ( .A(KEYINPUT88), .B(n804), .Z(n905) );
  XNOR2_X1 U888 ( .A(G2067), .B(KEYINPUT37), .ZN(n839) );
  NOR2_X1 U889 ( .A1(n905), .A2(n839), .ZN(n929) );
  NAND2_X1 U890 ( .A1(n841), .A2(n929), .ZN(n837) );
  XOR2_X1 U891 ( .A(KEYINPUT90), .B(G1991), .Z(n956) );
  NAND2_X1 U892 ( .A1(n896), .A2(G95), .ZN(n807) );
  NAND2_X1 U893 ( .A1(n897), .A2(G131), .ZN(n805) );
  XOR2_X1 U894 ( .A(KEYINPUT89), .B(n805), .Z(n806) );
  NAND2_X1 U895 ( .A1(n807), .A2(n806), .ZN(n811) );
  NAND2_X1 U896 ( .A1(G107), .A2(n893), .ZN(n809) );
  NAND2_X1 U897 ( .A1(G119), .A2(n617), .ZN(n808) );
  NAND2_X1 U898 ( .A1(n809), .A2(n808), .ZN(n810) );
  NOR2_X1 U899 ( .A1(n811), .A2(n810), .ZN(n904) );
  NOR2_X1 U900 ( .A1(n956), .A2(n904), .ZN(n822) );
  XOR2_X1 U901 ( .A(KEYINPUT92), .B(KEYINPUT38), .Z(n813) );
  NAND2_X1 U902 ( .A1(G105), .A2(n896), .ZN(n812) );
  XNOR2_X1 U903 ( .A(n813), .B(n812), .ZN(n818) );
  NAND2_X1 U904 ( .A1(G117), .A2(n893), .ZN(n815) );
  NAND2_X1 U905 ( .A1(G129), .A2(n617), .ZN(n814) );
  NAND2_X1 U906 ( .A1(n815), .A2(n814), .ZN(n816) );
  XOR2_X1 U907 ( .A(KEYINPUT91), .B(n816), .Z(n817) );
  NOR2_X1 U908 ( .A1(n818), .A2(n817), .ZN(n820) );
  NAND2_X1 U909 ( .A1(G141), .A2(n897), .ZN(n819) );
  NAND2_X1 U910 ( .A1(n820), .A2(n819), .ZN(n911) );
  AND2_X1 U911 ( .A1(n911), .A2(G1996), .ZN(n821) );
  NOR2_X1 U912 ( .A1(n822), .A2(n821), .ZN(n931) );
  INV_X1 U913 ( .A(n931), .ZN(n823) );
  NAND2_X1 U914 ( .A1(n823), .A2(n841), .ZN(n830) );
  NAND2_X1 U915 ( .A1(n837), .A2(n830), .ZN(n824) );
  NOR2_X1 U916 ( .A1(n825), .A2(n824), .ZN(n828) );
  XOR2_X1 U917 ( .A(G1986), .B(G290), .Z(n826) );
  XNOR2_X1 U918 ( .A(KEYINPUT87), .B(n826), .ZN(n987) );
  NAND2_X1 U919 ( .A1(n987), .A2(n841), .ZN(n827) );
  NAND2_X1 U920 ( .A1(n828), .A2(n827), .ZN(n844) );
  NOR2_X1 U921 ( .A1(n911), .A2(G1996), .ZN(n829) );
  XNOR2_X1 U922 ( .A(n829), .B(KEYINPUT104), .ZN(n926) );
  INV_X1 U923 ( .A(n830), .ZN(n833) );
  NOR2_X1 U924 ( .A1(G1986), .A2(G290), .ZN(n831) );
  AND2_X1 U925 ( .A1(n956), .A2(n904), .ZN(n936) );
  NOR2_X1 U926 ( .A1(n831), .A2(n936), .ZN(n832) );
  NOR2_X1 U927 ( .A1(n833), .A2(n832), .ZN(n834) );
  XOR2_X1 U928 ( .A(KEYINPUT105), .B(n834), .Z(n835) );
  NOR2_X1 U929 ( .A1(n926), .A2(n835), .ZN(n836) );
  XNOR2_X1 U930 ( .A(KEYINPUT39), .B(n836), .ZN(n838) );
  NAND2_X1 U931 ( .A1(n838), .A2(n837), .ZN(n840) );
  NAND2_X1 U932 ( .A1(n905), .A2(n839), .ZN(n930) );
  NAND2_X1 U933 ( .A1(n840), .A2(n930), .ZN(n842) );
  NAND2_X1 U934 ( .A1(n842), .A2(n841), .ZN(n843) );
  NAND2_X1 U935 ( .A1(n844), .A2(n843), .ZN(n845) );
  XNOR2_X1 U936 ( .A(n845), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U937 ( .A1(G2106), .A2(n846), .ZN(G217) );
  INV_X1 U938 ( .A(n846), .ZN(G223) );
  AND2_X1 U939 ( .A1(G15), .A2(G2), .ZN(n847) );
  NAND2_X1 U940 ( .A1(G661), .A2(n847), .ZN(G259) );
  NAND2_X1 U941 ( .A1(G3), .A2(G1), .ZN(n848) );
  NAND2_X1 U942 ( .A1(n849), .A2(n848), .ZN(G188) );
  XOR2_X1 U943 ( .A(G120), .B(KEYINPUT108), .Z(G236) );
  INV_X1 U945 ( .A(G108), .ZN(G238) );
  INV_X1 U946 ( .A(G96), .ZN(G221) );
  NOR2_X1 U947 ( .A1(n851), .A2(n850), .ZN(G325) );
  INV_X1 U948 ( .A(G325), .ZN(G261) );
  XOR2_X1 U949 ( .A(G286), .B(G171), .Z(n852) );
  XOR2_X1 U950 ( .A(n852), .B(n991), .Z(n854) );
  XNOR2_X1 U951 ( .A(n854), .B(n853), .ZN(n855) );
  NOR2_X1 U952 ( .A1(G37), .A2(n855), .ZN(G397) );
  XOR2_X1 U953 ( .A(G2100), .B(G2096), .Z(n857) );
  XNOR2_X1 U954 ( .A(KEYINPUT42), .B(G2678), .ZN(n856) );
  XNOR2_X1 U955 ( .A(n857), .B(n856), .ZN(n861) );
  XOR2_X1 U956 ( .A(KEYINPUT43), .B(G2090), .Z(n859) );
  XNOR2_X1 U957 ( .A(G2067), .B(G2072), .ZN(n858) );
  XNOR2_X1 U958 ( .A(n859), .B(n858), .ZN(n860) );
  XOR2_X1 U959 ( .A(n861), .B(n860), .Z(n863) );
  XNOR2_X1 U960 ( .A(G2084), .B(G2078), .ZN(n862) );
  XNOR2_X1 U961 ( .A(n863), .B(n862), .ZN(G227) );
  XNOR2_X1 U962 ( .A(G1981), .B(n864), .ZN(n866) );
  XNOR2_X1 U963 ( .A(G1996), .B(G1966), .ZN(n865) );
  XNOR2_X1 U964 ( .A(n866), .B(n865), .ZN(n870) );
  XOR2_X1 U965 ( .A(G1976), .B(G1971), .Z(n868) );
  XNOR2_X1 U966 ( .A(G1986), .B(G1956), .ZN(n867) );
  XNOR2_X1 U967 ( .A(n868), .B(n867), .ZN(n869) );
  XOR2_X1 U968 ( .A(n870), .B(n869), .Z(n872) );
  XNOR2_X1 U969 ( .A(KEYINPUT109), .B(KEYINPUT41), .ZN(n871) );
  XNOR2_X1 U970 ( .A(n872), .B(n871), .ZN(n874) );
  XOR2_X1 U971 ( .A(G1991), .B(G2474), .Z(n873) );
  XNOR2_X1 U972 ( .A(n874), .B(n873), .ZN(G229) );
  NAND2_X1 U973 ( .A1(G124), .A2(n617), .ZN(n875) );
  XNOR2_X1 U974 ( .A(n875), .B(KEYINPUT44), .ZN(n876) );
  XNOR2_X1 U975 ( .A(KEYINPUT110), .B(n876), .ZN(n879) );
  NAND2_X1 U976 ( .A1(n897), .A2(G136), .ZN(n877) );
  XOR2_X1 U977 ( .A(KEYINPUT111), .B(n877), .Z(n878) );
  NAND2_X1 U978 ( .A1(n879), .A2(n878), .ZN(n883) );
  NAND2_X1 U979 ( .A1(G112), .A2(n893), .ZN(n881) );
  NAND2_X1 U980 ( .A1(G100), .A2(n896), .ZN(n880) );
  NAND2_X1 U981 ( .A1(n881), .A2(n880), .ZN(n882) );
  NOR2_X1 U982 ( .A1(n883), .A2(n882), .ZN(G162) );
  NAND2_X1 U983 ( .A1(G115), .A2(n893), .ZN(n885) );
  NAND2_X1 U984 ( .A1(G127), .A2(n617), .ZN(n884) );
  NAND2_X1 U985 ( .A1(n885), .A2(n884), .ZN(n886) );
  XNOR2_X1 U986 ( .A(KEYINPUT47), .B(n886), .ZN(n892) );
  NAND2_X1 U987 ( .A1(n897), .A2(G139), .ZN(n887) );
  XOR2_X1 U988 ( .A(KEYINPUT114), .B(n887), .Z(n890) );
  NAND2_X1 U989 ( .A1(G103), .A2(n896), .ZN(n888) );
  XNOR2_X1 U990 ( .A(KEYINPUT113), .B(n888), .ZN(n889) );
  NOR2_X1 U991 ( .A1(n890), .A2(n889), .ZN(n891) );
  NAND2_X1 U992 ( .A1(n892), .A2(n891), .ZN(n942) );
  NAND2_X1 U993 ( .A1(G118), .A2(n893), .ZN(n895) );
  NAND2_X1 U994 ( .A1(G130), .A2(n617), .ZN(n894) );
  NAND2_X1 U995 ( .A1(n895), .A2(n894), .ZN(n903) );
  NAND2_X1 U996 ( .A1(n896), .A2(G106), .ZN(n899) );
  NAND2_X1 U997 ( .A1(G142), .A2(n897), .ZN(n898) );
  NAND2_X1 U998 ( .A1(n899), .A2(n898), .ZN(n900) );
  XOR2_X1 U999 ( .A(KEYINPUT112), .B(n900), .Z(n901) );
  XNOR2_X1 U1000 ( .A(KEYINPUT45), .B(n901), .ZN(n902) );
  NOR2_X1 U1001 ( .A1(n903), .A2(n902), .ZN(n909) );
  XOR2_X1 U1002 ( .A(G162), .B(n904), .Z(n907) );
  XNOR2_X1 U1003 ( .A(G160), .B(n905), .ZN(n906) );
  XNOR2_X1 U1004 ( .A(n907), .B(n906), .ZN(n908) );
  XOR2_X1 U1005 ( .A(n909), .B(n908), .Z(n910) );
  XNOR2_X1 U1006 ( .A(n942), .B(n910), .ZN(n916) );
  XOR2_X1 U1007 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n913) );
  XOR2_X1 U1008 ( .A(G164), .B(n911), .Z(n912) );
  XNOR2_X1 U1009 ( .A(n913), .B(n912), .ZN(n914) );
  XOR2_X1 U1010 ( .A(n933), .B(n914), .Z(n915) );
  XNOR2_X1 U1011 ( .A(n916), .B(n915), .ZN(n917) );
  NOR2_X1 U1012 ( .A1(G37), .A2(n917), .ZN(G395) );
  NOR2_X1 U1013 ( .A1(G401), .A2(n924), .ZN(n921) );
  NOR2_X1 U1014 ( .A1(G227), .A2(G229), .ZN(n918) );
  XNOR2_X1 U1015 ( .A(KEYINPUT49), .B(n918), .ZN(n919) );
  NOR2_X1 U1016 ( .A1(G397), .A2(n919), .ZN(n920) );
  NAND2_X1 U1017 ( .A1(n921), .A2(n920), .ZN(n922) );
  NOR2_X1 U1018 ( .A1(n922), .A2(G395), .ZN(n923) );
  XOR2_X1 U1019 ( .A(n923), .B(KEYINPUT115), .Z(G308) );
  INV_X1 U1020 ( .A(G308), .ZN(G225) );
  INV_X1 U1021 ( .A(n924), .ZN(G319) );
  INV_X1 U1022 ( .A(G69), .ZN(G235) );
  XOR2_X1 U1023 ( .A(G2090), .B(G162), .Z(n925) );
  NOR2_X1 U1024 ( .A1(n926), .A2(n925), .ZN(n927) );
  XNOR2_X1 U1025 ( .A(n927), .B(KEYINPUT51), .ZN(n928) );
  NOR2_X1 U1026 ( .A1(n929), .A2(n928), .ZN(n941) );
  NAND2_X1 U1027 ( .A1(n931), .A2(n930), .ZN(n939) );
  XNOR2_X1 U1028 ( .A(G160), .B(G2084), .ZN(n932) );
  XNOR2_X1 U1029 ( .A(n932), .B(KEYINPUT116), .ZN(n934) );
  NAND2_X1 U1030 ( .A1(n934), .A2(n933), .ZN(n935) );
  NOR2_X1 U1031 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1032 ( .A(KEYINPUT117), .B(n937), .ZN(n938) );
  NOR2_X1 U1033 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1034 ( .A1(n941), .A2(n940), .ZN(n948) );
  XOR2_X1 U1035 ( .A(G164), .B(G2078), .Z(n945) );
  XNOR2_X1 U1036 ( .A(KEYINPUT118), .B(n942), .ZN(n943) );
  XNOR2_X1 U1037 ( .A(G2072), .B(n943), .ZN(n944) );
  NOR2_X1 U1038 ( .A1(n945), .A2(n944), .ZN(n946) );
  XOR2_X1 U1039 ( .A(KEYINPUT50), .B(n946), .Z(n947) );
  NOR2_X1 U1040 ( .A1(n948), .A2(n947), .ZN(n949) );
  XOR2_X1 U1041 ( .A(KEYINPUT52), .B(n949), .Z(n950) );
  NOR2_X1 U1042 ( .A1(KEYINPUT55), .A2(n950), .ZN(n951) );
  XNOR2_X1 U1043 ( .A(KEYINPUT119), .B(n951), .ZN(n952) );
  NAND2_X1 U1044 ( .A1(n952), .A2(G29), .ZN(n1033) );
  XNOR2_X1 U1045 ( .A(G2067), .B(G26), .ZN(n954) );
  XNOR2_X1 U1046 ( .A(G33), .B(G2072), .ZN(n953) );
  NOR2_X1 U1047 ( .A1(n954), .A2(n953), .ZN(n963) );
  XOR2_X1 U1048 ( .A(G32), .B(G1996), .Z(n955) );
  NAND2_X1 U1049 ( .A1(n955), .A2(G28), .ZN(n961) );
  XNOR2_X1 U1050 ( .A(n956), .B(G25), .ZN(n959) );
  XNOR2_X1 U1051 ( .A(n957), .B(G27), .ZN(n958) );
  NAND2_X1 U1052 ( .A1(n959), .A2(n958), .ZN(n960) );
  NOR2_X1 U1053 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1054 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1055 ( .A(n964), .B(KEYINPUT53), .ZN(n967) );
  XOR2_X1 U1056 ( .A(G2084), .B(G34), .Z(n965) );
  XNOR2_X1 U1057 ( .A(KEYINPUT54), .B(n965), .ZN(n966) );
  NAND2_X1 U1058 ( .A1(n967), .A2(n966), .ZN(n969) );
  XNOR2_X1 U1059 ( .A(G35), .B(G2090), .ZN(n968) );
  NOR2_X1 U1060 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1061 ( .A(KEYINPUT55), .B(n970), .ZN(n972) );
  INV_X1 U1062 ( .A(G29), .ZN(n971) );
  NAND2_X1 U1063 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1064 ( .A1(n973), .A2(G11), .ZN(n1031) );
  INV_X1 U1065 ( .A(G16), .ZN(n1027) );
  XOR2_X1 U1066 ( .A(n1027), .B(KEYINPUT56), .Z(n1002) );
  XOR2_X1 U1067 ( .A(n974), .B(G1341), .Z(n976) );
  XNOR2_X1 U1068 ( .A(G301), .B(G1961), .ZN(n975) );
  NOR2_X1 U1069 ( .A1(n976), .A2(n975), .ZN(n990) );
  XOR2_X1 U1070 ( .A(G1971), .B(G303), .Z(n977) );
  XNOR2_X1 U1071 ( .A(n977), .B(KEYINPUT122), .ZN(n985) );
  INV_X1 U1072 ( .A(n978), .ZN(n979) );
  NAND2_X1 U1073 ( .A1(n980), .A2(n979), .ZN(n981) );
  XOR2_X1 U1074 ( .A(KEYINPUT121), .B(n981), .Z(n983) );
  XNOR2_X1 U1075 ( .A(G1956), .B(G299), .ZN(n982) );
  NOR2_X1 U1076 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1077 ( .A1(n985), .A2(n984), .ZN(n986) );
  NOR2_X1 U1078 ( .A1(n987), .A2(n986), .ZN(n988) );
  XOR2_X1 U1079 ( .A(KEYINPUT123), .B(n988), .Z(n989) );
  NAND2_X1 U1080 ( .A1(n990), .A2(n989), .ZN(n994) );
  XOR2_X1 U1081 ( .A(G1348), .B(n991), .Z(n992) );
  XNOR2_X1 U1082 ( .A(KEYINPUT120), .B(n992), .ZN(n993) );
  NOR2_X1 U1083 ( .A1(n994), .A2(n993), .ZN(n999) );
  XNOR2_X1 U1084 ( .A(G1966), .B(G168), .ZN(n996) );
  NAND2_X1 U1085 ( .A1(n996), .A2(n995), .ZN(n997) );
  XNOR2_X1 U1086 ( .A(n997), .B(KEYINPUT57), .ZN(n998) );
  NAND2_X1 U1087 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XNOR2_X1 U1088 ( .A(n1000), .B(KEYINPUT124), .ZN(n1001) );
  NAND2_X1 U1089 ( .A1(n1002), .A2(n1001), .ZN(n1029) );
  XOR2_X1 U1090 ( .A(KEYINPUT127), .B(KEYINPUT58), .Z(n1009) );
  XNOR2_X1 U1091 ( .A(G1986), .B(G24), .ZN(n1004) );
  XNOR2_X1 U1092 ( .A(G23), .B(G1976), .ZN(n1003) );
  NOR2_X1 U1093 ( .A1(n1004), .A2(n1003), .ZN(n1007) );
  XOR2_X1 U1094 ( .A(G1971), .B(KEYINPUT126), .Z(n1005) );
  XNOR2_X1 U1095 ( .A(G22), .B(n1005), .ZN(n1006) );
  NAND2_X1 U1096 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1097 ( .A(n1009), .B(n1008), .ZN(n1024) );
  XOR2_X1 U1098 ( .A(G5), .B(G1961), .Z(n1022) );
  XNOR2_X1 U1099 ( .A(G1348), .B(KEYINPUT59), .ZN(n1010) );
  XNOR2_X1 U1100 ( .A(n1010), .B(G4), .ZN(n1014) );
  XNOR2_X1 U1101 ( .A(G1341), .B(G19), .ZN(n1012) );
  XNOR2_X1 U1102 ( .A(G20), .B(G1956), .ZN(n1011) );
  NOR2_X1 U1103 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1104 ( .A1(n1014), .A2(n1013), .ZN(n1017) );
  XOR2_X1 U1105 ( .A(KEYINPUT125), .B(G1981), .Z(n1015) );
  XNOR2_X1 U1106 ( .A(G6), .B(n1015), .ZN(n1016) );
  NOR2_X1 U1107 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XOR2_X1 U1108 ( .A(KEYINPUT60), .B(n1018), .Z(n1020) );
  XNOR2_X1 U1109 ( .A(G1966), .B(G21), .ZN(n1019) );
  NOR2_X1 U1110 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1111 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NOR2_X1 U1112 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XNOR2_X1 U1113 ( .A(KEYINPUT61), .B(n1025), .ZN(n1026) );
  NAND2_X1 U1114 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NAND2_X1 U1115 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NOR2_X1 U1116 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  NAND2_X1 U1117 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  XNOR2_X1 U1118 ( .A(KEYINPUT62), .B(n1034), .ZN(G150) );
  INV_X1 U1119 ( .A(G150), .ZN(G311) );
endmodule

