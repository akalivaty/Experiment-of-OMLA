//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 1 1 0 0 0 0 0 0 0 0 0 1 1 1 1 1 1 1 0 0 0 0 0 1 0 0 1 0 1 0 1 0 0 0 0 0 1 0 1 1 1 0 0 0 1 0 0 1 0 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:16 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n682,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n699, new_n701, new_n702, new_n703, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n713, new_n714, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n919,
    new_n920, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001;
  NOR2_X1   g000(.A1(G237), .A2(G953), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G210), .ZN(new_n188));
  XOR2_X1   g002(.A(new_n188), .B(KEYINPUT27), .Z(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT26), .B(G101), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n189), .B(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT2), .B(G113), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  XNOR2_X1  g007(.A(G116), .B(G119), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(new_n194), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(new_n192), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G137), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n199), .A2(KEYINPUT11), .A3(G134), .ZN(new_n200));
  INV_X1    g014(.A(G134), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G137), .ZN(new_n202));
  AND2_X1   g016(.A1(new_n200), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT64), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n199), .A2(G134), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT11), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n204), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  AOI211_X1 g021(.A(KEYINPUT64), .B(KEYINPUT11), .C1(new_n199), .C2(G134), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n203), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G131), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT65), .ZN(new_n211));
  INV_X1    g025(.A(G131), .ZN(new_n212));
  OAI211_X1 g026(.A(new_n203), .B(new_n212), .C1(new_n207), .C2(new_n208), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n210), .A2(new_n211), .A3(new_n213), .ZN(new_n214));
  XNOR2_X1  g028(.A(G143), .B(G146), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n215), .A2(KEYINPUT0), .A3(G128), .ZN(new_n216));
  XNOR2_X1  g030(.A(KEYINPUT0), .B(G128), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n216), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n209), .A2(KEYINPUT65), .A3(G131), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n214), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT30), .ZN(new_n222));
  INV_X1    g036(.A(G146), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(G143), .ZN(new_n224));
  INV_X1    g038(.A(G143), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(G146), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n224), .A2(KEYINPUT1), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n227), .A2(new_n228), .A3(G128), .ZN(new_n229));
  INV_X1    g043(.A(G128), .ZN(new_n230));
  OAI211_X1 g044(.A(new_n224), .B(new_n226), .C1(KEYINPUT1), .C2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n205), .A2(new_n202), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(G131), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n233), .A2(new_n213), .A3(new_n235), .ZN(new_n236));
  AND3_X1   g050(.A1(new_n221), .A2(new_n222), .A3(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n213), .A2(new_n235), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT66), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n213), .A2(KEYINPUT66), .A3(new_n235), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n240), .A2(new_n241), .A3(new_n233), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n222), .B1(new_n242), .B2(new_n221), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n198), .B1(new_n237), .B2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(new_n198), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n242), .A2(new_n221), .A3(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(KEYINPUT67), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n244), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT67), .ZN(new_n250));
  OAI211_X1 g064(.A(new_n250), .B(new_n198), .C1(new_n237), .C2(new_n243), .ZN(new_n251));
  AOI211_X1 g065(.A(KEYINPUT31), .B(new_n191), .C1(new_n249), .C2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT31), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n242), .A2(new_n221), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(KEYINPUT30), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n221), .A2(new_n222), .A3(new_n236), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n245), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n251), .B1(new_n257), .B2(new_n247), .ZN(new_n258));
  INV_X1    g072(.A(new_n191), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n253), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n252), .A2(new_n260), .ZN(new_n261));
  AND3_X1   g075(.A1(new_n242), .A2(new_n221), .A3(new_n245), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n245), .B1(new_n221), .B2(new_n236), .ZN(new_n263));
  OAI21_X1  g077(.A(KEYINPUT28), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  OAI21_X1  g078(.A(KEYINPUT68), .B1(new_n262), .B2(KEYINPUT28), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT68), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT28), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n246), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n264), .A2(new_n265), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(new_n191), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT69), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n269), .A2(KEYINPUT69), .A3(new_n191), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  AOI21_X1  g088(.A(G902), .B1(new_n261), .B2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(G472), .ZN(new_n276));
  AOI21_X1  g090(.A(KEYINPUT32), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT29), .ZN(new_n278));
  AND3_X1   g092(.A1(new_n246), .A2(new_n266), .A3(new_n267), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n266), .B1(new_n246), .B2(new_n267), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n191), .B1(new_n281), .B2(new_n264), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n259), .B1(new_n249), .B2(new_n251), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n278), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n245), .B1(new_n242), .B2(new_n221), .ZN(new_n285));
  OAI21_X1  g099(.A(KEYINPUT28), .B1(new_n262), .B2(new_n285), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n191), .A2(new_n278), .ZN(new_n287));
  NAND4_X1  g101(.A1(new_n286), .A2(new_n265), .A3(new_n268), .A4(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT70), .ZN(new_n289));
  INV_X1    g103(.A(G902), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n288), .A2(new_n290), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(KEYINPUT70), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n284), .A2(new_n291), .A3(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(G472), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT32), .ZN(new_n296));
  NOR3_X1   g110(.A1(new_n296), .A2(G472), .A3(G902), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n258), .A2(new_n259), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(KEYINPUT31), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n258), .A2(new_n253), .A3(new_n259), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  AND3_X1   g115(.A1(new_n269), .A2(KEYINPUT69), .A3(new_n191), .ZN(new_n302));
  AOI21_X1  g116(.A(KEYINPUT69), .B1(new_n269), .B2(new_n191), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n297), .B1(new_n301), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n295), .A2(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(KEYINPUT71), .B1(new_n277), .B2(new_n306), .ZN(new_n307));
  OAI211_X1 g121(.A(new_n276), .B(new_n290), .C1(new_n301), .C2(new_n304), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(new_n296), .ZN(new_n309));
  OAI211_X1 g123(.A(new_n299), .B(new_n300), .C1(new_n303), .C2(new_n302), .ZN(new_n310));
  AOI22_X1  g124(.A1(G472), .A2(new_n294), .B1(new_n310), .B2(new_n297), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT71), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n309), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(G140), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(G125), .ZN(new_n315));
  INV_X1    g129(.A(G125), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(G140), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT74), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n315), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n316), .A2(G140), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(KEYINPUT74), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(KEYINPUT16), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT75), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n324), .B1(new_n315), .B2(KEYINPUT16), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n323), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n322), .A2(KEYINPUT75), .A3(KEYINPUT16), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n327), .A2(new_n223), .A3(new_n328), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n325), .B1(new_n322), .B2(KEYINPUT16), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT16), .ZN(new_n331));
  AOI211_X1 g145(.A(new_n324), .B(new_n331), .C1(new_n319), .C2(new_n321), .ZN(new_n332));
  OAI21_X1  g146(.A(G146), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n329), .A2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(G110), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n230), .A2(G119), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n230), .A2(G119), .ZN(new_n337));
  NAND2_X1  g151(.A1(KEYINPUT72), .A2(KEYINPUT23), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n336), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(new_n338), .ZN(new_n340));
  NOR2_X1   g154(.A1(KEYINPUT72), .A2(KEYINPUT23), .ZN(new_n341));
  OAI211_X1 g155(.A(G119), .B(new_n230), .C1(new_n340), .C2(new_n341), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n335), .B1(new_n339), .B2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(new_n336), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(new_n337), .ZN(new_n345));
  XNOR2_X1  g159(.A(KEYINPUT24), .B(G110), .ZN(new_n346));
  OAI22_X1  g160(.A1(new_n343), .A2(KEYINPUT73), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  AND2_X1   g161(.A1(new_n343), .A2(KEYINPUT73), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n334), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(G953), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n351), .A2(G221), .A3(G234), .ZN(new_n352));
  XNOR2_X1  g166(.A(new_n352), .B(KEYINPUT77), .ZN(new_n353));
  XOR2_X1   g167(.A(KEYINPUT22), .B(G137), .Z(new_n354));
  XNOR2_X1  g168(.A(new_n353), .B(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n339), .A2(new_n342), .A3(new_n335), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n345), .A2(new_n346), .ZN(new_n357));
  XNOR2_X1  g171(.A(G125), .B(G140), .ZN(new_n358));
  AOI22_X1  g172(.A1(new_n356), .A2(new_n357), .B1(new_n223), .B2(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n333), .A2(KEYINPUT76), .A3(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  AOI21_X1  g175(.A(KEYINPUT76), .B1(new_n333), .B2(new_n359), .ZN(new_n362));
  OAI211_X1 g176(.A(new_n350), .B(new_n355), .C1(new_n361), .C2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n362), .ZN(new_n364));
  AOI22_X1  g178(.A1(new_n364), .A2(new_n360), .B1(new_n334), .B2(new_n349), .ZN(new_n365));
  XNOR2_X1  g179(.A(new_n355), .B(KEYINPUT78), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  OAI211_X1 g181(.A(new_n363), .B(new_n290), .C1(new_n365), .C2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT25), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n350), .B1(new_n361), .B2(new_n362), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(new_n366), .ZN(new_n372));
  NAND4_X1  g186(.A1(new_n372), .A2(KEYINPUT25), .A3(new_n290), .A4(new_n363), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n370), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(G217), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n375), .B1(G234), .B2(new_n290), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(KEYINPUT79), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT79), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n374), .A2(new_n379), .A3(new_n376), .ZN(new_n380));
  AND2_X1   g194(.A1(new_n372), .A2(new_n363), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n376), .A2(G902), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n378), .A2(new_n380), .A3(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  NOR2_X1   g199(.A1(G475), .A2(G902), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(G237), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n388), .A2(new_n351), .A3(G214), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n389), .A2(KEYINPUT87), .A3(new_n225), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n225), .A2(KEYINPUT87), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n391), .A2(G214), .A3(new_n187), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n393), .A2(KEYINPUT18), .A3(G131), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n358), .A2(new_n223), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n395), .B1(new_n322), .B2(new_n223), .ZN(new_n396));
  NAND2_X1  g210(.A1(KEYINPUT18), .A2(G131), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n390), .A2(new_n397), .A3(new_n392), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n394), .A2(new_n396), .A3(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  XNOR2_X1  g214(.A(new_n393), .B(G131), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n401), .A2(KEYINPUT17), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n393), .A2(KEYINPUT17), .A3(G131), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n329), .A2(new_n333), .A3(new_n403), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n402), .B1(new_n404), .B2(KEYINPUT89), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT89), .ZN(new_n406));
  NAND4_X1  g220(.A1(new_n329), .A2(new_n333), .A3(new_n406), .A4(new_n403), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n400), .B1(new_n405), .B2(new_n407), .ZN(new_n408));
  XNOR2_X1  g222(.A(G113), .B(G122), .ZN(new_n409));
  XNOR2_X1  g223(.A(KEYINPUT88), .B(G104), .ZN(new_n410));
  XOR2_X1   g224(.A(new_n409), .B(new_n410), .Z(new_n411));
  NAND2_X1  g225(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n358), .A2(KEYINPUT19), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n413), .B1(new_n322), .B2(KEYINPUT19), .ZN(new_n414));
  OAI211_X1 g228(.A(new_n333), .B(new_n401), .C1(G146), .C2(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n411), .B1(new_n415), .B2(new_n399), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  AOI211_X1 g231(.A(KEYINPUT20), .B(new_n387), .C1(new_n412), .C2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT90), .ZN(new_n420));
  INV_X1    g234(.A(new_n411), .ZN(new_n421));
  AOI211_X1 g235(.A(new_n400), .B(new_n421), .C1(new_n405), .C2(new_n407), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n420), .B1(new_n422), .B2(new_n416), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n412), .A2(KEYINPUT90), .A3(new_n417), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n387), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT20), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n419), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n408), .A2(new_n411), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n290), .B1(new_n428), .B2(new_n422), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(G475), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n225), .A2(G128), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n230), .A2(G143), .ZN(new_n432));
  AND2_X1   g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  XNOR2_X1  g247(.A(new_n433), .B(new_n201), .ZN(new_n434));
  INV_X1    g248(.A(G116), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n435), .A2(KEYINPUT14), .A3(G122), .ZN(new_n436));
  XNOR2_X1  g250(.A(G116), .B(G122), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  OAI211_X1 g252(.A(G107), .B(new_n436), .C1(new_n438), .C2(KEYINPUT14), .ZN(new_n439));
  OAI211_X1 g253(.A(new_n434), .B(new_n439), .C1(G107), .C2(new_n438), .ZN(new_n440));
  INV_X1    g254(.A(new_n431), .ZN(new_n441));
  AND2_X1   g255(.A1(new_n441), .A2(KEYINPUT13), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n432), .B1(new_n441), .B2(KEYINPUT13), .ZN(new_n443));
  OAI21_X1  g257(.A(G134), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n433), .A2(new_n201), .ZN(new_n445));
  INV_X1    g259(.A(G107), .ZN(new_n446));
  XNOR2_X1  g260(.A(new_n437), .B(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n444), .A2(new_n445), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n440), .A2(new_n448), .ZN(new_n449));
  XNOR2_X1  g263(.A(KEYINPUT9), .B(G234), .ZN(new_n450));
  NOR3_X1   g264(.A1(new_n450), .A2(new_n375), .A3(G953), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n449), .B(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(new_n290), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(KEYINPUT91), .ZN(new_n455));
  INV_X1    g269(.A(G478), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n456), .A2(KEYINPUT15), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT91), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n453), .A2(new_n458), .A3(new_n290), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n455), .A2(new_n457), .A3(new_n459), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n457), .B(KEYINPUT92), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n453), .A2(new_n290), .A3(new_n461), .ZN(new_n462));
  OR2_X1    g276(.A1(new_n462), .A2(KEYINPUT93), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(KEYINPUT93), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n460), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(G234), .A2(G237), .ZN(new_n467));
  AND3_X1   g281(.A1(new_n467), .A2(G952), .A3(new_n351), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n467), .A2(G902), .A3(G953), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n469), .B(KEYINPUT94), .ZN(new_n470));
  XNOR2_X1  g284(.A(KEYINPUT21), .B(G898), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n468), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n427), .A2(new_n430), .A3(new_n466), .A4(new_n473), .ZN(new_n474));
  OAI21_X1  g288(.A(G221), .B1(new_n450), .B2(G902), .ZN(new_n475));
  OAI21_X1  g289(.A(G214), .B1(G237), .B2(G902), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  OAI21_X1  g291(.A(G210), .B1(G237), .B2(G902), .ZN(new_n478));
  XNOR2_X1  g292(.A(G110), .B(G122), .ZN(new_n479));
  XOR2_X1   g293(.A(new_n479), .B(KEYINPUT8), .Z(new_n480));
  INV_X1    g294(.A(G104), .ZN(new_n481));
  OAI21_X1  g295(.A(KEYINPUT3), .B1(new_n481), .B2(G107), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT3), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n483), .A2(new_n446), .A3(G104), .ZN(new_n484));
  INV_X1    g298(.A(G101), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n481), .A2(G107), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n482), .A2(new_n484), .A3(new_n485), .A4(new_n486), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n446), .A2(G104), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n481), .A2(G107), .ZN(new_n489));
  OAI21_X1  g303(.A(G101), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n487), .A2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n194), .A2(KEYINPUT5), .ZN(new_n493));
  INV_X1    g307(.A(G119), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(G116), .ZN(new_n495));
  OAI211_X1 g309(.A(new_n493), .B(G113), .C1(KEYINPUT5), .C2(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n492), .B1(new_n195), .B2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT86), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n480), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n496), .A2(new_n195), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(new_n491), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n492), .A2(new_n496), .A3(new_n195), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n501), .A2(new_n502), .A3(KEYINPUT86), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n499), .A2(new_n503), .ZN(new_n504));
  OAI211_X1 g318(.A(new_n216), .B(G125), .C1(new_n215), .C2(new_n217), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n505), .B1(G125), .B2(new_n232), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n351), .A2(G224), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(KEYINPUT7), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n506), .B(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n482), .A2(new_n484), .A3(new_n486), .ZN(new_n510));
  AND2_X1   g324(.A1(new_n510), .A2(G101), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT4), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n487), .A2(KEYINPUT4), .ZN(new_n514));
  OAI211_X1 g328(.A(new_n513), .B(new_n198), .C1(new_n511), .C2(new_n514), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n491), .A2(KEYINPUT81), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT81), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n517), .B1(new_n487), .B2(new_n490), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  OAI211_X1 g333(.A(new_n515), .B(new_n479), .C1(new_n519), .C2(new_n500), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n504), .A2(new_n509), .A3(new_n520), .ZN(new_n521));
  AND2_X1   g335(.A1(new_n521), .A2(new_n290), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n515), .B1(new_n519), .B2(new_n500), .ZN(new_n523));
  INV_X1    g337(.A(new_n479), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n525), .A2(KEYINPUT6), .A3(new_n520), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n507), .B(KEYINPUT85), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n506), .B(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT6), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n523), .A2(new_n529), .A3(new_n524), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n526), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n478), .B1(new_n522), .B2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n522), .A2(new_n531), .A3(new_n478), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n477), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  XOR2_X1   g349(.A(G110), .B(G140), .Z(new_n536));
  XNOR2_X1  g350(.A(new_n536), .B(KEYINPUT80), .ZN(new_n537));
  AND2_X1   g351(.A1(new_n351), .A2(G227), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n537), .B(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n214), .A2(new_n220), .ZN(new_n541));
  OAI211_X1 g355(.A(new_n219), .B(new_n513), .C1(new_n511), .C2(new_n514), .ZN(new_n542));
  OAI211_X1 g356(.A(KEYINPUT10), .B(new_n233), .C1(new_n516), .C2(new_n518), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT10), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n544), .B1(new_n232), .B2(new_n491), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n541), .A2(new_n542), .A3(new_n543), .A4(new_n545), .ZN(new_n546));
  AND2_X1   g360(.A1(new_n214), .A2(new_n220), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT82), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n548), .B1(new_n232), .B2(new_n491), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n232), .A2(new_n491), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n232), .A2(new_n491), .A3(new_n548), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n547), .A2(new_n553), .A3(KEYINPUT12), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(KEYINPUT12), .B1(new_n547), .B2(new_n553), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n546), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(KEYINPUT83), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n547), .A2(new_n553), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT12), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(new_n554), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT83), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n562), .A2(new_n563), .A3(new_n546), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n540), .B1(new_n558), .B2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(G469), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n542), .A2(new_n543), .A3(new_n545), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(new_n547), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n568), .A2(new_n540), .A3(new_n546), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  NOR3_X1   g384(.A1(new_n565), .A2(new_n566), .A3(new_n570), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n540), .B1(new_n568), .B2(new_n546), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(KEYINPUT84), .ZN(new_n573));
  OAI211_X1 g387(.A(new_n540), .B(new_n546), .C1(new_n555), .C2(new_n556), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n572), .A2(KEYINPUT84), .ZN(new_n576));
  OAI211_X1 g390(.A(new_n566), .B(new_n290), .C1(new_n575), .C2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(G469), .A2(G902), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  OAI211_X1 g393(.A(new_n475), .B(new_n535), .C1(new_n571), .C2(new_n579), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n474), .A2(new_n580), .ZN(new_n581));
  NAND4_X1  g395(.A1(new_n307), .A2(new_n313), .A3(new_n385), .A4(new_n581), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n582), .B(G101), .ZN(G3));
  OAI21_X1  g397(.A(new_n475), .B1(new_n571), .B2(new_n579), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n584), .A2(new_n384), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n310), .A2(new_n290), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(G472), .ZN(new_n587));
  AND2_X1   g401(.A1(new_n453), .A2(KEYINPUT33), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n453), .A2(KEYINPUT33), .ZN(new_n589));
  OAI211_X1 g403(.A(G478), .B(new_n290), .C1(new_n588), .C2(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n455), .A2(new_n456), .A3(new_n459), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n593), .B1(new_n427), .B2(new_n430), .ZN(new_n594));
  NAND4_X1  g408(.A1(new_n585), .A2(new_n587), .A3(new_n308), .A4(new_n594), .ZN(new_n595));
  AND3_X1   g409(.A1(new_n522), .A2(new_n531), .A3(new_n478), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n476), .B1(new_n596), .B2(new_n532), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT95), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  OAI211_X1 g413(.A(KEYINPUT95), .B(new_n476), .C1(new_n596), .C2(new_n532), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(new_n473), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n595), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(KEYINPUT34), .B(G104), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n603), .B(new_n604), .ZN(G6));
  AOI21_X1  g419(.A(new_n379), .B1(new_n374), .B2(new_n376), .ZN(new_n606));
  INV_X1    g420(.A(new_n376), .ZN(new_n607));
  AOI211_X1 g421(.A(KEYINPUT79), .B(new_n607), .C1(new_n370), .C2(new_n373), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n557), .A2(KEYINPUT83), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n563), .B1(new_n562), .B2(new_n546), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n539), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n612), .A2(G469), .A3(new_n569), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n613), .A2(new_n577), .A3(new_n578), .ZN(new_n614));
  NAND4_X1  g428(.A1(new_n609), .A2(new_n614), .A3(new_n383), .A4(new_n475), .ZN(new_n615));
  AOI211_X1 g429(.A(G472), .B(G902), .C1(new_n261), .C2(new_n274), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n276), .B1(new_n310), .B2(new_n290), .ZN(new_n617));
  NOR3_X1   g431(.A1(new_n615), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT96), .ZN(new_n620));
  AND2_X1   g434(.A1(new_n405), .A2(new_n407), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n421), .B1(new_n621), .B2(new_n400), .ZN(new_n622));
  AOI21_X1  g436(.A(G902), .B1(new_n622), .B2(new_n412), .ZN(new_n623));
  INV_X1    g437(.A(G475), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n620), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n429), .A2(KEYINPUT96), .A3(G475), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NOR3_X1   g441(.A1(new_n422), .A2(new_n420), .A3(new_n416), .ZN(new_n628));
  AOI21_X1  g442(.A(KEYINPUT90), .B1(new_n412), .B2(new_n417), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n386), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n630), .A2(KEYINPUT20), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n423), .A2(new_n424), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n426), .B1(new_n632), .B2(new_n386), .ZN(new_n633));
  OAI211_X1 g447(.A(new_n627), .B(new_n465), .C1(new_n631), .C2(new_n633), .ZN(new_n634));
  NOR3_X1   g448(.A1(new_n619), .A2(new_n602), .A3(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(KEYINPUT35), .B(G107), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G9));
  INV_X1    g451(.A(KEYINPUT36), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n365), .A2(new_n367), .A3(new_n638), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n371), .B1(KEYINPUT36), .B2(new_n366), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n639), .A2(new_n382), .A3(new_n640), .ZN(new_n641));
  XOR2_X1   g455(.A(new_n641), .B(KEYINPUT97), .Z(new_n642));
  NAND3_X1  g456(.A1(new_n378), .A2(new_n642), .A3(new_n380), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n581), .A2(new_n308), .A3(new_n587), .A4(new_n643), .ZN(new_n644));
  XOR2_X1   g458(.A(KEYINPUT37), .B(G110), .Z(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(KEYINPUT98), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n644), .B(new_n646), .ZN(G12));
  NAND4_X1  g461(.A1(new_n643), .A2(new_n601), .A3(new_n475), .A4(new_n614), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n425), .B(new_n426), .ZN(new_n649));
  INV_X1    g463(.A(G900), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n470), .A2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n468), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n649), .A2(new_n465), .A3(new_n627), .A4(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n648), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n655), .A2(new_n307), .A3(new_n313), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(G128), .ZN(G30));
  NOR2_X1   g471(.A1(new_n596), .A2(new_n532), .ZN(new_n658));
  XNOR2_X1  g472(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n659));
  XOR2_X1   g473(.A(new_n658), .B(new_n659), .Z(new_n660));
  AND3_X1   g474(.A1(new_n378), .A2(new_n642), .A3(new_n380), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n427), .A2(new_n430), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n466), .A2(new_n477), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n661), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n660), .B1(new_n664), .B2(KEYINPUT100), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n249), .A2(new_n259), .A3(new_n251), .ZN(new_n666));
  OR2_X1    g480(.A1(new_n262), .A2(new_n285), .ZN(new_n667));
  OAI211_X1 g481(.A(new_n666), .B(new_n290), .C1(new_n259), .C2(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(G472), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n309), .A2(new_n305), .A3(new_n669), .ZN(new_n670));
  OAI211_X1 g484(.A(new_n665), .B(new_n670), .C1(KEYINPUT100), .C2(new_n664), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT101), .ZN(new_n672));
  OR2_X1    g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n671), .A2(new_n672), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n653), .B(KEYINPUT39), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n584), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(KEYINPUT102), .B(KEYINPUT40), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n677), .B(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n673), .A2(new_n674), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G143), .ZN(G45));
  NAND2_X1  g495(.A1(new_n594), .A2(new_n653), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n648), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n683), .A2(new_n307), .A3(new_n313), .ZN(new_n684));
  XOR2_X1   g498(.A(KEYINPUT103), .B(G146), .Z(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(G48));
  INV_X1    g500(.A(new_n594), .ZN(new_n687));
  INV_X1    g501(.A(new_n577), .ZN(new_n688));
  OR2_X1    g502(.A1(new_n572), .A2(KEYINPUT84), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n689), .A2(new_n574), .A3(new_n573), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n566), .B1(new_n690), .B2(new_n290), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(new_n475), .ZN(new_n693));
  NOR3_X1   g507(.A1(new_n687), .A2(new_n602), .A3(new_n693), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n694), .A2(new_n307), .A3(new_n313), .A4(new_n385), .ZN(new_n695));
  XNOR2_X1  g509(.A(KEYINPUT41), .B(G113), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n695), .B(new_n696), .ZN(G15));
  NOR3_X1   g511(.A1(new_n602), .A2(new_n634), .A3(new_n693), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n307), .A2(new_n698), .A3(new_n313), .A4(new_n385), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G116), .ZN(G18));
  NAND3_X1  g514(.A1(new_n601), .A2(new_n475), .A3(new_n692), .ZN(new_n701));
  NOR3_X1   g515(.A1(new_n701), .A2(new_n661), .A3(new_n474), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n307), .A2(new_n702), .A3(new_n313), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G119), .ZN(G21));
  NAND3_X1  g518(.A1(new_n662), .A2(new_n601), .A3(new_n465), .ZN(new_n705));
  NOR3_X1   g519(.A1(new_n705), .A2(new_n472), .A3(new_n693), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n259), .B1(new_n281), .B2(new_n286), .ZN(new_n707));
  OAI211_X1 g521(.A(new_n276), .B(new_n290), .C1(new_n301), .C2(new_n707), .ZN(new_n708));
  AND2_X1   g522(.A1(new_n587), .A2(new_n708), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n706), .A2(new_n385), .A3(new_n709), .ZN(new_n710));
  XOR2_X1   g524(.A(KEYINPUT104), .B(G122), .Z(new_n711));
  XNOR2_X1  g525(.A(new_n710), .B(new_n711), .ZN(G24));
  NAND3_X1  g526(.A1(new_n587), .A2(new_n643), .A3(new_n708), .ZN(new_n713));
  NOR3_X1   g527(.A1(new_n713), .A2(new_n682), .A3(new_n701), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(new_n316), .ZN(G27));
  INV_X1    g529(.A(KEYINPUT106), .ZN(new_n716));
  XOR2_X1   g530(.A(new_n578), .B(KEYINPUT105), .Z(new_n717));
  NAND2_X1  g531(.A1(new_n577), .A2(new_n717), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n716), .B1(new_n571), .B2(new_n718), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n613), .A2(KEYINPUT106), .A3(new_n577), .A4(new_n717), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n658), .A2(new_n475), .A3(new_n476), .ZN(new_n722));
  INV_X1    g536(.A(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n724), .A2(new_n682), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n725), .A2(new_n307), .A3(new_n313), .A4(new_n385), .ZN(new_n726));
  XNOR2_X1  g540(.A(KEYINPUT107), .B(KEYINPUT42), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n722), .B1(new_n719), .B2(new_n720), .ZN(new_n729));
  INV_X1    g543(.A(new_n653), .ZN(new_n730));
  AOI211_X1 g544(.A(new_n730), .B(new_n593), .C1(new_n427), .C2(new_n430), .ZN(new_n731));
  AND3_X1   g545(.A1(new_n729), .A2(new_n731), .A3(KEYINPUT42), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n384), .B1(new_n309), .B2(new_n311), .ZN(new_n733));
  AOI21_X1  g547(.A(KEYINPUT108), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(new_n734), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n732), .A2(KEYINPUT108), .A3(new_n733), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n728), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G131), .ZN(G33));
  NOR2_X1   g552(.A1(new_n724), .A2(new_n654), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n739), .A2(new_n307), .A3(new_n313), .A4(new_n385), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT109), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  AND3_X1   g556(.A1(new_n309), .A2(new_n311), .A3(new_n312), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n312), .B1(new_n309), .B2(new_n311), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n745), .A2(KEYINPUT109), .A3(new_n385), .A4(new_n739), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n742), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G134), .ZN(G36));
  NOR2_X1   g562(.A1(new_n662), .A2(new_n593), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(KEYINPUT43), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n661), .B1(new_n587), .B2(new_n308), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n750), .A2(KEYINPUT44), .A3(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(KEYINPUT110), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n565), .A2(new_n570), .ZN(new_n754));
  OR2_X1    g568(.A1(new_n754), .A2(KEYINPUT45), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(KEYINPUT45), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n755), .A2(G469), .A3(new_n756), .ZN(new_n757));
  AOI21_X1  g571(.A(KEYINPUT46), .B1(new_n757), .B2(new_n717), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n758), .A2(new_n688), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n757), .A2(KEYINPUT46), .A3(new_n717), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n761), .A2(new_n475), .A3(new_n675), .ZN(new_n762));
  AOI21_X1  g576(.A(KEYINPUT44), .B1(new_n750), .B2(new_n751), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n658), .A2(new_n476), .ZN(new_n764));
  NOR3_X1   g578(.A1(new_n762), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n753), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G137), .ZN(G39));
  NAND2_X1  g581(.A1(new_n761), .A2(new_n475), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT47), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n761), .A2(KEYINPUT47), .A3(new_n475), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NOR4_X1   g586(.A1(new_n745), .A2(new_n385), .A3(new_n682), .A4(new_n764), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G140), .ZN(G42));
  INV_X1    g589(.A(new_n692), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(KEYINPUT49), .ZN(new_n777));
  AND3_X1   g591(.A1(new_n592), .A2(new_n475), .A3(new_n476), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n777), .A2(new_n660), .A3(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT49), .ZN(new_n780));
  AOI211_X1 g594(.A(new_n662), .B(new_n779), .C1(new_n780), .C2(new_n692), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n670), .A2(new_n384), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(new_n693), .ZN(new_n784));
  INV_X1    g598(.A(new_n764), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n782), .A2(new_n468), .A3(new_n784), .A4(new_n785), .ZN(new_n786));
  NOR3_X1   g600(.A1(new_n786), .A2(new_n662), .A3(new_n592), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n784), .A2(new_n785), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n750), .A2(new_n468), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(KEYINPUT115), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT115), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n750), .A2(new_n791), .A3(new_n468), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n788), .B1(new_n790), .B2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(new_n713), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n787), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n709), .A2(new_n385), .ZN(new_n796));
  INV_X1    g610(.A(new_n796), .ZN(new_n797));
  AND3_X1   g611(.A1(new_n784), .A2(new_n477), .A3(new_n660), .ZN(new_n798));
  INV_X1    g612(.A(new_n792), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n791), .B1(new_n750), .B2(new_n468), .ZN(new_n800));
  OAI211_X1 g614(.A(new_n797), .B(new_n798), .C1(new_n799), .C2(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(KEYINPUT50), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n796), .B1(new_n790), .B2(new_n792), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT50), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n803), .A2(new_n804), .A3(new_n798), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n795), .A2(new_n802), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n806), .A2(KEYINPUT116), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT116), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n795), .A2(new_n802), .A3(new_n805), .A4(new_n808), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n776), .A2(new_n475), .ZN(new_n810));
  INV_X1    g624(.A(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n770), .A2(new_n771), .A3(new_n811), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n812), .A2(new_n785), .A3(new_n803), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n807), .A2(new_n809), .A3(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT51), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n813), .A2(KEYINPUT51), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n817), .A2(new_n806), .ZN(new_n818));
  OAI211_X1 g632(.A(G952), .B(new_n351), .C1(new_n786), .C2(new_n687), .ZN(new_n819));
  INV_X1    g633(.A(new_n701), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n819), .B1(new_n803), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n793), .A2(new_n733), .ZN(new_n822));
  AND2_X1   g636(.A1(new_n822), .A2(KEYINPUT48), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n822), .A2(KEYINPUT48), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n821), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n818), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n816), .A2(KEYINPUT117), .A3(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT117), .ZN(new_n828));
  AND3_X1   g642(.A1(new_n812), .A2(new_n785), .A3(new_n803), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n829), .B1(new_n806), .B2(KEYINPUT116), .ZN(new_n830));
  AOI21_X1  g644(.A(KEYINPUT51), .B1(new_n830), .B2(new_n809), .ZN(new_n831));
  OAI221_X1 g645(.A(new_n821), .B1(new_n823), .B2(new_n824), .C1(new_n817), .C2(new_n806), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n828), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n827), .A2(new_n833), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n714), .B1(new_n745), .B2(new_n655), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n653), .A2(new_n475), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n705), .A2(new_n643), .A3(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n837), .A2(new_n670), .A3(new_n721), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n835), .A2(KEYINPUT52), .A3(new_n684), .A4(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n794), .A2(new_n731), .A3(new_n820), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n840), .A2(new_n684), .A3(new_n656), .A4(new_n838), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT52), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n839), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n535), .A2(new_n473), .ZN(new_n845));
  INV_X1    g659(.A(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n618), .A2(new_n594), .A3(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n582), .A2(new_n644), .A3(new_n847), .ZN(new_n848));
  OAI211_X1 g662(.A(new_n430), .B(new_n465), .C1(new_n633), .C2(new_n418), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT111), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n427), .A2(KEYINPUT111), .A3(new_n430), .A4(new_n465), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n845), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT112), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n618), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  AOI211_X1 g669(.A(KEYINPUT112), .B(new_n845), .C1(new_n851), .C2(new_n852), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  OAI21_X1  g671(.A(KEYINPUT113), .B1(new_n848), .B2(new_n857), .ZN(new_n858));
  AND2_X1   g672(.A1(new_n849), .A2(new_n850), .ZN(new_n859));
  INV_X1    g673(.A(new_n852), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n846), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(KEYINPUT112), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n853), .A2(new_n854), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n862), .A2(new_n618), .A3(new_n863), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n644), .B1(new_n595), .B2(new_n845), .ZN(new_n865));
  INV_X1    g679(.A(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT113), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n864), .A2(new_n866), .A3(new_n867), .A4(new_n582), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n858), .A2(new_n868), .ZN(new_n869));
  AND3_X1   g683(.A1(new_n732), .A2(KEYINPUT108), .A3(new_n733), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n870), .A2(new_n734), .ZN(new_n871));
  AOI22_X1  g685(.A1(new_n871), .A2(new_n728), .B1(new_n746), .B2(new_n742), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n695), .A2(new_n699), .A3(new_n703), .A4(new_n710), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n725), .A2(new_n709), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n307), .A2(new_n313), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n649), .A2(new_n627), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n723), .A2(new_n614), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n466), .A2(new_n653), .ZN(new_n878));
  OR3_X1    g692(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n874), .B1(new_n875), .B2(new_n879), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n873), .B1(new_n643), .B2(new_n880), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n844), .A2(new_n869), .A3(new_n872), .A4(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT53), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AND4_X1   g698(.A1(new_n695), .A2(new_n699), .A3(new_n703), .A4(new_n710), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n880), .A2(new_n643), .ZN(new_n886));
  AND4_X1   g700(.A1(new_n737), .A2(new_n747), .A3(new_n885), .A4(new_n886), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n887), .A2(KEYINPUT53), .A3(new_n844), .A4(new_n869), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT54), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n884), .A2(new_n888), .A3(KEYINPUT114), .A4(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n884), .A2(new_n888), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n891), .A2(KEYINPUT54), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT114), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n884), .A2(new_n889), .A3(new_n888), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n834), .B1(new_n890), .B2(new_n895), .ZN(new_n896));
  NOR2_X1   g710(.A1(G952), .A2(G953), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n783), .B1(new_n896), .B2(new_n897), .ZN(G75));
  NOR2_X1   g712(.A1(new_n351), .A2(G952), .ZN(new_n899));
  INV_X1    g713(.A(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n290), .B1(new_n884), .B2(new_n888), .ZN(new_n901));
  AOI21_X1  g715(.A(KEYINPUT56), .B1(new_n901), .B2(G210), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n526), .A2(new_n530), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(new_n528), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(KEYINPUT55), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n900), .B1(new_n902), .B2(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n906), .B1(new_n902), .B2(new_n905), .ZN(G51));
  INV_X1    g721(.A(KEYINPUT118), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n892), .A2(new_n908), .A3(new_n894), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n891), .A2(KEYINPUT118), .A3(KEYINPUT54), .ZN(new_n910));
  XOR2_X1   g724(.A(new_n717), .B(KEYINPUT57), .Z(new_n911));
  NAND3_X1  g725(.A1(new_n909), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(new_n690), .ZN(new_n913));
  INV_X1    g727(.A(new_n757), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n901), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n899), .B1(new_n913), .B2(new_n915), .ZN(G54));
  NAND2_X1  g730(.A1(KEYINPUT58), .A2(G475), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n917), .B(KEYINPUT119), .Z(new_n918));
  AND3_X1   g732(.A1(new_n901), .A2(new_n632), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n632), .B1(new_n901), .B2(new_n918), .ZN(new_n920));
  NOR3_X1   g734(.A1(new_n919), .A2(new_n920), .A3(new_n899), .ZN(G60));
  NOR2_X1   g735(.A1(new_n588), .A2(new_n589), .ZN(new_n922));
  XOR2_X1   g736(.A(new_n922), .B(KEYINPUT120), .Z(new_n923));
  NAND2_X1  g737(.A1(G478), .A2(G902), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n924), .B(KEYINPUT59), .Z(new_n925));
  NOR2_X1   g739(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n909), .A2(new_n910), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(KEYINPUT121), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT121), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n909), .A2(new_n929), .A3(new_n910), .A4(new_n926), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(new_n925), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n895), .A2(new_n890), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n899), .B1(new_n933), .B2(new_n923), .ZN(new_n934));
  AND2_X1   g748(.A1(new_n931), .A2(new_n934), .ZN(G63));
  NAND2_X1  g749(.A1(G217), .A2(G902), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n936), .B(KEYINPUT60), .Z(new_n937));
  NAND4_X1  g751(.A1(new_n891), .A2(new_n639), .A3(new_n640), .A4(new_n937), .ZN(new_n938));
  AND2_X1   g752(.A1(new_n891), .A2(new_n937), .ZN(new_n939));
  OAI211_X1 g753(.A(new_n900), .B(new_n938), .C1(new_n939), .C2(new_n381), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT122), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(KEYINPUT61), .ZN(G66));
  INV_X1    g757(.A(G224), .ZN(new_n944));
  OAI21_X1  g758(.A(G953), .B1(new_n471), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n869), .A2(new_n885), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n946), .B(KEYINPUT123), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n945), .B1(new_n947), .B2(G953), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n903), .B1(G898), .B2(new_n351), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n948), .B(new_n949), .ZN(G69));
  AOI21_X1  g764(.A(new_n351), .B1(G227), .B2(G900), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n951), .A2(KEYINPUT126), .ZN(new_n952));
  AND2_X1   g766(.A1(new_n835), .A2(new_n684), .ZN(new_n953));
  AND2_X1   g767(.A1(new_n680), .A2(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT62), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT124), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n954), .A2(KEYINPUT124), .A3(new_n955), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  OR2_X1    g774(.A1(new_n954), .A2(new_n955), .ZN(new_n961));
  NOR3_X1   g775(.A1(new_n859), .A2(new_n860), .A3(new_n594), .ZN(new_n962));
  NOR3_X1   g776(.A1(new_n962), .A2(new_n676), .A3(new_n877), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n963), .A2(new_n745), .A3(new_n385), .ZN(new_n964));
  AND2_X1   g778(.A1(new_n774), .A2(new_n964), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n960), .A2(new_n766), .A3(new_n961), .A4(new_n965), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n237), .A2(new_n243), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n967), .B(new_n414), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n968), .A2(G953), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n952), .B1(new_n966), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n951), .A2(KEYINPUT126), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n385), .B1(new_n277), .B2(new_n306), .ZN(new_n972));
  NOR3_X1   g786(.A1(new_n762), .A2(new_n705), .A3(new_n972), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n973), .B1(new_n772), .B2(new_n773), .ZN(new_n974));
  AND2_X1   g788(.A1(new_n974), .A2(new_n953), .ZN(new_n975));
  NAND4_X1  g789(.A1(new_n975), .A2(KEYINPUT125), .A3(new_n766), .A4(new_n872), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT125), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n974), .A2(new_n766), .A3(new_n953), .ZN(new_n978));
  INV_X1    g792(.A(new_n872), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n977), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  AOI21_X1  g794(.A(G953), .B1(new_n976), .B2(new_n980), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n968), .B1(G900), .B2(new_n351), .ZN(new_n982));
  OAI211_X1 g796(.A(new_n970), .B(new_n971), .C1(new_n981), .C2(new_n982), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n981), .A2(new_n982), .ZN(new_n984));
  OAI211_X1 g798(.A(new_n965), .B(new_n766), .C1(new_n954), .C2(new_n955), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n985), .B1(new_n958), .B2(new_n959), .ZN(new_n986));
  INV_X1    g800(.A(new_n969), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  OAI211_X1 g802(.A(KEYINPUT126), .B(new_n951), .C1(new_n984), .C2(new_n988), .ZN(new_n989));
  AND2_X1   g803(.A1(new_n983), .A2(new_n989), .ZN(G72));
  INV_X1    g804(.A(new_n283), .ZN(new_n991));
  NAND2_X1  g805(.A1(G472), .A2(G902), .ZN(new_n992));
  XOR2_X1   g806(.A(new_n992), .B(KEYINPUT63), .Z(new_n993));
  NAND4_X1  g807(.A1(new_n891), .A2(new_n991), .A3(new_n666), .A4(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(new_n993), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n995), .B1(new_n986), .B2(new_n947), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n994), .B1(new_n996), .B2(new_n666), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n976), .A2(new_n947), .A3(new_n980), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n991), .B1(new_n998), .B2(new_n993), .ZN(new_n999));
  OR3_X1    g813(.A1(new_n999), .A2(KEYINPUT127), .A3(new_n899), .ZN(new_n1000));
  OAI21_X1  g814(.A(KEYINPUT127), .B1(new_n999), .B2(new_n899), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n997), .B1(new_n1000), .B2(new_n1001), .ZN(G57));
endmodule


