//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 0 0 0 0 1 1 1 1 0 0 0 1 1 0 0 1 0 0 1 0 1 0 1 1 1 0 1 1 0 1 1 1 0 1 1 0 0 1 1 0 1 1 0 0 0 0 0 1 1 1 0 1 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:26 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n449, new_n450, new_n452, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n461, new_n462, new_n463, new_n464,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n547, new_n549, new_n550,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n564, new_n565, new_n566, new_n567, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n594, new_n595,
    new_n596, new_n597, new_n600, new_n602, new_n603, new_n604, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1117, new_n1118;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT64), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT65), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XOR2_X1   g017(.A(new_n442), .B(KEYINPUT66), .Z(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  INV_X1    g023(.A(G567), .ZN(new_n449));
  NOR2_X1   g024(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT67), .Z(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT68), .ZN(G217));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT2), .ZN(new_n455));
  NAND4_X1  g030(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT69), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G325));
  XOR2_X1   g034(.A(new_n458), .B(KEYINPUT70), .Z(G261));
  INV_X1    g035(.A(new_n455), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G2106), .ZN(new_n462));
  OR2_X1    g037(.A1(new_n457), .A2(new_n449), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(G319));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  XNOR2_X1  g041(.A(KEYINPUT3), .B(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G125), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT71), .ZN(new_n470));
  XNOR2_X1  g045(.A(new_n469), .B(new_n470), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n466), .B1(new_n468), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n466), .A2(G2104), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT72), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n466), .A2(KEYINPUT72), .A3(G2104), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n475), .A2(G101), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n467), .A2(new_n466), .ZN(new_n478));
  INV_X1    g053(.A(G137), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n472), .A2(new_n480), .ZN(G160));
  INV_X1    g056(.A(new_n478), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G136), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n483), .B(KEYINPUT73), .ZN(new_n484));
  INV_X1    g059(.A(new_n467), .ZN(new_n485));
  OAI21_X1  g060(.A(KEYINPUT74), .B1(new_n485), .B2(new_n466), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT74), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n467), .A2(new_n487), .A3(G2105), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G124), .ZN(new_n491));
  MUX2_X1   g066(.A(G100), .B(G112), .S(G2105), .Z(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G2104), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n484), .A2(new_n491), .A3(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(G162));
  AND2_X1   g070(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n496));
  NOR2_X1   g071(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n497));
  OAI211_X1 g072(.A(G138), .B(new_n466), .C1(new_n496), .C2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n467), .A2(KEYINPUT4), .A3(G138), .A4(new_n466), .ZN(new_n501));
  OAI21_X1  g076(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT75), .ZN(new_n504));
  INV_X1    g079(.A(G114), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n504), .B1(new_n505), .B2(G2105), .ZN(new_n506));
  NOR3_X1   g081(.A1(new_n466), .A2(KEYINPUT75), .A3(G114), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n503), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n467), .A2(G126), .A3(G2105), .ZN(new_n509));
  NAND4_X1  g084(.A1(new_n500), .A2(new_n501), .A3(new_n508), .A4(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(G164));
  XNOR2_X1  g086(.A(KEYINPUT6), .B(G651), .ZN(new_n512));
  XNOR2_X1  g087(.A(KEYINPUT5), .B(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(G88), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n512), .A2(G543), .ZN(new_n516));
  INV_X1    g091(.A(G50), .ZN(new_n517));
  OAI22_X1  g092(.A1(new_n514), .A2(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n513), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n519));
  INV_X1    g094(.A(G651), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n518), .A2(new_n521), .ZN(G166));
  NAND3_X1  g097(.A1(new_n513), .A2(G63), .A3(G651), .ZN(new_n523));
  INV_X1    g098(.A(G51), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n523), .B1(new_n516), .B2(new_n524), .ZN(new_n525));
  AND2_X1   g100(.A1(new_n525), .A2(KEYINPUT76), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n525), .A2(KEYINPUT76), .ZN(new_n527));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n528), .B(KEYINPUT7), .ZN(new_n529));
  INV_X1    g104(.A(G89), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n529), .B1(new_n514), .B2(new_n530), .ZN(new_n531));
  NOR3_X1   g106(.A1(new_n526), .A2(new_n527), .A3(new_n531), .ZN(G168));
  INV_X1    g107(.A(G90), .ZN(new_n533));
  INV_X1    g108(.A(G52), .ZN(new_n534));
  OAI22_X1  g109(.A1(new_n514), .A2(new_n533), .B1(new_n516), .B2(new_n534), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n513), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n536), .A2(new_n520), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n535), .A2(new_n537), .ZN(G171));
  INV_X1    g113(.A(G81), .ZN(new_n539));
  INV_X1    g114(.A(G43), .ZN(new_n540));
  OAI22_X1  g115(.A1(new_n514), .A2(new_n539), .B1(new_n516), .B2(new_n540), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n513), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n542), .A2(new_n520), .ZN(new_n543));
  OR2_X1    g118(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G860), .ZN(G153));
  AND3_X1   g121(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G36), .ZN(G176));
  NAND2_X1  g123(.A1(G1), .A2(G3), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT8), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n547), .A2(new_n550), .ZN(G188));
  INV_X1    g126(.A(new_n516), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G53), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT9), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n553), .B(new_n554), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n513), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n556));
  INV_X1    g131(.A(G91), .ZN(new_n557));
  OAI22_X1  g132(.A1(new_n556), .A2(new_n520), .B1(new_n514), .B2(new_n557), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(new_n559), .ZN(G299));
  INV_X1    g135(.A(G171), .ZN(G301));
  OR3_X1    g136(.A1(new_n526), .A2(new_n527), .A3(new_n531), .ZN(G286));
  INV_X1    g137(.A(G166), .ZN(G303));
  NAND2_X1  g138(.A1(new_n552), .A2(G49), .ZN(new_n564));
  AND2_X1   g139(.A1(new_n512), .A2(new_n513), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G87), .ZN(new_n566));
  OAI21_X1  g141(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n564), .A2(new_n566), .A3(new_n567), .ZN(G288));
  AOI22_X1  g143(.A1(new_n513), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n569));
  OR2_X1    g144(.A1(new_n569), .A2(new_n520), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n565), .A2(G86), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n552), .A2(G48), .ZN(new_n572));
  AND3_X1   g147(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(G305));
  INV_X1    g149(.A(G85), .ZN(new_n575));
  INV_X1    g150(.A(G47), .ZN(new_n576));
  OAI22_X1  g151(.A1(new_n514), .A2(new_n575), .B1(new_n516), .B2(new_n576), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n513), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n578));
  NOR2_X1   g153(.A1(new_n578), .A2(new_n520), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(G290));
  INV_X1    g156(.A(G868), .ZN(new_n582));
  NOR2_X1   g157(.A1(G301), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n565), .A2(G92), .ZN(new_n584));
  XOR2_X1   g159(.A(new_n584), .B(KEYINPUT10), .Z(new_n585));
  XNOR2_X1  g160(.A(new_n516), .B(KEYINPUT77), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n586), .A2(G54), .ZN(new_n587));
  AND2_X1   g162(.A1(new_n513), .A2(G66), .ZN(new_n588));
  AND2_X1   g163(.A1(G79), .A2(G543), .ZN(new_n589));
  OAI21_X1  g164(.A(G651), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  AND3_X1   g165(.A1(new_n585), .A2(new_n587), .A3(new_n590), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n583), .B1(new_n591), .B2(new_n582), .ZN(G284));
  AOI21_X1  g167(.A(new_n583), .B1(new_n591), .B2(new_n582), .ZN(G321));
  NOR2_X1   g168(.A1(G168), .A2(new_n582), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT78), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  AOI21_X1  g171(.A(KEYINPUT78), .B1(G299), .B2(new_n582), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n597), .B2(new_n594), .ZN(G297));
  OAI21_X1  g173(.A(new_n596), .B1(new_n597), .B2(new_n594), .ZN(G280));
  INV_X1    g174(.A(G559), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n591), .B1(new_n600), .B2(G860), .ZN(G148));
  NAND2_X1  g176(.A1(new_n545), .A2(new_n582), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n591), .A2(new_n600), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n603), .B2(new_n582), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n604), .B(KEYINPUT79), .ZN(G323));
  XNOR2_X1  g180(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND2_X1   g181(.A1(new_n475), .A2(new_n476), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n607), .A2(new_n467), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT12), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT13), .ZN(new_n610));
  INV_X1    g185(.A(G2100), .ZN(new_n611));
  OR2_X1    g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n610), .A2(new_n611), .ZN(new_n613));
  MUX2_X1   g188(.A(G99), .B(G111), .S(G2105), .Z(new_n614));
  AOI22_X1  g189(.A1(new_n482), .A2(G135), .B1(G2104), .B2(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(G123), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n489), .B2(new_n616), .ZN(new_n617));
  INV_X1    g192(.A(G2096), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n617), .B(new_n618), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n612), .A2(new_n613), .A3(new_n619), .ZN(G156));
  INV_X1    g195(.A(KEYINPUT14), .ZN(new_n621));
  XOR2_X1   g196(.A(KEYINPUT15), .B(G2435), .Z(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(G2438), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(G2427), .ZN(new_n624));
  INV_X1    g199(.A(G2430), .ZN(new_n625));
  AOI21_X1  g200(.A(new_n621), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n626), .B1(new_n625), .B2(new_n624), .ZN(new_n627));
  XNOR2_X1  g202(.A(G2451), .B(G2454), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT16), .ZN(new_n629));
  XNOR2_X1  g204(.A(G2443), .B(G2446), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(G1341), .B(G1348), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n627), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n627), .A2(new_n633), .ZN(new_n635));
  AND3_X1   g210(.A1(new_n634), .A2(G14), .A3(new_n635), .ZN(G401));
  XOR2_X1   g211(.A(G2084), .B(G2090), .Z(new_n637));
  INV_X1    g212(.A(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(G2072), .B(G2078), .Z(new_n639));
  XNOR2_X1  g214(.A(G2067), .B(G2678), .ZN(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(new_n641));
  NOR3_X1   g216(.A1(new_n638), .A2(new_n639), .A3(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT18), .ZN(new_n643));
  INV_X1    g218(.A(new_n639), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n644), .A2(KEYINPUT17), .ZN(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n640), .B1(new_n646), .B2(new_n637), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n647), .B1(new_n638), .B2(new_n645), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n638), .A2(new_n641), .ZN(new_n649));
  AOI21_X1  g224(.A(new_n644), .B1(new_n649), .B2(KEYINPUT17), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n643), .B1(new_n648), .B2(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(new_n618), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(new_n611), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(G227));
  XOR2_X1   g229(.A(G1971), .B(G1976), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT19), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1956), .B(G2474), .ZN(new_n657));
  XNOR2_X1  g232(.A(G1961), .B(G1966), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  AND2_X1   g234(.A1(new_n657), .A2(new_n658), .ZN(new_n660));
  NOR3_X1   g235(.A1(new_n656), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n656), .A2(new_n659), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n662), .B(KEYINPUT20), .Z(new_n663));
  AOI211_X1 g238(.A(new_n661), .B(new_n663), .C1(new_n656), .C2(new_n660), .ZN(new_n664));
  XOR2_X1   g239(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n665));
  XOR2_X1   g240(.A(new_n664), .B(new_n665), .Z(new_n666));
  XNOR2_X1  g241(.A(G1991), .B(G1996), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1981), .B(G1986), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n666), .B(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(G229));
  NOR2_X1   g246(.A1(G25), .A2(G29), .ZN(new_n672));
  MUX2_X1   g247(.A(G95), .B(G107), .S(G2105), .Z(new_n673));
  AOI22_X1  g248(.A1(new_n482), .A2(G131), .B1(G2104), .B2(new_n673), .ZN(new_n674));
  INV_X1    g249(.A(G119), .ZN(new_n675));
  OAI21_X1  g250(.A(new_n674), .B1(new_n489), .B2(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n676), .B(KEYINPUT80), .Z(new_n677));
  AOI21_X1  g252(.A(new_n672), .B1(new_n677), .B2(G29), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT81), .ZN(new_n679));
  XOR2_X1   g254(.A(KEYINPUT35), .B(G1991), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  NOR2_X1   g256(.A1(G16), .A2(G24), .ZN(new_n682));
  AOI21_X1  g257(.A(new_n682), .B1(new_n580), .B2(G16), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(G1986), .ZN(new_n684));
  NOR2_X1   g259(.A1(G6), .A2(G16), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n685), .B1(new_n573), .B2(G16), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT32), .B(G1981), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT82), .ZN(new_n688));
  XOR2_X1   g263(.A(new_n686), .B(new_n688), .Z(new_n689));
  INV_X1    g264(.A(G16), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n690), .A2(G23), .ZN(new_n691));
  INV_X1    g266(.A(G288), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n691), .B1(new_n692), .B2(new_n690), .ZN(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT33), .B(G1976), .ZN(new_n694));
  XOR2_X1   g269(.A(new_n693), .B(new_n694), .Z(new_n695));
  NOR2_X1   g270(.A1(G16), .A2(G22), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(G166), .B2(G16), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(G1971), .ZN(new_n698));
  NOR3_X1   g273(.A1(new_n689), .A2(new_n695), .A3(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(KEYINPUT34), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n684), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  OAI211_X1 g276(.A(new_n681), .B(new_n701), .C1(new_n700), .C2(new_n699), .ZN(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT83), .B(KEYINPUT36), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  NOR2_X1   g279(.A1(G29), .A2(G32), .ZN(new_n705));
  NAND3_X1  g280(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT26), .ZN(new_n707));
  AND2_X1   g282(.A1(new_n607), .A2(G105), .ZN(new_n708));
  AOI211_X1 g283(.A(new_n707), .B(new_n708), .C1(G141), .C2(new_n482), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n490), .A2(G129), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n705), .B1(new_n712), .B2(G29), .ZN(new_n713));
  XOR2_X1   g288(.A(new_n713), .B(KEYINPUT89), .Z(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT27), .B(G1996), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NOR2_X1   g291(.A1(G4), .A2(G16), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(KEYINPUT84), .Z(new_n718));
  NAND3_X1  g293(.A1(new_n585), .A2(new_n587), .A3(new_n590), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n718), .B1(new_n719), .B2(new_n690), .ZN(new_n720));
  XOR2_X1   g295(.A(KEYINPUT85), .B(G1348), .Z(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT86), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n720), .B(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(KEYINPUT25), .ZN(new_n724));
  INV_X1    g299(.A(G103), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n724), .B1(new_n473), .B2(new_n725), .ZN(new_n726));
  NAND4_X1  g301(.A1(new_n466), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n727));
  AOI22_X1  g302(.A1(new_n482), .A2(G139), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  AND2_X1   g303(.A1(new_n467), .A2(G127), .ZN(new_n729));
  AND2_X1   g304(.A1(G115), .A2(G2104), .ZN(new_n730));
  OAI21_X1  g305(.A(G2105), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n728), .A2(new_n731), .ZN(new_n732));
  MUX2_X1   g307(.A(G33), .B(new_n732), .S(G29), .Z(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(G2072), .Z(new_n734));
  INV_X1    g309(.A(G29), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n617), .A2(new_n735), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT91), .Z(new_n737));
  NOR2_X1   g312(.A1(G27), .A2(G29), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(G164), .B2(G29), .ZN(new_n739));
  XOR2_X1   g314(.A(KEYINPUT94), .B(G2078), .Z(new_n740));
  NAND2_X1  g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n734), .A2(new_n737), .A3(new_n741), .ZN(new_n742));
  NOR3_X1   g317(.A1(new_n716), .A2(new_n723), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n690), .A2(G5), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G171), .B2(new_n690), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n745), .A2(G1961), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT93), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n690), .A2(G21), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G168), .B2(new_n690), .ZN(new_n749));
  INV_X1    g324(.A(G1966), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(KEYINPUT30), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n735), .B1(new_n752), .B2(G28), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n753), .A2(KEYINPUT92), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(new_n752), .B2(G28), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n753), .A2(KEYINPUT92), .ZN(new_n756));
  AND2_X1   g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  XOR2_X1   g332(.A(KEYINPUT31), .B(G11), .Z(new_n758));
  AND2_X1   g333(.A1(KEYINPUT24), .A2(G34), .ZN(new_n759));
  NOR2_X1   g334(.A1(KEYINPUT24), .A2(G34), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n735), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(G160), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n761), .B1(new_n762), .B2(new_n735), .ZN(new_n763));
  INV_X1    g338(.A(G2084), .ZN(new_n764));
  AOI211_X1 g339(.A(new_n757), .B(new_n758), .C1(new_n763), .C2(new_n764), .ZN(new_n765));
  OAI221_X1 g340(.A(new_n765), .B1(G1961), .B2(new_n745), .C1(new_n764), .C2(new_n763), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n690), .A2(G20), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT95), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT23), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(new_n559), .B2(new_n690), .ZN(new_n770));
  XNOR2_X1  g345(.A(KEYINPUT96), .B(G1956), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n735), .A2(G26), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(KEYINPUT28), .Z(new_n774));
  MUX2_X1   g349(.A(G104), .B(G116), .S(G2105), .Z(new_n775));
  AOI22_X1  g350(.A1(new_n482), .A2(G140), .B1(G2104), .B2(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(G128), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n776), .B1(new_n489), .B2(new_n777), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n774), .B1(new_n778), .B2(G29), .ZN(new_n779));
  XOR2_X1   g354(.A(KEYINPUT88), .B(G2067), .Z(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  OAI211_X1 g356(.A(new_n772), .B(new_n781), .C1(new_n739), .C2(new_n740), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n690), .A2(G19), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(KEYINPUT87), .Z(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(new_n544), .B2(G16), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(G1341), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(new_n770), .B2(new_n771), .ZN(new_n787));
  NOR3_X1   g362(.A1(new_n766), .A2(new_n782), .A3(new_n787), .ZN(new_n788));
  NAND4_X1  g363(.A1(new_n743), .A2(new_n747), .A3(new_n751), .A4(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n714), .A2(new_n715), .ZN(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(KEYINPUT90), .Z(new_n791));
  NOR2_X1   g366(.A1(G29), .A2(G35), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(G162), .B2(G29), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT29), .ZN(new_n794));
  INV_X1    g369(.A(G2090), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n791), .A2(new_n796), .ZN(new_n797));
  NOR3_X1   g372(.A1(new_n704), .A2(new_n789), .A3(new_n797), .ZN(G311));
  INV_X1    g373(.A(G311), .ZN(G150));
  NAND2_X1  g374(.A1(new_n552), .A2(G55), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n565), .A2(G93), .ZN(new_n801));
  AOI22_X1  g376(.A1(new_n513), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n802));
  OAI211_X1 g377(.A(new_n800), .B(new_n801), .C1(new_n520), .C2(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n803), .A2(G860), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(KEYINPUT37), .Z(new_n805));
  AND2_X1   g380(.A1(new_n544), .A2(new_n803), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n544), .A2(new_n803), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT38), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n719), .A2(new_n600), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(new_n811), .ZN(new_n812));
  AND2_X1   g387(.A1(new_n812), .A2(KEYINPUT39), .ZN(new_n813));
  INV_X1    g388(.A(G860), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n814), .B1(new_n812), .B2(KEYINPUT39), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n805), .B1(new_n813), .B2(new_n815), .ZN(G145));
  XNOR2_X1  g391(.A(new_n617), .B(new_n762), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(new_n494), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n677), .B(KEYINPUT98), .ZN(new_n819));
  MUX2_X1   g394(.A(G106), .B(G118), .S(G2105), .Z(new_n820));
  AOI22_X1  g395(.A1(new_n482), .A2(G142), .B1(G2104), .B2(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(G130), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n821), .B1(new_n489), .B2(new_n822), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n609), .B(new_n823), .Z(new_n824));
  XNOR2_X1  g399(.A(new_n819), .B(new_n824), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n732), .A2(KEYINPUT97), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n711), .B(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n778), .B(G164), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n825), .A2(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT99), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  OR2_X1    g407(.A1(new_n825), .A2(new_n829), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n830), .A2(new_n831), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n818), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n818), .B(KEYINPUT100), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n837), .B1(new_n825), .B2(new_n829), .ZN(new_n838));
  AOI21_X1  g413(.A(G37), .B1(new_n833), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n836), .A2(new_n839), .ZN(new_n840));
  XOR2_X1   g415(.A(KEYINPUT101), .B(KEYINPUT40), .Z(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(G395));
  NOR2_X1   g417(.A1(new_n803), .A2(G868), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT102), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n591), .A2(new_n844), .A3(G299), .ZN(new_n845));
  OAI21_X1  g420(.A(KEYINPUT102), .B1(new_n719), .B2(new_n559), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n845), .A2(KEYINPUT103), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n719), .A2(new_n559), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n845), .A2(new_n846), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT103), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  NAND4_X1  g429(.A1(new_n853), .A2(KEYINPUT41), .A3(new_n848), .A4(new_n847), .ZN(new_n855));
  AOI22_X1  g430(.A1(new_n845), .A2(new_n846), .B1(new_n559), .B2(new_n719), .ZN(new_n856));
  OR2_X1    g431(.A1(new_n856), .A2(KEYINPUT41), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n603), .B(new_n808), .ZN(new_n859));
  MUX2_X1   g434(.A(new_n854), .B(new_n858), .S(new_n859), .Z(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT42), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n573), .B(G166), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n692), .B(new_n580), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n862), .B(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n861), .B(new_n864), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n843), .B1(new_n865), .B2(G868), .ZN(G295));
  AOI21_X1  g441(.A(new_n843), .B1(new_n865), .B2(G868), .ZN(G331));
  INV_X1    g442(.A(KEYINPUT44), .ZN(new_n868));
  NAND2_X1  g443(.A1(G168), .A2(G171), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  NOR2_X1   g445(.A1(G168), .A2(G171), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  XOR2_X1   g447(.A(new_n872), .B(new_n808), .Z(new_n873));
  NAND2_X1  g448(.A1(new_n854), .A2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n871), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n875), .A2(new_n808), .A3(new_n869), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n876), .A2(KEYINPUT104), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT104), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n872), .A2(new_n878), .A3(new_n808), .ZN(new_n879));
  OAI211_X1 g454(.A(new_n877), .B(new_n879), .C1(new_n808), .C2(new_n872), .ZN(new_n880));
  AND3_X1   g455(.A1(new_n858), .A2(KEYINPUT105), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(KEYINPUT105), .B1(new_n858), .B2(new_n880), .ZN(new_n882));
  OAI211_X1 g457(.A(new_n864), .B(new_n874), .C1(new_n881), .C2(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n880), .B1(new_n853), .B2(new_n850), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT41), .ZN(new_n885));
  AOI21_X1  g460(.A(KEYINPUT103), .B1(new_n845), .B2(new_n846), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n885), .B1(new_n849), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n856), .A2(KEYINPUT41), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT107), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n856), .A2(KEYINPUT107), .A3(KEYINPUT41), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n887), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n873), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n884), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  XOR2_X1   g469(.A(new_n864), .B(KEYINPUT106), .Z(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  OAI21_X1  g471(.A(KEYINPUT108), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT108), .ZN(new_n898));
  AND3_X1   g473(.A1(new_n856), .A2(KEYINPUT107), .A3(KEYINPUT41), .ZN(new_n899));
  AOI21_X1  g474(.A(KEYINPUT107), .B1(new_n856), .B2(KEYINPUT41), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n873), .B1(new_n901), .B2(new_n887), .ZN(new_n902));
  OAI211_X1 g477(.A(new_n898), .B(new_n895), .C1(new_n902), .C2(new_n884), .ZN(new_n903));
  INV_X1    g478(.A(G37), .ZN(new_n904));
  NAND4_X1  g479(.A1(new_n883), .A2(new_n897), .A3(new_n903), .A4(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(KEYINPUT43), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n874), .B1(new_n881), .B2(new_n882), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(new_n895), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT43), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n908), .A2(new_n909), .A3(new_n904), .A4(new_n883), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n868), .B1(new_n906), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n905), .A2(new_n909), .ZN(new_n912));
  NAND4_X1  g487(.A1(new_n908), .A2(KEYINPUT43), .A3(new_n904), .A4(new_n883), .ZN(new_n913));
  AOI21_X1  g488(.A(KEYINPUT44), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n911), .A2(new_n914), .ZN(G397));
  OR2_X1    g490(.A1(new_n677), .A2(new_n680), .ZN(new_n916));
  INV_X1    g491(.A(G1996), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n711), .B(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(G2067), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n778), .B(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n677), .A2(new_n680), .ZN(new_n921));
  NAND4_X1  g496(.A1(new_n916), .A2(new_n918), .A3(new_n920), .A4(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(G1384), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n510), .A2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT45), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(G160), .A2(G40), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n922), .A2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(G1986), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n928), .A2(new_n930), .A3(new_n580), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n931), .B(KEYINPUT48), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n918), .A2(new_n920), .ZN(new_n933));
  OAI22_X1  g508(.A1(new_n933), .A2(new_n921), .B1(G2067), .B2(new_n778), .ZN(new_n934));
  AOI22_X1  g509(.A1(new_n929), .A2(new_n932), .B1(new_n934), .B2(new_n928), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n928), .A2(new_n917), .ZN(new_n936));
  OR2_X1    g511(.A1(new_n936), .A2(KEYINPUT46), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(KEYINPUT46), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n712), .A2(new_n920), .ZN(new_n939));
  AOI22_X1  g514(.A1(new_n937), .A2(new_n938), .B1(new_n939), .B2(new_n928), .ZN(new_n940));
  XOR2_X1   g515(.A(new_n940), .B(KEYINPUT47), .Z(new_n941));
  NAND2_X1  g516(.A1(new_n935), .A2(new_n941), .ZN(new_n942));
  XOR2_X1   g517(.A(new_n942), .B(KEYINPUT127), .Z(new_n943));
  NAND2_X1  g518(.A1(G303), .A2(G8), .ZN(new_n944));
  XOR2_X1   g519(.A(new_n944), .B(KEYINPUT55), .Z(new_n945));
  INV_X1    g520(.A(G40), .ZN(new_n946));
  NOR3_X1   g521(.A1(new_n472), .A2(new_n480), .A3(new_n946), .ZN(new_n947));
  AND3_X1   g522(.A1(new_n510), .A2(KEYINPUT50), .A3(new_n923), .ZN(new_n948));
  AOI21_X1  g523(.A(KEYINPUT50), .B1(new_n510), .B2(new_n923), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n947), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  OR2_X1    g525(.A1(new_n950), .A2(G2090), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT109), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n924), .A2(new_n952), .A3(new_n925), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n510), .A2(KEYINPUT45), .A3(new_n923), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(KEYINPUT109), .ZN(new_n955));
  AOI21_X1  g530(.A(KEYINPUT45), .B1(new_n510), .B2(new_n923), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n953), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  AOI21_X1  g532(.A(G1971), .B1(new_n957), .B2(new_n947), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n951), .B1(new_n958), .B2(KEYINPUT110), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n926), .A2(KEYINPUT109), .A3(new_n954), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n927), .B1(new_n960), .B2(new_n953), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT110), .ZN(new_n962));
  NOR3_X1   g537(.A1(new_n961), .A2(new_n962), .A3(G1971), .ZN(new_n963));
  OAI211_X1 g538(.A(G8), .B(new_n945), .C1(new_n959), .C2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT111), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n962), .B1(new_n961), .B2(G1971), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n958), .A2(KEYINPUT110), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n967), .A2(new_n968), .A3(new_n951), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n969), .A2(KEYINPUT111), .A3(G8), .A4(new_n945), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n966), .A2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(G1981), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n573), .A2(KEYINPUT113), .A3(new_n972), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n570), .A2(new_n972), .A3(new_n571), .A4(new_n572), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT113), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n973), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n572), .A2(new_n571), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT114), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n572), .A2(new_n571), .A3(KEYINPUT114), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n980), .A2(new_n981), .A3(new_n570), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(G1981), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n977), .A2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT116), .ZN(new_n985));
  XNOR2_X1  g560(.A(KEYINPUT115), .B(KEYINPUT49), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n984), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  AOI22_X1  g562(.A1(new_n973), .A2(new_n976), .B1(new_n982), .B2(G1981), .ZN(new_n988));
  INV_X1    g563(.A(new_n986), .ZN(new_n989));
  OAI21_X1  g564(.A(KEYINPUT116), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n987), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(G8), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n927), .A2(new_n924), .ZN(new_n993));
  AOI211_X1 g568(.A(new_n992), .B(new_n993), .C1(new_n988), .C2(KEYINPUT49), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n991), .A2(new_n994), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n993), .A2(new_n992), .ZN(new_n996));
  INV_X1    g571(.A(G1976), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n996), .B1(new_n997), .B2(G288), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(KEYINPUT52), .ZN(new_n999));
  XNOR2_X1  g574(.A(KEYINPUT112), .B(G1976), .ZN(new_n1000));
  AOI21_X1  g575(.A(KEYINPUT52), .B1(G288), .B2(new_n1000), .ZN(new_n1001));
  OAI211_X1 g576(.A(new_n996), .B(new_n1001), .C1(new_n997), .C2(G288), .ZN(new_n1002));
  AND2_X1   g577(.A1(new_n999), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n995), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(new_n958), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n992), .B1(new_n1006), .B2(new_n951), .ZN(new_n1007));
  OR2_X1    g582(.A1(new_n1007), .A2(new_n945), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n971), .A2(new_n1005), .A3(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(G2078), .ZN(new_n1010));
  AOI21_X1  g585(.A(KEYINPUT53), .B1(new_n961), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT123), .ZN(new_n1012));
  INV_X1    g587(.A(G1961), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n950), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT53), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1015), .A2(G2078), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n926), .A2(new_n954), .A3(new_n947), .A4(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1012), .B1(new_n1014), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1018), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1014), .A2(new_n1012), .A3(new_n1017), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1011), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  XNOR2_X1  g596(.A(G171), .B(KEYINPUT54), .ZN(new_n1022));
  OR2_X1    g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1017), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1024), .B1(KEYINPUT124), .B2(new_n1014), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n957), .A2(new_n947), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1015), .B1(new_n1026), .B2(G2078), .ZN(new_n1027));
  OAI211_X1 g602(.A(new_n1025), .B(new_n1027), .C1(KEYINPUT124), .C2(new_n1014), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT121), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n947), .A2(new_n954), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n750), .B1(new_n1030), .B2(new_n956), .ZN(new_n1031));
  OAI211_X1 g606(.A(new_n764), .B(new_n947), .C1(new_n948), .C2(new_n949), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  OAI211_X1 g608(.A(new_n1029), .B(G8), .C1(new_n1033), .C2(G286), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT122), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT51), .ZN(new_n1037));
  OAI211_X1 g612(.A(KEYINPUT122), .B(G8), .C1(new_n1033), .C2(G286), .ZN(new_n1038));
  AND3_X1   g613(.A1(new_n1036), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(G8), .B1(new_n1033), .B2(G286), .ZN(new_n1040));
  OAI211_X1 g615(.A(new_n1035), .B(KEYINPUT51), .C1(new_n1040), .C2(KEYINPUT121), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n992), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(G286), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1041), .A2(new_n1043), .ZN(new_n1044));
  OAI211_X1 g619(.A(new_n1023), .B(new_n1028), .C1(new_n1039), .C2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g620(.A(KEYINPUT125), .B1(new_n1009), .B2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1028), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1044), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1036), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1047), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1004), .B1(new_n966), .B2(new_n970), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT125), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1050), .A2(new_n1051), .A3(new_n1052), .A4(new_n1008), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT61), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT118), .ZN(new_n1055));
  INV_X1    g630(.A(new_n950), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1055), .B1(new_n1056), .B2(G1956), .ZN(new_n1057));
  INV_X1    g632(.A(G1956), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n950), .A2(KEYINPUT118), .A3(new_n1058), .ZN(new_n1059));
  XOR2_X1   g634(.A(KEYINPUT56), .B(G2072), .Z(new_n1060));
  OAI211_X1 g635(.A(new_n1057), .B(new_n1059), .C1(new_n1026), .C2(new_n1060), .ZN(new_n1061));
  XNOR2_X1  g636(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n1062));
  XNOR2_X1  g637(.A(new_n559), .B(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1064), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1054), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  OR2_X1    g642(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1068), .A2(KEYINPUT61), .A3(new_n1064), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n993), .A2(KEYINPUT120), .A3(new_n919), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT120), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n947), .A2(new_n923), .A3(new_n510), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1071), .B1(new_n1072), .B2(G2067), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1070), .B(new_n1073), .C1(new_n1056), .C2(G1348), .ZN(new_n1074));
  NOR3_X1   g649(.A1(new_n1074), .A2(KEYINPUT60), .A3(new_n719), .ZN(new_n1075));
  XNOR2_X1  g650(.A(new_n1074), .B(new_n591), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1075), .B1(new_n1076), .B2(KEYINPUT60), .ZN(new_n1077));
  XNOR2_X1  g652(.A(KEYINPUT58), .B(G1341), .ZN(new_n1078));
  OAI22_X1  g653(.A1(new_n1026), .A2(G1996), .B1(new_n993), .B2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(new_n545), .ZN(new_n1080));
  XNOR2_X1  g655(.A(new_n1080), .B(KEYINPUT59), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1067), .A2(new_n1069), .A3(new_n1077), .A4(new_n1081), .ZN(new_n1082));
  AND2_X1   g657(.A1(new_n1074), .A2(new_n591), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1065), .B1(new_n1068), .B2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1082), .A2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1046), .A2(new_n1053), .A3(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n692), .A2(new_n997), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1087), .B1(new_n991), .B2(new_n994), .ZN(new_n1088));
  INV_X1    g663(.A(new_n977), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n996), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1090), .B1(new_n971), .B2(new_n1004), .ZN(new_n1091));
  OAI21_X1  g666(.A(KEYINPUT62), .B1(new_n1039), .B2(new_n1044), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT62), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1049), .A2(new_n1093), .A3(new_n1041), .A4(new_n1043), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1021), .A2(G301), .ZN(new_n1095));
  AND3_X1   g670(.A1(new_n1092), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1009), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1091), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1042), .A2(G168), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1099), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n971), .A2(new_n1005), .A3(new_n1100), .A4(new_n1008), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT63), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1101), .A2(KEYINPUT117), .A3(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n945), .B1(new_n969), .B2(G8), .ZN(new_n1104));
  NOR3_X1   g679(.A1(new_n1104), .A2(new_n1102), .A3(new_n1099), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1051), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1103), .A2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(KEYINPUT117), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1108));
  OAI211_X1 g683(.A(new_n1086), .B(new_n1098), .C1(new_n1107), .C2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT126), .ZN(new_n1110));
  XNOR2_X1  g685(.A(new_n580), .B(new_n930), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n928), .B1(new_n922), .B2(new_n1111), .ZN(new_n1112));
  AND3_X1   g687(.A1(new_n1109), .A2(new_n1110), .A3(new_n1112), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1110), .B1(new_n1109), .B2(new_n1112), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n943), .B1(new_n1113), .B2(new_n1114), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g690(.A1(G401), .A2(new_n464), .ZN(new_n1117));
  AND4_X1   g691(.A1(new_n653), .A2(new_n840), .A3(new_n670), .A4(new_n1117), .ZN(new_n1118));
  AND3_X1   g692(.A1(new_n1118), .A2(new_n912), .A3(new_n913), .ZN(G308));
  NAND3_X1  g693(.A1(new_n1118), .A2(new_n912), .A3(new_n913), .ZN(G225));
endmodule


