//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 0 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 1 1 0 1 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 0 0 1 1 0 1 0 0 0 0 0 0 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:43 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n450, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n554, new_n555, new_n556, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n566, new_n567, new_n568, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n602,
    new_n605, new_n607, new_n608, new_n609, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n827, new_n828, new_n829,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1217, new_n1218;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(G234));
  NAND2_X1  g024(.A1(new_n447), .A2(G2106), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT66), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT67), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  AND2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n462), .A2(G2105), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G137), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  AND2_X1   g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G101), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  XNOR2_X1  g043(.A(KEYINPUT3), .B(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G125), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n465), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n468), .A2(new_n472), .ZN(G160));
  NOR2_X1   g048(.A1(new_n462), .A2(new_n465), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G124), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(new_n476));
  OAI21_X1  g051(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n477));
  INV_X1    g052(.A(G112), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n477), .B1(new_n478), .B2(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n463), .A2(KEYINPUT68), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT68), .ZN(new_n481));
  OAI21_X1  g056(.A(new_n481), .B1(new_n462), .B2(G2105), .ZN(new_n482));
  AND2_X1   g057(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  AOI211_X1 g058(.A(new_n476), .B(new_n479), .C1(new_n483), .C2(G136), .ZN(G162));
  OAI21_X1  g059(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n485));
  INV_X1    g060(.A(G114), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n485), .B1(new_n486), .B2(G2105), .ZN(new_n487));
  AND2_X1   g062(.A1(G126), .A2(G2105), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n488), .B1(new_n460), .B2(new_n461), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT69), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  OAI211_X1 g066(.A(KEYINPUT69), .B(new_n488), .C1(new_n460), .C2(new_n461), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n487), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT70), .ZN(new_n494));
  OAI211_X1 g069(.A(G138), .B(new_n465), .C1(new_n460), .C2(new_n461), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT4), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n469), .A2(new_n497), .A3(G138), .A4(new_n465), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  AND3_X1   g074(.A1(new_n493), .A2(new_n494), .A3(new_n499), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n494), .B1(new_n493), .B2(new_n499), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n500), .A2(new_n501), .ZN(G164));
  NAND2_X1  g077(.A1(G75), .A2(G543), .ZN(new_n503));
  INV_X1    g078(.A(G543), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT5), .ZN(new_n505));
  OAI21_X1  g080(.A(new_n504), .B1(new_n505), .B2(KEYINPUT72), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT72), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n507), .A2(KEYINPUT5), .A3(G543), .ZN(new_n508));
  AND2_X1   g083(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(G62), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n503), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G651), .ZN(new_n512));
  INV_X1    g087(.A(G651), .ZN(new_n513));
  OAI21_X1  g088(.A(KEYINPUT71), .B1(new_n513), .B2(KEYINPUT6), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT71), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT6), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n515), .A2(new_n516), .A3(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n514), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n513), .A2(KEYINPUT6), .ZN(new_n519));
  AND2_X1   g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n506), .A2(new_n508), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(G88), .ZN(new_n523));
  INV_X1    g098(.A(G50), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n520), .A2(G543), .ZN(new_n525));
  OAI221_X1 g100(.A(new_n512), .B1(new_n522), .B2(new_n523), .C1(new_n524), .C2(new_n525), .ZN(G303));
  INV_X1    g101(.A(G303), .ZN(G166));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n528), .B(KEYINPUT73), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n529), .B(KEYINPUT7), .ZN(new_n530));
  INV_X1    g105(.A(G89), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n530), .B1(new_n531), .B2(new_n522), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n521), .A2(G63), .A3(G651), .ZN(new_n533));
  INV_X1    g108(.A(G51), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n533), .B1(new_n525), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n532), .A2(new_n535), .ZN(G168));
  AOI22_X1  g111(.A1(new_n521), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  OR2_X1    g112(.A1(new_n537), .A2(new_n513), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n518), .A2(new_n519), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n539), .A2(new_n504), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G52), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n539), .A2(new_n509), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G90), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n538), .A2(new_n541), .A3(new_n543), .ZN(G301));
  INV_X1    g119(.A(G301), .ZN(G171));
  AOI22_X1  g120(.A1(new_n521), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n546));
  OR2_X1    g121(.A1(new_n546), .A2(new_n513), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n540), .A2(G43), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n542), .A2(G81), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  NAND4_X1  g127(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g128(.A(KEYINPUT74), .B(KEYINPUT8), .Z(new_n554));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n554), .B(new_n555), .ZN(new_n556));
  NAND4_X1  g131(.A1(G319), .A2(G483), .A3(G661), .A4(new_n556), .ZN(G188));
  NAND2_X1  g132(.A1(G78), .A2(G543), .ZN(new_n558));
  INV_X1    g133(.A(G65), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n558), .B1(new_n509), .B2(new_n559), .ZN(new_n560));
  AOI22_X1  g135(.A1(G91), .A2(new_n542), .B1(new_n560), .B2(G651), .ZN(new_n561));
  NAND4_X1  g136(.A1(new_n518), .A2(G53), .A3(G543), .A4(new_n519), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT9), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n561), .A2(new_n563), .ZN(G299));
  OR2_X1    g139(.A1(new_n532), .A2(new_n535), .ZN(G286));
  NAND2_X1  g140(.A1(new_n540), .A2(G49), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n542), .A2(G87), .ZN(new_n567));
  OAI21_X1  g142(.A(G651), .B1(new_n521), .B2(G74), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(G288));
  NAND2_X1  g144(.A1(new_n521), .A2(G61), .ZN(new_n570));
  NAND2_X1  g145(.A1(G73), .A2(G543), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(G651), .ZN(new_n573));
  NAND4_X1  g148(.A1(new_n518), .A2(new_n521), .A3(G86), .A4(new_n519), .ZN(new_n574));
  NAND4_X1  g149(.A1(new_n518), .A2(G48), .A3(G543), .A4(new_n519), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(G305));
  AOI22_X1  g151(.A1(new_n521), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n577));
  OR2_X1    g152(.A1(new_n577), .A2(new_n513), .ZN(new_n578));
  XNOR2_X1  g153(.A(KEYINPUT75), .B(G85), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n542), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n540), .A2(G47), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n578), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT76), .ZN(new_n583));
  OR2_X1    g158(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n582), .A2(new_n583), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(new_n585), .ZN(G290));
  INV_X1    g161(.A(G868), .ZN(new_n587));
  NOR2_X1   g162(.A1(G301), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n542), .A2(G92), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT10), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n589), .B(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(G79), .A2(G543), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n592), .B(KEYINPUT77), .ZN(new_n593));
  INV_X1    g168(.A(G66), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n509), .B2(new_n594), .ZN(new_n595));
  AOI22_X1  g170(.A1(G54), .A2(new_n540), .B1(new_n595), .B2(G651), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n591), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT78), .ZN(new_n598));
  XNOR2_X1  g173(.A(new_n597), .B(new_n598), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n588), .B1(new_n599), .B2(new_n587), .ZN(G284));
  XOR2_X1   g175(.A(G284), .B(KEYINPUT79), .Z(G321));
  NAND2_X1  g176(.A1(G299), .A2(new_n587), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n602), .B1(G168), .B2(new_n587), .ZN(G297));
  OAI21_X1  g178(.A(new_n602), .B1(G168), .B2(new_n587), .ZN(G280));
  INV_X1    g179(.A(G559), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n599), .B1(new_n605), .B2(G860), .ZN(G148));
  NAND2_X1  g181(.A1(new_n550), .A2(new_n587), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n597), .B(KEYINPUT78), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n608), .A2(G559), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n607), .B1(new_n609), .B2(new_n587), .ZN(G323));
  XOR2_X1   g185(.A(KEYINPUT80), .B(KEYINPUT11), .Z(new_n611));
  XNOR2_X1  g186(.A(G323), .B(new_n611), .ZN(G282));
  NAND2_X1  g187(.A1(new_n483), .A2(G135), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n474), .A2(G123), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n465), .A2(G111), .ZN(new_n615));
  OAI21_X1  g190(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n616));
  OAI211_X1 g191(.A(new_n613), .B(new_n614), .C1(new_n615), .C2(new_n616), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT82), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(G2096), .ZN(new_n619));
  NAND2_X1  g194(.A1(KEYINPUT81), .A2(G2100), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n469), .A2(new_n466), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT12), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT13), .ZN(new_n623));
  NOR2_X1   g198(.A1(KEYINPUT81), .A2(G2100), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n620), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  OAI211_X1 g200(.A(new_n619), .B(new_n625), .C1(new_n623), .C2(new_n620), .ZN(G156));
  INV_X1    g201(.A(G14), .ZN(new_n627));
  XNOR2_X1  g202(.A(G2427), .B(G2438), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2430), .ZN(new_n629));
  XNOR2_X1  g204(.A(KEYINPUT15), .B(G2435), .ZN(new_n630));
  OR2_X1    g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n629), .A2(new_n630), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n631), .A2(KEYINPUT14), .A3(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2451), .B(G2454), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT16), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n633), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2443), .B(G2446), .ZN(new_n637));
  OR2_X1    g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n636), .A2(new_n637), .ZN(new_n639));
  AND2_X1   g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(G1341), .B(G1348), .ZN(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n627), .B1(new_n640), .B2(new_n642), .ZN(new_n643));
  INV_X1    g218(.A(KEYINPUT83), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n638), .A2(new_n639), .ZN(new_n645));
  AOI21_X1  g220(.A(new_n644), .B1(new_n645), .B2(new_n641), .ZN(new_n646));
  AOI211_X1 g221(.A(KEYINPUT83), .B(new_n642), .C1(new_n638), .C2(new_n639), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n643), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(G401));
  XOR2_X1   g224(.A(KEYINPUT84), .B(KEYINPUT18), .Z(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(G2084), .B(G2090), .Z(new_n652));
  XNOR2_X1  g227(.A(G2067), .B(G2678), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n654), .A2(KEYINPUT17), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n652), .A2(new_n653), .ZN(new_n656));
  OAI21_X1  g231(.A(new_n651), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G2072), .B(G2078), .Z(new_n658));
  AOI21_X1  g233(.A(new_n658), .B1(new_n654), .B2(new_n650), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n657), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2096), .B(G2100), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n660), .B(new_n661), .Z(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(G227));
  XNOR2_X1  g238(.A(G1981), .B(G1986), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1956), .B(G2474), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1961), .B(G1966), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n666), .A2(new_n667), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(KEYINPUT85), .B(KEYINPUT19), .Z(new_n671));
  XNOR2_X1  g246(.A(G1971), .B(G1976), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  MUX2_X1   g248(.A(new_n670), .B(new_n669), .S(new_n673), .Z(new_n674));
  NAND2_X1  g249(.A1(new_n668), .A2(KEYINPUT86), .ZN(new_n675));
  OR3_X1    g250(.A1(new_n666), .A2(new_n667), .A3(KEYINPUT86), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n673), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(KEYINPUT87), .B(KEYINPUT20), .Z(new_n678));
  OR2_X1    g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n677), .A2(new_n678), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n674), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT88), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n681), .B(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(G1991), .B(G1996), .Z(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  AND2_X1   g261(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n684), .A2(new_n686), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n665), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  OR2_X1    g264(.A1(new_n684), .A2(new_n686), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n684), .A2(new_n686), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n690), .A2(new_n664), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(G229));
  INV_X1    g269(.A(G29), .ZN(new_n695));
  AND2_X1   g270(.A1(new_n695), .A2(G32), .ZN(new_n696));
  AND2_X1   g271(.A1(new_n483), .A2(G141), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n466), .A2(G105), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT93), .ZN(new_n699));
  NAND3_X1  g274(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n700));
  XOR2_X1   g275(.A(new_n700), .B(KEYINPUT26), .Z(new_n701));
  NAND2_X1  g276(.A1(new_n474), .A2(G129), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n699), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  OR2_X1    g278(.A1(new_n697), .A2(new_n703), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n696), .B1(new_n704), .B2(G29), .ZN(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT27), .B(G1996), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT94), .ZN(new_n707));
  INV_X1    g282(.A(KEYINPUT24), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n695), .B1(new_n708), .B2(G34), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n709), .B1(new_n708), .B2(G34), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n710), .B1(G160), .B2(G29), .ZN(new_n711));
  AOI22_X1  g286(.A1(new_n705), .A2(new_n707), .B1(G2084), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n695), .A2(G33), .ZN(new_n713));
  AND3_X1   g288(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT25), .ZN(new_n715));
  AOI22_X1  g290(.A1(new_n469), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n715), .B1(new_n716), .B2(new_n465), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(new_n483), .B2(G139), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n713), .B1(new_n718), .B2(new_n695), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(G2072), .Z(new_n720));
  NAND2_X1  g295(.A1(new_n712), .A2(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(KEYINPUT95), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(G1961), .ZN(new_n724));
  INV_X1    g299(.A(G16), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n725), .A2(G5), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G171), .B2(new_n725), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(KEYINPUT97), .Z(new_n728));
  AOI21_X1  g303(.A(new_n723), .B1(new_n724), .B2(new_n728), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n617), .A2(new_n695), .ZN(new_n730));
  INV_X1    g305(.A(G28), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n731), .A2(KEYINPUT30), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT96), .Z(new_n733));
  AOI211_X1 g308(.A(G29), .B(new_n733), .C1(KEYINPUT30), .C2(new_n731), .ZN(new_n734));
  XOR2_X1   g309(.A(KEYINPUT31), .B(G11), .Z(new_n735));
  NOR3_X1   g310(.A1(new_n730), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  OAI221_X1 g311(.A(new_n736), .B1(G2084), .B2(new_n711), .C1(new_n705), .C2(new_n707), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n725), .A2(G21), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(G168), .B2(new_n725), .ZN(new_n739));
  AND2_X1   g314(.A1(new_n739), .A2(G1966), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n695), .A2(G27), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(G164), .B2(new_n695), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(G2078), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n739), .A2(G1966), .ZN(new_n744));
  NOR4_X1   g319(.A1(new_n737), .A2(new_n740), .A3(new_n743), .A4(new_n744), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n728), .A2(new_n724), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(new_n722), .B2(new_n721), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n729), .A2(new_n745), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n748), .A2(KEYINPUT98), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT90), .ZN(new_n750));
  OR3_X1    g325(.A1(new_n750), .A2(G4), .A3(G16), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n750), .B1(G4), .B2(G16), .ZN(new_n752));
  OAI211_X1 g327(.A(new_n751), .B(new_n752), .C1(new_n608), .C2(new_n725), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(G1348), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n725), .A2(G20), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT23), .Z(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(G299), .B2(G16), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(G1956), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n695), .A2(G35), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G162), .B2(new_n695), .ZN(new_n760));
  XNOR2_X1  g335(.A(KEYINPUT29), .B(G2090), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  NOR2_X1   g337(.A1(G16), .A2(G19), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(new_n551), .B2(G16), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n762), .B1(G1341), .B2(new_n764), .ZN(new_n765));
  AND3_X1   g340(.A1(new_n695), .A2(KEYINPUT28), .A3(G26), .ZN(new_n766));
  AOI21_X1  g341(.A(KEYINPUT28), .B1(new_n695), .B2(G26), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n474), .A2(G128), .ZN(new_n768));
  OR2_X1    g343(.A1(new_n768), .A2(KEYINPUT91), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n768), .A2(KEYINPUT91), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n483), .A2(G140), .ZN(new_n772));
  OAI21_X1  g347(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n773));
  INV_X1    g348(.A(G116), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n773), .B1(new_n774), .B2(G2105), .ZN(new_n775));
  INV_X1    g350(.A(new_n775), .ZN(new_n776));
  NAND3_X1  g351(.A1(new_n771), .A2(new_n772), .A3(new_n776), .ZN(new_n777));
  AOI211_X1 g352(.A(new_n766), .B(new_n767), .C1(new_n777), .C2(G29), .ZN(new_n778));
  XOR2_X1   g353(.A(KEYINPUT92), .B(G2067), .Z(new_n779));
  INV_X1    g354(.A(new_n779), .ZN(new_n780));
  AND2_X1   g355(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n778), .A2(new_n780), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n764), .A2(G1341), .ZN(new_n783));
  NOR3_X1   g358(.A1(new_n781), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  AND4_X1   g359(.A1(new_n754), .A2(new_n758), .A3(new_n765), .A4(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(KEYINPUT98), .ZN(new_n786));
  NAND4_X1  g361(.A1(new_n729), .A2(new_n786), .A3(new_n745), .A4(new_n747), .ZN(new_n787));
  AND3_X1   g362(.A1(new_n749), .A2(new_n785), .A3(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n725), .A2(G24), .ZN(new_n789));
  AND2_X1   g364(.A1(new_n584), .A2(new_n585), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n789), .B1(new_n790), .B2(new_n725), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT89), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n792), .A2(G1986), .ZN(new_n793));
  OR2_X1    g368(.A1(new_n791), .A2(KEYINPUT89), .ZN(new_n794));
  INV_X1    g369(.A(G1986), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n791), .A2(KEYINPUT89), .ZN(new_n796));
  NAND3_X1  g371(.A1(new_n794), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n483), .A2(G131), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n474), .A2(G119), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n465), .A2(G107), .ZN(new_n800));
  OAI21_X1  g375(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n801));
  OAI211_X1 g376(.A(new_n798), .B(new_n799), .C1(new_n800), .C2(new_n801), .ZN(new_n802));
  MUX2_X1   g377(.A(G25), .B(new_n802), .S(G29), .Z(new_n803));
  XOR2_X1   g378(.A(KEYINPUT35), .B(G1991), .Z(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  NAND3_X1  g380(.A1(new_n793), .A2(new_n797), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n725), .A2(G22), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(G166), .B2(new_n725), .ZN(new_n808));
  INV_X1    g383(.A(G1971), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  NOR2_X1   g385(.A1(G6), .A2(G16), .ZN(new_n811));
  INV_X1    g386(.A(G305), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n811), .B1(new_n812), .B2(G16), .ZN(new_n813));
  XOR2_X1   g388(.A(KEYINPUT32), .B(G1981), .Z(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n725), .A2(G23), .ZN(new_n816));
  AND3_X1   g391(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n816), .B1(new_n817), .B2(new_n725), .ZN(new_n818));
  XNOR2_X1  g393(.A(KEYINPUT33), .B(G1976), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n810), .A2(new_n815), .A3(new_n820), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT34), .ZN(new_n822));
  OR3_X1    g397(.A1(new_n806), .A2(new_n822), .A3(KEYINPUT36), .ZN(new_n823));
  OAI21_X1  g398(.A(KEYINPUT36), .B1(new_n806), .B2(new_n822), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  AND2_X1   g400(.A1(new_n788), .A2(new_n825), .ZN(G311));
  INV_X1    g401(.A(KEYINPUT99), .ZN(new_n827));
  AND3_X1   g402(.A1(new_n788), .A2(new_n827), .A3(new_n825), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n827), .B1(new_n788), .B2(new_n825), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n828), .A2(new_n829), .ZN(G150));
  NAND2_X1  g405(.A1(new_n599), .A2(G559), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT38), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  AOI22_X1  g408(.A1(new_n521), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n834));
  OR2_X1    g409(.A1(new_n834), .A2(new_n513), .ZN(new_n835));
  AOI22_X1  g410(.A1(G55), .A2(new_n540), .B1(new_n542), .B2(G93), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n836), .A2(KEYINPUT100), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n540), .A2(G55), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n542), .A2(G93), .ZN(new_n839));
  AND3_X1   g414(.A1(new_n838), .A2(new_n839), .A3(KEYINPUT100), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n835), .B1(new_n837), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n841), .A2(new_n550), .ZN(new_n842));
  OAI211_X1 g417(.A(new_n551), .B(new_n835), .C1(new_n837), .C2(new_n840), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n833), .B(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT39), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(G860), .ZN(new_n849));
  OR2_X1    g424(.A1(new_n833), .A2(new_n845), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n833), .A2(new_n845), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n850), .A2(KEYINPUT39), .A3(new_n851), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n848), .A2(new_n849), .A3(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n841), .A2(G860), .ZN(new_n854));
  XOR2_X1   g429(.A(KEYINPUT101), .B(KEYINPUT37), .Z(new_n855));
  XNOR2_X1  g430(.A(new_n854), .B(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n853), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n857), .A2(KEYINPUT102), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT102), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n853), .A2(new_n859), .A3(new_n856), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n858), .A2(new_n860), .ZN(G145));
  XNOR2_X1  g436(.A(new_n617), .B(G160), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(G162), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n474), .A2(G130), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT104), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n864), .B(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n483), .A2(G142), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n465), .A2(G118), .ZN(new_n868));
  OAI21_X1  g443(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n869));
  OAI211_X1 g444(.A(new_n866), .B(new_n867), .C1(new_n868), .C2(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n718), .A2(KEYINPUT103), .ZN(new_n871));
  XOR2_X1   g446(.A(new_n870), .B(new_n871), .Z(new_n872));
  NAND2_X1  g447(.A1(new_n493), .A2(new_n499), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n777), .A2(new_n873), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n697), .A2(new_n703), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n775), .B1(new_n769), .B2(new_n770), .ZN(new_n876));
  INV_X1    g451(.A(new_n873), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n876), .A2(new_n877), .A3(new_n772), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n874), .A2(new_n875), .A3(new_n878), .ZN(new_n879));
  OR2_X1    g454(.A1(new_n718), .A2(KEYINPUT103), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n875), .B1(new_n874), .B2(new_n878), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n872), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n802), .B(new_n622), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n870), .B(new_n871), .ZN(new_n885));
  INV_X1    g460(.A(new_n878), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n877), .B1(new_n876), .B2(new_n772), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n704), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND4_X1  g463(.A1(new_n885), .A2(new_n888), .A3(new_n880), .A4(new_n879), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n883), .A2(new_n884), .A3(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT105), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n884), .B1(new_n883), .B2(new_n889), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n863), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(G37), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n883), .A2(new_n889), .ZN(new_n896));
  INV_X1    g471(.A(new_n884), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n863), .ZN(new_n899));
  NAND4_X1  g474(.A1(new_n898), .A2(new_n891), .A3(new_n899), .A4(new_n890), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n894), .A2(new_n895), .A3(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g477(.A1(new_n790), .A2(G305), .ZN(new_n903));
  XNOR2_X1  g478(.A(G303), .B(G288), .ZN(new_n904));
  AOI21_X1  g479(.A(G305), .B1(new_n584), .B2(new_n585), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n903), .A2(new_n904), .A3(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(new_n904), .ZN(new_n908));
  NOR2_X1   g483(.A1(G290), .A2(new_n812), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n908), .B1(new_n909), .B2(new_n905), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n907), .A2(new_n910), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n609), .A2(new_n844), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n599), .A2(new_n605), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n913), .A2(new_n845), .ZN(new_n914));
  INV_X1    g489(.A(G299), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n591), .A2(new_n915), .A3(new_n596), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n915), .B1(new_n591), .B2(new_n596), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NOR3_X1   g494(.A1(new_n912), .A2(new_n914), .A3(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT41), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n921), .B1(new_n917), .B2(new_n918), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n597), .A2(G299), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n923), .A2(KEYINPUT41), .A3(new_n916), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n609), .A2(new_n844), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n913), .A2(new_n845), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n926), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NOR3_X1   g504(.A1(new_n920), .A2(new_n929), .A3(KEYINPUT42), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT42), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n925), .B1(new_n912), .B2(new_n914), .ZN(new_n932));
  OAI211_X1 g507(.A(new_n927), .B(new_n928), .C1(new_n918), .C2(new_n917), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n931), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n911), .B1(new_n930), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g510(.A(KEYINPUT42), .B1(new_n920), .B2(new_n929), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n932), .A2(new_n933), .A3(new_n931), .ZN(new_n937));
  INV_X1    g512(.A(new_n911), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n936), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n587), .B1(new_n935), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n841), .A2(new_n587), .ZN(new_n941));
  INV_X1    g516(.A(new_n941), .ZN(new_n942));
  OAI21_X1  g517(.A(KEYINPUT106), .B1(new_n940), .B2(new_n942), .ZN(new_n943));
  NOR3_X1   g518(.A1(new_n930), .A2(new_n934), .A3(new_n911), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n938), .B1(new_n936), .B2(new_n937), .ZN(new_n945));
  OAI21_X1  g520(.A(G868), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT106), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n946), .A2(new_n947), .A3(new_n941), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n943), .A2(new_n948), .ZN(G295));
  NAND2_X1  g524(.A1(new_n946), .A2(new_n941), .ZN(G331));
  NAND2_X1  g525(.A1(G286), .A2(G301), .ZN(new_n951));
  NAND2_X1  g526(.A1(G168), .A2(G171), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n844), .A2(new_n953), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n842), .A2(new_n843), .A3(new_n951), .A4(new_n952), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n954), .A2(new_n919), .A3(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(new_n955), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT107), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n954), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n844), .A2(new_n953), .A3(KEYINPUT107), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n957), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n956), .B1(new_n961), .B2(new_n925), .ZN(new_n962));
  AOI21_X1  g537(.A(G37), .B1(new_n962), .B2(new_n938), .ZN(new_n963));
  OAI211_X1 g538(.A(new_n911), .B(new_n956), .C1(new_n961), .C2(new_n925), .ZN(new_n964));
  AOI21_X1  g539(.A(KEYINPUT43), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n955), .A2(new_n919), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n966), .B1(new_n959), .B2(new_n960), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n925), .B1(new_n955), .B2(new_n954), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n938), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n964), .A2(new_n969), .A3(new_n895), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT43), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  OAI21_X1  g547(.A(KEYINPUT44), .B1(new_n965), .B2(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n971), .B1(new_n963), .B2(new_n964), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n964), .A2(new_n969), .A3(new_n971), .A4(new_n895), .ZN(new_n975));
  INV_X1    g550(.A(new_n975), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n973), .B1(new_n977), .B2(KEYINPUT44), .ZN(G397));
  AOI21_X1  g553(.A(G1384), .B1(new_n493), .B2(new_n499), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n979), .A2(KEYINPUT45), .ZN(new_n980));
  INV_X1    g555(.A(G40), .ZN(new_n981));
  NOR3_X1   g556(.A1(new_n468), .A2(new_n472), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n983), .A2(G1996), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(new_n875), .ZN(new_n985));
  OR2_X1    g560(.A1(new_n985), .A2(KEYINPUT108), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(KEYINPUT108), .ZN(new_n987));
  INV_X1    g562(.A(G2067), .ZN(new_n988));
  XNOR2_X1  g563(.A(new_n777), .B(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(G1996), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n989), .B1(new_n990), .B2(new_n875), .ZN(new_n991));
  INV_X1    g566(.A(new_n983), .ZN(new_n992));
  AOI22_X1  g567(.A1(new_n986), .A2(new_n987), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(new_n804), .ZN(new_n994));
  AND2_X1   g569(.A1(new_n802), .A2(new_n994), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n802), .A2(new_n994), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n992), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  AND2_X1   g572(.A1(new_n993), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n790), .A2(new_n795), .A3(new_n992), .ZN(new_n999));
  XNOR2_X1  g574(.A(new_n999), .B(KEYINPUT48), .ZN(new_n1000));
  AND2_X1   g575(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n984), .A2(KEYINPUT46), .ZN(new_n1002));
  XNOR2_X1  g577(.A(new_n1002), .B(KEYINPUT124), .ZN(new_n1003));
  AND2_X1   g578(.A1(new_n989), .A2(new_n875), .ZN(new_n1004));
  OAI221_X1 g579(.A(new_n1003), .B1(KEYINPUT46), .B2(new_n984), .C1(new_n983), .C2(new_n1004), .ZN(new_n1005));
  XOR2_X1   g580(.A(KEYINPUT125), .B(KEYINPUT47), .Z(new_n1006));
  XNOR2_X1  g581(.A(new_n1005), .B(new_n1006), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n777), .A2(G2067), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1008), .B1(new_n993), .B2(new_n996), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT123), .ZN(new_n1010));
  OR2_X1    g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n983), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1012));
  AOI211_X1 g587(.A(new_n1001), .B(new_n1007), .C1(new_n1011), .C2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n574), .A2(new_n575), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n513), .B1(new_n570), .B2(new_n571), .ZN(new_n1015));
  OAI21_X1  g590(.A(G1981), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  OR2_X1    g591(.A1(new_n1016), .A2(KEYINPUT111), .ZN(new_n1017));
  XNOR2_X1  g592(.A(KEYINPUT110), .B(G1981), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n573), .A2(new_n574), .A3(new_n575), .A4(new_n1018), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1019), .A2(KEYINPUT111), .A3(new_n1016), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT49), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1017), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(G1384), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n873), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n470), .A2(new_n471), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(G2105), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n1026), .A2(G40), .A3(new_n467), .A4(new_n464), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1024), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(G8), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1022), .A2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1021), .B1(new_n1017), .B2(new_n1020), .ZN(new_n1032));
  OR2_X1    g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NOR2_X1   g608(.A1(G288), .A2(G1976), .ZN(new_n1034));
  AOI22_X1  g609(.A1(new_n1033), .A2(new_n1034), .B1(new_n812), .B2(new_n1018), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT113), .ZN(new_n1036));
  AND2_X1   g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1030), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n817), .A2(G1976), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n982), .A2(new_n979), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1039), .A2(new_n1040), .A3(G8), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(KEYINPUT52), .ZN(new_n1042));
  INV_X1    g617(.A(G1976), .ZN(new_n1043));
  AOI21_X1  g618(.A(KEYINPUT52), .B1(G288), .B2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1030), .A2(new_n1039), .A3(new_n1044), .ZN(new_n1045));
  OAI211_X1 g620(.A(new_n1042), .B(new_n1045), .C1(new_n1031), .C2(new_n1032), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT112), .ZN(new_n1047));
  AND2_X1   g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1023), .B1(new_n500), .B2(new_n501), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT45), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1027), .B1(new_n979), .B2(KEYINPUT45), .ZN(new_n1054));
  AOI21_X1  g629(.A(G1971), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1055), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n982), .B1(new_n1024), .B2(KEYINPUT50), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1057), .B1(KEYINPUT50), .B2(new_n1051), .ZN(new_n1058));
  XNOR2_X1  g633(.A(KEYINPUT109), .B(G2090), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1029), .B1(new_n1056), .B2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(G303), .A2(G8), .ZN(new_n1062));
  XNOR2_X1  g637(.A(new_n1062), .B(KEYINPUT55), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1061), .A2(new_n1064), .ZN(new_n1065));
  OAI22_X1  g640(.A1(new_n1037), .A2(new_n1038), .B1(new_n1050), .B2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1046), .B1(new_n1061), .B2(new_n1064), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT50), .ZN(new_n1068));
  OAI211_X1 g643(.A(new_n1068), .B(new_n1023), .C1(new_n500), .C2(new_n501), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1027), .B1(new_n1024), .B2(KEYINPUT50), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1069), .A2(new_n1070), .A3(new_n1059), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n873), .A2(KEYINPUT45), .A3(new_n1023), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(new_n982), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1073), .B1(new_n1052), .B2(new_n1051), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1071), .B1(new_n1074), .B2(G1971), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT114), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1029), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  OAI211_X1 g652(.A(new_n1071), .B(KEYINPUT114), .C1(new_n1074), .C2(G1971), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1064), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT115), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1067), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  AND3_X1   g656(.A1(new_n1069), .A2(new_n1070), .A3(new_n1059), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1076), .B1(new_n1055), .B2(new_n1082), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1083), .A2(G8), .A3(new_n1078), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(new_n1063), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1085), .A2(KEYINPUT115), .ZN(new_n1086));
  XNOR2_X1  g661(.A(KEYINPUT122), .B(KEYINPUT53), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1074), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1087), .B1(new_n1088), .B2(G2078), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1027), .B1(new_n1024), .B2(new_n1052), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1090), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT53), .ZN(new_n1092));
  OR3_X1    g667(.A1(new_n1091), .A2(new_n1092), .A3(G2078), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1027), .B1(new_n979), .B2(new_n1068), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n873), .A2(KEYINPUT70), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n493), .A2(new_n494), .A3(new_n499), .ZN(new_n1096));
  AOI21_X1  g671(.A(G1384), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1094), .B1(new_n1097), .B2(new_n1068), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(KEYINPUT116), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT116), .ZN(new_n1100));
  OAI211_X1 g675(.A(new_n1100), .B(new_n1094), .C1(new_n1097), .C2(new_n1068), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1102));
  OAI211_X1 g677(.A(new_n1089), .B(new_n1093), .C1(new_n1102), .C2(G1961), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(G171), .ZN(new_n1104));
  NOR3_X1   g679(.A1(new_n1081), .A2(new_n1086), .A3(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT62), .ZN(new_n1106));
  INV_X1    g681(.A(G2084), .ZN(new_n1107));
  INV_X1    g682(.A(G1966), .ZN(new_n1108));
  AOI22_X1  g683(.A1(new_n1058), .A2(new_n1107), .B1(new_n1091), .B2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1029), .B1(new_n1109), .B2(G168), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT51), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1091), .A2(new_n1108), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1114), .B1(G2084), .B2(new_n1098), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(G286), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1111), .B1(new_n1110), .B2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1106), .B1(new_n1113), .B2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g693(.A(G8), .B1(new_n1115), .B2(G286), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1109), .A2(G168), .ZN(new_n1120));
  OAI21_X1  g695(.A(KEYINPUT51), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1121), .A2(KEYINPUT62), .A3(new_n1112), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1118), .A2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1066), .B1(new_n1105), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1085), .A2(KEYINPUT115), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1126));
  NOR3_X1   g701(.A1(new_n1109), .A2(new_n1029), .A3(G286), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1125), .A2(new_n1126), .A3(new_n1067), .A4(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT63), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1050), .ZN(new_n1131));
  OR2_X1    g706(.A1(new_n1061), .A2(new_n1064), .ZN(new_n1132));
  AND2_X1   g707(.A1(new_n1127), .A2(KEYINPUT63), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1131), .A2(new_n1065), .A3(new_n1132), .A4(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1130), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1124), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1137));
  INV_X1    g712(.A(G1956), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT57), .ZN(new_n1140));
  XNOR2_X1  g715(.A(G299), .B(new_n1140), .ZN(new_n1141));
  XNOR2_X1  g716(.A(KEYINPUT56), .B(G2072), .ZN(new_n1142));
  OAI211_X1 g717(.A(new_n1054), .B(new_n1142), .C1(new_n1097), .C2(KEYINPUT45), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1139), .A2(new_n1141), .A3(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(G1348), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1099), .A2(new_n1145), .A3(new_n1101), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1028), .A2(new_n988), .ZN(new_n1147));
  AND2_X1   g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g723(.A(KEYINPUT117), .B1(new_n1148), .B2(new_n597), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1139), .A2(new_n1143), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1141), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1149), .A2(new_n1152), .ZN(new_n1153));
  NOR3_X1   g728(.A1(new_n1148), .A2(KEYINPUT117), .A3(new_n597), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1144), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1148), .A2(KEYINPUT120), .A3(KEYINPUT60), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1146), .A2(KEYINPUT60), .A3(new_n1147), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT120), .ZN(new_n1158));
  AND3_X1   g733(.A1(new_n1157), .A2(new_n1158), .A3(new_n597), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n597), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1156), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT121), .ZN(new_n1162));
  OR2_X1    g737(.A1(new_n1148), .A2(KEYINPUT60), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1161), .A2(new_n1162), .A3(new_n1163), .ZN(new_n1164));
  NOR2_X1   g739(.A1(KEYINPUT118), .A2(KEYINPUT59), .ZN(new_n1165));
  INV_X1    g740(.A(new_n1165), .ZN(new_n1166));
  OAI211_X1 g741(.A(new_n990), .B(new_n1054), .C1(new_n1097), .C2(KEYINPUT45), .ZN(new_n1167));
  XOR2_X1   g742(.A(KEYINPUT58), .B(G1341), .Z(new_n1168));
  NAND2_X1  g743(.A1(new_n1040), .A2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1167), .A2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(KEYINPUT118), .A2(KEYINPUT59), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n551), .A2(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1172), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1166), .B1(new_n1170), .B2(new_n1173), .ZN(new_n1174));
  AOI211_X1 g749(.A(new_n1165), .B(new_n1172), .C1(new_n1167), .C2(new_n1169), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT61), .ZN(new_n1177));
  AND3_X1   g752(.A1(new_n1139), .A2(new_n1141), .A3(new_n1143), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1141), .B1(new_n1139), .B2(new_n1143), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1177), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1152), .A2(KEYINPUT61), .A3(new_n1144), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1176), .A2(new_n1180), .A3(new_n1181), .ZN(new_n1182));
  XNOR2_X1  g757(.A(new_n1182), .B(KEYINPUT119), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1164), .A2(new_n1183), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1162), .B1(new_n1161), .B2(new_n1163), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1155), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  XNOR2_X1  g761(.A(G301), .B(KEYINPUT54), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1103), .A2(new_n1187), .ZN(new_n1188));
  AOI211_X1 g763(.A(new_n1092), .B(G2078), .C1(new_n979), .C2(KEYINPUT45), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n1187), .B1(new_n1090), .B2(new_n1189), .ZN(new_n1190));
  OAI211_X1 g765(.A(new_n1089), .B(new_n1190), .C1(new_n1102), .C2(G1961), .ZN(new_n1191));
  OAI211_X1 g766(.A(new_n1188), .B(new_n1191), .C1(new_n1113), .C2(new_n1117), .ZN(new_n1192));
  NOR3_X1   g767(.A1(new_n1192), .A2(new_n1086), .A3(new_n1081), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1136), .B1(new_n1186), .B2(new_n1193), .ZN(new_n1194));
  XNOR2_X1  g769(.A(G290), .B(new_n795), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n998), .B1(new_n983), .B2(new_n1195), .ZN(new_n1196));
  OAI21_X1  g771(.A(new_n1013), .B1(new_n1194), .B2(new_n1196), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g772(.A1(new_n662), .A2(G319), .ZN(new_n1199));
  XOR2_X1   g773(.A(new_n1199), .B(KEYINPUT126), .Z(new_n1200));
  AND3_X1   g774(.A1(new_n648), .A2(new_n693), .A3(new_n1200), .ZN(new_n1201));
  NAND2_X1  g775(.A1(new_n1201), .A2(new_n901), .ZN(new_n1202));
  INV_X1    g776(.A(new_n956), .ZN(new_n1203));
  INV_X1    g777(.A(new_n960), .ZN(new_n1204));
  AOI21_X1  g778(.A(KEYINPUT107), .B1(new_n844), .B2(new_n953), .ZN(new_n1205));
  OAI21_X1  g779(.A(new_n955), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  AOI21_X1  g780(.A(new_n1203), .B1(new_n1206), .B2(new_n926), .ZN(new_n1207));
  OAI21_X1  g781(.A(new_n895), .B1(new_n1207), .B2(new_n911), .ZN(new_n1208));
  INV_X1    g782(.A(new_n964), .ZN(new_n1209));
  OAI21_X1  g783(.A(KEYINPUT43), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  AOI211_X1 g784(.A(KEYINPUT127), .B(new_n1202), .C1(new_n1210), .C2(new_n975), .ZN(new_n1211));
  INV_X1    g785(.A(KEYINPUT127), .ZN(new_n1212));
  NAND2_X1  g786(.A1(new_n1210), .A2(new_n975), .ZN(new_n1213));
  INV_X1    g787(.A(new_n1202), .ZN(new_n1214));
  AOI21_X1  g788(.A(new_n1212), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  NOR2_X1   g789(.A1(new_n1211), .A2(new_n1215), .ZN(G308));
  OAI21_X1  g790(.A(KEYINPUT127), .B1(new_n977), .B2(new_n1202), .ZN(new_n1217));
  NAND3_X1  g791(.A1(new_n1213), .A2(new_n1212), .A3(new_n1214), .ZN(new_n1218));
  NAND2_X1  g792(.A1(new_n1217), .A2(new_n1218), .ZN(G225));
endmodule


