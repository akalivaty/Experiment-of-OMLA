//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 0 1 1 0 1 0 1 1 0 1 0 0 0 0 0 0 0 1 0 1 1 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 1 1 0 0 1 1 1 0 1 1 0 0 0 0 0 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n718, new_n719, new_n720, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n748, new_n749, new_n750, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n811, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n880, new_n882, new_n883, new_n885,
    new_n886, new_n887, new_n888, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n947, new_n948, new_n950, new_n951, new_n953,
    new_n954, new_n955, new_n957, new_n959, new_n960, new_n961, new_n963,
    new_n964, new_n965, new_n966, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n995,
    new_n996;
  INV_X1    g000(.A(KEYINPUT72), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT36), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(KEYINPUT72), .A2(KEYINPUT36), .ZN(new_n205));
  NOR2_X1   g004(.A1(G169gat), .A2(G176gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT66), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  OAI21_X1  g007(.A(KEYINPUT66), .B1(G169gat), .B2(G176gat), .ZN(new_n209));
  AOI21_X1  g008(.A(KEYINPUT26), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(G169gat), .A2(G176gat), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT26), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n211), .B1(new_n206), .B2(new_n212), .ZN(new_n213));
  OR2_X1    g012(.A1(new_n210), .A2(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(KEYINPUT68), .B(KEYINPUT28), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(G190gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n218));
  INV_X1    g017(.A(new_n218), .ZN(new_n219));
  NOR2_X1   g018(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n217), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n216), .A2(new_n221), .A3(KEYINPUT67), .ZN(new_n222));
  NAND2_X1  g021(.A1(G183gat), .A2(G190gat), .ZN(new_n223));
  OR2_X1    g022(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n224));
  AOI21_X1  g023(.A(G190gat), .B1(new_n224), .B2(new_n218), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT67), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n215), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND4_X1  g026(.A1(new_n214), .A2(new_n222), .A3(new_n223), .A4(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n211), .A2(KEYINPUT23), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n229), .B1(G169gat), .B2(G176gat), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT24), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n223), .A2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(G183gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(new_n217), .ZN(new_n234));
  NAND3_X1  g033(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n232), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n230), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT23), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n238), .B1(new_n208), .B2(new_n209), .ZN(new_n239));
  OAI21_X1  g038(.A(KEYINPUT25), .B1(new_n237), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n235), .A2(KEYINPUT64), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(new_n232), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT65), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n234), .A2(new_n243), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n233), .A2(new_n217), .A3(KEYINPUT65), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n223), .A2(KEYINPUT64), .A3(new_n231), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n242), .A2(new_n244), .A3(new_n245), .A4(new_n246), .ZN(new_n247));
  AOI21_X1  g046(.A(KEYINPUT25), .B1(new_n206), .B2(KEYINPUT23), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n247), .A2(new_n230), .A3(new_n248), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n228), .A2(new_n240), .A3(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(G134gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(G127gat), .ZN(new_n252));
  INV_X1    g051(.A(G127gat), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(G134gat), .ZN(new_n254));
  AOI21_X1  g053(.A(KEYINPUT69), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT69), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n256), .B1(G127gat), .B2(new_n251), .ZN(new_n257));
  OAI21_X1  g056(.A(KEYINPUT70), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  XOR2_X1   g057(.A(G113gat), .B(G120gat), .Z(new_n259));
  INV_X1    g058(.A(KEYINPUT1), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT70), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n252), .A2(KEYINPUT69), .ZN(new_n263));
  XNOR2_X1  g062(.A(G127gat), .B(G134gat), .ZN(new_n264));
  OAI211_X1 g063(.A(new_n262), .B(new_n263), .C1(new_n264), .C2(KEYINPUT69), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n258), .A2(new_n261), .A3(new_n265), .ZN(new_n266));
  OR2_X1    g065(.A1(new_n261), .A2(new_n264), .ZN(new_n267));
  AND2_X1   g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n250), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(G227gat), .A2(G233gat), .ZN(new_n270));
  AND2_X1   g069(.A1(new_n249), .A2(new_n240), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n266), .A2(new_n267), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n271), .A2(new_n272), .A3(new_n228), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n269), .A2(new_n270), .A3(new_n273), .ZN(new_n274));
  XOR2_X1   g073(.A(new_n274), .B(KEYINPUT34), .Z(new_n275));
  XNOR2_X1  g074(.A(G15gat), .B(G43gat), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n276), .B(G71gat), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n277), .B(G99gat), .ZN(new_n278));
  AND2_X1   g077(.A1(new_n278), .A2(KEYINPUT71), .ZN(new_n279));
  OAI21_X1  g078(.A(KEYINPUT33), .B1(new_n278), .B2(KEYINPUT71), .ZN(new_n280));
  AND2_X1   g079(.A1(new_n269), .A2(new_n273), .ZN(new_n281));
  OAI221_X1 g080(.A(KEYINPUT32), .B1(new_n279), .B2(new_n280), .C1(new_n281), .C2(new_n270), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT33), .ZN(new_n283));
  OAI22_X1  g082(.A1(new_n281), .A2(new_n270), .B1(KEYINPUT32), .B2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n278), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n275), .A2(new_n282), .A3(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n275), .B1(new_n282), .B2(new_n286), .ZN(new_n289));
  OAI211_X1 g088(.A(new_n204), .B(new_n205), .C1(new_n288), .C2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n275), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n286), .A2(new_n282), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND4_X1  g092(.A1(new_n293), .A2(new_n202), .A3(new_n203), .A4(new_n287), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n290), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(G218gat), .ZN(new_n296));
  INV_X1    g095(.A(G211gat), .ZN(new_n297));
  XNOR2_X1  g096(.A(KEYINPUT73), .B(G211gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(G218gat), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT22), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  XOR2_X1   g100(.A(G197gat), .B(G204gat), .Z(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n297), .B1(new_n301), .B2(new_n303), .ZN(new_n304));
  AOI21_X1  g103(.A(KEYINPUT22), .B1(new_n298), .B2(G218gat), .ZN(new_n305));
  NOR3_X1   g104(.A1(new_n305), .A2(G211gat), .A3(new_n302), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n296), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n301), .A2(new_n297), .A3(new_n303), .ZN(new_n308));
  OAI21_X1  g107(.A(G211gat), .B1(new_n305), .B2(new_n302), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n308), .A2(G218gat), .A3(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n307), .A2(KEYINPUT74), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n307), .A2(new_n310), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT74), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(G226gat), .A2(G233gat), .ZN(new_n315));
  XNOR2_X1  g114(.A(new_n315), .B(KEYINPUT75), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n316), .B(KEYINPUT76), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT29), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n318), .B1(new_n250), .B2(new_n319), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n316), .B1(new_n271), .B2(new_n228), .ZN(new_n321));
  OAI211_X1 g120(.A(new_n311), .B(new_n314), .C1(new_n320), .C2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n249), .A2(new_n240), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n227), .A2(new_n222), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n223), .B1(new_n210), .B2(new_n213), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n319), .B1(new_n323), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(new_n316), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n250), .A2(new_n318), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n328), .A2(new_n312), .A3(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(G8gat), .B(G36gat), .ZN(new_n331));
  INV_X1    g130(.A(G64gat), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n331), .B(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(G92gat), .ZN(new_n334));
  XNOR2_X1  g133(.A(new_n333), .B(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  NAND4_X1  g135(.A1(new_n322), .A2(new_n330), .A3(KEYINPUT30), .A4(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT78), .ZN(new_n338));
  XNOR2_X1  g137(.A(new_n337), .B(new_n338), .ZN(new_n339));
  AND3_X1   g138(.A1(new_n322), .A2(KEYINPUT77), .A3(new_n330), .ZN(new_n340));
  AOI21_X1  g139(.A(KEYINPUT77), .B1(new_n322), .B2(new_n330), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n335), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(KEYINPUT30), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n322), .A2(new_n330), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n344), .A2(new_n335), .ZN(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n339), .B1(new_n343), .B2(new_n346), .ZN(new_n347));
  XNOR2_X1  g146(.A(KEYINPUT0), .B(G57gat), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n348), .B(G85gat), .ZN(new_n349));
  XNOR2_X1  g148(.A(G1gat), .B(G29gat), .ZN(new_n350));
  XOR2_X1   g149(.A(new_n349), .B(new_n350), .Z(new_n351));
  XOR2_X1   g150(.A(G141gat), .B(G148gat), .Z(new_n352));
  INV_X1    g151(.A(G155gat), .ZN(new_n353));
  INV_X1    g152(.A(G162gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(G155gat), .A2(G162gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(KEYINPUT2), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n352), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(G141gat), .B(G148gat), .ZN(new_n360));
  OAI211_X1 g159(.A(new_n356), .B(new_n355), .C1(new_n360), .C2(KEYINPUT2), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n272), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(KEYINPUT80), .ZN(new_n365));
  AOI21_X1  g164(.A(KEYINPUT79), .B1(new_n359), .B2(new_n361), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n359), .A2(new_n361), .A3(KEYINPUT79), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(new_n268), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n362), .B1(new_n266), .B2(new_n267), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT80), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n365), .A2(new_n370), .A3(new_n373), .ZN(new_n374));
  AND2_X1   g173(.A1(G225gat), .A2(G233gat), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n371), .A2(new_n372), .ZN(new_n377));
  AOI211_X1 g176(.A(KEYINPUT80), .B(new_n362), .C1(new_n266), .C2(new_n267), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT4), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n375), .A2(new_n379), .ZN(new_n380));
  NOR3_X1   g179(.A1(new_n377), .A2(new_n378), .A3(new_n380), .ZN(new_n381));
  AND3_X1   g180(.A1(new_n359), .A2(new_n361), .A3(KEYINPUT79), .ZN(new_n382));
  OAI21_X1  g181(.A(KEYINPUT3), .B1(new_n382), .B2(new_n366), .ZN(new_n383));
  OR2_X1    g182(.A1(new_n362), .A2(KEYINPUT3), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n383), .A2(new_n268), .A3(new_n384), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n385), .B1(new_n379), .B2(new_n364), .ZN(new_n386));
  OAI211_X1 g185(.A(new_n376), .B(KEYINPUT5), .C1(new_n381), .C2(new_n386), .ZN(new_n387));
  OAI21_X1  g186(.A(KEYINPUT4), .B1(new_n377), .B2(new_n378), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n375), .A2(KEYINPUT5), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n364), .A2(new_n379), .ZN(new_n390));
  NAND4_X1  g189(.A1(new_n388), .A2(new_n389), .A3(new_n390), .A4(new_n385), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n351), .B1(new_n387), .B2(new_n391), .ZN(new_n392));
  XOR2_X1   g191(.A(KEYINPUT81), .B(KEYINPUT6), .Z(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n387), .A2(new_n391), .A3(new_n351), .ZN(new_n395));
  INV_X1    g194(.A(new_n393), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n394), .B1(new_n397), .B2(new_n392), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n347), .A2(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(KEYINPUT29), .B1(new_n307), .B2(new_n310), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n362), .B1(new_n400), .B2(KEYINPUT3), .ZN(new_n401));
  INV_X1    g200(.A(new_n312), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n384), .A2(new_n319), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(G228gat), .A2(G233gat), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT82), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n384), .A2(new_n408), .A3(new_n319), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n403), .A2(KEYINPUT82), .ZN(new_n410));
  NAND4_X1  g209(.A1(new_n314), .A2(new_n409), .A3(new_n311), .A4(new_n410), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n369), .B1(new_n400), .B2(KEYINPUT3), .ZN(new_n412));
  INV_X1    g211(.A(new_n406), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(G22gat), .ZN(new_n415));
  AND3_X1   g214(.A1(new_n407), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n415), .B1(new_n407), .B2(new_n414), .ZN(new_n417));
  OAI21_X1  g216(.A(KEYINPUT83), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  AND3_X1   g217(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n413), .B1(new_n401), .B2(new_n404), .ZN(new_n420));
  OAI21_X1  g219(.A(G22gat), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT83), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n407), .A2(new_n414), .A3(new_n415), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n421), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  XNOR2_X1  g223(.A(G78gat), .B(G106gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(KEYINPUT31), .B(G50gat), .ZN(new_n426));
  XOR2_X1   g225(.A(new_n425), .B(new_n426), .Z(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n418), .A2(new_n424), .A3(new_n428), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n421), .A2(new_n422), .A3(new_n423), .A4(new_n427), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n295), .B1(new_n399), .B2(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n388), .A2(new_n390), .A3(new_n385), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(new_n375), .ZN(new_n434));
  OR2_X1    g233(.A1(new_n374), .A2(new_n375), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n434), .A2(KEYINPUT39), .A3(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT39), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n433), .A2(new_n437), .A3(new_n375), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n436), .A2(KEYINPUT40), .A3(new_n351), .A4(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT84), .ZN(new_n440));
  AOI211_X1 g239(.A(new_n440), .B(new_n351), .C1(new_n387), .C2(new_n391), .ZN(new_n441));
  OAI21_X1  g240(.A(KEYINPUT5), .B1(new_n381), .B2(new_n386), .ZN(new_n442));
  AND2_X1   g241(.A1(new_n374), .A2(new_n375), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n391), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n351), .ZN(new_n445));
  AOI21_X1  g244(.A(KEYINPUT84), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n439), .B1(new_n441), .B2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  XNOR2_X1  g247(.A(new_n337), .B(KEYINPUT78), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT30), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT77), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n344), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n322), .A2(KEYINPUT77), .A3(new_n330), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n450), .B1(new_n454), .B2(new_n335), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n449), .B1(new_n455), .B2(new_n345), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT85), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT40), .ZN(new_n458));
  AND3_X1   g257(.A1(new_n434), .A2(KEYINPUT39), .A3(new_n435), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n438), .A2(new_n351), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n458), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND4_X1  g260(.A1(new_n448), .A2(new_n456), .A3(new_n457), .A4(new_n461), .ZN(new_n462));
  OAI211_X1 g261(.A(new_n461), .B(new_n439), .C1(new_n446), .C2(new_n441), .ZN(new_n463));
  OAI21_X1  g262(.A(KEYINPUT85), .B1(new_n463), .B2(new_n347), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  OAI211_X1 g264(.A(new_n396), .B(new_n395), .C1(new_n441), .C2(new_n446), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(new_n394), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT38), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n468), .B1(new_n344), .B2(KEYINPUT37), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT37), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n320), .A2(new_n321), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n314), .A2(new_n311), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n328), .A2(new_n329), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(new_n402), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n470), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n335), .B1(new_n469), .B2(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n344), .A2(new_n468), .A3(new_n336), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n470), .B1(new_n452), .B2(new_n453), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n344), .A2(KEYINPUT37), .ZN(new_n481));
  OAI21_X1  g280(.A(KEYINPUT38), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n479), .A2(new_n482), .ZN(new_n483));
  OAI211_X1 g282(.A(new_n430), .B(new_n429), .C1(new_n467), .C2(new_n483), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n432), .B1(new_n465), .B2(new_n484), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n288), .A2(new_n289), .ZN(new_n486));
  AND3_X1   g285(.A1(new_n429), .A2(new_n430), .A3(new_n486), .ZN(new_n487));
  XOR2_X1   g286(.A(KEYINPUT86), .B(KEYINPUT35), .Z(new_n488));
  NAND4_X1  g287(.A1(new_n487), .A2(new_n467), .A3(new_n347), .A4(new_n488), .ZN(new_n489));
  NAND4_X1  g288(.A1(new_n347), .A2(new_n429), .A3(new_n430), .A4(new_n486), .ZN(new_n490));
  INV_X1    g289(.A(new_n398), .ZN(new_n491));
  OAI21_X1  g290(.A(KEYINPUT35), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n485), .A2(new_n493), .ZN(new_n494));
  XOR2_X1   g293(.A(KEYINPUT89), .B(KEYINPUT17), .Z(new_n495));
  INV_X1    g294(.A(KEYINPUT88), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT87), .ZN(new_n497));
  INV_X1    g296(.A(G29gat), .ZN(new_n498));
  INV_X1    g297(.A(G36gat), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n498), .A2(new_n499), .A3(KEYINPUT14), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT14), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n501), .B1(G29gat), .B2(G36gat), .ZN(new_n502));
  NAND2_X1  g301(.A1(G29gat), .A2(G36gat), .ZN(new_n503));
  AND3_X1   g302(.A1(new_n500), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(G50gat), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(G43gat), .ZN(new_n506));
  INV_X1    g305(.A(G43gat), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(G50gat), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n506), .A2(new_n508), .A3(KEYINPUT15), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n497), .B1(new_n504), .B2(new_n509), .ZN(new_n510));
  AND3_X1   g309(.A1(new_n506), .A2(new_n508), .A3(KEYINPUT15), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n500), .A2(new_n502), .A3(new_n503), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n511), .A2(new_n512), .A3(KEYINPUT87), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n506), .A2(new_n508), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT15), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n504), .A2(new_n517), .A3(new_n509), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n496), .B1(new_n514), .B2(new_n518), .ZN(new_n519));
  AND3_X1   g318(.A1(new_n511), .A2(KEYINPUT87), .A3(new_n512), .ZN(new_n520));
  AOI21_X1  g319(.A(KEYINPUT87), .B1(new_n511), .B2(new_n512), .ZN(new_n521));
  OAI211_X1 g320(.A(new_n496), .B(new_n518), .C1(new_n520), .C2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n495), .B1(new_n519), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n514), .A2(KEYINPUT17), .A3(new_n518), .ZN(new_n525));
  AND2_X1   g324(.A1(KEYINPUT98), .A2(KEYINPUT7), .ZN(new_n526));
  NOR2_X1   g325(.A1(KEYINPUT98), .A2(KEYINPUT7), .ZN(new_n527));
  INV_X1    g326(.A(G85gat), .ZN(new_n528));
  OAI22_X1  g327(.A1(new_n526), .A2(new_n527), .B1(new_n528), .B2(new_n334), .ZN(new_n529));
  OR2_X1    g328(.A1(KEYINPUT98), .A2(KEYINPUT7), .ZN(new_n530));
  AND2_X1   g329(.A1(G85gat), .A2(G92gat), .ZN(new_n531));
  NAND2_X1  g330(.A1(KEYINPUT98), .A2(KEYINPUT7), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  AND2_X1   g332(.A1(new_n529), .A2(new_n533), .ZN(new_n534));
  NOR2_X1   g333(.A1(G85gat), .A2(G92gat), .ZN(new_n535));
  AND3_X1   g334(.A1(KEYINPUT99), .A2(G99gat), .A3(G106gat), .ZN(new_n536));
  AOI21_X1  g335(.A(KEYINPUT99), .B1(G99gat), .B2(G106gat), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n535), .B1(new_n538), .B2(KEYINPUT8), .ZN(new_n539));
  XOR2_X1   g338(.A(G99gat), .B(G106gat), .Z(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n534), .A2(new_n539), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(G99gat), .A2(G106gat), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT99), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(KEYINPUT99), .A2(G99gat), .A3(G106gat), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n545), .A2(KEYINPUT8), .A3(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(new_n535), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n547), .A2(new_n529), .A3(new_n533), .A4(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(new_n540), .ZN(new_n550));
  AND3_X1   g349(.A1(new_n542), .A2(new_n550), .A3(KEYINPUT100), .ZN(new_n551));
  AOI21_X1  g350(.A(KEYINPUT100), .B1(new_n542), .B2(new_n550), .ZN(new_n552));
  OAI21_X1  g351(.A(KEYINPUT101), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n542), .A2(new_n550), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT100), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT101), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n542), .A2(new_n550), .A3(KEYINPUT100), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  NAND4_X1  g358(.A1(new_n524), .A2(new_n525), .A3(new_n553), .A4(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n514), .A2(new_n518), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(KEYINPUT88), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n562), .A2(new_n522), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n563), .A2(new_n558), .A3(new_n556), .ZN(new_n564));
  AND3_X1   g363(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n560), .A2(new_n564), .A3(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(G190gat), .B(G218gat), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  NAND4_X1  g369(.A1(new_n560), .A2(new_n564), .A3(new_n568), .A4(new_n566), .ZN(new_n571));
  XNOR2_X1  g370(.A(G134gat), .B(G162gat), .ZN(new_n572));
  AOI21_X1  g371(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n572), .B(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n570), .A2(new_n571), .A3(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT102), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n570), .A2(KEYINPUT102), .A3(new_n571), .A4(new_n575), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n570), .A2(new_n571), .ZN(new_n581));
  AOI21_X1  g380(.A(KEYINPUT103), .B1(new_n581), .B2(new_n574), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT103), .ZN(new_n583));
  AOI211_X1 g382(.A(new_n583), .B(new_n575), .C1(new_n570), .C2(new_n571), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n580), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n587), .B(KEYINPUT20), .ZN(new_n588));
  XNOR2_X1  g387(.A(G183gat), .B(G211gat), .ZN(new_n589));
  XOR2_X1   g388(.A(new_n588), .B(new_n589), .Z(new_n590));
  XNOR2_X1  g389(.A(G15gat), .B(G22gat), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT16), .ZN(new_n592));
  AOI21_X1  g391(.A(G1gat), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(G8gat), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT90), .ZN(new_n595));
  AND2_X1   g394(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n594), .B(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(G57gat), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n598), .A2(new_n332), .ZN(new_n599));
  NAND2_X1  g398(.A1(G57gat), .A2(G64gat), .ZN(new_n600));
  AND2_X1   g399(.A1(G71gat), .A2(G78gat), .ZN(new_n601));
  OAI211_X1 g400(.A(new_n599), .B(new_n600), .C1(new_n601), .C2(KEYINPUT9), .ZN(new_n602));
  OAI21_X1  g401(.A(KEYINPUT93), .B1(G71gat), .B2(G78gat), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NOR2_X1   g403(.A1(G71gat), .A2(G78gat), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n601), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  OAI211_X1 g406(.A(new_n602), .B(new_n603), .C1(new_n601), .C2(new_n605), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT96), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n607), .A2(new_n608), .A3(KEYINPUT96), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT21), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n597), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(KEYINPUT97), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n607), .A2(new_n608), .A3(new_n615), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n618), .B(KEYINPUT95), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT97), .ZN(new_n620));
  OAI211_X1 g419(.A(new_n597), .B(new_n620), .C1(new_n614), .C2(new_n615), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n617), .A2(new_n619), .A3(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n619), .B1(new_n617), .B2(new_n621), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n590), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n624), .ZN(new_n626));
  INV_X1    g425(.A(new_n590), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n626), .A2(new_n627), .A3(new_n622), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n625), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(G127gat), .B(G155gat), .ZN(new_n630));
  NAND2_X1  g429(.A1(G231gat), .A2(G233gat), .ZN(new_n631));
  XOR2_X1   g430(.A(new_n630), .B(new_n631), .Z(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n629), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n625), .A2(new_n628), .A3(new_n632), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT105), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n549), .A2(KEYINPUT104), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n609), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n639), .A2(new_n554), .ZN(new_n640));
  NAND4_X1  g439(.A1(new_n609), .A2(new_n542), .A3(new_n550), .A4(new_n638), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(G230gat), .A2(G233gat), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n637), .B1(new_n642), .B2(new_n644), .ZN(new_n645));
  AOI211_X1 g444(.A(KEYINPUT105), .B(new_n643), .C1(new_n640), .C2(new_n641), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND4_X1  g446(.A1(new_n613), .A2(new_n556), .A3(KEYINPUT10), .A4(new_n558), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT10), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n640), .A2(new_n649), .A3(new_n641), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n651), .A2(new_n643), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n647), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(G120gat), .B(G148gat), .ZN(new_n654));
  INV_X1    g453(.A(G176gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(G204gat), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n653), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n653), .A2(new_n658), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n586), .A2(new_n636), .A3(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(KEYINPUT106), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT106), .ZN(new_n666));
  NAND4_X1  g465(.A1(new_n586), .A2(new_n666), .A3(new_n636), .A4(new_n663), .ZN(new_n667));
  AND3_X1   g466(.A1(new_n494), .A2(new_n665), .A3(new_n667), .ZN(new_n668));
  XNOR2_X1  g467(.A(KEYINPUT11), .B(G169gat), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(G197gat), .ZN(new_n670));
  XOR2_X1   g469(.A(G113gat), .B(G141gat), .Z(new_n671));
  XNOR2_X1  g470(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(KEYINPUT12), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n524), .A2(new_n597), .A3(new_n525), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n594), .A2(new_n596), .ZN(new_n675));
  OR2_X1    g474(.A1(new_n594), .A2(new_n596), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n563), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(G229gat), .A2(G233gat), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n678), .B(KEYINPUT91), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n674), .A2(new_n677), .A3(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT92), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT18), .ZN(new_n683));
  AND3_X1   g482(.A1(new_n681), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n683), .B1(new_n681), .B2(new_n682), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  XOR2_X1   g485(.A(new_n679), .B(KEYINPUT13), .Z(new_n687));
  NAND3_X1  g486(.A1(new_n597), .A2(new_n562), .A3(new_n522), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n687), .B1(new_n677), .B2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n673), .B1(new_n686), .B2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n673), .ZN(new_n692));
  NOR4_X1   g491(.A1(new_n684), .A2(new_n685), .A3(new_n692), .A4(new_n689), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n668), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n398), .B(KEYINPUT107), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  XOR2_X1   g497(.A(KEYINPUT108), .B(G1gat), .Z(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(KEYINPUT109), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n698), .B(new_n700), .ZN(G1324gat));
  NOR2_X1   g500(.A1(new_n696), .A2(new_n347), .ZN(new_n702));
  INV_X1    g501(.A(G8gat), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n592), .A2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n592), .A2(new_n703), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n702), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT42), .ZN(new_n708));
  OR2_X1    g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n707), .A2(new_n708), .ZN(new_n710));
  OAI211_X1 g509(.A(new_n709), .B(new_n710), .C1(new_n703), .C2(new_n702), .ZN(G1325gat));
  INV_X1    g510(.A(G15gat), .ZN(new_n712));
  NAND4_X1  g511(.A1(new_n668), .A2(new_n712), .A3(new_n695), .A4(new_n486), .ZN(new_n713));
  INV_X1    g512(.A(new_n295), .ZN(new_n714));
  OAI21_X1  g513(.A(G15gat), .B1(new_n696), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(KEYINPUT110), .ZN(G1326gat));
  INV_X1    g516(.A(new_n431), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n696), .A2(new_n718), .ZN(new_n719));
  XOR2_X1   g518(.A(KEYINPUT43), .B(G22gat), .Z(new_n720));
  XNOR2_X1  g519(.A(new_n719), .B(new_n720), .ZN(G1327gat));
  AOI21_X1  g520(.A(new_n586), .B1(new_n485), .B2(new_n493), .ZN(new_n722));
  NOR3_X1   g521(.A1(new_n636), .A2(new_n694), .A3(new_n662), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(new_n697), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n725), .A2(new_n498), .A3(new_n726), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(KEYINPUT45), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n581), .A2(new_n574), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(new_n583), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n581), .A2(KEYINPUT103), .A3(new_n574), .ZN(new_n731));
  AOI221_X4 g530(.A(KEYINPUT112), .B1(new_n578), .B2(new_n579), .C1(new_n730), .C2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT112), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n730), .A2(new_n731), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n733), .B1(new_n734), .B2(new_n580), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n736), .A2(KEYINPUT44), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT111), .ZN(new_n738));
  AND3_X1   g537(.A1(new_n485), .A2(new_n738), .A3(new_n493), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n738), .B1(new_n485), .B2(new_n493), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n737), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n494), .A2(new_n585), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(KEYINPUT44), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(new_n723), .ZN(new_n745));
  OAI21_X1  g544(.A(G29gat), .B1(new_n745), .B2(new_n697), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n728), .A2(new_n746), .ZN(G1328gat));
  OAI21_X1  g546(.A(G36gat), .B1(new_n745), .B2(new_n347), .ZN(new_n748));
  NOR3_X1   g547(.A1(new_n724), .A2(G36gat), .A3(new_n347), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(KEYINPUT46), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n748), .A2(new_n750), .ZN(G1329gat));
  NAND3_X1  g550(.A1(new_n744), .A2(new_n295), .A3(new_n723), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(KEYINPUT113), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT113), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n744), .A2(new_n754), .A3(new_n295), .A4(new_n723), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n753), .A2(G43gat), .A3(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(new_n486), .ZN(new_n757));
  NOR3_X1   g556(.A1(new_n724), .A2(G43gat), .A3(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(new_n758), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n756), .A2(KEYINPUT47), .A3(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT47), .ZN(new_n761));
  AND2_X1   g560(.A1(new_n752), .A2(G43gat), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n761), .B1(new_n762), .B2(new_n758), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n760), .A2(new_n763), .ZN(G1330gat));
  INV_X1    g563(.A(new_n723), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n431), .A2(G50gat), .ZN(new_n766));
  AOI211_X1 g565(.A(new_n765), .B(new_n766), .C1(new_n741), .C2(new_n743), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n505), .B1(new_n724), .B2(new_n718), .ZN(new_n768));
  INV_X1    g567(.A(new_n768), .ZN(new_n769));
  OAI21_X1  g568(.A(KEYINPUT114), .B1(new_n767), .B2(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT114), .ZN(new_n771));
  OAI211_X1 g570(.A(new_n771), .B(new_n768), .C1(new_n745), .C2(new_n766), .ZN(new_n772));
  AND3_X1   g571(.A1(new_n770), .A2(new_n772), .A3(KEYINPUT48), .ZN(new_n773));
  AOI21_X1  g572(.A(KEYINPUT48), .B1(new_n770), .B2(new_n772), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n773), .A2(new_n774), .ZN(G1331gat));
  INV_X1    g574(.A(new_n636), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n776), .A2(new_n585), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n695), .A2(new_n663), .ZN(new_n778));
  OAI211_X1 g577(.A(new_n777), .B(new_n778), .C1(new_n739), .C2(new_n740), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n779), .A2(new_n697), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n780), .B(new_n598), .ZN(G1332gat));
  INV_X1    g580(.A(KEYINPUT115), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n779), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n494), .A2(KEYINPUT111), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n485), .A2(new_n493), .A3(new_n738), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND4_X1  g585(.A1(new_n786), .A2(KEYINPUT115), .A3(new_n777), .A4(new_n778), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n347), .B1(new_n783), .B2(new_n787), .ZN(new_n788));
  NOR2_X1   g587(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n789));
  AND2_X1   g588(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n788), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n791), .B1(new_n788), .B2(new_n789), .ZN(G1333gat));
  INV_X1    g591(.A(KEYINPUT50), .ZN(new_n793));
  INV_X1    g592(.A(new_n777), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n794), .B1(new_n784), .B2(new_n785), .ZN(new_n795));
  AOI21_X1  g594(.A(KEYINPUT115), .B1(new_n795), .B2(new_n778), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n779), .A2(new_n782), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n295), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(G71gat), .ZN(new_n799));
  OAI21_X1  g598(.A(KEYINPUT116), .B1(new_n779), .B2(new_n757), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT116), .ZN(new_n801));
  NAND4_X1  g600(.A1(new_n795), .A2(new_n801), .A3(new_n486), .A4(new_n778), .ZN(new_n802));
  AOI21_X1  g601(.A(G71gat), .B1(new_n800), .B2(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(new_n803), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n793), .B1(new_n799), .B2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(G71gat), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n783), .A2(new_n787), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n806), .B1(new_n807), .B2(new_n295), .ZN(new_n808));
  NOR3_X1   g607(.A1(new_n808), .A2(new_n803), .A3(KEYINPUT50), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n805), .A2(new_n809), .ZN(G1334gat));
  NAND2_X1  g609(.A1(new_n807), .A2(new_n431), .ZN(new_n811));
  XNOR2_X1  g610(.A(new_n811), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g611(.A1(new_n695), .A2(new_n636), .A3(new_n663), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n744), .A2(new_n813), .ZN(new_n814));
  OR3_X1    g613(.A1(new_n814), .A2(KEYINPUT117), .A3(new_n697), .ZN(new_n815));
  OAI21_X1  g614(.A(KEYINPUT117), .B1(new_n814), .B2(new_n697), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n815), .A2(G85gat), .A3(new_n816), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n695), .A2(new_n636), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n494), .A2(new_n585), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(KEYINPUT51), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT51), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n722), .A2(new_n821), .A3(new_n818), .ZN(new_n822));
  AND2_X1   g621(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n823), .A2(new_n528), .A3(new_n726), .A4(new_n662), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n817), .A2(new_n824), .ZN(G1336gat));
  NAND4_X1  g624(.A1(new_n823), .A2(new_n334), .A3(new_n662), .A4(new_n456), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n814), .A2(new_n347), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n826), .B1(new_n827), .B2(new_n334), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(KEYINPUT52), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT52), .ZN(new_n830));
  OAI211_X1 g629(.A(new_n830), .B(new_n826), .C1(new_n827), .C2(new_n334), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n829), .A2(new_n831), .ZN(G1337gat));
  OAI21_X1  g631(.A(G99gat), .B1(new_n814), .B2(new_n714), .ZN(new_n833));
  INV_X1    g632(.A(G99gat), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n823), .A2(new_n834), .A3(new_n662), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n833), .B1(new_n757), .B2(new_n835), .ZN(G1338gat));
  NAND4_X1  g635(.A1(new_n744), .A2(G106gat), .A3(new_n431), .A4(new_n813), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n820), .A2(new_n662), .A3(new_n431), .A4(new_n822), .ZN(new_n838));
  INV_X1    g637(.A(G106gat), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n837), .A2(new_n840), .ZN(new_n841));
  XNOR2_X1  g640(.A(KEYINPUT118), .B(KEYINPUT53), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(KEYINPUT119), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n837), .A2(new_n840), .A3(KEYINPUT53), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT119), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n841), .A2(new_n846), .A3(new_n842), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n844), .A2(new_n845), .A3(new_n847), .ZN(G1339gat));
  NAND3_X1  g647(.A1(new_n648), .A2(new_n644), .A3(new_n650), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n652), .A2(KEYINPUT54), .A3(new_n849), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n644), .B1(new_n648), .B2(new_n650), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT54), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n657), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  AND3_X1   g652(.A1(new_n850), .A2(KEYINPUT55), .A3(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(KEYINPUT55), .B1(new_n850), .B2(new_n853), .ZN(new_n855));
  NOR3_X1   g654(.A1(new_n854), .A2(new_n855), .A3(new_n659), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n686), .A2(new_n673), .A3(new_n690), .ZN(new_n857));
  AND3_X1   g656(.A1(new_n677), .A2(new_n688), .A3(new_n687), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n680), .B1(new_n674), .B2(new_n677), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n672), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n856), .A2(new_n857), .A3(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(new_n861), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n862), .B1(new_n732), .B2(new_n735), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n856), .B1(new_n691), .B2(new_n693), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n857), .A2(new_n662), .A3(new_n860), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n585), .A2(KEYINPUT112), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n734), .A2(new_n733), .A3(new_n580), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n866), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n863), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(new_n776), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n777), .A2(new_n694), .A3(new_n663), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n697), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(new_n490), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  OR3_X1    g674(.A1(new_n875), .A2(G113gat), .A3(new_n694), .ZN(new_n876));
  OAI21_X1  g675(.A(G113gat), .B1(new_n875), .B2(new_n694), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  XOR2_X1   g677(.A(new_n878), .B(KEYINPUT120), .Z(G1340gat));
  NOR2_X1   g678(.A1(new_n875), .A2(new_n663), .ZN(new_n880));
  XOR2_X1   g679(.A(new_n880), .B(G120gat), .Z(G1341gat));
  NOR2_X1   g680(.A1(new_n875), .A2(new_n776), .ZN(new_n882));
  NOR2_X1   g681(.A1(KEYINPUT121), .A2(G127gat), .ZN(new_n883));
  XNOR2_X1  g682(.A(new_n882), .B(new_n883), .ZN(G1342gat));
  NAND2_X1  g683(.A1(new_n585), .A2(new_n347), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n873), .A2(new_n487), .ZN(new_n886));
  AOI211_X1 g685(.A(new_n885), .B(new_n886), .C1(KEYINPUT56), .C2(G134gat), .ZN(new_n887));
  NOR2_X1   g686(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n888));
  XNOR2_X1  g687(.A(new_n887), .B(new_n888), .ZN(G1343gat));
  XNOR2_X1  g688(.A(KEYINPUT123), .B(KEYINPUT58), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT122), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n295), .B1(new_n873), .B2(new_n891), .ZN(new_n892));
  INV_X1    g691(.A(G141gat), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n636), .B1(new_n863), .B2(new_n869), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n664), .A2(new_n695), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n726), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n718), .B1(new_n896), .B2(KEYINPUT122), .ZN(new_n897));
  NAND4_X1  g696(.A1(new_n892), .A2(new_n893), .A3(new_n347), .A4(new_n897), .ZN(new_n898));
  OR2_X1    g697(.A1(new_n898), .A2(new_n694), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT57), .ZN(new_n900));
  OAI211_X1 g699(.A(new_n900), .B(new_n431), .C1(new_n894), .C2(new_n895), .ZN(new_n901));
  NOR3_X1   g700(.A1(new_n697), .A2(new_n456), .A3(new_n295), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n861), .B1(new_n867), .B2(new_n868), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n585), .B1(new_n864), .B2(new_n865), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n776), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n718), .B1(new_n905), .B2(new_n872), .ZN(new_n906));
  OAI211_X1 g705(.A(new_n901), .B(new_n902), .C1(new_n900), .C2(new_n906), .ZN(new_n907));
  OAI21_X1  g706(.A(G141gat), .B1(new_n907), .B2(new_n694), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n890), .B1(new_n899), .B2(new_n908), .ZN(new_n909));
  OAI211_X1 g708(.A(new_n908), .B(new_n890), .C1(new_n898), .C2(new_n694), .ZN(new_n910));
  INV_X1    g709(.A(new_n910), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n909), .A2(new_n911), .ZN(G1344gat));
  INV_X1    g711(.A(KEYINPUT125), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT59), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n431), .B1(new_n894), .B2(new_n895), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(KEYINPUT57), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n665), .A2(new_n667), .A3(new_n694), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n586), .A2(new_n861), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n776), .B1(new_n918), .B2(new_n904), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n718), .A2(KEYINPUT57), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND4_X1  g721(.A1(new_n916), .A2(new_n662), .A3(new_n922), .A4(new_n902), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n914), .B1(new_n923), .B2(G148gat), .ZN(new_n924));
  INV_X1    g723(.A(G148gat), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n925), .A2(KEYINPUT59), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n926), .B1(new_n907), .B2(new_n663), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT124), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n866), .A2(new_n586), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n636), .B1(new_n863), .B2(new_n930), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n431), .B1(new_n931), .B2(new_n895), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(KEYINPUT57), .ZN(new_n933));
  NAND4_X1  g732(.A1(new_n933), .A2(new_n662), .A3(new_n902), .A4(new_n901), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n934), .A2(KEYINPUT124), .A3(new_n926), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n924), .B1(new_n929), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n892), .A2(new_n897), .ZN(new_n937));
  NOR4_X1   g736(.A1(new_n937), .A2(G148gat), .A3(new_n663), .A4(new_n456), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n913), .B1(new_n936), .B2(new_n938), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n937), .A2(new_n456), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n940), .A2(new_n925), .A3(new_n662), .ZN(new_n941));
  AND3_X1   g740(.A1(new_n934), .A2(KEYINPUT124), .A3(new_n926), .ZN(new_n942));
  AOI21_X1  g741(.A(KEYINPUT124), .B1(new_n934), .B2(new_n926), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  OAI211_X1 g743(.A(KEYINPUT125), .B(new_n941), .C1(new_n944), .C2(new_n924), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n939), .A2(new_n945), .ZN(G1345gat));
  NOR3_X1   g745(.A1(new_n907), .A2(new_n353), .A3(new_n776), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n940), .A2(new_n636), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n947), .B1(new_n948), .B2(new_n353), .ZN(G1346gat));
  OAI21_X1  g748(.A(G162gat), .B1(new_n907), .B2(new_n736), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n585), .A2(new_n354), .A3(new_n347), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n950), .B1(new_n937), .B2(new_n951), .ZN(G1347gat));
  NOR2_X1   g751(.A1(new_n726), .A2(new_n347), .ZN(new_n953));
  OAI211_X1 g752(.A(new_n487), .B(new_n953), .C1(new_n894), .C2(new_n895), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n954), .A2(new_n694), .ZN(new_n955));
  XOR2_X1   g754(.A(new_n955), .B(G169gat), .Z(G1348gat));
  NOR2_X1   g755(.A1(new_n954), .A2(new_n663), .ZN(new_n957));
  XNOR2_X1  g756(.A(new_n957), .B(new_n655), .ZN(G1349gat));
  NOR2_X1   g757(.A1(new_n954), .A2(new_n776), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n959), .B1(new_n220), .B2(new_n219), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n960), .B1(new_n233), .B2(new_n959), .ZN(new_n961));
  XNOR2_X1  g760(.A(new_n961), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g761(.A(G190gat), .B1(new_n954), .B2(new_n586), .ZN(new_n963));
  XNOR2_X1  g762(.A(new_n963), .B(KEYINPUT61), .ZN(new_n964));
  INV_X1    g763(.A(new_n736), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n965), .A2(new_n217), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n964), .B1(new_n954), .B2(new_n966), .ZN(G1351gat));
  INV_X1    g766(.A(KEYINPUT126), .ZN(new_n968));
  AOI22_X1  g767(.A1(new_n915), .A2(KEYINPUT57), .B1(new_n920), .B2(new_n921), .ZN(new_n969));
  NOR3_X1   g768(.A1(new_n726), .A2(new_n347), .A3(new_n295), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n968), .B1(new_n971), .B2(new_n694), .ZN(new_n972));
  NAND4_X1  g771(.A1(new_n969), .A2(KEYINPUT126), .A3(new_n695), .A4(new_n970), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n972), .A2(G197gat), .A3(new_n973), .ZN(new_n974));
  INV_X1    g773(.A(new_n915), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n975), .A2(new_n970), .ZN(new_n976));
  OR2_X1    g775(.A1(new_n694), .A2(G197gat), .ZN(new_n977));
  OAI21_X1  g776(.A(new_n974), .B1(new_n976), .B2(new_n977), .ZN(G1352gat));
  NOR3_X1   g777(.A1(new_n976), .A2(G204gat), .A3(new_n663), .ZN(new_n979));
  INV_X1    g778(.A(KEYINPUT62), .ZN(new_n980));
  OR2_X1    g779(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n969), .A2(new_n662), .A3(new_n970), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n982), .A2(G204gat), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n979), .A2(new_n980), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n981), .A2(new_n983), .A3(new_n984), .ZN(G1353gat));
  NAND4_X1  g784(.A1(new_n916), .A2(new_n636), .A3(new_n922), .A4(new_n970), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n986), .A2(KEYINPUT127), .ZN(new_n987));
  INV_X1    g786(.A(KEYINPUT127), .ZN(new_n988));
  NAND4_X1  g787(.A1(new_n969), .A2(new_n988), .A3(new_n636), .A4(new_n970), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n987), .A2(new_n989), .A3(G211gat), .ZN(new_n990));
  INV_X1    g789(.A(KEYINPUT63), .ZN(new_n991));
  XNOR2_X1  g790(.A(new_n990), .B(new_n991), .ZN(new_n992));
  OR3_X1    g791(.A1(new_n976), .A2(new_n776), .A3(new_n298), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n992), .A2(new_n993), .ZN(G1354gat));
  OAI21_X1  g793(.A(G218gat), .B1(new_n971), .B2(new_n586), .ZN(new_n995));
  NAND3_X1  g794(.A1(new_n975), .A2(new_n296), .A3(new_n970), .ZN(new_n996));
  OAI21_X1  g795(.A(new_n995), .B1(new_n736), .B2(new_n996), .ZN(G1355gat));
endmodule


