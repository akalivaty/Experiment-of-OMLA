//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 1 1 1 0 0 0 1 0 1 0 0 0 0 1 0 0 0 0 0 0 0 0 1 1 1 0 1 0 1 1 0 1 1 1 0 1 1 0 0 0 1 1 0 0 0 0 1 1 0 1 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:16 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n759, new_n760, new_n761, new_n762, new_n763, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n786, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016;
  INV_X1    g000(.A(KEYINPUT23), .ZN(new_n187));
  INV_X1    g001(.A(G119), .ZN(new_n188));
  OAI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G128), .ZN(new_n189));
  INV_X1    g003(.A(G128), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n190), .A2(KEYINPUT23), .A3(G119), .ZN(new_n191));
  OAI211_X1 g005(.A(new_n189), .B(new_n191), .C1(G119), .C2(new_n190), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G110), .ZN(new_n193));
  XOR2_X1   g007(.A(KEYINPUT24), .B(G110), .Z(new_n194));
  XNOR2_X1  g008(.A(G119), .B(G128), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n193), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G125), .ZN(new_n198));
  OR3_X1    g012(.A1(new_n198), .A2(KEYINPUT16), .A3(G140), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT72), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  XNOR2_X1  g015(.A(G125), .B(G140), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(KEYINPUT16), .ZN(new_n203));
  AND2_X1   g017(.A1(new_n203), .A2(new_n199), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n201), .B1(new_n204), .B2(new_n200), .ZN(new_n205));
  INV_X1    g019(.A(G146), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  OAI211_X1 g021(.A(G146), .B(new_n201), .C1(new_n204), .C2(new_n200), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n197), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(new_n209), .ZN(new_n210));
  OAI22_X1  g024(.A1(new_n192), .A2(G110), .B1(new_n195), .B2(new_n194), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n202), .A2(new_n206), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n208), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  XNOR2_X1  g027(.A(KEYINPUT22), .B(G137), .ZN(new_n214));
  INV_X1    g028(.A(G953), .ZN(new_n215));
  AND3_X1   g029(.A1(new_n215), .A2(G221), .A3(G234), .ZN(new_n216));
  XOR2_X1   g030(.A(new_n214), .B(new_n216), .Z(new_n217));
  NAND3_X1  g031(.A1(new_n210), .A2(new_n213), .A3(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(G902), .ZN(new_n219));
  INV_X1    g033(.A(new_n217), .ZN(new_n220));
  INV_X1    g034(.A(new_n213), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n220), .B1(new_n209), .B2(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n218), .A2(new_n219), .A3(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(KEYINPUT25), .ZN(new_n224));
  NAND2_X1  g038(.A1(G217), .A2(G902), .ZN(new_n225));
  INV_X1    g039(.A(G217), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n225), .B1(new_n226), .B2(G234), .ZN(new_n227));
  XNOR2_X1  g041(.A(new_n227), .B(KEYINPUT71), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT25), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n218), .A2(new_n222), .A3(new_n229), .A4(new_n219), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n224), .A2(new_n228), .A3(new_n230), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n228), .A2(G902), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n218), .A2(new_n222), .A3(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(G134), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G137), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n235), .A2(G137), .ZN(new_n238));
  OAI21_X1  g052(.A(G131), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT11), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n240), .B1(new_n235), .B2(G137), .ZN(new_n241));
  INV_X1    g055(.A(G137), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n242), .A2(KEYINPUT11), .A3(G134), .ZN(new_n243));
  INV_X1    g057(.A(G131), .ZN(new_n244));
  NAND4_X1  g058(.A1(new_n241), .A2(new_n243), .A3(new_n244), .A4(new_n236), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n239), .A2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT1), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(KEYINPUT64), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT64), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(KEYINPUT1), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n248), .A2(new_n250), .A3(G128), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n206), .A2(G143), .ZN(new_n252));
  INV_X1    g066(.A(G143), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G146), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  OAI21_X1  g069(.A(KEYINPUT65), .B1(new_n251), .B2(new_n255), .ZN(new_n256));
  XNOR2_X1  g070(.A(G143), .B(G146), .ZN(new_n257));
  XNOR2_X1  g071(.A(KEYINPUT64), .B(KEYINPUT1), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT65), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n257), .A2(new_n258), .A3(new_n259), .A4(G128), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n256), .A2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(new_n252), .ZN(new_n262));
  OAI21_X1  g076(.A(G128), .B1(new_n258), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(new_n255), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n246), .B1(new_n261), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(KEYINPUT0), .A2(G128), .ZN(new_n266));
  OR2_X1    g080(.A1(KEYINPUT0), .A2(G128), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n255), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n257), .A2(KEYINPUT0), .A3(G128), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n241), .A2(new_n236), .A3(new_n243), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(G131), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n270), .B1(new_n245), .B2(new_n272), .ZN(new_n273));
  OAI21_X1  g087(.A(KEYINPUT30), .B1(new_n265), .B2(new_n273), .ZN(new_n274));
  AND2_X1   g088(.A1(new_n268), .A2(new_n269), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n272), .A2(new_n245), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT30), .ZN(new_n278));
  AOI22_X1  g092(.A1(new_n256), .A2(new_n260), .B1(new_n263), .B2(new_n255), .ZN(new_n279));
  OAI211_X1 g093(.A(new_n277), .B(new_n278), .C1(new_n279), .C2(new_n246), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n274), .A2(new_n280), .ZN(new_n281));
  XOR2_X1   g095(.A(KEYINPUT2), .B(G113), .Z(new_n282));
  XNOR2_X1  g096(.A(G116), .B(G119), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n282), .B1(KEYINPUT66), .B2(new_n283), .ZN(new_n284));
  XNOR2_X1  g098(.A(KEYINPUT2), .B(G113), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT66), .ZN(new_n286));
  INV_X1    g100(.A(G116), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n287), .A2(G119), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n188), .A2(G116), .ZN(new_n289));
  OAI211_X1 g103(.A(new_n285), .B(new_n286), .C1(new_n288), .C2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n284), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n281), .A2(new_n291), .ZN(new_n292));
  AND2_X1   g106(.A1(new_n284), .A2(new_n290), .ZN(new_n293));
  AND2_X1   g107(.A1(new_n272), .A2(new_n245), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n293), .B1(new_n294), .B2(new_n270), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT67), .ZN(new_n296));
  NOR3_X1   g110(.A1(new_n295), .A2(new_n265), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n261), .A2(new_n264), .ZN(new_n298));
  INV_X1    g112(.A(new_n246), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n291), .B1(new_n276), .B2(new_n275), .ZN(new_n301));
  AOI21_X1  g115(.A(KEYINPUT67), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n297), .A2(new_n302), .ZN(new_n303));
  XOR2_X1   g117(.A(KEYINPUT68), .B(KEYINPUT27), .Z(new_n304));
  INV_X1    g118(.A(G237), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n305), .A2(new_n215), .A3(G210), .ZN(new_n306));
  XNOR2_X1  g120(.A(new_n304), .B(new_n306), .ZN(new_n307));
  XNOR2_X1  g121(.A(KEYINPUT26), .B(G101), .ZN(new_n308));
  XNOR2_X1  g122(.A(new_n307), .B(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n292), .A2(new_n303), .A3(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT31), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n293), .B1(new_n274), .B2(new_n280), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n296), .B1(new_n295), .B2(new_n265), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n300), .A2(KEYINPUT67), .A3(new_n301), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n314), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n318), .A2(KEYINPUT31), .A3(new_n310), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n313), .A2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT69), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n295), .A2(new_n265), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n322), .A2(KEYINPUT28), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n291), .B1(new_n265), .B2(new_n273), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n315), .A2(new_n316), .A3(new_n324), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n323), .B1(new_n325), .B2(KEYINPUT28), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n321), .B1(new_n326), .B2(new_n310), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n325), .A2(KEYINPUT28), .ZN(new_n328));
  INV_X1    g142(.A(new_n323), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n330), .A2(KEYINPUT69), .A3(new_n309), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n320), .A2(new_n327), .A3(new_n331), .ZN(new_n332));
  NOR2_X1   g146(.A1(G472), .A2(G902), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT32), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  AND3_X1   g150(.A1(new_n332), .A2(KEYINPUT70), .A3(new_n336), .ZN(new_n337));
  AOI21_X1  g151(.A(KEYINPUT70), .B1(new_n332), .B2(new_n336), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(G472), .ZN(new_n340));
  AND2_X1   g154(.A1(new_n326), .A2(new_n310), .ZN(new_n341));
  AOI21_X1  g155(.A(G902), .B1(new_n341), .B2(KEYINPUT29), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n326), .A2(new_n310), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT29), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n309), .B1(new_n314), .B2(new_n317), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n343), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n340), .B1(new_n342), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n332), .A2(new_n333), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n347), .B1(new_n335), .B2(new_n348), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n234), .B1(new_n339), .B2(new_n349), .ZN(new_n350));
  AND2_X1   g164(.A1(new_n215), .A2(G952), .ZN(new_n351));
  NAND2_X1  g165(.A1(G234), .A2(G237), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  XNOR2_X1  g167(.A(KEYINPUT21), .B(G898), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n352), .A2(G902), .A3(G953), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n353), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  XNOR2_X1  g171(.A(G128), .B(G143), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(KEYINPUT13), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n253), .A2(G128), .ZN(new_n360));
  OAI211_X1 g174(.A(new_n359), .B(G134), .C1(KEYINPUT13), .C2(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n358), .A2(KEYINPUT96), .A3(new_n235), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT96), .ZN(new_n363));
  INV_X1    g177(.A(new_n358), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n363), .B1(new_n364), .B2(G134), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n361), .A2(new_n362), .A3(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT95), .ZN(new_n367));
  AND2_X1   g181(.A1(KEYINPUT91), .A2(G122), .ZN(new_n368));
  NOR2_X1   g182(.A1(KEYINPUT91), .A2(G122), .ZN(new_n369));
  OAI21_X1  g183(.A(G116), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(KEYINPUT92), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT92), .ZN(new_n372));
  OAI211_X1 g186(.A(new_n372), .B(G116), .C1(new_n368), .C2(new_n369), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(G122), .ZN(new_n375));
  OAI21_X1  g189(.A(KEYINPUT93), .B1(new_n375), .B2(G116), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT93), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n377), .A2(new_n287), .A3(G122), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  AND3_X1   g193(.A1(new_n374), .A2(KEYINPUT94), .A3(new_n379), .ZN(new_n380));
  AOI21_X1  g194(.A(KEYINPUT94), .B1(new_n374), .B2(new_n379), .ZN(new_n381));
  INV_X1    g195(.A(G107), .ZN(new_n382));
  NOR3_X1   g196(.A1(new_n380), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  XNOR2_X1  g197(.A(KEYINPUT91), .B(G122), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n372), .B1(new_n384), .B2(G116), .ZN(new_n385));
  INV_X1    g199(.A(new_n373), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n379), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT94), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n374), .A2(KEYINPUT94), .A3(new_n379), .ZN(new_n390));
  AOI21_X1  g204(.A(G107), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n367), .B1(new_n383), .B2(new_n391), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n382), .B1(new_n380), .B2(new_n381), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n389), .A2(G107), .A3(new_n390), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n393), .A2(KEYINPUT95), .A3(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n366), .B1(new_n392), .B2(new_n395), .ZN(new_n396));
  XNOR2_X1  g210(.A(new_n358), .B(new_n235), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n393), .A2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT14), .ZN(new_n399));
  XNOR2_X1  g213(.A(new_n379), .B(new_n399), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n382), .B1(new_n400), .B2(new_n374), .ZN(new_n401));
  OR2_X1    g215(.A1(new_n401), .A2(KEYINPUT97), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(KEYINPUT97), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n398), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  XNOR2_X1  g218(.A(KEYINPUT9), .B(G234), .ZN(new_n405));
  NOR3_X1   g219(.A1(new_n405), .A2(new_n226), .A3(G953), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  NOR3_X1   g221(.A1(new_n396), .A2(new_n404), .A3(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n366), .ZN(new_n409));
  AND3_X1   g223(.A1(new_n393), .A2(KEYINPUT95), .A3(new_n394), .ZN(new_n410));
  AOI21_X1  g224(.A(KEYINPUT95), .B1(new_n393), .B2(new_n394), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n409), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n402), .A2(new_n403), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n413), .A2(new_n393), .A3(new_n397), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n406), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n219), .B1(new_n408), .B2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(G478), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n417), .A2(KEYINPUT15), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n407), .B1(new_n396), .B2(new_n404), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n412), .A2(new_n414), .A3(new_n406), .ZN(new_n421));
  AOI21_X1  g235(.A(G902), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n418), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  OR2_X1    g238(.A1(new_n253), .A2(KEYINPUT86), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n305), .A2(new_n215), .A3(G214), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  XNOR2_X1  g241(.A(KEYINPUT86), .B(G143), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n427), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  OR2_X1    g243(.A1(new_n429), .A2(G131), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT17), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n429), .A2(G131), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n430), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n429), .A2(KEYINPUT17), .A3(G131), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n207), .A2(new_n433), .A3(new_n208), .A4(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n429), .A2(KEYINPUT18), .A3(G131), .ZN(new_n436));
  NAND2_X1  g250(.A1(KEYINPUT18), .A2(G131), .ZN(new_n437));
  OAI211_X1 g251(.A(new_n427), .B(new_n437), .C1(new_n426), .C2(new_n428), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n202), .B(new_n206), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n436), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT87), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND4_X1  g256(.A1(new_n436), .A2(KEYINPUT87), .A3(new_n438), .A4(new_n439), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  XNOR2_X1  g258(.A(G113), .B(G122), .ZN(new_n445));
  XNOR2_X1  g259(.A(KEYINPUT89), .B(G104), .ZN(new_n446));
  XNOR2_X1  g260(.A(new_n445), .B(new_n446), .ZN(new_n447));
  AND3_X1   g261(.A1(new_n435), .A2(new_n444), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n430), .A2(new_n432), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT88), .ZN(new_n450));
  OR2_X1    g264(.A1(new_n450), .A2(KEYINPUT19), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(KEYINPUT19), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n202), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n453), .B1(new_n202), .B2(new_n452), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(new_n206), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n449), .A2(new_n208), .A3(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n447), .B1(new_n444), .B2(new_n456), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n448), .A2(new_n457), .ZN(new_n458));
  NOR2_X1   g272(.A1(G475), .A2(G902), .ZN(new_n459));
  XNOR2_X1  g273(.A(new_n459), .B(KEYINPUT90), .ZN(new_n460));
  OAI21_X1  g274(.A(KEYINPUT20), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT20), .ZN(new_n462));
  INV_X1    g276(.A(new_n460), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n462), .B(new_n463), .C1(new_n448), .C2(new_n457), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n447), .B1(new_n435), .B2(new_n444), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n219), .B1(new_n448), .B2(new_n465), .ZN(new_n466));
  AOI22_X1  g280(.A1(new_n461), .A2(new_n464), .B1(G475), .B2(new_n466), .ZN(new_n467));
  AND4_X1   g281(.A1(new_n357), .A2(new_n419), .A3(new_n424), .A4(new_n467), .ZN(new_n468));
  OAI21_X1  g282(.A(G214), .B1(G237), .B2(G902), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(G104), .ZN(new_n471));
  OAI21_X1  g285(.A(KEYINPUT3), .B1(new_n471), .B2(G107), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT3), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n473), .A2(new_n382), .A3(G104), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n471), .A2(G107), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n472), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(KEYINPUT73), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT73), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n472), .A2(new_n474), .A3(new_n478), .A4(new_n475), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n477), .A2(G101), .A3(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(G101), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n472), .A2(new_n474), .A3(new_n481), .A4(new_n475), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n480), .A2(KEYINPUT4), .A3(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT82), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT4), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n477), .A2(new_n485), .A3(G101), .A4(new_n479), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n483), .A2(new_n484), .A3(new_n291), .A4(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n291), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n482), .A2(KEYINPUT4), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n481), .B1(new_n476), .B2(KEYINPUT73), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n489), .B1(new_n490), .B2(new_n479), .ZN(new_n491));
  OAI21_X1  g305(.A(KEYINPUT82), .B1(new_n488), .B2(new_n491), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n471), .A2(G107), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n382), .A2(G104), .ZN(new_n494));
  OAI21_X1  g308(.A(G101), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n482), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(KEYINPUT75), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT75), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n482), .A2(new_n495), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n283), .A2(KEYINPUT5), .ZN(new_n501));
  INV_X1    g315(.A(G113), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT5), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n502), .B1(new_n288), .B2(new_n503), .ZN(new_n504));
  AOI22_X1  g318(.A1(new_n501), .A2(new_n504), .B1(new_n282), .B2(new_n283), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n500), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n487), .A2(new_n492), .A3(new_n506), .ZN(new_n507));
  XNOR2_X1  g321(.A(G110), .B(G122), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n487), .A2(new_n492), .A3(new_n508), .A4(new_n506), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n510), .A2(KEYINPUT6), .A3(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT6), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n507), .A2(new_n513), .A3(new_n509), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n198), .B1(new_n268), .B2(new_n269), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n515), .B1(new_n279), .B2(new_n198), .ZN(new_n516));
  INV_X1    g330(.A(G224), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n517), .A2(G953), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n516), .B(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n512), .A2(new_n514), .A3(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n261), .A2(new_n198), .A3(new_n264), .ZN(new_n522));
  INV_X1    g336(.A(new_n515), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT84), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n524), .A2(new_n525), .A3(KEYINPUT7), .A4(new_n519), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n519), .A2(KEYINPUT7), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n518), .A2(new_n525), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n527), .B1(new_n516), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n526), .A2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n496), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(KEYINPUT83), .ZN(new_n532));
  OR2_X1    g346(.A1(new_n532), .A2(new_n505), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n505), .ZN(new_n534));
  XNOR2_X1  g348(.A(new_n508), .B(KEYINPUT8), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n530), .A2(new_n511), .A3(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT85), .ZN(new_n538));
  AND3_X1   g352(.A1(new_n537), .A2(new_n538), .A3(new_n219), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n538), .B1(new_n537), .B2(new_n219), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n521), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  OAI21_X1  g355(.A(G210), .B1(G237), .B2(G902), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n542), .B(new_n521), .C1(new_n539), .C2(new_n540), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n470), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  AND2_X1   g360(.A1(new_n468), .A2(new_n546), .ZN(new_n547));
  XNOR2_X1  g361(.A(KEYINPUT79), .B(G469), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n483), .A2(new_n275), .A3(new_n486), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT10), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n550), .B1(new_n261), .B2(new_n264), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(new_n500), .ZN(new_n552));
  XNOR2_X1  g366(.A(KEYINPUT74), .B(KEYINPUT10), .ZN(new_n553));
  OAI22_X1  g367(.A1(new_n257), .A2(G128), .B1(new_n247), .B2(new_n254), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n554), .B1(new_n256), .B2(new_n260), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n553), .B1(new_n555), .B2(new_n496), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n549), .A2(new_n552), .A3(new_n294), .A4(new_n556), .ZN(new_n557));
  XNOR2_X1  g371(.A(G110), .B(G140), .ZN(new_n558));
  INV_X1    g372(.A(G227), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n559), .A2(G953), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n558), .B(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n557), .A2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT12), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n564), .A2(KEYINPUT76), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n565), .A2(KEYINPUT12), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  AND2_X1   g381(.A1(new_n276), .A2(KEYINPUT76), .ZN(new_n568));
  AND3_X1   g382(.A1(new_n261), .A2(new_n264), .A3(new_n496), .ZN(new_n569));
  INV_X1    g383(.A(new_n554), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n496), .B1(new_n261), .B2(new_n570), .ZN(new_n571));
  OAI211_X1 g385(.A(new_n567), .B(new_n568), .C1(new_n569), .C2(new_n571), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n568), .B1(new_n569), .B2(new_n571), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(new_n566), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n563), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n549), .A2(new_n552), .A3(new_n556), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(new_n276), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n562), .B1(new_n577), .B2(new_n557), .ZN(new_n578));
  OAI211_X1 g392(.A(new_n219), .B(new_n548), .C1(new_n575), .C2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT80), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n261), .A2(new_n570), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(new_n531), .ZN(new_n583));
  AOI22_X1  g397(.A1(new_n583), .A2(new_n553), .B1(new_n551), .B2(new_n500), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n294), .B1(new_n584), .B2(new_n549), .ZN(new_n585));
  INV_X1    g399(.A(new_n557), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n561), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n574), .A2(new_n572), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n588), .A2(new_n562), .A3(new_n557), .ZN(new_n589));
  AOI21_X1  g403(.A(G902), .B1(new_n587), .B2(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n590), .A2(KEYINPUT80), .A3(new_n548), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n581), .A2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(new_n572), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n261), .A2(new_n264), .A3(new_n496), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n594), .B1(new_n496), .B2(new_n555), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n567), .B1(new_n595), .B2(new_n568), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n557), .B1(new_n593), .B2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT77), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  OAI211_X1 g413(.A(KEYINPUT77), .B(new_n557), .C1(new_n593), .C2(new_n596), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n562), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n563), .A2(new_n585), .ZN(new_n602));
  OAI21_X1  g416(.A(KEYINPUT78), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n600), .ZN(new_n604));
  AOI21_X1  g418(.A(KEYINPUT77), .B1(new_n588), .B2(new_n557), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n561), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT78), .ZN(new_n607));
  INV_X1    g421(.A(new_n602), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  AOI21_X1  g423(.A(G902), .B1(new_n603), .B2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(G469), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n592), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT81), .ZN(new_n613));
  INV_X1    g427(.A(G221), .ZN(new_n614));
  INV_X1    g428(.A(new_n405), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n614), .B1(new_n615), .B2(new_n219), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  AND3_X1   g431(.A1(new_n612), .A2(new_n613), .A3(new_n617), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n613), .B1(new_n612), .B2(new_n617), .ZN(new_n619));
  OAI211_X1 g433(.A(new_n350), .B(new_n547), .C1(new_n618), .C2(new_n619), .ZN(new_n620));
  XNOR2_X1  g434(.A(KEYINPUT98), .B(G101), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n620), .B(new_n621), .ZN(G3));
  NAND2_X1  g436(.A1(new_n612), .A2(new_n617), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(KEYINPUT81), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n612), .A2(new_n613), .A3(new_n617), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n310), .B1(new_n328), .B2(new_n329), .ZN(new_n627));
  AOI22_X1  g441(.A1(new_n313), .A2(new_n319), .B1(new_n627), .B2(KEYINPUT69), .ZN(new_n628));
  AOI21_X1  g442(.A(G902), .B1(new_n628), .B2(new_n327), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n348), .B1(new_n629), .B2(new_n340), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n630), .A2(new_n234), .ZN(new_n631));
  AND2_X1   g445(.A1(new_n626), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n544), .A2(new_n545), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n633), .A2(new_n469), .A3(new_n357), .ZN(new_n634));
  OAI21_X1  g448(.A(KEYINPUT33), .B1(new_n406), .B2(KEYINPUT99), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n420), .A2(new_n421), .A3(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n636), .B1(new_n420), .B2(new_n421), .ZN(new_n639));
  OAI21_X1  g453(.A(G478), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n467), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n417), .A2(new_n219), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n642), .B1(new_n422), .B2(new_n417), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n640), .A2(new_n641), .A3(new_n643), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n634), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n632), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(G104), .ZN(new_n647));
  XNOR2_X1  g461(.A(KEYINPUT100), .B(KEYINPUT34), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G6));
  NAND2_X1  g463(.A1(new_n419), .A2(new_n424), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(new_n467), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n634), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n632), .A2(new_n652), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT35), .B(G107), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G9));
  NOR2_X1   g469(.A1(new_n220), .A2(KEYINPUT36), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n210), .A2(new_n213), .A3(new_n656), .ZN(new_n657));
  OAI22_X1  g471(.A1(new_n209), .A2(new_n221), .B1(KEYINPUT36), .B2(new_n220), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n657), .A2(new_n232), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n231), .A2(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n630), .A2(new_n661), .ZN(new_n662));
  OAI211_X1 g476(.A(new_n547), .B(new_n662), .C1(new_n618), .C2(new_n619), .ZN(new_n663));
  XOR2_X1   g477(.A(KEYINPUT37), .B(G110), .Z(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(KEYINPUT101), .B(KEYINPUT102), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(G12));
  NAND2_X1  g481(.A1(new_n348), .A2(new_n335), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n332), .A2(new_n336), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT70), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(new_n346), .ZN(new_n672));
  OAI21_X1  g486(.A(new_n219), .B1(new_n343), .B2(new_n344), .ZN(new_n673));
  OAI21_X1  g487(.A(G472), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n332), .A2(KEYINPUT70), .A3(new_n336), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n668), .A2(new_n671), .A3(new_n674), .A4(new_n675), .ZN(new_n676));
  OR2_X1    g490(.A1(new_n356), .A2(G900), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(new_n353), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n651), .A2(new_n679), .ZN(new_n680));
  AND4_X1   g494(.A1(new_n676), .A2(new_n680), .A3(new_n546), .A4(new_n660), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n626), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G128), .ZN(G30));
  INV_X1    g497(.A(KEYINPUT106), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n678), .B(KEYINPUT39), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n685), .B1(new_n618), .B2(new_n619), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT40), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  AOI21_X1  g502(.A(KEYINPUT40), .B1(new_n626), .B2(new_n685), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n684), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n467), .A2(new_n470), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n650), .A2(new_n691), .A3(new_n661), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(KEYINPUT104), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n633), .B(KEYINPUT38), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n318), .A2(new_n309), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n219), .B1(new_n325), .B2(new_n310), .ZN(new_n696));
  OAI21_X1  g510(.A(G472), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(KEYINPUT103), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n339), .A2(new_n668), .A3(new_n698), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n693), .A2(new_n694), .A3(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT105), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n700), .B(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n686), .A2(new_n687), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n626), .A2(KEYINPUT40), .A3(new_n685), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n703), .A2(new_n704), .A3(KEYINPUT106), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n690), .A2(new_n702), .A3(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G143), .ZN(G45));
  NAND2_X1  g521(.A1(new_n671), .A2(new_n675), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n334), .B1(new_n628), .B2(new_n327), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n674), .B1(new_n709), .B2(KEYINPUT32), .ZN(new_n710));
  OAI211_X1 g524(.A(new_n546), .B(new_n660), .C1(new_n708), .C2(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n644), .A2(new_n679), .ZN(new_n713));
  OAI211_X1 g527(.A(new_n712), .B(new_n713), .C1(new_n618), .C2(new_n619), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G146), .ZN(G48));
  INV_X1    g529(.A(KEYINPUT108), .ZN(new_n716));
  INV_X1    g530(.A(new_n234), .ZN(new_n717));
  OR2_X1    g531(.A1(new_n590), .A2(new_n611), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n579), .A2(new_n580), .ZN(new_n719));
  AOI21_X1  g533(.A(KEYINPUT80), .B1(new_n590), .B2(new_n548), .ZN(new_n720));
  OAI211_X1 g534(.A(new_n617), .B(new_n718), .C1(new_n719), .C2(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT107), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n592), .A2(KEYINPUT107), .A3(new_n617), .A4(new_n718), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n676), .A2(new_n717), .A3(new_n723), .A4(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(new_n642), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n726), .B1(new_n416), .B2(G478), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n635), .B1(new_n408), .B2(new_n415), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n417), .B1(new_n728), .B2(new_n637), .ZN(new_n729));
  NOR3_X1   g543(.A1(new_n727), .A2(new_n729), .A3(new_n467), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n730), .A2(new_n546), .A3(new_n357), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n716), .B1(new_n725), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n723), .A2(new_n724), .ZN(new_n733));
  INV_X1    g547(.A(new_n733), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n734), .A2(new_n350), .A3(KEYINPUT108), .A4(new_n645), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(KEYINPUT41), .B(G113), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n736), .B(new_n737), .ZN(G15));
  AND4_X1   g552(.A1(new_n676), .A2(new_n717), .A3(new_n723), .A4(new_n724), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(new_n652), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G116), .ZN(G18));
  AND3_X1   g555(.A1(new_n723), .A2(new_n468), .A3(new_n724), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n661), .B1(new_n339), .B2(new_n349), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n742), .A2(KEYINPUT109), .A3(new_n546), .A4(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT109), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n723), .A2(new_n468), .A3(new_n724), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n745), .B1(new_n711), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n744), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G119), .ZN(G21));
  INV_X1    g563(.A(new_n627), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n334), .B1(new_n320), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n332), .A2(new_n219), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n751), .B1(new_n752), .B2(G472), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(new_n717), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n633), .A2(new_n650), .A3(new_n691), .A4(new_n357), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n734), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G122), .ZN(G24));
  NAND3_X1  g572(.A1(new_n723), .A2(new_n546), .A3(new_n724), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n727), .A2(new_n729), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n760), .A2(new_n641), .A3(new_n678), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n753), .A2(new_n660), .ZN(new_n762));
  NOR3_X1   g576(.A1(new_n759), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(new_n198), .ZN(G27));
  NAND3_X1  g578(.A1(new_n544), .A2(new_n469), .A3(new_n545), .ZN(new_n765));
  INV_X1    g579(.A(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(G469), .A2(G902), .ZN(new_n767));
  XOR2_X1   g581(.A(new_n767), .B(KEYINPUT110), .Z(new_n768));
  NOR2_X1   g582(.A1(new_n601), .A2(new_n602), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n768), .B1(new_n769), .B2(G469), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n616), .B1(new_n770), .B2(new_n592), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n730), .A2(new_n766), .A3(new_n771), .A4(new_n678), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT111), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n669), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n332), .A2(KEYINPUT111), .A3(new_n336), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n717), .B1(new_n776), .B2(new_n710), .ZN(new_n777));
  OAI21_X1  g591(.A(KEYINPUT42), .B1(new_n772), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n770), .A2(new_n592), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(new_n617), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n780), .A2(new_n765), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT42), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n781), .A2(new_n350), .A3(new_n782), .A4(new_n713), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n778), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(new_n244), .ZN(G33));
  NAND3_X1  g599(.A1(new_n781), .A2(new_n350), .A3(new_n680), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G134), .ZN(G36));
  INV_X1    g601(.A(new_n768), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n769), .A2(KEYINPUT45), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(G469), .ZN(new_n790));
  AOI21_X1  g604(.A(KEYINPUT45), .B1(new_n603), .B2(new_n609), .ZN(new_n791));
  OAI211_X1 g605(.A(KEYINPUT46), .B(new_n788), .C1(new_n790), .C2(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n792), .A2(KEYINPUT112), .A3(new_n592), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT46), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n790), .A2(new_n791), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n794), .B1(new_n795), .B2(new_n768), .ZN(new_n796));
  AND2_X1   g610(.A1(new_n793), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n792), .A2(new_n592), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT112), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n616), .B1(new_n797), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n760), .A2(new_n467), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n802), .A2(KEYINPUT43), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n630), .A2(new_n660), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT43), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n760), .A2(new_n805), .A3(new_n467), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n803), .A2(new_n804), .A3(KEYINPUT44), .A4(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n803), .A2(new_n804), .A3(new_n806), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT44), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n765), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n801), .A2(new_n685), .A3(new_n807), .A4(new_n810), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n811), .B(G137), .ZN(G39));
  NAND2_X1  g626(.A1(new_n713), .A2(new_n766), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n813), .A2(new_n676), .A3(new_n717), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n797), .A2(new_n800), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n815), .A2(KEYINPUT47), .A3(new_n617), .ZN(new_n816));
  INV_X1    g630(.A(new_n816), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n801), .A2(KEYINPUT47), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n814), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(G140), .ZN(G42));
  NAND3_X1  g634(.A1(new_n717), .A2(new_n617), .A3(new_n469), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n592), .A2(new_n718), .ZN(new_n822));
  AOI211_X1 g636(.A(new_n821), .B(new_n802), .C1(KEYINPUT49), .C2(new_n822), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n823), .B(KEYINPUT113), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n822), .A2(KEYINPUT49), .ZN(new_n825));
  OR4_X1    g639(.A1(new_n694), .A2(new_n824), .A3(new_n699), .A4(new_n825), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n733), .A2(new_n765), .ZN(new_n827));
  INV_X1    g641(.A(new_n699), .ZN(new_n828));
  INV_X1    g642(.A(new_n353), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n827), .A2(new_n717), .A3(new_n828), .A4(new_n829), .ZN(new_n830));
  OR3_X1    g644(.A1(new_n830), .A2(new_n641), .A3(new_n760), .ZN(new_n831));
  AND2_X1   g645(.A1(new_n803), .A2(new_n806), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n832), .A2(new_n829), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n833), .A2(new_n827), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n831), .B1(new_n834), .B2(new_n762), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT114), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT51), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  OR2_X1    g653(.A1(new_n801), .A2(KEYINPUT47), .ZN(new_n840));
  OAI211_X1 g654(.A(new_n840), .B(new_n816), .C1(new_n617), .C2(new_n822), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n832), .A2(new_n717), .A3(new_n829), .A4(new_n753), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n842), .A2(new_n765), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  OR3_X1    g658(.A1(new_n694), .A2(new_n733), .A3(new_n469), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n842), .A2(new_n845), .ZN(new_n846));
  OR2_X1    g660(.A1(new_n846), .A2(KEYINPUT50), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(KEYINPUT50), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n835), .A2(new_n836), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n839), .A2(new_n844), .A3(new_n849), .A4(new_n850), .ZN(new_n851));
  OAI221_X1 g665(.A(new_n351), .B1(new_n644), .B2(new_n830), .C1(new_n842), .C2(new_n759), .ZN(new_n852));
  INV_X1    g666(.A(new_n777), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n833), .A2(new_n853), .A3(new_n827), .ZN(new_n854));
  XOR2_X1   g668(.A(KEYINPUT115), .B(KEYINPUT48), .Z(new_n855));
  OR2_X1    g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n854), .A2(new_n855), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n852), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  AOI221_X4 g672(.A(new_n835), .B1(new_n847), .B2(new_n848), .C1(new_n841), .C2(new_n843), .ZN(new_n859));
  OAI211_X1 g673(.A(new_n851), .B(new_n858), .C1(new_n859), .C2(KEYINPUT51), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT54), .ZN(new_n861));
  INV_X1    g675(.A(new_n763), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n780), .A2(new_n660), .A3(new_n679), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n650), .A2(new_n633), .A3(new_n691), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n863), .A2(new_n699), .A3(new_n864), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n682), .A2(new_n714), .A3(new_n862), .A4(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(KEYINPUT52), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n763), .B1(new_n626), .B2(new_n681), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT52), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n868), .A2(new_n869), .A3(new_n714), .A4(new_n865), .ZN(new_n870));
  AND2_X1   g684(.A1(new_n867), .A2(new_n870), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n778), .A2(new_n783), .A3(new_n786), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n679), .B1(new_n231), .B2(new_n659), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n873), .A2(new_n419), .A3(new_n424), .A4(new_n467), .ZN(new_n874));
  AOI211_X1 g688(.A(new_n765), .B(new_n874), .C1(new_n339), .C2(new_n349), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n761), .A2(new_n762), .ZN(new_n876));
  AOI22_X1  g690(.A1(new_n626), .A2(new_n875), .B1(new_n876), .B2(new_n781), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n872), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n736), .A2(new_n663), .A3(new_n748), .ZN(new_n879));
  OAI221_X1 g693(.A(new_n631), .B1(new_n645), .B2(new_n652), .C1(new_n618), .C2(new_n619), .ZN(new_n880));
  AOI22_X1  g694(.A1(new_n739), .A2(new_n652), .B1(new_n734), .B2(new_n756), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n880), .A2(new_n881), .A3(new_n620), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n878), .A2(new_n879), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n682), .A2(new_n862), .ZN(new_n884));
  AOI21_X1  g698(.A(KEYINPUT53), .B1(new_n884), .B2(KEYINPUT52), .ZN(new_n885));
  INV_X1    g699(.A(new_n885), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n871), .A2(new_n883), .A3(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT53), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n867), .A2(new_n870), .ZN(new_n889));
  AND3_X1   g703(.A1(new_n736), .A2(new_n663), .A3(new_n748), .ZN(new_n890));
  AND3_X1   g704(.A1(new_n880), .A2(new_n881), .A3(new_n620), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n875), .B1(new_n618), .B2(new_n619), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n876), .A2(new_n781), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n778), .A2(new_n783), .A3(new_n786), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n890), .A2(new_n891), .A3(new_n896), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n888), .B1(new_n889), .B2(new_n897), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n861), .B1(new_n887), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g713(.A(KEYINPUT53), .B1(new_n868), .B2(new_n869), .ZN(new_n900));
  INV_X1    g714(.A(new_n900), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n883), .A2(new_n867), .A3(new_n870), .A4(new_n901), .ZN(new_n902));
  AND3_X1   g716(.A1(new_n898), .A2(new_n902), .A3(new_n861), .ZN(new_n903));
  NOR3_X1   g717(.A1(new_n860), .A2(new_n899), .A3(new_n903), .ZN(new_n904));
  NOR2_X1   g718(.A1(G952), .A2(G953), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n826), .B1(new_n904), .B2(new_n905), .ZN(G75));
  AOI21_X1  g720(.A(new_n219), .B1(new_n898), .B2(new_n902), .ZN(new_n907));
  AOI21_X1  g721(.A(KEYINPUT56), .B1(new_n907), .B2(G210), .ZN(new_n908));
  AND2_X1   g722(.A1(new_n512), .A2(new_n514), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n909), .B(new_n520), .ZN(new_n910));
  XNOR2_X1  g724(.A(KEYINPUT116), .B(KEYINPUT55), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n910), .B(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(new_n912), .ZN(new_n913));
  OAI22_X1  g727(.A1(new_n908), .A2(new_n913), .B1(G952), .B2(new_n215), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n914), .B1(new_n908), .B2(new_n913), .ZN(G51));
  NOR2_X1   g729(.A1(new_n215), .A2(G952), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n898), .A2(new_n902), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(KEYINPUT54), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n898), .A2(new_n902), .A3(new_n861), .ZN(new_n919));
  AND2_X1   g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n768), .B(KEYINPUT57), .Z(new_n921));
  OAI22_X1  g735(.A1(new_n920), .A2(new_n921), .B1(new_n578), .B2(new_n575), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n907), .A2(new_n795), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n916), .B1(new_n922), .B2(new_n923), .ZN(G54));
  NAND2_X1  g738(.A1(KEYINPUT58), .A2(G475), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n925), .B(KEYINPUT117), .Z(new_n926));
  NAND2_X1  g740(.A1(new_n907), .A2(new_n926), .ZN(new_n927));
  AND2_X1   g741(.A1(new_n927), .A2(new_n458), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n927), .A2(new_n458), .ZN(new_n929));
  NOR3_X1   g743(.A1(new_n928), .A2(new_n929), .A3(new_n916), .ZN(G60));
  XNOR2_X1  g744(.A(new_n642), .B(KEYINPUT59), .ZN(new_n931));
  AOI21_X1  g745(.A(KEYINPUT53), .B1(new_n871), .B2(new_n883), .ZN(new_n932));
  NOR3_X1   g746(.A1(new_n889), .A2(new_n897), .A3(new_n885), .ZN(new_n933));
  OAI21_X1  g747(.A(KEYINPUT54), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n931), .B1(new_n934), .B2(new_n919), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n638), .A2(new_n639), .ZN(new_n936));
  OAI21_X1  g750(.A(KEYINPUT118), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT118), .ZN(new_n938));
  INV_X1    g752(.A(new_n936), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n903), .A2(new_n899), .ZN(new_n940));
  OAI211_X1 g754(.A(new_n938), .B(new_n939), .C1(new_n940), .C2(new_n931), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n918), .A2(new_n919), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n939), .A2(new_n931), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n916), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  AND3_X1   g758(.A1(new_n937), .A2(new_n941), .A3(new_n944), .ZN(G63));
  XNOR2_X1  g759(.A(new_n225), .B(KEYINPUT60), .ZN(new_n946));
  INV_X1    g760(.A(new_n946), .ZN(new_n947));
  NOR3_X1   g761(.A1(new_n889), .A2(new_n897), .A3(new_n900), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n947), .B1(new_n932), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n218), .A2(new_n222), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n916), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT120), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n657), .A2(new_n658), .ZN(new_n953));
  XOR2_X1   g767(.A(new_n953), .B(KEYINPUT119), .Z(new_n954));
  AND4_X1   g768(.A1(new_n952), .A2(new_n917), .A3(new_n947), .A4(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n946), .B1(new_n898), .B2(new_n902), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n952), .B1(new_n956), .B2(new_n954), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n951), .B1(new_n955), .B2(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT61), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  OAI211_X1 g774(.A(new_n951), .B(KEYINPUT61), .C1(new_n955), .C2(new_n957), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n960), .A2(new_n961), .ZN(G66));
  OAI21_X1  g776(.A(G953), .B1(new_n354), .B2(new_n517), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n879), .A2(new_n882), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n963), .B1(new_n964), .B2(G953), .ZN(new_n965));
  INV_X1    g779(.A(new_n909), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n966), .B1(G898), .B2(new_n215), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n965), .B(new_n967), .ZN(G69));
  XOR2_X1   g782(.A(new_n454), .B(KEYINPUT121), .Z(new_n969));
  XNOR2_X1  g783(.A(new_n281), .B(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n765), .B1(new_n651), .B2(new_n644), .ZN(new_n971));
  NAND4_X1  g785(.A1(new_n626), .A2(new_n350), .A3(new_n685), .A4(new_n971), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n819), .A2(new_n811), .A3(new_n972), .ZN(new_n973));
  AND2_X1   g787(.A1(new_n868), .A2(new_n714), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n706), .A2(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT62), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n706), .A2(KEYINPUT62), .A3(new_n974), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n973), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n970), .B1(new_n979), .B2(G953), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT123), .ZN(new_n981));
  INV_X1    g795(.A(new_n814), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n982), .B1(new_n840), .B2(new_n816), .ZN(new_n983));
  NAND4_X1  g797(.A1(new_n801), .A2(new_n685), .A3(new_n864), .A4(new_n853), .ZN(new_n984));
  NAND4_X1  g798(.A1(new_n811), .A2(new_n984), .A3(new_n872), .A4(new_n974), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n981), .B1(new_n983), .B2(new_n985), .ZN(new_n986));
  AND3_X1   g800(.A1(new_n811), .A2(new_n872), .A3(new_n974), .ZN(new_n987));
  NAND4_X1  g801(.A1(new_n987), .A2(new_n819), .A3(KEYINPUT123), .A4(new_n984), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n986), .A2(new_n988), .A3(new_n215), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n970), .B1(G900), .B2(G953), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n980), .A2(new_n991), .ZN(new_n992));
  INV_X1    g806(.A(KEYINPUT124), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n980), .A2(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(G900), .ZN(new_n995));
  OAI21_X1  g809(.A(G953), .B1(new_n559), .B2(new_n995), .ZN(new_n996));
  XNOR2_X1  g810(.A(new_n996), .B(KEYINPUT122), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n992), .A2(new_n994), .A3(new_n997), .ZN(new_n998));
  INV_X1    g812(.A(new_n997), .ZN(new_n999));
  OAI211_X1 g813(.A(new_n980), .B(new_n991), .C1(new_n993), .C2(new_n999), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n998), .A2(new_n1000), .ZN(G72));
  NOR3_X1   g815(.A1(new_n314), .A2(new_n317), .A3(new_n310), .ZN(new_n1002));
  AND3_X1   g816(.A1(new_n986), .A2(new_n988), .A3(new_n964), .ZN(new_n1003));
  XNOR2_X1  g817(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n1004));
  NOR2_X1   g818(.A1(new_n340), .A2(new_n219), .ZN(new_n1005));
  XOR2_X1   g819(.A(new_n1004), .B(new_n1005), .Z(new_n1006));
  OAI21_X1  g820(.A(new_n1002), .B1(new_n1003), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n887), .A2(new_n898), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n1006), .B1(new_n311), .B2(new_n345), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n916), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1007), .A2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n1006), .B1(new_n979), .B2(new_n964), .ZN(new_n1012));
  INV_X1    g826(.A(KEYINPUT126), .ZN(new_n1013));
  OR2_X1    g827(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g828(.A(new_n695), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n1015), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n1011), .B1(new_n1014), .B2(new_n1016), .ZN(G57));
endmodule


