//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 0 1 0 1 0 1 0 1 1 0 0 0 0 0 0 0 1 1 1 1 0 0 0 0 1 1 1 0 1 1 1 0 0 1 1 0 0 1 1 1 0 1 1 0 0 1 0 0 1 0 0 1 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:33 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n761, new_n762, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n782, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023;
  XNOR2_X1  g000(.A(G110), .B(G140), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  AND2_X1   g002(.A1(new_n188), .A2(G227), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n187), .B(new_n189), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT78), .B(G101), .ZN(new_n191));
  INV_X1    g005(.A(G104), .ZN(new_n192));
  OAI21_X1  g006(.A(KEYINPUT3), .B1(new_n192), .B2(G107), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT3), .ZN(new_n194));
  INV_X1    g008(.A(G107), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n194), .A2(new_n195), .A3(G104), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n192), .A2(G107), .ZN(new_n197));
  NAND4_X1  g011(.A1(new_n191), .A2(new_n193), .A3(new_n196), .A4(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G143), .ZN(new_n199));
  OAI21_X1  g013(.A(KEYINPUT1), .B1(new_n199), .B2(G146), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n199), .A2(G146), .ZN(new_n201));
  INV_X1    g015(.A(G146), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n202), .A2(G143), .ZN(new_n203));
  OAI211_X1 g017(.A(G128), .B(new_n200), .C1(new_n201), .C2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n202), .A2(G143), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n199), .A2(G146), .ZN(new_n206));
  INV_X1    g020(.A(G128), .ZN(new_n207));
  OAI211_X1 g021(.A(new_n205), .B(new_n206), .C1(KEYINPUT1), .C2(new_n207), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n192), .A2(G107), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n195), .A2(G104), .ZN(new_n210));
  OAI21_X1  g024(.A(G101), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n198), .A2(new_n204), .A3(new_n208), .A4(new_n211), .ZN(new_n212));
  XNOR2_X1  g026(.A(new_n212), .B(KEYINPUT10), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT64), .ZN(new_n214));
  XNOR2_X1  g028(.A(G143), .B(G146), .ZN(new_n215));
  XNOR2_X1  g029(.A(KEYINPUT0), .B(G128), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  AND2_X1   g031(.A1(KEYINPUT0), .A2(G128), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n205), .A2(new_n206), .ZN(new_n220));
  NOR2_X1   g034(.A1(KEYINPUT0), .A2(G128), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n218), .A2(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n220), .A2(new_n222), .A3(KEYINPUT64), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n217), .A2(new_n219), .A3(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT67), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND4_X1  g040(.A1(new_n217), .A2(new_n223), .A3(KEYINPUT67), .A4(new_n219), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n193), .A2(new_n196), .A3(new_n197), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(G101), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n229), .A2(KEYINPUT4), .A3(new_n198), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT4), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n228), .A2(new_n231), .A3(G101), .ZN(new_n232));
  NAND4_X1  g046(.A1(new_n226), .A2(new_n227), .A3(new_n230), .A4(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT11), .ZN(new_n234));
  INV_X1    g048(.A(G134), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n234), .B1(new_n235), .B2(G137), .ZN(new_n236));
  INV_X1    g050(.A(G137), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n237), .A2(KEYINPUT11), .A3(G134), .ZN(new_n238));
  AND2_X1   g052(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  AOI21_X1  g053(.A(G131), .B1(new_n235), .B2(G137), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n235), .A2(G137), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n236), .A2(new_n238), .A3(new_n241), .ZN(new_n242));
  AOI22_X1  g056(.A1(new_n239), .A2(new_n240), .B1(new_n242), .B2(G131), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n213), .A2(new_n233), .A3(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n243), .B1(new_n213), .B2(new_n233), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n190), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n190), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n198), .A2(new_n211), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n204), .A2(new_n208), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(new_n212), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n242), .A2(G131), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n236), .A2(new_n240), .A3(new_n238), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT12), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT79), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n256), .B1(new_n243), .B2(new_n257), .ZN(new_n258));
  AND3_X1   g072(.A1(new_n252), .A2(new_n255), .A3(new_n258), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n258), .B1(new_n252), .B2(new_n255), .ZN(new_n260));
  OAI211_X1 g074(.A(new_n244), .B(new_n248), .C1(new_n259), .C2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n247), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(G469), .ZN(new_n263));
  INV_X1    g077(.A(G902), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n262), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  AND2_X1   g079(.A1(new_n244), .A2(new_n248), .ZN(new_n266));
  INV_X1    g080(.A(new_n246), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n244), .B1(new_n259), .B2(new_n260), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(new_n190), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n268), .A2(G469), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(G469), .A2(G902), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n265), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(G221), .ZN(new_n274));
  XNOR2_X1  g088(.A(KEYINPUT9), .B(G234), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n274), .B1(new_n276), .B2(new_n264), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n273), .A2(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(G478), .B1(KEYINPUT94), .B2(KEYINPUT15), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n280), .B1(KEYINPUT94), .B2(KEYINPUT15), .ZN(new_n281));
  INV_X1    g095(.A(G217), .ZN(new_n282));
  NOR3_X1   g096(.A1(new_n275), .A2(new_n282), .A3(G953), .ZN(new_n283));
  INV_X1    g097(.A(G116), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(G122), .ZN(new_n285));
  XNOR2_X1  g099(.A(new_n285), .B(KEYINPUT93), .ZN(new_n286));
  OR2_X1    g100(.A1(new_n286), .A2(KEYINPUT14), .ZN(new_n287));
  INV_X1    g101(.A(G122), .ZN(new_n288));
  AOI22_X1  g102(.A1(new_n286), .A2(KEYINPUT14), .B1(G116), .B2(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n195), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n288), .A2(G116), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n286), .A2(new_n195), .A3(new_n291), .ZN(new_n292));
  XNOR2_X1  g106(.A(G128), .B(G143), .ZN(new_n293));
  XNOR2_X1  g107(.A(new_n293), .B(new_n235), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  OR2_X1    g109(.A1(new_n290), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n207), .A2(G143), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT13), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n297), .A2(new_n298), .A3(G134), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n294), .A2(new_n299), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n293), .A2(new_n298), .A3(G134), .A4(new_n297), .ZN(new_n301));
  INV_X1    g115(.A(new_n292), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n195), .B1(new_n286), .B2(new_n291), .ZN(new_n303));
  OAI211_X1 g117(.A(new_n300), .B(new_n301), .C1(new_n302), .C2(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n283), .B1(new_n296), .B2(new_n304), .ZN(new_n305));
  OAI211_X1 g119(.A(new_n304), .B(new_n283), .C1(new_n290), .C2(new_n295), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n264), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT95), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n304), .B1(new_n290), .B2(new_n295), .ZN(new_n311));
  INV_X1    g125(.A(new_n283), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  AOI21_X1  g127(.A(G902), .B1(new_n313), .B2(new_n306), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(KEYINPUT95), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n281), .B1(new_n310), .B2(new_n315), .ZN(new_n316));
  AND2_X1   g130(.A1(new_n315), .A2(new_n281), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  NOR2_X1   g133(.A1(G475), .A2(G902), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT89), .ZN(new_n322));
  INV_X1    g136(.A(G140), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G125), .ZN(new_n324));
  INV_X1    g138(.A(G125), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(G140), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n324), .A2(new_n326), .A3(KEYINPUT16), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT16), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n328), .A2(new_n323), .A3(G125), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n327), .A2(new_n329), .A3(G146), .ZN(new_n330));
  NAND2_X1  g144(.A1(KEYINPUT88), .A2(KEYINPUT19), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n324), .A2(new_n326), .A3(new_n331), .ZN(new_n332));
  XOR2_X1   g146(.A(KEYINPUT88), .B(KEYINPUT19), .Z(new_n333));
  XNOR2_X1  g147(.A(G125), .B(G140), .ZN(new_n334));
  OAI211_X1 g148(.A(new_n332), .B(new_n202), .C1(new_n333), .C2(new_n334), .ZN(new_n335));
  NOR2_X1   g149(.A1(G237), .A2(G953), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n336), .A2(G143), .A3(G214), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  AOI21_X1  g152(.A(G143), .B1(new_n336), .B2(G214), .ZN(new_n339));
  NOR3_X1   g153(.A1(new_n338), .A2(new_n339), .A3(G131), .ZN(new_n340));
  INV_X1    g154(.A(G131), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n336), .A2(G214), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(new_n199), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n341), .B1(new_n343), .B2(new_n337), .ZN(new_n344));
  OAI211_X1 g158(.A(new_n330), .B(new_n335), .C1(new_n340), .C2(new_n344), .ZN(new_n345));
  OAI211_X1 g159(.A(KEYINPUT18), .B(G131), .C1(new_n338), .C2(new_n339), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n324), .A2(new_n326), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(G146), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n334), .A2(new_n202), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(KEYINPUT18), .A2(G131), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n343), .A2(new_n337), .A3(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n346), .A2(new_n350), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n345), .A2(new_n353), .ZN(new_n354));
  XNOR2_X1  g168(.A(G113), .B(G122), .ZN(new_n355));
  XNOR2_X1  g169(.A(new_n355), .B(new_n192), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n322), .B1(new_n354), .B2(new_n357), .ZN(new_n358));
  AOI211_X1 g172(.A(KEYINPUT89), .B(new_n356), .C1(new_n345), .C2(new_n353), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT75), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n330), .A2(new_n361), .ZN(new_n362));
  AOI21_X1  g176(.A(G146), .B1(new_n327), .B2(new_n329), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  AOI211_X1 g178(.A(new_n361), .B(G146), .C1(new_n327), .C2(new_n329), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n344), .A2(KEYINPUT17), .ZN(new_n367));
  OAI21_X1  g181(.A(G131), .B1(new_n338), .B2(new_n339), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n343), .A2(new_n341), .A3(new_n337), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n367), .B1(new_n370), .B2(KEYINPUT17), .ZN(new_n371));
  OAI211_X1 g185(.A(new_n356), .B(new_n353), .C1(new_n366), .C2(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n321), .B1(new_n360), .B2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT20), .ZN(new_n374));
  OAI21_X1  g188(.A(KEYINPUT90), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  AND2_X1   g189(.A1(new_n335), .A2(new_n330), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n338), .A2(new_n339), .ZN(new_n377));
  AOI22_X1  g191(.A1(new_n377), .A2(new_n351), .B1(new_n349), .B2(new_n348), .ZN(new_n378));
  AOI22_X1  g192(.A1(new_n376), .A2(new_n370), .B1(new_n378), .B2(new_n346), .ZN(new_n379));
  OAI21_X1  g193(.A(KEYINPUT89), .B1(new_n379), .B2(new_n356), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n354), .A2(new_n322), .A3(new_n357), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n380), .A2(new_n372), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(new_n320), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT90), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n383), .A2(new_n384), .A3(KEYINPUT20), .ZN(new_n385));
  OAI211_X1 g199(.A(new_n375), .B(new_n385), .C1(KEYINPUT20), .C2(new_n383), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n353), .B1(new_n366), .B2(new_n371), .ZN(new_n387));
  OR2_X1    g201(.A1(new_n356), .A2(KEYINPUT92), .ZN(new_n388));
  OR2_X1    g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n387), .A2(new_n388), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n389), .A2(new_n264), .A3(new_n390), .ZN(new_n391));
  XOR2_X1   g205(.A(KEYINPUT91), .B(G475), .Z(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n386), .A2(new_n393), .ZN(new_n394));
  AND2_X1   g208(.A1(new_n188), .A2(G952), .ZN(new_n395));
  NAND2_X1  g209(.A1(G234), .A2(G237), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n396), .A2(G902), .A3(G953), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  XNOR2_X1  g214(.A(KEYINPUT21), .B(G898), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n398), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NOR4_X1   g216(.A1(new_n279), .A2(new_n319), .A3(new_n394), .A4(new_n402), .ZN(new_n403));
  XNOR2_X1  g217(.A(KEYINPUT22), .B(G137), .ZN(new_n404));
  AND3_X1   g218(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n405));
  XOR2_X1   g219(.A(new_n404), .B(new_n405), .Z(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n207), .A2(G119), .ZN(new_n408));
  INV_X1    g222(.A(G119), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(G128), .ZN(new_n410));
  AND3_X1   g224(.A1(new_n408), .A2(new_n410), .A3(KEYINPUT73), .ZN(new_n411));
  AOI21_X1  g225(.A(KEYINPUT73), .B1(new_n408), .B2(new_n410), .ZN(new_n412));
  XNOR2_X1  g226(.A(KEYINPUT24), .B(G110), .ZN(new_n413));
  NOR3_X1   g227(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(KEYINPUT74), .A2(KEYINPUT23), .ZN(new_n415));
  NOR2_X1   g229(.A1(KEYINPUT74), .A2(KEYINPUT23), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n415), .B1(new_n408), .B2(new_n416), .ZN(new_n417));
  XNOR2_X1  g231(.A(G119), .B(G128), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n417), .B1(new_n418), .B2(new_n415), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n414), .B1(G110), .B2(new_n419), .ZN(new_n420));
  OR2_X1    g234(.A1(new_n362), .A2(new_n363), .ZN(new_n421));
  INV_X1    g235(.A(new_n365), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n420), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n330), .A2(new_n349), .ZN(new_n424));
  INV_X1    g238(.A(new_n415), .ZN(new_n425));
  INV_X1    g239(.A(new_n416), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n409), .A2(G128), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n425), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n415), .B1(new_n408), .B2(new_n410), .ZN(new_n429));
  NOR3_X1   g243(.A1(new_n428), .A2(new_n429), .A3(G110), .ZN(new_n430));
  INV_X1    g244(.A(new_n413), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n408), .A2(new_n410), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT73), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n408), .A2(new_n410), .A3(KEYINPUT73), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n431), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  OAI21_X1  g250(.A(KEYINPUT76), .B1(new_n430), .B2(new_n436), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n413), .B1(new_n411), .B2(new_n412), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT76), .ZN(new_n439));
  INV_X1    g253(.A(G110), .ZN(new_n440));
  OAI211_X1 g254(.A(new_n417), .B(new_n440), .C1(new_n418), .C2(new_n415), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n438), .A2(new_n439), .A3(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n424), .B1(new_n437), .B2(new_n442), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n423), .B1(new_n443), .B2(KEYINPUT77), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT77), .ZN(new_n445));
  AOI211_X1 g259(.A(new_n445), .B(new_n424), .C1(new_n437), .C2(new_n442), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n407), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT25), .ZN(new_n448));
  AND3_X1   g262(.A1(new_n438), .A2(new_n439), .A3(new_n441), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n439), .B1(new_n438), .B2(new_n441), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n445), .B1(new_n451), .B2(new_n424), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n443), .A2(KEYINPUT77), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n452), .A2(new_n453), .A3(new_n423), .A4(new_n406), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n447), .A2(new_n448), .A3(new_n454), .A4(new_n264), .ZN(new_n455));
  NAND2_X1  g269(.A1(G217), .A2(G902), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n456), .B1(new_n282), .B2(G234), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n457), .B(KEYINPUT72), .ZN(new_n458));
  AND2_X1   g272(.A1(new_n455), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n447), .A2(new_n264), .A3(new_n454), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(KEYINPUT25), .ZN(new_n461));
  AND2_X1   g275(.A1(new_n447), .A2(new_n454), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n458), .A2(G902), .ZN(new_n463));
  AOI22_X1  g277(.A1(new_n459), .A2(new_n461), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n226), .A2(new_n255), .A3(new_n227), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n409), .A2(G116), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n284), .A2(G119), .ZN(new_n468));
  INV_X1    g282(.A(G113), .ZN(new_n469));
  AND2_X1   g283(.A1(new_n469), .A2(KEYINPUT2), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n469), .A2(KEYINPUT2), .ZN(new_n471));
  OAI211_X1 g285(.A(new_n467), .B(new_n468), .C1(new_n470), .C2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n467), .A2(new_n468), .ZN(new_n473));
  XNOR2_X1  g287(.A(KEYINPUT2), .B(G113), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n237), .A2(G134), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(new_n241), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(G131), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n204), .A2(new_n480), .A3(new_n254), .A4(new_n208), .ZN(new_n481));
  AND2_X1   g295(.A1(new_n477), .A2(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(KEYINPUT28), .B1(new_n466), .B2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT68), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n481), .B(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n485), .A2(new_n466), .A3(new_n477), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n255), .A2(new_n217), .A3(new_n219), .A4(new_n223), .ZN(new_n487));
  AND3_X1   g301(.A1(new_n236), .A2(new_n240), .A3(new_n238), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n341), .B1(new_n478), .B2(new_n241), .ZN(new_n489));
  OAI21_X1  g303(.A(KEYINPUT65), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  AND2_X1   g304(.A1(new_n204), .A2(new_n208), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT65), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n480), .A2(new_n254), .A3(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n490), .A2(new_n491), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n487), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(new_n476), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n486), .A2(new_n496), .ZN(new_n497));
  XOR2_X1   g311(.A(KEYINPUT69), .B(KEYINPUT28), .Z(new_n498));
  AOI21_X1  g312(.A(new_n483), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n336), .A2(G210), .ZN(new_n500));
  XNOR2_X1  g314(.A(new_n500), .B(KEYINPUT27), .ZN(new_n501));
  XNOR2_X1  g315(.A(KEYINPUT26), .B(G101), .ZN(new_n502));
  XNOR2_X1  g316(.A(new_n501), .B(new_n502), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n499), .A2(new_n503), .ZN(new_n504));
  AND2_X1   g318(.A1(new_n486), .A2(new_n503), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT30), .ZN(new_n506));
  AOI21_X1  g320(.A(KEYINPUT66), .B1(new_n495), .B2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT66), .ZN(new_n508));
  AOI211_X1 g322(.A(new_n508), .B(KEYINPUT30), .C1(new_n487), .C2(new_n494), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n485), .A2(new_n466), .A3(KEYINPUT30), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(new_n476), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n505), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT31), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  OAI211_X1 g329(.A(new_n476), .B(new_n511), .C1(new_n507), .C2(new_n509), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n516), .A2(KEYINPUT31), .A3(new_n505), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n504), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g332(.A1(G472), .A2(G902), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  OAI21_X1  g334(.A(KEYINPUT32), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  AND3_X1   g335(.A1(new_n516), .A2(KEYINPUT31), .A3(new_n505), .ZN(new_n522));
  AOI21_X1  g336(.A(KEYINPUT31), .B1(new_n516), .B2(new_n505), .ZN(new_n523));
  OAI22_X1  g337(.A1(new_n522), .A2(new_n523), .B1(new_n503), .B2(new_n499), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT32), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n524), .A2(new_n525), .A3(new_n519), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n521), .A2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT70), .ZN(new_n528));
  INV_X1    g342(.A(new_n486), .ZN(new_n529));
  AND2_X1   g343(.A1(new_n511), .A2(new_n476), .ZN(new_n530));
  AND3_X1   g344(.A1(new_n490), .A2(new_n491), .A3(new_n493), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n224), .A2(new_n243), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n506), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(new_n508), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n495), .A2(KEYINPUT66), .A3(new_n506), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n529), .B1(new_n530), .B2(new_n536), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n528), .B1(new_n537), .B2(new_n503), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n516), .A2(new_n486), .ZN(new_n539));
  INV_X1    g353(.A(new_n503), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n539), .A2(KEYINPUT70), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(KEYINPUT29), .B1(new_n499), .B2(new_n503), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n538), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n486), .A2(KEYINPUT71), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n485), .A2(new_n466), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(new_n476), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT71), .ZN(new_n547));
  NAND4_X1  g361(.A1(new_n485), .A2(new_n466), .A3(new_n547), .A4(new_n477), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n544), .A2(new_n546), .A3(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n483), .B1(new_n549), .B2(KEYINPUT28), .ZN(new_n550));
  AND2_X1   g364(.A1(new_n503), .A2(KEYINPUT29), .ZN(new_n551));
  AOI21_X1  g365(.A(G902), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n543), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(G472), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n465), .B1(new_n527), .B2(new_n554), .ZN(new_n555));
  OAI21_X1  g369(.A(G214), .B1(G237), .B2(G902), .ZN(new_n556));
  OR2_X1    g370(.A1(new_n224), .A2(new_n325), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n491), .A2(new_n325), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(G224), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n561), .A2(G953), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT7), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n562), .B1(KEYINPUT85), .B2(new_n563), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n564), .B1(KEYINPUT85), .B2(new_n563), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n560), .A2(new_n565), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n559), .B1(new_n561), .B2(G953), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n566), .B1(new_n567), .B2(new_n563), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n230), .A2(new_n476), .A3(new_n232), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n284), .A2(G119), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT5), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(KEYINPUT80), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT80), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(KEYINPUT5), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n570), .A2(new_n572), .A3(new_n574), .ZN(new_n575));
  XNOR2_X1  g389(.A(KEYINPUT80), .B(KEYINPUT5), .ZN(new_n576));
  OAI211_X1 g390(.A(new_n575), .B(G113), .C1(new_n473), .C2(new_n576), .ZN(new_n577));
  NAND4_X1  g391(.A1(new_n577), .A2(new_n472), .A3(new_n198), .A4(new_n211), .ZN(new_n578));
  XNOR2_X1  g392(.A(G110), .B(G122), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n569), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n473), .A2(new_n571), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n469), .B1(new_n576), .B2(new_n570), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT84), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n581), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n585), .B1(new_n584), .B2(new_n583), .ZN(new_n586));
  AND3_X1   g400(.A1(new_n198), .A2(new_n472), .A3(new_n211), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n577), .A2(new_n472), .ZN(new_n588));
  AOI22_X1  g402(.A1(new_n586), .A2(new_n587), .B1(new_n249), .B2(new_n588), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n579), .B(KEYINPUT8), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n580), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n264), .B1(new_n568), .B2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  OAI21_X1  g408(.A(G210), .B1(G237), .B2(G902), .ZN(new_n595));
  XOR2_X1   g409(.A(new_n595), .B(KEYINPUT86), .Z(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n560), .A2(new_n562), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(new_n567), .ZN(new_n599));
  AND3_X1   g413(.A1(new_n229), .A2(KEYINPUT4), .A3(new_n198), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n476), .A2(new_n232), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n578), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(KEYINPUT81), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT81), .ZN(new_n604));
  OAI211_X1 g418(.A(new_n604), .B(new_n578), .C1(new_n600), .C2(new_n601), .ZN(new_n605));
  INV_X1    g419(.A(new_n579), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n603), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  AND2_X1   g421(.A1(new_n580), .A2(KEYINPUT6), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n605), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n604), .B1(new_n569), .B2(new_n578), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n579), .A2(KEYINPUT6), .ZN(new_n613));
  AOI21_X1  g427(.A(KEYINPUT82), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND4_X1  g428(.A1(new_n603), .A2(KEYINPUT82), .A3(new_n605), .A4(new_n613), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  OAI211_X1 g430(.A(new_n599), .B(new_n609), .C1(new_n614), .C2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT83), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n603), .A2(new_n605), .A3(new_n613), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT82), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  AOI22_X1  g436(.A1(new_n622), .A2(new_n615), .B1(new_n607), .B2(new_n608), .ZN(new_n623));
  AOI21_X1  g437(.A(KEYINPUT83), .B1(new_n623), .B2(new_n599), .ZN(new_n624));
  OAI211_X1 g438(.A(new_n594), .B(new_n597), .C1(new_n619), .C2(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n617), .A2(new_n618), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n623), .A2(KEYINPUT83), .A3(new_n599), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n593), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  XOR2_X1   g442(.A(new_n596), .B(KEYINPUT87), .Z(new_n629));
  OAI21_X1  g443(.A(new_n625), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND4_X1  g444(.A1(new_n403), .A2(new_n555), .A3(new_n556), .A4(new_n630), .ZN(new_n631));
  XOR2_X1   g445(.A(new_n631), .B(new_n191), .Z(G3));
  NAND2_X1  g446(.A1(new_n524), .A2(new_n264), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(G472), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n524), .A2(new_n519), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NOR3_X1   g450(.A1(new_n636), .A2(new_n279), .A3(new_n465), .ZN(new_n637));
  XOR2_X1   g451(.A(new_n637), .B(KEYINPUT96), .Z(new_n638));
  NAND2_X1  g452(.A1(new_n626), .A2(new_n627), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n597), .B1(new_n639), .B2(new_n594), .ZN(new_n640));
  AOI211_X1 g454(.A(new_n593), .B(new_n596), .C1(new_n626), .C2(new_n627), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n556), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(KEYINPUT97), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT97), .ZN(new_n644));
  OAI211_X1 g458(.A(new_n644), .B(new_n556), .C1(new_n640), .C2(new_n641), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT33), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT98), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n646), .B1(new_n306), .B2(new_n647), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n648), .B1(new_n307), .B2(new_n305), .ZN(new_n649));
  OAI211_X1 g463(.A(new_n313), .B(new_n306), .C1(new_n647), .C2(new_n646), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n649), .A2(G478), .A3(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(G478), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n652), .A2(new_n264), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n653), .B1(new_n314), .B2(new_n652), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  AOI211_X1 g469(.A(new_n402), .B(new_n655), .C1(new_n386), .C2(new_n393), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n643), .A2(new_n645), .A3(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n638), .A2(new_n658), .ZN(new_n659));
  XOR2_X1   g473(.A(KEYINPUT34), .B(G104), .Z(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G6));
  NOR2_X1   g475(.A1(new_n383), .A2(KEYINPUT20), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT99), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n384), .B1(new_n383), .B2(KEYINPUT20), .ZN(new_n664));
  AOI211_X1 g478(.A(KEYINPUT90), .B(new_n374), .C1(new_n382), .C2(new_n320), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n663), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n375), .A2(KEYINPUT99), .A3(new_n385), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n662), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n393), .B1(new_n316), .B2(new_n317), .ZN(new_n669));
  NOR3_X1   g483(.A1(new_n668), .A2(new_n669), .A3(new_n402), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n643), .A2(new_n645), .A3(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n638), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G107), .ZN(new_n674));
  XNOR2_X1  g488(.A(KEYINPUT100), .B(KEYINPUT35), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G9));
  NAND3_X1  g490(.A1(new_n403), .A2(new_n556), .A3(new_n630), .ZN(new_n677));
  INV_X1    g491(.A(new_n636), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n452), .A2(new_n453), .A3(new_n423), .ZN(new_n679));
  OR2_X1    g493(.A1(new_n407), .A2(KEYINPUT36), .ZN(new_n680));
  OR2_X1    g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n679), .A2(new_n680), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n681), .A2(new_n463), .A3(new_n682), .ZN(new_n683));
  AND2_X1   g497(.A1(new_n460), .A2(KEYINPUT25), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n455), .A2(new_n458), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n683), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT101), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  OAI211_X1 g502(.A(KEYINPUT101), .B(new_n683), .C1(new_n684), .C2(new_n685), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n678), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n677), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(KEYINPUT37), .B(G110), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(KEYINPUT102), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n692), .B(new_n694), .ZN(G12));
  NAND2_X1  g509(.A1(new_n527), .A2(new_n554), .ZN(new_n696));
  XOR2_X1   g510(.A(KEYINPUT103), .B(G900), .Z(new_n697));
  AOI21_X1  g511(.A(new_n398), .B1(new_n400), .B2(new_n697), .ZN(new_n698));
  NOR3_X1   g512(.A1(new_n668), .A2(new_n669), .A3(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(new_n279), .ZN(new_n700));
  AND4_X1   g514(.A1(new_n696), .A2(new_n699), .A3(new_n700), .A4(new_n690), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n701), .A2(KEYINPUT104), .A3(new_n645), .A4(new_n643), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT104), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n643), .A2(new_n645), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n696), .A2(new_n699), .A3(new_n700), .A4(new_n690), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n703), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n702), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G128), .ZN(G30));
  XOR2_X1   g522(.A(new_n698), .B(KEYINPUT39), .Z(new_n709));
  NAND2_X1  g523(.A1(new_n700), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(KEYINPUT40), .ZN(new_n711));
  INV_X1    g525(.A(new_n394), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n712), .A2(new_n318), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n711), .A2(new_n556), .A3(new_n713), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n710), .A2(KEYINPUT40), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n630), .B(KEYINPUT38), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n539), .A2(new_n503), .ZN(new_n718));
  OR2_X1    g532(.A1(new_n549), .A2(new_n503), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n718), .A2(new_n719), .A3(KEYINPUT105), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(new_n264), .ZN(new_n721));
  AOI21_X1  g535(.A(KEYINPUT105), .B1(new_n718), .B2(new_n719), .ZN(new_n722));
  OAI21_X1  g536(.A(G472), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n527), .A2(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(new_n724), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n725), .A2(new_n690), .ZN(new_n726));
  AND3_X1   g540(.A1(new_n716), .A2(new_n717), .A3(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(new_n199), .ZN(G45));
  AOI21_X1  g542(.A(new_n279), .B1(new_n527), .B2(new_n554), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(new_n690), .ZN(new_n730));
  AOI211_X1 g544(.A(new_n698), .B(new_n655), .C1(new_n386), .C2(new_n393), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n643), .A2(new_n645), .A3(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT106), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n643), .A2(KEYINPUT106), .A3(new_n645), .A4(new_n731), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n730), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(new_n202), .ZN(G48));
  INV_X1    g551(.A(new_n555), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n263), .B1(new_n262), .B2(new_n264), .ZN(new_n739));
  AOI211_X1 g553(.A(G469), .B(G902), .C1(new_n247), .C2(new_n261), .ZN(new_n740));
  OR2_X1    g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n741), .A2(new_n277), .ZN(new_n742));
  INV_X1    g556(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n738), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n658), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(KEYINPUT41), .B(G113), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n745), .B(new_n746), .ZN(G15));
  NAND2_X1  g561(.A1(new_n672), .A2(new_n744), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G116), .ZN(G18));
  NAND3_X1  g563(.A1(new_n643), .A2(new_n645), .A3(new_n742), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n394), .A2(new_n402), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n696), .A2(new_n751), .A3(new_n318), .A4(new_n690), .ZN(new_n752));
  OR2_X1    g566(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G119), .ZN(G21));
  OAI22_X1  g568(.A1(new_n522), .A2(new_n523), .B1(new_n550), .B2(new_n503), .ZN(new_n755));
  AOI22_X1  g569(.A1(new_n633), .A2(G472), .B1(new_n519), .B2(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(new_n402), .ZN(new_n757));
  AND4_X1   g571(.A1(new_n464), .A2(new_n756), .A3(new_n742), .A4(new_n757), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n758), .A2(new_n645), .A3(new_n643), .A4(new_n713), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G122), .ZN(G24));
  AND3_X1   g574(.A1(new_n690), .A2(new_n731), .A3(new_n756), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n761), .A2(new_n643), .A3(new_n645), .A4(new_n742), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G125), .ZN(G27));
  INV_X1    g577(.A(KEYINPUT42), .ZN(new_n764));
  OAI211_X1 g578(.A(new_n625), .B(new_n556), .C1(new_n628), .C2(new_n629), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n272), .B(KEYINPUT107), .ZN(new_n766));
  INV_X1    g580(.A(new_n766), .ZN(new_n767));
  AOI22_X1  g581(.A1(new_n267), .A2(new_n266), .B1(new_n269), .B2(new_n190), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n767), .B1(new_n768), .B2(G469), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n277), .B1(new_n769), .B2(new_n265), .ZN(new_n770));
  INV_X1    g584(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n765), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n772), .A2(new_n555), .A3(new_n731), .ZN(new_n773));
  AOI211_X1 g587(.A(KEYINPUT109), .B(new_n764), .C1(new_n773), .C2(KEYINPUT108), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(KEYINPUT109), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(KEYINPUT42), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n773), .A2(KEYINPUT108), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT109), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n774), .B1(new_n776), .B2(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(new_n341), .ZN(G33));
  NAND3_X1  g595(.A1(new_n772), .A2(new_n555), .A3(new_n699), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G134), .ZN(G36));
  INV_X1    g597(.A(new_n655), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n712), .A2(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(KEYINPUT43), .ZN(new_n786));
  OR2_X1    g600(.A1(new_n786), .A2(KEYINPUT110), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(KEYINPUT110), .ZN(new_n788));
  INV_X1    g602(.A(new_n690), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n678), .A2(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n787), .A2(new_n788), .A3(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT44), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n787), .A2(new_n788), .A3(KEYINPUT44), .A4(new_n790), .ZN(new_n794));
  OR2_X1    g608(.A1(new_n768), .A2(KEYINPUT45), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n768), .A2(KEYINPUT45), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n795), .A2(G469), .A3(new_n796), .ZN(new_n797));
  AOI21_X1  g611(.A(KEYINPUT46), .B1(new_n797), .B2(new_n766), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n798), .A2(new_n740), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n797), .A2(KEYINPUT46), .A3(new_n766), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n277), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(new_n709), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n802), .A2(new_n765), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n793), .A2(new_n794), .A3(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(KEYINPUT111), .B(G137), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n804), .B(new_n805), .ZN(G39));
  XNOR2_X1  g620(.A(new_n801), .B(KEYINPUT47), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n731), .A2(new_n465), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n808), .A2(new_n696), .A3(new_n765), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  XOR2_X1   g624(.A(KEYINPUT112), .B(G140), .Z(new_n811));
  XNOR2_X1  g625(.A(new_n810), .B(new_n811), .ZN(G42));
  NOR2_X1   g626(.A1(new_n786), .A2(new_n397), .ZN(new_n813));
  INV_X1    g627(.A(new_n756), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n814), .A2(new_n465), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  NOR4_X1   g630(.A1(new_n816), .A2(new_n556), .A3(new_n717), .A4(new_n743), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(KEYINPUT50), .ZN(new_n818));
  INV_X1    g632(.A(new_n816), .ZN(new_n819));
  INV_X1    g633(.A(new_n765), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n741), .A2(new_n278), .ZN(new_n821));
  OAI211_X1 g635(.A(new_n819), .B(new_n820), .C1(new_n807), .C2(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n820), .A2(new_n742), .ZN(new_n823));
  OR4_X1    g637(.A1(new_n465), .A2(new_n823), .A3(new_n397), .A4(new_n724), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n824), .A2(new_n394), .A3(new_n784), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n789), .A2(new_n814), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n786), .A2(new_n397), .A3(new_n823), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n825), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n818), .A2(new_n822), .A3(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT51), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n827), .A2(new_n555), .ZN(new_n832));
  XOR2_X1   g646(.A(new_n832), .B(KEYINPUT48), .Z(new_n833));
  NOR2_X1   g647(.A1(new_n712), .A2(new_n655), .ZN(new_n834));
  INV_X1    g648(.A(new_n834), .ZN(new_n835));
  OAI221_X1 g649(.A(new_n395), .B1(new_n824), .B2(new_n835), .C1(new_n750), .C2(new_n816), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n831), .A2(new_n833), .A3(new_n836), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n837), .B1(new_n830), .B2(new_n829), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT54), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n681), .A2(new_n682), .ZN(new_n840));
  AOI22_X1  g654(.A1(new_n459), .A2(new_n461), .B1(new_n840), .B2(new_n463), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT115), .ZN(new_n842));
  INV_X1    g656(.A(new_n698), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n841), .A2(new_n770), .A3(new_n842), .A4(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n271), .A2(new_n766), .ZN(new_n845));
  OAI211_X1 g659(.A(new_n278), .B(new_n843), .C1(new_n845), .C2(new_n740), .ZN(new_n846));
  OAI21_X1  g660(.A(KEYINPUT115), .B1(new_n846), .B2(new_n686), .ZN(new_n847));
  AOI22_X1  g661(.A1(new_n844), .A2(new_n847), .B1(new_n527), .B2(new_n723), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n848), .A2(new_n643), .A3(new_n645), .A4(new_n713), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n762), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n707), .A2(new_n850), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n851), .A2(KEYINPUT52), .A3(new_n736), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT52), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n762), .A2(new_n849), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n854), .B1(new_n706), .B2(new_n702), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n734), .A2(new_n735), .ZN(new_n856));
  INV_X1    g670(.A(new_n730), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n853), .B1(new_n855), .B2(new_n858), .ZN(new_n859));
  OAI21_X1  g673(.A(KEYINPUT116), .B1(new_n852), .B2(new_n859), .ZN(new_n860));
  OAI21_X1  g674(.A(KEYINPUT52), .B1(new_n851), .B2(new_n736), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT116), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n855), .A2(new_n853), .A3(new_n858), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n860), .A2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT113), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n630), .A2(new_n556), .ZN(new_n867));
  INV_X1    g681(.A(new_n656), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n866), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n656), .A2(new_n630), .A3(KEYINPUT113), .A4(new_n556), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n869), .A2(new_n637), .A3(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT114), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n871), .A2(new_n631), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n872), .B1(new_n871), .B2(new_n631), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n637), .A2(new_n751), .A3(new_n319), .ZN(new_n875));
  OAI22_X1  g689(.A1(new_n875), .A2(new_n867), .B1(new_n677), .B2(new_n691), .ZN(new_n876));
  NOR3_X1   g690(.A1(new_n873), .A2(new_n874), .A3(new_n876), .ZN(new_n877));
  AOI211_X1 g691(.A(new_n738), .B(new_n743), .C1(new_n657), .C2(new_n671), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n759), .B1(new_n750), .B2(new_n752), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n318), .A2(new_n393), .A3(new_n843), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n765), .A2(new_n668), .A3(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n881), .A2(new_n690), .A3(new_n729), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n761), .A2(new_n772), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n882), .A2(new_n883), .A3(new_n782), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n878), .A2(new_n879), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n779), .A2(new_n776), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n886), .B1(new_n764), .B2(new_n779), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n877), .A2(new_n885), .A3(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(new_n888), .ZN(new_n889));
  XOR2_X1   g703(.A(KEYINPUT117), .B(KEYINPUT53), .Z(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n865), .A2(new_n889), .A3(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(new_n884), .ZN(new_n893));
  INV_X1    g707(.A(new_n704), .ZN(new_n894));
  OAI211_X1 g708(.A(new_n894), .B(new_n744), .C1(new_n656), .C2(new_n670), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n893), .A2(new_n895), .A3(new_n753), .A4(new_n759), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n780), .A2(new_n896), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n897), .A2(new_n861), .A3(new_n863), .A4(new_n877), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT53), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n839), .B1(new_n892), .B2(new_n900), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n839), .B1(new_n898), .B2(new_n899), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n865), .A2(new_n889), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n902), .B1(new_n903), .B2(new_n890), .ZN(new_n904));
  NOR3_X1   g718(.A1(new_n838), .A2(new_n901), .A3(new_n904), .ZN(new_n905));
  NOR2_X1   g719(.A1(G952), .A2(G953), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n741), .B(KEYINPUT49), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n712), .A2(new_n556), .A3(new_n278), .A4(new_n784), .ZN(new_n908));
  OR4_X1    g722(.A1(new_n465), .A2(new_n907), .A3(new_n724), .A4(new_n908), .ZN(new_n909));
  OAI22_X1  g723(.A1(new_n905), .A2(new_n906), .B1(new_n717), .B2(new_n909), .ZN(G75));
  XOR2_X1   g724(.A(new_n623), .B(new_n599), .Z(new_n911));
  XNOR2_X1  g725(.A(new_n911), .B(KEYINPUT55), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n861), .A2(new_n863), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n913), .A2(new_n888), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(KEYINPUT53), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n888), .B1(new_n860), .B2(new_n864), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n915), .B1(new_n916), .B2(new_n891), .ZN(new_n917));
  INV_X1    g731(.A(new_n917), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n918), .A2(new_n264), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(new_n596), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT56), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n912), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n188), .A2(G952), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n912), .A2(new_n921), .ZN(new_n924));
  INV_X1    g738(.A(new_n629), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n924), .B1(new_n919), .B2(new_n925), .ZN(new_n926));
  NOR3_X1   g740(.A1(new_n922), .A2(new_n923), .A3(new_n926), .ZN(G51));
  NOR3_X1   g741(.A1(new_n918), .A2(new_n264), .A3(new_n797), .ZN(new_n928));
  INV_X1    g742(.A(new_n262), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n891), .B1(new_n865), .B2(new_n889), .ZN(new_n930));
  OAI21_X1  g744(.A(KEYINPUT119), .B1(new_n930), .B2(new_n902), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n917), .A2(KEYINPUT54), .ZN(new_n932));
  AOI21_X1  g746(.A(KEYINPUT54), .B1(new_n914), .B2(KEYINPUT53), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT119), .ZN(new_n934));
  OAI211_X1 g748(.A(new_n933), .B(new_n934), .C1(new_n891), .C2(new_n916), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n931), .A2(new_n932), .A3(new_n935), .ZN(new_n936));
  XNOR2_X1  g750(.A(KEYINPUT118), .B(KEYINPUT57), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n766), .B(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n929), .B1(new_n936), .B2(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n928), .B1(new_n939), .B2(KEYINPUT120), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT120), .ZN(new_n941));
  INV_X1    g755(.A(new_n938), .ZN(new_n942));
  AOI22_X1  g756(.A1(new_n904), .A2(new_n934), .B1(new_n917), .B2(KEYINPUT54), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n942), .B1(new_n943), .B2(new_n931), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n941), .B1(new_n944), .B2(new_n929), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n923), .B1(new_n940), .B2(new_n945), .ZN(G54));
  AND2_X1   g760(.A1(KEYINPUT58), .A2(G475), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n917), .A2(G902), .A3(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(new_n382), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n923), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n950), .B1(new_n949), .B2(new_n948), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n951), .B(KEYINPUT121), .ZN(G60));
  AND2_X1   g766(.A1(new_n649), .A2(new_n650), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n653), .B(KEYINPUT59), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n936), .A2(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(new_n954), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n957), .B1(new_n901), .B2(new_n904), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n958), .A2(new_n953), .ZN(new_n959));
  INV_X1    g773(.A(new_n923), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n956), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(KEYINPUT122), .ZN(new_n962));
  INV_X1    g776(.A(KEYINPUT122), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n956), .A2(new_n959), .A3(new_n963), .A4(new_n960), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n962), .A2(new_n964), .ZN(G63));
  XOR2_X1   g779(.A(new_n456), .B(KEYINPUT124), .Z(new_n966));
  XOR2_X1   g780(.A(new_n966), .B(KEYINPUT60), .Z(new_n967));
  NAND3_X1  g781(.A1(new_n917), .A2(new_n840), .A3(new_n967), .ZN(new_n968));
  AND2_X1   g782(.A1(new_n917), .A2(new_n967), .ZN(new_n969));
  OAI211_X1 g783(.A(new_n960), .B(new_n968), .C1(new_n969), .C2(new_n462), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT123), .ZN(new_n971));
  AND3_X1   g785(.A1(new_n970), .A2(new_n971), .A3(KEYINPUT61), .ZN(new_n972));
  AOI21_X1  g786(.A(KEYINPUT61), .B1(new_n970), .B2(new_n971), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n972), .A2(new_n973), .ZN(G66));
  OAI21_X1  g788(.A(G953), .B1(new_n401), .B2(new_n561), .ZN(new_n975));
  INV_X1    g789(.A(new_n877), .ZN(new_n976));
  NOR3_X1   g790(.A1(new_n976), .A2(new_n878), .A3(new_n879), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n975), .B1(new_n977), .B2(G953), .ZN(new_n978));
  INV_X1    g792(.A(new_n623), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n979), .B1(G898), .B2(new_n188), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n980), .B(KEYINPUT125), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n978), .B(new_n981), .ZN(G69));
  INV_X1    g796(.A(new_n782), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n802), .A2(new_n738), .ZN(new_n984));
  NOR3_X1   g798(.A1(new_n704), .A2(new_n712), .A3(new_n318), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n983), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  AND3_X1   g800(.A1(new_n804), .A2(new_n986), .A3(new_n810), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n858), .A2(new_n707), .A3(new_n762), .ZN(new_n988));
  INV_X1    g802(.A(new_n988), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n987), .A2(new_n887), .A3(new_n989), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n990), .A2(KEYINPUT126), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n536), .A2(new_n511), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n332), .B1(new_n333), .B2(new_n334), .ZN(new_n993));
  XNOR2_X1  g807(.A(new_n992), .B(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT126), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n987), .A2(new_n995), .A3(new_n887), .A4(new_n989), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n991), .A2(new_n994), .A3(new_n996), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n804), .A2(new_n810), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n834), .B1(new_n712), .B2(new_n319), .ZN(new_n999));
  NOR3_X1   g813(.A1(new_n999), .A2(new_n738), .A3(new_n710), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n998), .B1(new_n820), .B2(new_n1000), .ZN(new_n1001));
  OR2_X1    g815(.A1(new_n988), .A2(new_n727), .ZN(new_n1002));
  OR2_X1    g816(.A1(new_n1002), .A2(KEYINPUT62), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1002), .A2(KEYINPUT62), .ZN(new_n1004));
  AND3_X1   g818(.A1(new_n1001), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  OAI211_X1 g819(.A(new_n997), .B(new_n188), .C1(new_n994), .C2(new_n1005), .ZN(new_n1006));
  OR2_X1    g820(.A1(new_n994), .A2(G227), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n994), .A2(G227), .ZN(new_n1008));
  NAND4_X1  g822(.A1(new_n1007), .A2(G900), .A3(G953), .A4(new_n1008), .ZN(new_n1009));
  AND2_X1   g823(.A1(new_n1006), .A2(new_n1009), .ZN(G72));
  NAND3_X1  g824(.A1(new_n991), .A2(new_n977), .A3(new_n996), .ZN(new_n1011));
  NAND2_X1  g825(.A1(G472), .A2(G902), .ZN(new_n1012));
  XOR2_X1   g826(.A(new_n1012), .B(KEYINPUT63), .Z(new_n1013));
  NAND2_X1  g827(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g828(.A1(new_n539), .A2(new_n503), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n892), .A2(new_n900), .ZN(new_n1017));
  NAND3_X1  g831(.A1(new_n538), .A2(new_n541), .A3(new_n513), .ZN(new_n1018));
  NAND3_X1  g832(.A1(new_n1017), .A2(new_n1013), .A3(new_n1018), .ZN(new_n1019));
  NAND4_X1  g833(.A1(new_n1001), .A2(new_n1003), .A3(new_n977), .A4(new_n1004), .ZN(new_n1020));
  AOI21_X1  g834(.A(new_n718), .B1(new_n1020), .B2(new_n1013), .ZN(new_n1021));
  NOR2_X1   g835(.A1(new_n1021), .A2(new_n923), .ZN(new_n1022));
  NAND3_X1  g836(.A1(new_n1016), .A2(new_n1019), .A3(new_n1022), .ZN(new_n1023));
  XNOR2_X1  g837(.A(new_n1023), .B(KEYINPUT127), .ZN(G57));
endmodule


