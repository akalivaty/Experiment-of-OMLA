//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 0 1 0 0 1 1 1 0 1 1 1 0 0 1 0 0 0 1 1 1 1 0 0 0 1 1 1 1 0 1 0 0 0 0 1 0 0 1 0 0 0 0 1 1 1 0 0 0 0 1 0 0 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:30 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n490, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n557, new_n558, new_n559, new_n560, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n571, new_n572, new_n573, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n582, new_n583,
    new_n584, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n613, new_n614, new_n617, new_n619,
    new_n620, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1152, new_n1153, new_n1155;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT64), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  INV_X1    g023(.A(new_n447), .ZN(new_n449));
  NAND2_X1  g024(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n449), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  XOR2_X1   g030(.A(KEYINPUT66), .B(KEYINPUT67), .Z(new_n456));
  XNOR2_X1  g031(.A(new_n455), .B(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n454), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n454), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n457), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  AND2_X1   g038(.A1(KEYINPUT68), .A2(G2105), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT68), .A2(G2105), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  XNOR2_X1  g041(.A(KEYINPUT3), .B(G2104), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n466), .A2(new_n467), .A3(G137), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  AND3_X1   g044(.A1(new_n469), .A2(KEYINPUT70), .A3(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(KEYINPUT70), .B1(new_n469), .B2(G2104), .ZN(new_n471));
  OAI21_X1  g046(.A(G101), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n468), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(KEYINPUT71), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT71), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n468), .A2(new_n472), .A3(new_n475), .ZN(new_n476));
  AND2_X1   g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  NOR2_X1   g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(G125), .ZN(new_n480));
  OAI21_X1  g055(.A(KEYINPUT69), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT69), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n482), .B(G125), .C1(new_n477), .C2(new_n478), .ZN(new_n483));
  NAND2_X1  g058(.A1(G113), .A2(G2104), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n481), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT68), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(new_n469), .ZN(new_n487));
  NAND2_X1  g062(.A1(KEYINPUT68), .A2(G2105), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  AOI22_X1  g064(.A1(new_n474), .A2(new_n476), .B1(new_n485), .B2(new_n489), .ZN(new_n490));
  XOR2_X1   g065(.A(new_n490), .B(KEYINPUT72), .Z(G160));
  NAND2_X1  g066(.A1(new_n489), .A2(new_n467), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n467), .A2(new_n469), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  AOI22_X1  g070(.A1(G124), .A2(new_n493), .B1(new_n495), .B2(G136), .ZN(new_n496));
  OAI221_X1 g071(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n466), .C2(G112), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  XOR2_X1   g073(.A(new_n498), .B(KEYINPUT73), .Z(G162));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n500), .A2(KEYINPUT76), .ZN(new_n501));
  OAI211_X1 g076(.A(new_n487), .B(new_n488), .C1(new_n477), .C2(new_n478), .ZN(new_n502));
  INV_X1    g077(.A(G138), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n501), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n466), .A2(new_n467), .A3(new_n505), .A4(G138), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT75), .ZN(new_n508));
  NAND2_X1  g083(.A1(G126), .A2(G2105), .ZN(new_n509));
  OAI21_X1  g084(.A(G2105), .B1(KEYINPUT74), .B2(G114), .ZN(new_n510));
  AND2_X1   g085(.A1(KEYINPUT74), .A2(G114), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  OAI21_X1  g087(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n513));
  OAI221_X1 g088(.A(new_n508), .B1(new_n479), .B2(new_n509), .C1(new_n512), .C2(new_n513), .ZN(new_n514));
  OAI22_X1  g089(.A1(new_n512), .A2(new_n513), .B1(new_n479), .B2(new_n509), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(KEYINPUT75), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n507), .A2(new_n514), .A3(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(new_n517), .ZN(G164));
  NAND2_X1  g093(.A1(G75), .A2(G543), .ZN(new_n519));
  OR2_X1    g094(.A1(KEYINPUT5), .A2(G543), .ZN(new_n520));
  NAND2_X1  g095(.A1(KEYINPUT5), .A2(G543), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(G62), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n519), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G651), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT6), .ZN(new_n527));
  OAI21_X1  g102(.A(KEYINPUT77), .B1(new_n527), .B2(G651), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT77), .ZN(new_n529));
  INV_X1    g104(.A(G651), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n529), .A2(new_n530), .A3(KEYINPUT6), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  OAI21_X1  g107(.A(KEYINPUT78), .B1(new_n530), .B2(KEYINPUT6), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT78), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n534), .A2(new_n527), .A3(G651), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  NAND4_X1  g111(.A1(new_n532), .A2(new_n536), .A3(G88), .A4(new_n522), .ZN(new_n537));
  NAND4_X1  g112(.A1(new_n532), .A2(new_n536), .A3(G50), .A4(G543), .ZN(new_n538));
  AND3_X1   g113(.A1(new_n537), .A2(new_n538), .A3(KEYINPUT79), .ZN(new_n539));
  AOI21_X1  g114(.A(KEYINPUT79), .B1(new_n537), .B2(new_n538), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n526), .B1(new_n539), .B2(new_n540), .ZN(G303));
  INV_X1    g116(.A(G303), .ZN(G166));
  NAND2_X1  g117(.A1(new_n532), .A2(new_n536), .ZN(new_n543));
  INV_X1    g118(.A(G543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G51), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n543), .A2(new_n523), .ZN(new_n547));
  XOR2_X1   g122(.A(KEYINPUT80), .B(G89), .Z(new_n548));
  NAND2_X1  g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g124(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n550));
  OR2_X1    g125(.A1(new_n550), .A2(KEYINPUT7), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n550), .A2(KEYINPUT7), .ZN(new_n552));
  AND2_X1   g127(.A1(G63), .A2(G651), .ZN(new_n553));
  AOI22_X1  g128(.A1(new_n551), .A2(new_n552), .B1(new_n522), .B2(new_n553), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n546), .A2(new_n549), .A3(new_n554), .ZN(G286));
  INV_X1    g130(.A(G286), .ZN(G168));
  NAND2_X1  g131(.A1(new_n545), .A2(G52), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n547), .A2(G90), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n522), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n559));
  OR2_X1    g134(.A1(new_n559), .A2(new_n530), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n557), .A2(new_n558), .A3(new_n560), .ZN(G301));
  INV_X1    g136(.A(G301), .ZN(G171));
  NAND2_X1  g137(.A1(new_n545), .A2(G43), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n547), .A2(G81), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n522), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n565));
  OR2_X1    g140(.A1(new_n565), .A2(new_n530), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n563), .A2(new_n564), .A3(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G860), .ZN(G153));
  NAND4_X1  g144(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g145(.A1(G1), .A2(G3), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n571), .B(KEYINPUT8), .ZN(new_n572));
  NAND4_X1  g147(.A1(G319), .A2(G483), .A3(G661), .A4(new_n572), .ZN(new_n573));
  XOR2_X1   g148(.A(new_n573), .B(KEYINPUT81), .Z(G188));
  NAND4_X1  g149(.A1(new_n532), .A2(new_n536), .A3(G53), .A4(G543), .ZN(new_n575));
  XNOR2_X1  g150(.A(new_n575), .B(KEYINPUT9), .ZN(new_n576));
  NAND2_X1  g151(.A1(G78), .A2(G543), .ZN(new_n577));
  INV_X1    g152(.A(G65), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n523), .B2(new_n578), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n547), .A2(G91), .B1(new_n579), .B2(G651), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n576), .A2(new_n580), .ZN(G299));
  NAND4_X1  g156(.A1(new_n532), .A2(new_n536), .A3(G49), .A4(G543), .ZN(new_n582));
  NAND4_X1  g157(.A1(new_n532), .A2(new_n536), .A3(G87), .A4(new_n522), .ZN(new_n583));
  OAI21_X1  g158(.A(G651), .B1(new_n522), .B2(G74), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(G288));
  INV_X1    g160(.A(new_n543), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n586), .A2(G48), .A3(G543), .ZN(new_n587));
  NAND4_X1  g162(.A1(new_n532), .A2(new_n536), .A3(G86), .A4(new_n522), .ZN(new_n588));
  INV_X1    g163(.A(G61), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n589), .B1(new_n520), .B2(new_n521), .ZN(new_n590));
  AND2_X1   g165(.A1(G73), .A2(G543), .ZN(new_n591));
  OAI21_X1  g166(.A(G651), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n587), .A2(new_n588), .A3(new_n592), .ZN(G305));
  NAND2_X1  g168(.A1(new_n545), .A2(G47), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n547), .A2(G85), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n522), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n596));
  OAI211_X1 g171(.A(new_n594), .B(new_n595), .C1(new_n530), .C2(new_n596), .ZN(G290));
  NAND2_X1  g172(.A1(G301), .A2(G868), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n547), .A2(G92), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT10), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n547), .A2(KEYINPUT10), .A3(G92), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(G79), .A2(G543), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n604), .B(KEYINPUT82), .ZN(new_n605));
  INV_X1    g180(.A(G66), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n523), .B2(new_n606), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n545), .A2(G54), .B1(new_n607), .B2(G651), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n603), .A2(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n598), .B1(new_n610), .B2(G868), .ZN(G284));
  OAI21_X1  g186(.A(new_n598), .B1(new_n610), .B2(G868), .ZN(G321));
  INV_X1    g187(.A(G868), .ZN(new_n613));
  NAND2_X1  g188(.A1(G299), .A2(new_n613), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n614), .B1(new_n613), .B2(G168), .ZN(G297));
  OAI21_X1  g190(.A(new_n614), .B1(new_n613), .B2(G168), .ZN(G280));
  INV_X1    g191(.A(G559), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n610), .B1(new_n617), .B2(G860), .ZN(G148));
  NAND2_X1  g193(.A1(new_n567), .A2(new_n613), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n609), .A2(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n620), .B2(new_n613), .ZN(G323));
  XNOR2_X1  g196(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OR2_X1    g197(.A1(new_n470), .A2(new_n471), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n623), .A2(new_n467), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(KEYINPUT12), .Z(new_n625));
  XOR2_X1   g200(.A(new_n625), .B(KEYINPUT13), .Z(new_n626));
  XNOR2_X1  g201(.A(KEYINPUT83), .B(G2100), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n628), .B(KEYINPUT84), .Z(new_n629));
  AOI22_X1  g204(.A1(G123), .A2(new_n493), .B1(new_n495), .B2(G135), .ZN(new_n630));
  OAI221_X1 g205(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n466), .C2(G111), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  XOR2_X1   g207(.A(new_n632), .B(G2096), .Z(new_n633));
  OAI211_X1 g208(.A(new_n629), .B(new_n633), .C1(new_n627), .C2(new_n626), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(KEYINPUT85), .Z(G156));
  XNOR2_X1  g210(.A(G2427), .B(G2438), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2430), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT15), .B(G2435), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n637), .A2(new_n638), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n639), .A2(KEYINPUT14), .A3(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2443), .B(G2446), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(G2451), .B(G2454), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT16), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n645), .B(KEYINPUT86), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n643), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G1341), .B(G1348), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT87), .ZN(new_n650));
  OAI211_X1 g225(.A(new_n650), .B(G14), .C1(new_n648), .C2(new_n647), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(G401));
  XOR2_X1   g227(.A(G2072), .B(G2078), .Z(new_n653));
  XOR2_X1   g228(.A(G2084), .B(G2090), .Z(new_n654));
  XNOR2_X1  g229(.A(G2067), .B(G2678), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  AOI21_X1  g231(.A(new_n653), .B1(new_n656), .B2(KEYINPUT18), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT88), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(G2100), .ZN(new_n659));
  INV_X1    g234(.A(KEYINPUT18), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n656), .A2(KEYINPUT17), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n654), .A2(new_n655), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n660), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(G2096), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n659), .B(new_n664), .ZN(G227));
  XOR2_X1   g240(.A(KEYINPUT89), .B(KEYINPUT19), .Z(new_n666));
  XNOR2_X1  g241(.A(G1971), .B(G1976), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1956), .B(G2474), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1961), .B(G1966), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT20), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n669), .A2(new_n670), .ZN(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n668), .A2(new_n675), .ZN(new_n676));
  OR2_X1    g251(.A1(new_n675), .A2(new_n671), .ZN(new_n677));
  OAI211_X1 g252(.A(new_n673), .B(new_n676), .C1(new_n668), .C2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(G1991), .B(G1996), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1981), .B(G1986), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(G229));
  INV_X1    g260(.A(G16), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n686), .A2(G22), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n687), .B1(G166), .B2(new_n686), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(G1971), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n686), .A2(G23), .ZN(new_n690));
  INV_X1    g265(.A(G288), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n690), .B1(new_n691), .B2(new_n686), .ZN(new_n692));
  XOR2_X1   g267(.A(new_n692), .B(KEYINPUT93), .Z(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT33), .B(G1976), .ZN(new_n694));
  AND2_X1   g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  MUX2_X1   g270(.A(G6), .B(G305), .S(G16), .Z(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT32), .B(G1981), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT92), .ZN(new_n698));
  XOR2_X1   g273(.A(new_n696), .B(new_n698), .Z(new_n699));
  NOR2_X1   g274(.A1(new_n693), .A2(new_n694), .ZN(new_n700));
  NOR4_X1   g275(.A1(new_n689), .A2(new_n695), .A3(new_n699), .A4(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(KEYINPUT34), .ZN(new_n702));
  OR2_X1    g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  MUX2_X1   g278(.A(G24), .B(G290), .S(G16), .Z(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(G1986), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  AND2_X1   g281(.A1(new_n706), .A2(KEYINPUT91), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n706), .A2(KEYINPUT91), .ZN(new_n708));
  INV_X1    g283(.A(G29), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G25), .ZN(new_n710));
  AOI22_X1  g285(.A1(G119), .A2(new_n493), .B1(new_n495), .B2(G131), .ZN(new_n711));
  OAI221_X1 g286(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n466), .C2(G107), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n710), .B1(new_n714), .B2(new_n709), .ZN(new_n715));
  XOR2_X1   g290(.A(KEYINPUT35), .B(G1991), .Z(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT90), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n715), .B(new_n717), .ZN(new_n718));
  NOR3_X1   g293(.A1(new_n707), .A2(new_n708), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n701), .A2(new_n702), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n703), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n721), .B(KEYINPUT36), .Z(new_n722));
  NAND2_X1  g297(.A1(new_n623), .A2(G105), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(KEYINPUT96), .Z(new_n724));
  NAND3_X1  g299(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n725), .B(KEYINPUT26), .Z(new_n726));
  INV_X1    g301(.A(G141), .ZN(new_n727));
  INV_X1    g302(.A(G129), .ZN(new_n728));
  OAI221_X1 g303(.A(new_n726), .B1(new_n494), .B2(new_n727), .C1(new_n728), .C2(new_n492), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n724), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n730), .A2(new_n709), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(new_n709), .B2(G32), .ZN(new_n732));
  XNOR2_X1  g307(.A(KEYINPUT27), .B(G1996), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n709), .A2(G33), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT25), .Z(new_n737));
  AOI22_X1  g312(.A1(new_n467), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n738));
  OR2_X1    g313(.A1(new_n738), .A2(new_n466), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n495), .A2(G139), .ZN(new_n740));
  NAND3_X1  g315(.A1(new_n737), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(new_n741), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n735), .B1(new_n742), .B2(new_n709), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n734), .B1(G2072), .B2(new_n743), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n743), .A2(G2072), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(KEYINPUT95), .Z(new_n746));
  NAND2_X1  g321(.A1(new_n732), .A2(new_n733), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n744), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  XNOR2_X1  g323(.A(KEYINPUT31), .B(G11), .ZN(new_n749));
  XNOR2_X1  g324(.A(KEYINPUT97), .B(G28), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n750), .A2(KEYINPUT30), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n750), .A2(KEYINPUT30), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n752), .A2(new_n709), .ZN(new_n753));
  OAI221_X1 g328(.A(new_n749), .B1(new_n751), .B2(new_n753), .C1(new_n632), .C2(new_n709), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n709), .A2(G26), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT28), .Z(new_n756));
  NAND2_X1  g331(.A1(new_n493), .A2(G128), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n495), .A2(G140), .ZN(new_n758));
  OAI21_X1  g333(.A(KEYINPUT94), .B1(G104), .B2(G2105), .ZN(new_n759));
  INV_X1    g334(.A(new_n759), .ZN(new_n760));
  NOR3_X1   g335(.A1(KEYINPUT94), .A2(G104), .A3(G2105), .ZN(new_n761));
  OAI221_X1 g336(.A(G2104), .B1(new_n760), .B2(new_n761), .C1(new_n466), .C2(G116), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n757), .A2(new_n758), .A3(new_n762), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n756), .B1(new_n763), .B2(G29), .ZN(new_n764));
  INV_X1    g339(.A(G2067), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n764), .B(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n686), .A2(G21), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(G168), .B2(new_n686), .ZN(new_n768));
  AOI211_X1 g343(.A(new_n754), .B(new_n766), .C1(G1966), .C2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n686), .A2(G5), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G171), .B2(new_n686), .ZN(new_n771));
  INV_X1    g346(.A(G1961), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n769), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g349(.A(KEYINPUT101), .B(KEYINPUT23), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n686), .A2(G20), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(G299), .B2(G16), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(G1956), .ZN(new_n779));
  NAND2_X1  g354(.A1(G160), .A2(G29), .ZN(new_n780));
  INV_X1    g355(.A(G34), .ZN(new_n781));
  AOI21_X1  g356(.A(G29), .B1(new_n781), .B2(KEYINPUT24), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(KEYINPUT24), .B2(new_n781), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n780), .A2(new_n783), .ZN(new_n784));
  INV_X1    g359(.A(G2084), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n779), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NOR3_X1   g361(.A1(new_n748), .A2(new_n774), .A3(new_n786), .ZN(new_n787));
  NOR2_X1   g362(.A1(G29), .A2(G35), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(G162), .B2(G29), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT29), .ZN(new_n790));
  INV_X1    g365(.A(G2090), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n686), .A2(G19), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(new_n568), .B2(new_n686), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(G1341), .Z(new_n795));
  NOR2_X1   g370(.A1(G4), .A2(G16), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(new_n610), .B2(G16), .ZN(new_n797));
  INV_X1    g372(.A(G1348), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  NAND4_X1  g374(.A1(new_n787), .A2(new_n792), .A3(new_n795), .A4(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n784), .A2(new_n785), .ZN(new_n801));
  XOR2_X1   g376(.A(new_n801), .B(KEYINPUT99), .Z(new_n802));
  NAND2_X1  g377(.A1(new_n709), .A2(G27), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(G164), .B2(new_n709), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT100), .ZN(new_n805));
  INV_X1    g380(.A(G2078), .ZN(new_n806));
  OR2_X1    g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n768), .A2(G1966), .ZN(new_n808));
  XOR2_X1   g383(.A(new_n808), .B(KEYINPUT98), .Z(new_n809));
  NAND2_X1  g384(.A1(new_n805), .A2(new_n806), .ZN(new_n810));
  NAND4_X1  g385(.A1(new_n802), .A2(new_n807), .A3(new_n809), .A4(new_n810), .ZN(new_n811));
  NOR3_X1   g386(.A1(new_n722), .A2(new_n800), .A3(new_n811), .ZN(G311));
  INV_X1    g387(.A(G311), .ZN(G150));
  NAND2_X1  g388(.A1(new_n545), .A2(G55), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n547), .A2(G93), .ZN(new_n815));
  AOI22_X1  g390(.A1(new_n522), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n816));
  OAI211_X1 g391(.A(new_n814), .B(new_n815), .C1(new_n530), .C2(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT102), .ZN(new_n818));
  OR2_X1    g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n817), .A2(new_n818), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n819), .A2(new_n568), .A3(new_n820), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n817), .A2(new_n818), .A3(new_n567), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n823), .B(KEYINPUT38), .Z(new_n824));
  NAND2_X1  g399(.A1(new_n610), .A2(G559), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  AND2_X1   g401(.A1(new_n826), .A2(KEYINPUT39), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n826), .A2(KEYINPUT39), .ZN(new_n828));
  NOR3_X1   g403(.A1(new_n827), .A2(new_n828), .A3(G860), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n817), .A2(G860), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT37), .ZN(new_n831));
  OR2_X1    g406(.A1(new_n829), .A2(new_n831), .ZN(G145));
  AOI22_X1  g407(.A1(G130), .A2(new_n493), .B1(new_n495), .B2(G142), .ZN(new_n833));
  OR3_X1    g408(.A1(new_n466), .A2(KEYINPUT105), .A3(G118), .ZN(new_n834));
  OAI21_X1  g409(.A(KEYINPUT105), .B1(new_n466), .B2(G118), .ZN(new_n835));
  OR2_X1    g410(.A1(G106), .A2(G2105), .ZN(new_n836));
  NAND4_X1  g411(.A1(new_n834), .A2(G2104), .A3(new_n835), .A4(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n833), .A2(new_n837), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(KEYINPUT107), .Z(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(new_n714), .ZN(new_n840));
  INV_X1    g415(.A(new_n840), .ZN(new_n841));
  OR2_X1    g416(.A1(new_n724), .A2(new_n729), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n515), .B1(new_n504), .B2(new_n506), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n763), .B(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(new_n515), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n507), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(new_n763), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(new_n730), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n845), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n850), .A2(new_n742), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT103), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n851), .B(new_n852), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n845), .A2(new_n741), .A3(new_n849), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT104), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n625), .B(KEYINPUT106), .ZN(new_n856));
  NOR3_X1   g431(.A1(new_n853), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(new_n856), .ZN(new_n858));
  INV_X1    g433(.A(new_n855), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n851), .B(KEYINPUT103), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n858), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n841), .B1(new_n857), .B2(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(G160), .B(new_n632), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(G162), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n856), .B1(new_n853), .B2(new_n855), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n859), .A2(new_n860), .A3(new_n858), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n865), .A2(new_n866), .A3(new_n840), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n862), .A2(new_n864), .A3(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT108), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND4_X1  g445(.A1(new_n862), .A2(new_n867), .A3(KEYINPUT108), .A4(new_n864), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n864), .B1(new_n862), .B2(new_n867), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n873), .A2(G37), .ZN(new_n874));
  AND3_X1   g449(.A1(new_n872), .A2(KEYINPUT40), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(KEYINPUT40), .B1(new_n872), .B2(new_n874), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n875), .A2(new_n876), .ZN(G395));
  XNOR2_X1  g452(.A(new_n823), .B(new_n620), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n609), .B(G299), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  XOR2_X1   g456(.A(new_n879), .B(KEYINPUT41), .Z(new_n882));
  AOI21_X1  g457(.A(new_n881), .B1(new_n878), .B2(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(KEYINPUT42), .ZN(new_n884));
  XNOR2_X1  g459(.A(G303), .B(G290), .ZN(new_n885));
  XNOR2_X1  g460(.A(G305), .B(G288), .ZN(new_n886));
  XOR2_X1   g461(.A(new_n885), .B(new_n886), .Z(new_n887));
  AND2_X1   g462(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n884), .A2(new_n887), .ZN(new_n889));
  OAI21_X1  g464(.A(G868), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n817), .A2(new_n613), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(G295));
  NAND2_X1  g467(.A1(new_n890), .A2(new_n891), .ZN(G331));
  INV_X1    g468(.A(KEYINPUT44), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT43), .ZN(new_n895));
  XOR2_X1   g470(.A(G286), .B(G301), .Z(new_n896));
  XNOR2_X1  g471(.A(new_n823), .B(new_n896), .ZN(new_n897));
  OR2_X1    g472(.A1(new_n882), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n880), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n900), .A2(KEYINPUT109), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT109), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n898), .A2(new_n902), .A3(new_n899), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n901), .A2(new_n887), .A3(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n887), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n898), .A2(new_n905), .A3(new_n899), .ZN(new_n906));
  INV_X1    g481(.A(G37), .ZN(new_n907));
  AND2_X1   g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n895), .B1(new_n904), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n900), .A2(new_n887), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n910), .A2(new_n907), .A3(new_n906), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n911), .A2(KEYINPUT43), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n894), .B1(new_n909), .B2(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n894), .B1(new_n911), .B2(KEYINPUT43), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n904), .A2(new_n908), .A3(new_n895), .ZN(new_n915));
  AND3_X1   g490(.A1(new_n914), .A2(KEYINPUT110), .A3(new_n915), .ZN(new_n916));
  AOI21_X1  g491(.A(KEYINPUT110), .B1(new_n914), .B2(new_n915), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n913), .B1(new_n916), .B2(new_n917), .ZN(G397));
  INV_X1    g493(.A(KEYINPUT45), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n919), .A2(G1384), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n847), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n921), .A2(new_n490), .A3(G40), .ZN(new_n922));
  INV_X1    g497(.A(G1384), .ZN(new_n923));
  AOI21_X1  g498(.A(KEYINPUT45), .B1(new_n517), .B2(new_n923), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  XNOR2_X1  g500(.A(KEYINPUT56), .B(G2072), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT3), .ZN(new_n927));
  INV_X1    g502(.A(G2104), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n480), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n484), .B1(new_n931), .B2(new_n482), .ZN(new_n932));
  INV_X1    g507(.A(new_n483), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n489), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n475), .B1(new_n468), .B2(new_n472), .ZN(new_n935));
  AND3_X1   g510(.A1(new_n468), .A2(new_n472), .A3(new_n475), .ZN(new_n936));
  OAI211_X1 g511(.A(new_n934), .B(G40), .C1(new_n935), .C2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT50), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n517), .A2(new_n939), .A3(new_n923), .ZN(new_n940));
  OAI21_X1  g515(.A(KEYINPUT50), .B1(new_n843), .B2(G1384), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n938), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(G1956), .ZN(new_n943));
  AOI22_X1  g518(.A1(new_n925), .A2(new_n926), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT57), .ZN(new_n945));
  AND3_X1   g520(.A1(new_n576), .A2(new_n945), .A3(new_n580), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n945), .B1(new_n576), .B2(new_n580), .ZN(new_n947));
  OAI21_X1  g522(.A(KEYINPUT119), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(G299), .A2(KEYINPUT57), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT119), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n576), .A2(new_n945), .A3(new_n580), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n949), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n948), .A2(new_n952), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n944), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n941), .A2(new_n490), .A3(G40), .ZN(new_n955));
  AND3_X1   g530(.A1(new_n517), .A2(new_n939), .A3(new_n923), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n943), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n517), .A2(new_n923), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(new_n919), .ZN(new_n959));
  INV_X1    g534(.A(new_n920), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n843), .A2(new_n960), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n937), .A2(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n959), .A2(new_n962), .A3(new_n926), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n946), .A2(new_n947), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n957), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  NOR3_X1   g540(.A1(new_n843), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n966), .A2(new_n937), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n958), .A2(KEYINPUT50), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(new_n798), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n847), .A2(new_n923), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n971), .A2(new_n937), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(new_n765), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n609), .B1(new_n970), .B2(new_n973), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n954), .B1(new_n965), .B2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT60), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n609), .A2(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n939), .B1(new_n517), .B2(new_n923), .ZN(new_n978));
  NOR3_X1   g553(.A1(new_n978), .A2(new_n937), .A3(new_n966), .ZN(new_n979));
  OAI211_X1 g554(.A(new_n977), .B(new_n973), .C1(new_n979), .C2(G1348), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n610), .A2(KEYINPUT60), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n970), .A2(KEYINPUT60), .A3(new_n610), .A4(new_n973), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT61), .ZN(new_n985));
  AND3_X1   g560(.A1(new_n957), .A2(new_n964), .A3(new_n963), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n964), .B1(new_n957), .B2(new_n963), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n985), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NOR3_X1   g563(.A1(new_n922), .A2(G1996), .A3(new_n924), .ZN(new_n989));
  XNOR2_X1  g564(.A(KEYINPUT120), .B(KEYINPUT58), .ZN(new_n990));
  XNOR2_X1  g565(.A(new_n990), .B(G1341), .ZN(new_n991));
  INV_X1    g566(.A(new_n991), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n972), .A2(new_n992), .ZN(new_n993));
  OAI211_X1 g568(.A(KEYINPUT122), .B(new_n568), .C1(new_n989), .C2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT59), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  OAI211_X1 g571(.A(KEYINPUT61), .B(new_n965), .C1(new_n944), .C2(new_n953), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n984), .A2(new_n988), .A3(new_n996), .A4(new_n997), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n989), .A2(new_n993), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n999), .A2(new_n567), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT121), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(KEYINPUT59), .ZN(new_n1002));
  AOI22_X1  g577(.A1(new_n1000), .A2(new_n1002), .B1(new_n1001), .B2(new_n994), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n975), .B1(new_n998), .B2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g579(.A(KEYINPUT114), .B1(new_n922), .B2(new_n924), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT114), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n959), .A2(new_n962), .A3(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(G1971), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1005), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n979), .A2(new_n791), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(G303), .A2(G8), .ZN(new_n1012));
  AND2_X1   g587(.A1(KEYINPUT115), .A2(KEYINPUT55), .ZN(new_n1013));
  NOR2_X1   g588(.A1(KEYINPUT115), .A2(KEYINPUT55), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1012), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1015), .B1(new_n1012), .B2(new_n1014), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1011), .A2(G8), .A3(new_n1016), .ZN(new_n1017));
  OAI21_X1  g592(.A(G8), .B1(new_n971), .B2(new_n937), .ZN(new_n1018));
  NAND2_X1  g593(.A1(G305), .A2(G1981), .ZN(new_n1019));
  INV_X1    g594(.A(G1981), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n587), .A2(new_n588), .A3(new_n592), .A4(new_n1020), .ZN(new_n1021));
  AND2_X1   g596(.A1(new_n1021), .A2(KEYINPUT118), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1021), .A2(KEYINPUT118), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1019), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT49), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1018), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  OAI211_X1 g601(.A(new_n1019), .B(KEYINPUT49), .C1(new_n1022), .C2(new_n1023), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1018), .ZN(new_n1028));
  AOI21_X1  g603(.A(KEYINPUT117), .B1(new_n691), .B2(G1976), .ZN(new_n1029));
  XOR2_X1   g604(.A(KEYINPUT116), .B(G1976), .Z(new_n1030));
  NOR2_X1   g605(.A1(new_n691), .A2(new_n1030), .ZN(new_n1031));
  OAI211_X1 g606(.A(new_n1028), .B(new_n1029), .C1(KEYINPUT52), .C2(new_n1031), .ZN(new_n1032));
  OAI211_X1 g607(.A(new_n1029), .B(G8), .C1(new_n937), .C2(new_n971), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT52), .ZN(new_n1034));
  OAI211_X1 g609(.A(new_n1031), .B(G8), .C1(new_n971), .C2(new_n937), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1033), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  AOI22_X1  g611(.A1(new_n1026), .A2(new_n1027), .B1(new_n1032), .B2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1017), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(G8), .ZN(new_n1039));
  OR2_X1    g614(.A1(new_n942), .A2(G2090), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1039), .B1(new_n1009), .B2(new_n1040), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1041), .A2(new_n1016), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1038), .A2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n969), .A2(new_n772), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n919), .B1(new_n843), .B2(G1384), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n517), .A2(new_n920), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n938), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n806), .A2(KEYINPUT53), .ZN(new_n1048));
  OAI211_X1 g623(.A(new_n1044), .B(KEYINPUT123), .C1(new_n1047), .C2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT123), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1051));
  AOI21_X1  g626(.A(G1961), .B1(new_n967), .B2(new_n968), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1050), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1049), .A2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(G2078), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1055));
  OR2_X1    g630(.A1(new_n1055), .A2(KEYINPUT53), .ZN(new_n1056));
  XNOR2_X1  g631(.A(G301), .B(KEYINPUT54), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1054), .A2(new_n1056), .A3(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1057), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT124), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1044), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1052), .A2(KEYINPUT124), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1045), .ZN(new_n1063));
  OR4_X1    g638(.A1(new_n937), .A2(new_n1063), .A3(new_n961), .A4(new_n1048), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1061), .A2(new_n1062), .A3(new_n1064), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1055), .A2(KEYINPUT53), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1059), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(G1966), .ZN(new_n1068));
  AOI22_X1  g643(.A1(new_n979), .A2(new_n785), .B1(new_n1047), .B2(new_n1068), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1069), .A2(G168), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1047), .A2(new_n1068), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n967), .A2(new_n968), .A3(new_n785), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1071), .A2(G168), .A3(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(G8), .ZN(new_n1074));
  OAI21_X1  g649(.A(KEYINPUT51), .B1(new_n1070), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT51), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1073), .A2(new_n1076), .A3(G8), .ZN(new_n1077));
  AOI22_X1  g652(.A1(new_n1058), .A2(new_n1067), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1004), .A2(new_n1043), .A3(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT63), .ZN(new_n1080));
  OAI211_X1 g655(.A(new_n1017), .B(new_n1037), .C1(new_n1041), .C2(new_n1016), .ZN(new_n1081));
  OR3_X1    g656(.A1(new_n1069), .A2(new_n1039), .A3(G286), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1080), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1082), .A2(new_n1080), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1039), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1085));
  OR2_X1    g660(.A1(new_n1085), .A2(new_n1016), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1084), .A2(new_n1086), .A3(new_n1017), .A4(new_n1037), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1083), .A2(new_n1087), .ZN(new_n1088));
  AOI211_X1 g663(.A(G1976), .B(G288), .C1(new_n1026), .C2(new_n1027), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1090));
  OR2_X1    g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1017), .ZN(new_n1092));
  AOI22_X1  g667(.A1(new_n1091), .A2(new_n1028), .B1(new_n1092), .B2(new_n1037), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1079), .A2(new_n1088), .A3(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT125), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1079), .A2(new_n1088), .A3(KEYINPUT125), .A4(new_n1093), .ZN(new_n1097));
  AOI21_X1  g672(.A(G301), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1043), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1075), .A2(new_n1077), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT62), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1075), .A2(KEYINPUT62), .A3(new_n1077), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1099), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1096), .A2(new_n1097), .A3(new_n1105), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1045), .A2(new_n937), .ZN(new_n1107));
  INV_X1    g682(.A(G1996), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1109), .A2(new_n842), .ZN(new_n1110));
  XOR2_X1   g685(.A(new_n1110), .B(KEYINPUT111), .Z(new_n1111));
  INV_X1    g686(.A(KEYINPUT112), .ZN(new_n1112));
  XNOR2_X1  g687(.A(new_n763), .B(new_n765), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1113), .B1(new_n730), .B2(new_n1108), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(new_n1107), .ZN(new_n1115));
  AND3_X1   g690(.A1(new_n1111), .A2(new_n1112), .A3(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1112), .B1(new_n1111), .B2(new_n1115), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  XNOR2_X1  g693(.A(new_n713), .B(new_n716), .ZN(new_n1119));
  OR2_X1    g694(.A1(new_n1119), .A2(KEYINPUT113), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(KEYINPUT113), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1120), .A2(new_n1107), .A3(new_n1121), .ZN(new_n1122));
  AND2_X1   g697(.A1(new_n1118), .A2(new_n1122), .ZN(new_n1123));
  XNOR2_X1  g698(.A(G290), .B(G1986), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(new_n1107), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1106), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT127), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1107), .ZN(new_n1130));
  NOR3_X1   g705(.A1(new_n1130), .A2(G1986), .A3(G290), .ZN(new_n1131));
  XOR2_X1   g706(.A(new_n1131), .B(KEYINPUT48), .Z(new_n1132));
  NAND3_X1  g707(.A1(new_n1118), .A2(new_n1122), .A3(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1130), .B1(new_n730), .B2(new_n1113), .ZN(new_n1134));
  XNOR2_X1  g709(.A(new_n1134), .B(KEYINPUT126), .ZN(new_n1135));
  XNOR2_X1  g710(.A(new_n1109), .B(KEYINPUT46), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  XNOR2_X1  g712(.A(new_n1137), .B(KEYINPUT47), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1133), .A2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1118), .A2(new_n714), .A3(new_n716), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1140), .B1(G2067), .B2(new_n763), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1139), .B1(new_n1141), .B2(new_n1107), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1128), .A2(new_n1129), .A3(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1104), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1126), .B1(new_n1144), .B2(new_n1097), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1141), .A2(new_n1107), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1139), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g723(.A(KEYINPUT127), .B1(new_n1145), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1143), .A2(new_n1149), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g725(.A1(G229), .A2(G401), .A3(new_n462), .A4(G227), .ZN(new_n1152));
  OAI21_X1  g726(.A(new_n1152), .B1(new_n909), .B2(new_n912), .ZN(new_n1153));
  AOI21_X1  g727(.A(new_n1153), .B1(new_n872), .B2(new_n874), .ZN(G308));
  NAND2_X1  g728(.A1(new_n872), .A2(new_n874), .ZN(new_n1155));
  OAI211_X1 g729(.A(new_n1155), .B(new_n1152), .C1(new_n909), .C2(new_n912), .ZN(G225));
endmodule


