//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 1 0 1 0 1 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 0 1 0 0 0 0 1 1 0 0 0 1 1 1 0 1 0 0 0 1 0 1 0 0 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:32 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n753, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n778, new_n779, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n911, new_n912, new_n913,
    new_n914, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960;
  XNOR2_X1  g000(.A(KEYINPUT2), .B(G113), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT68), .ZN(new_n188));
  INV_X1    g002(.A(G116), .ZN(new_n189));
  OAI21_X1  g003(.A(new_n188), .B1(new_n189), .B2(G119), .ZN(new_n190));
  INV_X1    g004(.A(G119), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n191), .A2(KEYINPUT68), .A3(G116), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT69), .B(G116), .ZN(new_n193));
  OAI211_X1 g007(.A(new_n190), .B(new_n192), .C1(new_n193), .C2(new_n191), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT67), .ZN(new_n195));
  AOI21_X1  g009(.A(new_n187), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n189), .A2(KEYINPUT69), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT69), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G116), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n191), .B1(new_n197), .B2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n190), .A2(new_n192), .ZN(new_n201));
  OAI211_X1 g015(.A(new_n195), .B(new_n187), .C1(new_n200), .C2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(new_n202), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n196), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT11), .ZN(new_n205));
  INV_X1    g019(.A(G134), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n205), .B1(new_n206), .B2(G137), .ZN(new_n207));
  INV_X1    g021(.A(G137), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n208), .A2(KEYINPUT11), .A3(G134), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n206), .A2(G137), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n207), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT66), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n207), .A2(new_n209), .A3(KEYINPUT66), .A4(new_n210), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n213), .A2(G131), .A3(new_n214), .ZN(new_n215));
  XOR2_X1   g029(.A(KEYINPUT65), .B(G131), .Z(new_n216));
  NOR2_X1   g030(.A1(new_n211), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(G143), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G146), .ZN(new_n221));
  INV_X1    g035(.A(G146), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G143), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(G128), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g040(.A(KEYINPUT64), .B1(new_n220), .B2(G146), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT64), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n228), .A2(new_n222), .A3(G143), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n227), .A2(new_n229), .A3(new_n221), .ZN(new_n230));
  XOR2_X1   g044(.A(KEYINPUT0), .B(G128), .Z(new_n231));
  AOI22_X1  g045(.A1(new_n226), .A2(KEYINPUT0), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n219), .A2(new_n232), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n206), .A2(G137), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n208), .A2(G134), .ZN(new_n235));
  OAI21_X1  g049(.A(G131), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n236), .B1(new_n211), .B2(new_n216), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT1), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n221), .A2(new_n223), .A3(new_n238), .A4(G128), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n223), .A2(KEYINPUT1), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G128), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(new_n230), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n237), .B1(new_n239), .B2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n204), .B1(new_n233), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n230), .A2(new_n231), .ZN(new_n246));
  NAND4_X1  g060(.A1(new_n221), .A2(new_n223), .A3(KEYINPUT0), .A4(G128), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n248), .B1(new_n215), .B2(new_n218), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n195), .B1(new_n200), .B2(new_n201), .ZN(new_n250));
  INV_X1    g064(.A(new_n187), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(new_n202), .ZN(new_n253));
  NOR3_X1   g067(.A1(new_n249), .A2(new_n253), .A3(new_n243), .ZN(new_n254));
  OAI21_X1  g068(.A(KEYINPUT28), .B1(new_n245), .B2(new_n254), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n233), .A2(new_n244), .A3(new_n204), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT28), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(G953), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(KEYINPUT70), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT70), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G953), .ZN(new_n262));
  AOI21_X1  g076(.A(G237), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G210), .ZN(new_n264));
  XNOR2_X1  g078(.A(new_n264), .B(G101), .ZN(new_n265));
  XNOR2_X1  g079(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n266));
  XNOR2_X1  g080(.A(new_n265), .B(new_n266), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n255), .A2(KEYINPUT29), .A3(new_n258), .A4(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT72), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n242), .A2(new_n239), .ZN(new_n271));
  INV_X1    g085(.A(new_n237), .ZN(new_n272));
  AOI22_X1  g086(.A1(new_n219), .A2(new_n232), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  AOI21_X1  g087(.A(KEYINPUT28), .B1(new_n273), .B2(new_n204), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n253), .B1(new_n249), .B2(new_n243), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n256), .A2(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n274), .B1(new_n276), .B2(KEYINPUT28), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n277), .A2(KEYINPUT72), .A3(KEYINPUT29), .A4(new_n267), .ZN(new_n278));
  INV_X1    g092(.A(G902), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n270), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT73), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND4_X1  g096(.A1(new_n270), .A2(new_n278), .A3(KEYINPUT73), .A4(new_n279), .ZN(new_n283));
  AOI21_X1  g097(.A(KEYINPUT29), .B1(new_n277), .B2(new_n267), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT30), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n233), .A2(new_n244), .A3(new_n285), .ZN(new_n286));
  OAI21_X1  g100(.A(KEYINPUT30), .B1(new_n249), .B2(new_n243), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n254), .B1(new_n288), .B2(new_n253), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n284), .B1(new_n267), .B2(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n282), .A2(new_n283), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(G472), .ZN(new_n292));
  INV_X1    g106(.A(G472), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n285), .B1(new_n233), .B2(new_n244), .ZN(new_n294));
  NOR3_X1   g108(.A1(new_n249), .A2(KEYINPUT30), .A3(new_n243), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n253), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT31), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n296), .A2(new_n297), .A3(new_n256), .A4(new_n267), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(KEYINPUT71), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT71), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n289), .A2(new_n300), .A3(new_n297), .A4(new_n267), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(new_n267), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n257), .B1(new_n256), .B2(new_n275), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n303), .B1(new_n304), .B2(new_n274), .ZN(new_n305));
  AOI22_X1  g119(.A1(new_n305), .A2(new_n297), .B1(new_n289), .B2(new_n267), .ZN(new_n306));
  OAI211_X1 g120(.A(new_n293), .B(new_n279), .C1(new_n302), .C2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT32), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  AND2_X1   g123(.A1(new_n305), .A2(new_n297), .ZN(new_n310));
  INV_X1    g124(.A(new_n289), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n311), .A2(new_n303), .ZN(new_n312));
  OAI211_X1 g126(.A(new_n299), .B(new_n301), .C1(new_n310), .C2(new_n312), .ZN(new_n313));
  NAND4_X1  g127(.A1(new_n313), .A2(KEYINPUT32), .A3(new_n293), .A4(new_n279), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n292), .A2(new_n309), .A3(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT76), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n316), .B1(new_n191), .B2(G128), .ZN(new_n317));
  OR2_X1    g131(.A1(new_n317), .A2(KEYINPUT23), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(KEYINPUT23), .ZN(new_n319));
  OAI211_X1 g133(.A(new_n318), .B(new_n319), .C1(G119), .C2(new_n225), .ZN(new_n320));
  XNOR2_X1  g134(.A(G119), .B(G128), .ZN(new_n321));
  XOR2_X1   g135(.A(KEYINPUT24), .B(G110), .Z(new_n322));
  OAI22_X1  g136(.A1(new_n320), .A2(G110), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  XNOR2_X1  g137(.A(G125), .B(G140), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(new_n222), .ZN(new_n325));
  XNOR2_X1  g139(.A(KEYINPUT77), .B(G125), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT16), .ZN(new_n327));
  INV_X1    g141(.A(G140), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n326), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  NOR2_X1   g143(.A1(G125), .A2(G140), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n330), .B1(new_n326), .B2(G140), .ZN(new_n331));
  OAI211_X1 g145(.A(G146), .B(new_n329), .C1(new_n331), .C2(new_n327), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n323), .A2(new_n325), .A3(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(G125), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(KEYINPUT77), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT77), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(G125), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n335), .A2(new_n337), .A3(G140), .ZN(new_n338));
  INV_X1    g152(.A(new_n330), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n327), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  AND4_X1   g154(.A1(new_n327), .A2(new_n335), .A3(new_n337), .A4(new_n328), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n222), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(new_n332), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n320), .A2(G110), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n322), .A2(new_n321), .ZN(new_n345));
  XNOR2_X1  g159(.A(new_n345), .B(KEYINPUT75), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n343), .A2(new_n344), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n333), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n260), .A2(new_n262), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n349), .A2(G221), .A3(G234), .ZN(new_n350));
  XNOR2_X1  g164(.A(KEYINPUT22), .B(G137), .ZN(new_n351));
  XNOR2_X1  g165(.A(new_n350), .B(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n348), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n333), .A2(new_n347), .A3(new_n352), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n357), .A2(KEYINPUT25), .A3(new_n279), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT25), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n359), .B1(new_n356), .B2(G902), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  XOR2_X1   g175(.A(KEYINPUT74), .B(G217), .Z(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n363), .B1(G234), .B2(new_n279), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n364), .A2(G902), .ZN(new_n365));
  AOI22_X1  g179(.A1(new_n361), .A2(new_n364), .B1(new_n357), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n315), .A2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT78), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  XNOR2_X1  g183(.A(KEYINPUT70), .B(G953), .ZN(new_n370));
  INV_X1    g184(.A(G214), .ZN(new_n371));
  NOR2_X1   g185(.A1(KEYINPUT90), .A2(G143), .ZN(new_n372));
  NOR4_X1   g186(.A1(new_n370), .A2(new_n371), .A3(G237), .A4(new_n372), .ZN(new_n373));
  AND2_X1   g187(.A1(KEYINPUT90), .A2(G143), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n374), .A2(new_n372), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n375), .B1(new_n263), .B2(G214), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n216), .B1(new_n373), .B2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT17), .ZN(new_n378));
  INV_X1    g192(.A(new_n372), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n263), .A2(G214), .A3(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(new_n216), .ZN(new_n381));
  NOR3_X1   g195(.A1(new_n370), .A2(new_n371), .A3(G237), .ZN(new_n382));
  OAI211_X1 g196(.A(new_n380), .B(new_n381), .C1(new_n382), .C2(new_n375), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n377), .A2(new_n378), .A3(new_n383), .ZN(new_n384));
  AND2_X1   g198(.A1(new_n342), .A2(new_n332), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n380), .B1(new_n382), .B2(new_n375), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n386), .A2(KEYINPUT17), .A3(new_n216), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n384), .A2(new_n385), .A3(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT91), .ZN(new_n389));
  NAND2_X1  g203(.A1(KEYINPUT18), .A2(G131), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n389), .B1(new_n386), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n386), .A2(new_n391), .ZN(new_n393));
  INV_X1    g207(.A(new_n331), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n325), .B1(new_n394), .B2(new_n222), .ZN(new_n395));
  INV_X1    g209(.A(new_n376), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n396), .A2(KEYINPUT91), .A3(new_n390), .A4(new_n380), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n392), .A2(new_n393), .A3(new_n395), .A4(new_n397), .ZN(new_n398));
  XNOR2_X1  g212(.A(G113), .B(G122), .ZN(new_n399));
  XNOR2_X1  g213(.A(KEYINPUT93), .B(G104), .ZN(new_n400));
  XNOR2_X1  g214(.A(new_n399), .B(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n388), .A2(new_n398), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(KEYINPUT94), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT94), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n388), .A2(new_n398), .A3(new_n404), .A4(new_n401), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n324), .A2(KEYINPUT19), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n407), .B1(new_n394), .B2(KEYINPUT19), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT92), .ZN(new_n409));
  OR3_X1    g223(.A1(new_n408), .A2(new_n409), .A3(G146), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n377), .A2(new_n383), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n409), .B1(new_n408), .B2(G146), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n410), .A2(new_n332), .A3(new_n411), .A4(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(new_n398), .ZN(new_n414));
  INV_X1    g228(.A(new_n401), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n406), .A2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(G475), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n417), .A2(new_n418), .A3(new_n279), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(KEYINPUT20), .ZN(new_n420));
  AOI21_X1  g234(.A(G475), .B1(new_n406), .B2(new_n416), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT20), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n421), .A2(new_n422), .A3(new_n279), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n420), .A2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(G122), .ZN(new_n425));
  OR3_X1    g239(.A1(new_n193), .A2(KEYINPUT14), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(G116), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT96), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n427), .B(new_n428), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n198), .A2(G116), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n189), .A2(KEYINPUT69), .ZN(new_n431));
  OAI21_X1  g245(.A(G122), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(KEYINPUT14), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n426), .A2(new_n429), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(G107), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(KEYINPUT100), .ZN(new_n436));
  INV_X1    g250(.A(G107), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(KEYINPUT79), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT79), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(G107), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n429), .A2(new_n432), .A3(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT99), .ZN(new_n443));
  XNOR2_X1  g257(.A(new_n442), .B(new_n443), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n220), .A2(G128), .ZN(new_n445));
  XNOR2_X1  g259(.A(new_n445), .B(KEYINPUT98), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n220), .A2(G128), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(new_n206), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n446), .A2(G134), .A3(new_n447), .ZN(new_n450));
  AND2_X1   g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT100), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n434), .A2(new_n452), .A3(G107), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n436), .A2(new_n444), .A3(new_n451), .A4(new_n453), .ZN(new_n454));
  XOR2_X1   g268(.A(KEYINPUT97), .B(KEYINPUT13), .Z(new_n455));
  NAND3_X1  g269(.A1(new_n446), .A2(G134), .A3(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n449), .A2(new_n450), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n429), .A2(new_n432), .ZN(new_n458));
  XNOR2_X1  g272(.A(KEYINPUT79), .B(G107), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(new_n442), .ZN(new_n461));
  OAI211_X1 g275(.A(new_n457), .B(new_n461), .C1(new_n448), .C2(new_n456), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n454), .A2(new_n462), .ZN(new_n463));
  XOR2_X1   g277(.A(KEYINPUT9), .B(G234), .Z(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  NOR3_X1   g279(.A1(new_n363), .A2(new_n465), .A3(G953), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n463), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n454), .A2(new_n466), .A3(new_n462), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(new_n279), .ZN(new_n471));
  INV_X1    g285(.A(G478), .ZN(new_n472));
  NOR2_X1   g286(.A1(KEYINPUT101), .A2(KEYINPUT15), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(KEYINPUT101), .A2(KEYINPUT15), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n472), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n471), .A2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(new_n476), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n470), .A2(new_n279), .A3(new_n478), .ZN(new_n479));
  AND2_X1   g293(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(G952), .ZN(new_n481));
  AOI211_X1 g295(.A(G953), .B(new_n481), .C1(G234), .C2(G237), .ZN(new_n482));
  AOI211_X1 g296(.A(new_n279), .B(new_n349), .C1(G234), .C2(G237), .ZN(new_n483));
  XOR2_X1   g297(.A(KEYINPUT21), .B(G898), .Z(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n482), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n388), .A2(new_n398), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(new_n415), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n406), .A2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT95), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n490), .A2(new_n491), .A3(new_n279), .ZN(new_n492));
  AOI22_X1  g306(.A1(new_n403), .A2(new_n405), .B1(new_n415), .B2(new_n488), .ZN(new_n493));
  OAI21_X1  g307(.A(KEYINPUT95), .B1(new_n493), .B2(G902), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n492), .A2(new_n494), .A3(G475), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n424), .A2(new_n480), .A3(new_n487), .A4(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT102), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n496), .B(new_n497), .ZN(new_n498));
  OAI21_X1  g312(.A(G221), .B1(new_n465), .B2(G902), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  OAI21_X1  g314(.A(G210), .B1(G237), .B2(G902), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(G104), .ZN(new_n503));
  AOI211_X1 g317(.A(KEYINPUT3), .B(new_n503), .C1(new_n438), .C2(new_n440), .ZN(new_n504));
  AOI21_X1  g318(.A(KEYINPUT3), .B1(new_n503), .B2(G107), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n503), .A2(G107), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  OAI21_X1  g321(.A(G101), .B1(new_n504), .B2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT3), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n441), .A2(new_n509), .A3(G104), .ZN(new_n510));
  OR2_X1    g324(.A1(new_n505), .A2(new_n506), .ZN(new_n511));
  INV_X1    g325(.A(G101), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n508), .A2(KEYINPUT4), .A3(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT4), .ZN(new_n515));
  OAI211_X1 g329(.A(new_n515), .B(G101), .C1(new_n504), .C2(new_n507), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n514), .A2(new_n253), .A3(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n438), .A2(new_n440), .A3(new_n503), .ZN(new_n518));
  INV_X1    g332(.A(new_n506), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(KEYINPUT80), .B1(new_n520), .B2(G101), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT80), .ZN(new_n522));
  AOI211_X1 g336(.A(new_n522), .B(new_n512), .C1(new_n518), .C2(new_n519), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  OAI21_X1  g338(.A(G119), .B1(new_n430), .B2(new_n431), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n525), .A2(KEYINPUT5), .A3(new_n190), .A4(new_n192), .ZN(new_n526));
  NOR3_X1   g340(.A1(new_n189), .A2(KEYINPUT5), .A3(G119), .ZN(new_n527));
  INV_X1    g341(.A(G113), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n200), .A2(new_n201), .ZN(new_n530));
  AOI22_X1  g344(.A1(new_n526), .A2(new_n529), .B1(new_n530), .B2(new_n251), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n524), .A2(new_n531), .A3(new_n513), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n517), .A2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT6), .ZN(new_n534));
  XOR2_X1   g348(.A(G110), .B(G122), .Z(new_n535));
  NAND4_X1  g349(.A1(new_n533), .A2(KEYINPUT87), .A3(new_n534), .A4(new_n535), .ZN(new_n536));
  AND2_X1   g350(.A1(new_n242), .A2(new_n239), .ZN(new_n537));
  INV_X1    g351(.A(new_n326), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  OAI21_X1  g353(.A(KEYINPUT88), .B1(new_n232), .B2(new_n538), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT88), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n248), .A2(new_n541), .A3(new_n326), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n539), .A2(new_n540), .A3(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(G224), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n544), .A2(G953), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(new_n545), .ZN(new_n547));
  NAND4_X1  g361(.A1(new_n539), .A2(new_n540), .A3(new_n547), .A4(new_n542), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT87), .ZN(new_n550));
  INV_X1    g364(.A(new_n535), .ZN(new_n551));
  AOI211_X1 g365(.A(new_n550), .B(new_n551), .C1(new_n517), .C2(new_n532), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n517), .A2(new_n532), .A3(new_n551), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(KEYINPUT6), .ZN(new_n554));
  OAI211_X1 g368(.A(new_n536), .B(new_n549), .C1(new_n552), .C2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(new_n279), .ZN(new_n556));
  INV_X1    g370(.A(new_n531), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n506), .B1(new_n459), .B2(new_n503), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n522), .B1(new_n558), .B2(new_n512), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n520), .A2(KEYINPUT80), .A3(G101), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n559), .A2(new_n513), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n557), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(new_n532), .ZN(new_n563));
  XNOR2_X1  g377(.A(new_n535), .B(KEYINPUT8), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT7), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n543), .B1(new_n567), .B2(new_n545), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n566), .A2(new_n568), .A3(new_n553), .ZN(new_n569));
  AND3_X1   g383(.A1(new_n539), .A2(new_n540), .A3(new_n542), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT89), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n570), .A2(new_n571), .A3(KEYINPUT7), .A4(new_n547), .ZN(new_n572));
  OAI21_X1  g386(.A(KEYINPUT89), .B1(new_n548), .B2(new_n567), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n569), .A2(new_n574), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n502), .B1(new_n556), .B2(new_n575), .ZN(new_n576));
  OR2_X1    g390(.A1(new_n569), .A2(new_n574), .ZN(new_n577));
  NAND4_X1  g391(.A1(new_n577), .A2(new_n279), .A3(new_n501), .A4(new_n555), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  OAI21_X1  g393(.A(G214), .B1(G237), .B2(G902), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n271), .A2(KEYINPUT10), .ZN(new_n582));
  OAI21_X1  g396(.A(KEYINPUT81), .B1(new_n561), .B2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT81), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT10), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n585), .B1(new_n242), .B2(new_n239), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n524), .A2(new_n584), .A3(new_n513), .A4(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n514), .A2(new_n516), .A3(new_n232), .ZN(new_n588));
  INV_X1    g402(.A(new_n224), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n225), .B1(new_n223), .B2(KEYINPUT1), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n239), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n559), .A2(new_n591), .A3(new_n513), .A4(new_n560), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(new_n585), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n583), .A2(new_n587), .A3(new_n588), .A4(new_n593), .ZN(new_n594));
  XOR2_X1   g408(.A(new_n219), .B(KEYINPUT82), .Z(new_n595));
  NOR2_X1   g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n594), .A2(new_n219), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT84), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n594), .A2(KEYINPUT84), .A3(new_n219), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n596), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n349), .A2(G227), .ZN(new_n602));
  XNOR2_X1  g416(.A(G110), .B(G140), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n602), .B(new_n603), .ZN(new_n604));
  OAI21_X1  g418(.A(KEYINPUT86), .B1(new_n601), .B2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n596), .ZN(new_n606));
  INV_X1    g420(.A(new_n600), .ZN(new_n607));
  AOI21_X1  g421(.A(KEYINPUT84), .B1(new_n594), .B2(new_n219), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n606), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT86), .ZN(new_n610));
  INV_X1    g424(.A(new_n604), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n561), .A2(new_n537), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(new_n592), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(new_n219), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT12), .ZN(new_n616));
  OAI21_X1  g430(.A(KEYINPUT83), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n615), .A2(new_n616), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT83), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n614), .A2(new_n619), .A3(KEYINPUT12), .A4(new_n219), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n617), .A2(new_n618), .A3(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n621), .A2(new_n606), .A3(new_n604), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n605), .A2(new_n612), .A3(new_n622), .ZN(new_n623));
  XOR2_X1   g437(.A(KEYINPUT85), .B(G469), .Z(new_n624));
  NAND3_X1  g438(.A1(new_n623), .A2(new_n279), .A3(new_n624), .ZN(new_n625));
  AOI211_X1 g439(.A(new_n596), .B(new_n611), .C1(new_n599), .C2(new_n600), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n604), .B1(new_n621), .B2(new_n606), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  OAI21_X1  g442(.A(G469), .B1(new_n628), .B2(G902), .ZN(new_n629));
  AOI211_X1 g443(.A(new_n500), .B(new_n581), .C1(new_n625), .C2(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n315), .A2(KEYINPUT78), .A3(new_n366), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n369), .A2(new_n498), .A3(new_n630), .A4(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(G101), .ZN(G3));
  NAND2_X1  g447(.A1(new_n625), .A2(new_n629), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n279), .B1(new_n302), .B2(new_n306), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(G472), .ZN(new_n636));
  AND2_X1   g450(.A1(new_n636), .A2(new_n307), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n634), .A2(new_n499), .A3(new_n637), .A4(new_n366), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(KEYINPUT103), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n500), .B1(new_n625), .B2(new_n629), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT103), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n640), .A2(new_n641), .A3(new_n366), .A4(new_n637), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n639), .A2(new_n642), .ZN(new_n643));
  AND2_X1   g457(.A1(new_n492), .A2(new_n494), .ZN(new_n644));
  AOI22_X1  g458(.A1(new_n644), .A2(G475), .B1(new_n420), .B2(new_n423), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n468), .A2(KEYINPUT104), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n470), .A2(new_n646), .A3(KEYINPUT33), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT33), .ZN(new_n648));
  OAI211_X1 g462(.A(new_n468), .B(new_n469), .C1(KEYINPUT104), .C2(new_n648), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n647), .A2(G478), .A3(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n470), .A2(new_n472), .A3(new_n279), .ZN(new_n651));
  NAND2_X1  g465(.A1(G478), .A2(G902), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n650), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n645), .A2(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n579), .A2(new_n487), .A3(new_n580), .ZN(new_n656));
  NOR3_X1   g470(.A1(new_n643), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(KEYINPUT34), .B(G104), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G6));
  INV_X1    g473(.A(new_n580), .ZN(new_n660));
  AOI211_X1 g474(.A(new_n486), .B(new_n660), .C1(new_n576), .C2(new_n578), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT105), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n477), .A2(new_n479), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n645), .A2(new_n661), .A3(new_n662), .A4(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n423), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n422), .B1(new_n421), .B2(new_n279), .ZN(new_n666));
  OAI211_X1 g480(.A(new_n495), .B(new_n663), .C1(new_n665), .C2(new_n666), .ZN(new_n667));
  OAI21_X1  g481(.A(KEYINPUT105), .B1(new_n667), .B2(new_n656), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n664), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n639), .A2(new_n642), .A3(new_n669), .ZN(new_n670));
  XOR2_X1   g484(.A(KEYINPUT35), .B(G107), .Z(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G9));
  NAND2_X1  g486(.A1(new_n361), .A2(new_n364), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n353), .A2(KEYINPUT36), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n348), .B(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(new_n365), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n498), .A2(new_n630), .A3(new_n637), .A4(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G110), .ZN(new_n679));
  XNOR2_X1  g493(.A(KEYINPUT106), .B(KEYINPUT37), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(G12));
  INV_X1    g495(.A(new_n677), .ZN(new_n682));
  AND2_X1   g496(.A1(new_n314), .A2(new_n309), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n682), .B1(new_n683), .B2(new_n292), .ZN(new_n684));
  INV_X1    g498(.A(G900), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n482), .B1(new_n483), .B2(new_n685), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n667), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n630), .A2(new_n684), .A3(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G128), .ZN(G30));
  XNOR2_X1  g503(.A(new_n686), .B(KEYINPUT39), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n640), .A2(new_n691), .ZN(new_n692));
  XOR2_X1   g506(.A(KEYINPUT107), .B(KEYINPUT40), .Z(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n579), .B(KEYINPUT38), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n289), .A2(new_n303), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n279), .B1(new_n276), .B2(new_n267), .ZN(new_n697));
  OAI21_X1  g511(.A(G472), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n314), .A2(new_n309), .A3(new_n698), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n480), .B1(new_n424), .B2(new_n495), .ZN(new_n700));
  AND3_X1   g514(.A1(new_n699), .A2(new_n700), .A3(new_n682), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n694), .A2(new_n580), .A3(new_n695), .A4(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G143), .ZN(G45));
  NOR3_X1   g517(.A1(new_n645), .A2(new_n653), .A3(new_n686), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n630), .A2(new_n684), .A3(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G146), .ZN(G48));
  NAND2_X1  g520(.A1(new_n357), .A2(new_n365), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n673), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n708), .B1(new_n683), .B2(new_n292), .ZN(new_n709));
  AND3_X1   g523(.A1(new_n623), .A2(new_n279), .A3(new_n624), .ZN(new_n710));
  INV_X1    g524(.A(G469), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n711), .B1(new_n623), .B2(new_n279), .ZN(new_n712));
  NOR3_X1   g526(.A1(new_n710), .A2(new_n712), .A3(new_n500), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n709), .A2(new_n713), .A3(new_n654), .A4(new_n661), .ZN(new_n714));
  XNOR2_X1  g528(.A(KEYINPUT41), .B(G113), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n714), .B(new_n715), .ZN(G15));
  NAND3_X1  g530(.A1(new_n669), .A2(new_n709), .A3(new_n713), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G116), .ZN(G18));
  NAND2_X1  g532(.A1(new_n623), .A2(new_n279), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(G469), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(new_n625), .ZN(new_n721));
  NOR3_X1   g535(.A1(new_n721), .A2(new_n500), .A3(new_n581), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n722), .A2(new_n498), .A3(new_n684), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G119), .ZN(G21));
  NAND2_X1  g538(.A1(new_n708), .A2(KEYINPUT108), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT108), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n366), .A2(new_n726), .ZN(new_n727));
  AND4_X1   g541(.A1(new_n307), .A2(new_n725), .A3(new_n636), .A4(new_n727), .ZN(new_n728));
  NOR3_X1   g542(.A1(new_n645), .A2(new_n480), .A3(new_n581), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n713), .A2(new_n728), .A3(new_n487), .A4(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G122), .ZN(G24));
  NAND3_X1  g545(.A1(new_n636), .A2(new_n677), .A3(new_n307), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT109), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n636), .A2(new_n677), .A3(KEYINPUT109), .A4(new_n307), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(new_n581), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n736), .A2(new_n713), .A3(new_n737), .A4(new_n704), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G125), .ZN(G27));
  AOI211_X1 g553(.A(new_n500), .B(new_n708), .C1(new_n625), .C2(new_n629), .ZN(new_n740));
  AND2_X1   g554(.A1(new_n740), .A2(new_n315), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n424), .A2(new_n495), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n579), .A2(new_n660), .ZN(new_n743));
  AND3_X1   g557(.A1(new_n650), .A2(new_n651), .A3(new_n652), .ZN(new_n744));
  INV_X1    g558(.A(new_n686), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n742), .A2(new_n743), .A3(new_n744), .A4(new_n745), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n746), .A2(KEYINPUT42), .ZN(new_n747));
  AND4_X1   g561(.A1(new_n742), .A2(new_n743), .A3(new_n744), .A4(new_n745), .ZN(new_n748));
  AND2_X1   g562(.A1(new_n725), .A2(new_n727), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n748), .A2(new_n640), .A3(new_n315), .A4(new_n749), .ZN(new_n750));
  AOI22_X1  g564(.A1(new_n741), .A2(new_n747), .B1(new_n750), .B2(KEYINPUT42), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G131), .ZN(G33));
  NAND4_X1  g566(.A1(new_n740), .A2(new_n315), .A3(new_n687), .A4(new_n743), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G134), .ZN(G36));
  NAND2_X1  g568(.A1(new_n628), .A2(KEYINPUT45), .ZN(new_n755));
  XOR2_X1   g569(.A(new_n755), .B(KEYINPUT110), .Z(new_n756));
  OR2_X1    g570(.A1(new_n628), .A2(KEYINPUT45), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n756), .A2(G469), .A3(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(G469), .A2(G902), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT46), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n758), .A2(KEYINPUT46), .A3(new_n759), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n762), .A2(new_n625), .A3(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n764), .A2(new_n499), .A3(new_n691), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(KEYINPUT111), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT111), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n764), .A2(new_n767), .A3(new_n499), .A4(new_n691), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n743), .B(KEYINPUT112), .ZN(new_n769));
  INV_X1    g583(.A(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n645), .A2(new_n744), .ZN(new_n771));
  XOR2_X1   g585(.A(new_n771), .B(KEYINPUT43), .Z(new_n772));
  INV_X1    g586(.A(new_n637), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n772), .A2(new_n773), .A3(new_n677), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(KEYINPUT44), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n766), .A2(new_n768), .A3(new_n770), .A4(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G137), .ZN(G39));
  NOR2_X1   g591(.A1(new_n315), .A2(new_n366), .ZN(new_n778));
  AND3_X1   g592(.A1(new_n764), .A2(KEYINPUT47), .A3(new_n499), .ZN(new_n779));
  AOI21_X1  g593(.A(KEYINPUT47), .B1(new_n764), .B2(new_n499), .ZN(new_n780));
  OAI211_X1 g594(.A(new_n748), .B(new_n778), .C1(new_n779), .C2(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G140), .ZN(G42));
  OAI211_X1 g596(.A(new_n630), .B(new_n684), .C1(new_n687), .C2(new_n704), .ZN(new_n783));
  AOI211_X1 g597(.A(new_n500), .B(new_n686), .C1(new_n625), .C2(new_n629), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n701), .A2(new_n784), .A3(new_n737), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n783), .A2(new_n738), .A3(new_n785), .ZN(new_n786));
  AND2_X1   g600(.A1(new_n786), .A2(KEYINPUT52), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT52), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n783), .A2(new_n738), .A3(new_n785), .A4(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(new_n751), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n723), .A2(new_n714), .A3(new_n717), .A4(new_n730), .ZN(new_n791));
  NOR3_X1   g605(.A1(new_n787), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n655), .A2(new_n667), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n639), .A2(new_n793), .A3(new_n642), .A4(new_n661), .ZN(new_n794));
  AND3_X1   g608(.A1(new_n794), .A2(new_n632), .A3(new_n678), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT115), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT113), .ZN(new_n797));
  AND4_X1   g611(.A1(new_n640), .A2(new_n315), .A3(new_n366), .A4(new_n687), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n634), .A2(new_n499), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n799), .A2(new_n746), .ZN(new_n800));
  AOI22_X1  g614(.A1(new_n798), .A2(new_n743), .B1(new_n800), .B2(new_n736), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n645), .A2(new_n480), .ZN(new_n802));
  INV_X1    g616(.A(new_n802), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n684), .A2(new_n784), .A3(new_n803), .A4(new_n743), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n797), .B1(new_n801), .B2(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n736), .A2(new_n640), .A3(new_n748), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n804), .A2(new_n753), .A3(new_n806), .A4(new_n797), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  OAI211_X1 g622(.A(new_n795), .B(new_n796), .C1(new_n805), .C2(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n792), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n794), .A2(new_n632), .A3(new_n678), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n804), .A2(new_n753), .A3(new_n806), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n812), .A2(KEYINPUT113), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n811), .B1(new_n813), .B2(new_n807), .ZN(new_n814));
  OAI21_X1  g628(.A(KEYINPUT53), .B1(new_n814), .B2(new_n796), .ZN(new_n815));
  OAI21_X1  g629(.A(KEYINPUT116), .B1(new_n810), .B2(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n717), .A2(new_n714), .A3(new_n730), .ZN(new_n817));
  AND3_X1   g631(.A1(new_n722), .A2(new_n498), .A3(new_n684), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n786), .A2(KEYINPUT52), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n819), .A2(new_n820), .A3(new_n751), .A4(new_n789), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n821), .B1(new_n796), .B2(new_n814), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT53), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n795), .B1(new_n805), .B2(new_n808), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n823), .B1(new_n824), .B2(KEYINPUT115), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT116), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n822), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT54), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n792), .A2(new_n814), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n829), .A2(new_n823), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n816), .A2(new_n827), .A3(new_n828), .A4(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  AOI21_X1  g646(.A(KEYINPUT114), .B1(new_n829), .B2(new_n823), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n829), .A2(new_n823), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n833), .B(new_n834), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n832), .B1(new_n835), .B2(KEYINPUT54), .ZN(new_n836));
  AND3_X1   g650(.A1(new_n713), .A2(new_n482), .A3(new_n743), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n772), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n749), .A2(new_n315), .ZN(new_n839));
  INV_X1    g653(.A(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  XOR2_X1   g655(.A(KEYINPUT119), .B(KEYINPUT48), .Z(new_n842));
  XNOR2_X1  g656(.A(new_n841), .B(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n772), .A2(new_n482), .A3(new_n728), .ZN(new_n844));
  INV_X1    g658(.A(new_n713), .ZN(new_n845));
  NOR3_X1   g659(.A1(new_n844), .A2(new_n581), .A3(new_n845), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n846), .A2(new_n481), .A3(G953), .ZN(new_n847));
  INV_X1    g661(.A(new_n699), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n837), .A2(new_n366), .A3(new_n848), .ZN(new_n849));
  OAI211_X1 g663(.A(new_n843), .B(new_n847), .C1(new_n655), .C2(new_n849), .ZN(new_n850));
  XOR2_X1   g664(.A(new_n850), .B(KEYINPUT120), .Z(new_n851));
  NOR4_X1   g665(.A1(new_n844), .A2(new_n580), .A3(new_n695), .A4(new_n845), .ZN(new_n852));
  XNOR2_X1  g666(.A(new_n852), .B(KEYINPUT50), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n838), .A2(new_n736), .ZN(new_n854));
  OR3_X1    g668(.A1(new_n849), .A2(new_n742), .A3(new_n744), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n853), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT51), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n844), .A2(new_n769), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n779), .A2(new_n780), .ZN(new_n860));
  INV_X1    g674(.A(new_n721), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(new_n500), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n859), .B1(new_n863), .B2(KEYINPUT118), .ZN(new_n864));
  AND2_X1   g678(.A1(new_n863), .A2(KEYINPUT118), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n858), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n836), .A2(new_n851), .A3(new_n866), .ZN(new_n867));
  AND2_X1   g681(.A1(new_n863), .A2(new_n859), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n857), .B1(new_n868), .B2(new_n856), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT117), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n869), .B(new_n870), .ZN(new_n871));
  OAI22_X1  g685(.A1(new_n867), .A2(new_n871), .B1(G952), .B2(G953), .ZN(new_n872));
  XOR2_X1   g686(.A(new_n721), .B(KEYINPUT49), .Z(new_n873));
  NOR4_X1   g687(.A1(new_n771), .A2(new_n695), .A3(new_n500), .A4(new_n660), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n873), .A2(new_n848), .A3(new_n749), .A4(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n872), .A2(new_n875), .ZN(G75));
  OAI21_X1  g690(.A(new_n536), .B1(new_n552), .B2(new_n554), .ZN(new_n877));
  XNOR2_X1  g691(.A(new_n877), .B(new_n549), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n878), .B(KEYINPUT55), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT56), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n879), .B1(KEYINPUT121), .B2(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n816), .A2(new_n827), .A3(new_n830), .ZN(new_n883));
  AND2_X1   g697(.A1(new_n883), .A2(G902), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(G210), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n882), .B1(new_n885), .B2(new_n880), .ZN(new_n886));
  AOI211_X1 g700(.A(KEYINPUT56), .B(new_n881), .C1(new_n884), .C2(G210), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n349), .A2(G952), .ZN(new_n888));
  XOR2_X1   g702(.A(new_n888), .B(KEYINPUT122), .Z(new_n889));
  NOR3_X1   g703(.A1(new_n886), .A2(new_n887), .A3(new_n889), .ZN(G51));
  INV_X1    g704(.A(new_n888), .ZN(new_n891));
  INV_X1    g705(.A(new_n623), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n883), .A2(KEYINPUT54), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n893), .A2(new_n831), .ZN(new_n894));
  XOR2_X1   g708(.A(new_n759), .B(KEYINPUT57), .Z(new_n895));
  AOI21_X1  g709(.A(new_n892), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(new_n758), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n883), .A2(G902), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(KEYINPUT123), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT123), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n883), .A2(new_n900), .A3(G902), .A4(new_n897), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n891), .B1(new_n896), .B2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT124), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  OAI211_X1 g719(.A(KEYINPUT124), .B(new_n891), .C1(new_n896), .C2(new_n902), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(G54));
  NAND3_X1  g721(.A1(new_n884), .A2(KEYINPUT58), .A3(G475), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n908), .B(new_n417), .ZN(new_n909));
  AND2_X1   g723(.A1(new_n909), .A2(new_n891), .ZN(G60));
  AND2_X1   g724(.A1(new_n647), .A2(new_n649), .ZN(new_n911));
  XOR2_X1   g725(.A(new_n652), .B(KEYINPUT59), .Z(new_n912));
  AOI211_X1 g726(.A(new_n911), .B(new_n912), .C1(new_n893), .C2(new_n831), .ZN(new_n913));
  OR2_X1    g727(.A1(new_n836), .A2(new_n912), .ZN(new_n914));
  AOI211_X1 g728(.A(new_n889), .B(new_n913), .C1(new_n914), .C2(new_n911), .ZN(G63));
  INV_X1    g729(.A(new_n889), .ZN(new_n916));
  NAND2_X1  g730(.A1(G217), .A2(G902), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n917), .B(KEYINPUT60), .Z(new_n918));
  NAND3_X1  g732(.A1(new_n883), .A2(new_n675), .A3(new_n918), .ZN(new_n919));
  AND2_X1   g733(.A1(new_n883), .A2(new_n918), .ZN(new_n920));
  OAI211_X1 g734(.A(new_n916), .B(new_n919), .C1(new_n920), .C2(new_n357), .ZN(new_n921));
  XOR2_X1   g735(.A(new_n921), .B(KEYINPUT61), .Z(G66));
  OAI21_X1  g736(.A(G953), .B1(new_n485), .B2(new_n544), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n811), .A2(new_n791), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n923), .B1(new_n924), .B2(new_n370), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n877), .B1(G898), .B2(new_n349), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n925), .B(new_n926), .ZN(G69));
  XNOR2_X1  g741(.A(new_n288), .B(new_n408), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n776), .A2(new_n781), .A3(new_n753), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n766), .A2(new_n729), .A3(new_n840), .A4(new_n768), .ZN(new_n930));
  AND2_X1   g744(.A1(new_n783), .A2(new_n738), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n930), .A2(new_n751), .A3(new_n931), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n349), .B1(new_n929), .B2(new_n932), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n349), .B1(G227), .B2(G900), .ZN(new_n934));
  XNOR2_X1  g748(.A(KEYINPUT125), .B(G900), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n928), .B1(new_n933), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n702), .A2(new_n931), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n938), .B(KEYINPUT62), .Z(new_n939));
  NAND2_X1  g753(.A1(new_n369), .A2(new_n631), .ZN(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(new_n692), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n941), .A2(new_n942), .A3(new_n743), .A4(new_n793), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n939), .A2(new_n776), .A3(new_n781), .A4(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n934), .B1(new_n944), .B2(new_n349), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n937), .B1(new_n928), .B2(new_n945), .ZN(G72));
  INV_X1    g760(.A(new_n924), .ZN(new_n947));
  NOR3_X1   g761(.A1(new_n929), .A2(new_n932), .A3(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT126), .ZN(new_n949));
  NAND2_X1  g763(.A1(G472), .A2(G902), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n950), .B(KEYINPUT63), .Z(new_n951));
  INV_X1    g765(.A(new_n951), .ZN(new_n952));
  OR3_X1    g766(.A1(new_n948), .A2(new_n949), .A3(new_n952), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n311), .A2(new_n267), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n949), .B1(new_n948), .B2(new_n952), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n953), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n951), .B1(new_n944), .B2(new_n947), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n888), .B1(new_n957), .B2(new_n696), .ZN(new_n958));
  NOR3_X1   g772(.A1(new_n954), .A2(new_n696), .A3(new_n952), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n835), .A2(new_n959), .ZN(new_n960));
  AND3_X1   g774(.A1(new_n956), .A2(new_n958), .A3(new_n960), .ZN(G57));
endmodule


