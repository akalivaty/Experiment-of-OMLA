

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803;

  INV_X1 U382 ( .A(n777), .ZN(n362) );
  INV_X1 U383 ( .A(n777), .ZN(n365) );
  AND2_X1 U384 ( .A1(n721), .A2(n437), .ZN(n436) );
  XNOR2_X1 U385 ( .A(n478), .B(KEYINPUT68), .ZN(n740) );
  BUF_X1 U386 ( .A(G116), .Z(n361) );
  XNOR2_X1 U387 ( .A(n783), .B(n466), .ZN(n507) );
  XNOR2_X1 U388 ( .A(n785), .B(n507), .ZN(n509) );
  XNOR2_X2 U389 ( .A(n462), .B(n506), .ZN(n785) );
  NAND2_X1 U390 ( .A1(n739), .A2(n740), .ZN(n490) );
  INV_X4 U391 ( .A(G146), .ZN(n426) );
  AND2_X2 U392 ( .A1(n363), .A2(n362), .ZN(n680) );
  XNOR2_X1 U393 ( .A(n676), .B(n364), .ZN(n363) );
  INV_X1 U394 ( .A(n675), .ZN(n364) );
  AND2_X2 U395 ( .A1(n366), .A2(n365), .ZN(n688) );
  XNOR2_X1 U396 ( .A(n686), .B(n367), .ZN(n366) );
  INV_X1 U397 ( .A(n685), .ZN(n367) );
  NAND2_X1 U398 ( .A1(n368), .A2(n592), .ZN(n595) );
  NAND2_X1 U399 ( .A1(n689), .A2(n387), .ZN(n368) );
  XNOR2_X1 U400 ( .A(G113), .B(G116), .ZN(n491) );
  INV_X2 U401 ( .A(G953), .ZN(n794) );
  NOR2_X2 U402 ( .A1(n698), .A2(n801), .ZN(n387) );
  AND2_X1 U403 ( .A1(n613), .A2(n612), .ZN(n642) );
  INV_X1 U404 ( .A(n710), .ZN(n700) );
  INV_X2 U405 ( .A(G122), .ZN(n465) );
  INV_X2 U406 ( .A(G143), .ZN(n479) );
  AND2_X1 U407 ( .A1(n561), .A2(n560), .ZN(n690) );
  AND2_X1 U408 ( .A1(n391), .A2(n502), .ZN(n584) );
  XNOR2_X1 U409 ( .A(n558), .B(n395), .ZN(n391) );
  XNOR2_X1 U410 ( .A(n563), .B(n404), .ZN(n390) );
  NAND2_X1 U411 ( .A1(n571), .A2(n572), .ZN(n710) );
  XNOR2_X1 U412 ( .A(G119), .B(G128), .ZN(n471) );
  NAND2_X1 U413 ( .A1(n399), .A2(n396), .ZN(n756) );
  XNOR2_X1 U414 ( .A(n406), .B(n538), .ZN(n674) );
  XNOR2_X1 U415 ( .A(n410), .B(n791), .ZN(n774) );
  XNOR2_X1 U416 ( .A(n461), .B(G110), .ZN(n506) );
  INV_X1 U417 ( .A(n491), .ZN(n493) );
  XNOR2_X1 U418 ( .A(KEYINPUT67), .B(G101), .ZN(n494) );
  XNOR2_X2 U419 ( .A(n499), .B(n457), .ZN(n668) );
  NAND2_X1 U420 ( .A1(n430), .A2(n719), .ZN(n369) );
  XNOR2_X1 U421 ( .A(n512), .B(n511), .ZN(n370) );
  NAND2_X1 U422 ( .A1(n430), .A2(n719), .ZN(n666) );
  XNOR2_X1 U423 ( .A(n512), .B(n511), .ZN(n402) );
  XNOR2_X1 U424 ( .A(n412), .B(n411), .ZN(n410) );
  BUF_X1 U425 ( .A(n563), .Z(n371) );
  NOR2_X1 U426 ( .A1(G953), .A2(G237), .ZN(n526) );
  XNOR2_X1 U427 ( .A(n392), .B(KEYINPUT10), .ZN(n535) );
  INV_X1 U428 ( .A(n494), .ZN(n466) );
  NOR2_X1 U429 ( .A1(n418), .A2(n417), .ZN(n416) );
  OR2_X2 U430 ( .A1(n774), .A2(G902), .ZN(n389) );
  XNOR2_X1 U431 ( .A(n548), .B(n463), .ZN(n462) );
  XNOR2_X1 U432 ( .A(n464), .B(KEYINPUT75), .ZN(n463) );
  INV_X1 U433 ( .A(KEYINPUT16), .ZN(n464) );
  XOR2_X1 U434 ( .A(KEYINPUT64), .B(KEYINPUT46), .Z(n628) );
  NAND2_X1 U435 ( .A1(n455), .A2(n454), .ZN(n444) );
  NAND2_X1 U436 ( .A1(n489), .A2(G902), .ZN(n454) );
  XNOR2_X1 U437 ( .A(n392), .B(n425), .ZN(n424) );
  XNOR2_X1 U438 ( .A(KEYINPUT81), .B(KEYINPUT18), .ZN(n425) );
  XNOR2_X1 U439 ( .A(n423), .B(KEYINPUT17), .ZN(n422) );
  XNOR2_X1 U440 ( .A(KEYINPUT70), .B(KEYINPUT4), .ZN(n427) );
  INV_X1 U441 ( .A(KEYINPUT22), .ZN(n395) );
  XNOR2_X1 U442 ( .A(n497), .B(n498), .ZN(n458) );
  XNOR2_X1 U443 ( .A(n535), .B(n414), .ZN(n791) );
  INV_X1 U444 ( .A(n484), .ZN(n414) );
  XNOR2_X1 U445 ( .A(n468), .B(n467), .ZN(n543) );
  INV_X1 U446 ( .A(KEYINPUT8), .ZN(n467) );
  XNOR2_X1 U447 ( .A(n471), .B(n469), .ZN(n413) );
  XNOR2_X1 U448 ( .A(n536), .B(n537), .ZN(n406) );
  XNOR2_X1 U449 ( .A(G104), .B(KEYINPUT92), .ZN(n461) );
  XNOR2_X1 U450 ( .A(n655), .B(n456), .ZN(n428) );
  INV_X1 U451 ( .A(KEYINPUT86), .ZN(n456) );
  NAND2_X1 U452 ( .A1(n398), .A2(n397), .ZN(n396) );
  AND2_X1 U453 ( .A1(n401), .A2(n400), .ZN(n399) );
  NOR2_X1 U454 ( .A1(n725), .A2(n378), .ZN(n397) );
  XNOR2_X1 U455 ( .A(n615), .B(KEYINPUT39), .ZN(n658) );
  NAND2_X1 U456 ( .A1(n705), .A2(n408), .ZN(n649) );
  XNOR2_X1 U457 ( .A(n554), .B(G478), .ZN(n572) );
  NAND2_X1 U458 ( .A1(n452), .A2(n451), .ZN(n450) );
  NAND2_X1 U459 ( .A1(G953), .A2(G902), .ZN(n602) );
  NOR2_X1 U460 ( .A1(G237), .A2(G902), .ZN(n510) );
  OR2_X1 U461 ( .A1(n450), .A2(n448), .ZN(n442) );
  XOR2_X1 U462 ( .A(G134), .B(KEYINPUT7), .Z(n545) );
  XNOR2_X1 U463 ( .A(G113), .B(G143), .ZN(n530) );
  INV_X1 U464 ( .A(G140), .ZN(n529) );
  XNOR2_X1 U465 ( .A(G122), .B(G104), .ZN(n533) );
  XOR2_X1 U466 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n534) );
  XOR2_X1 U467 ( .A(KEYINPUT101), .B(G131), .Z(n528) );
  NAND2_X1 U468 ( .A1(G234), .A2(G237), .ZN(n517) );
  XNOR2_X1 U469 ( .A(n542), .B(n541), .ZN(n570) );
  INV_X1 U470 ( .A(KEYINPUT95), .ZN(n404) );
  AND2_X1 U471 ( .A1(n449), .A2(n448), .ZN(n446) );
  XNOR2_X1 U472 ( .A(n439), .B(n792), .ZN(n796) );
  XNOR2_X1 U473 ( .A(KEYINPUT97), .B(KEYINPUT80), .ZN(n480) );
  XNOR2_X1 U474 ( .A(G107), .B(KEYINPUT96), .ZN(n483) );
  XNOR2_X1 U475 ( .A(n424), .B(n422), .ZN(n403) );
  NAND2_X1 U476 ( .A1(n428), .A2(n802), .ZN(n460) );
  BUF_X1 U477 ( .A(n721), .Z(n757) );
  XOR2_X1 U478 ( .A(KEYINPUT106), .B(n700), .Z(n656) );
  XNOR2_X1 U479 ( .A(n470), .B(n413), .ZN(n412) );
  NAND2_X1 U480 ( .A1(n543), .A2(G221), .ZN(n411) );
  XNOR2_X1 U481 ( .A(n553), .B(n552), .ZN(n771) );
  XNOR2_X1 U482 ( .A(n674), .B(n673), .ZN(n675) );
  NAND2_X1 U483 ( .A1(n756), .A2(n634), .ZN(n627) );
  XNOR2_X1 U484 ( .A(n617), .B(n616), .ZN(n672) );
  OR2_X1 U485 ( .A1(n633), .A2(n394), .ZN(n714) );
  INV_X1 U486 ( .A(KEYINPUT36), .ZN(n407) );
  XNOR2_X1 U487 ( .A(n586), .B(n585), .ZN(n801) );
  XNOR2_X1 U488 ( .A(n565), .B(n564), .ZN(n711) );
  INV_X1 U489 ( .A(n708), .ZN(n705) );
  OR2_X1 U490 ( .A1(n572), .A2(n571), .ZN(n708) );
  XNOR2_X1 U491 ( .A(n379), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U492 ( .A1(n380), .A2(n671), .ZN(n379) );
  XNOR2_X1 U493 ( .A(n669), .B(n372), .ZN(n380) );
  XOR2_X1 U494 ( .A(n668), .B(n667), .Z(n372) );
  XOR2_X1 U495 ( .A(n474), .B(n473), .Z(n373) );
  INV_X1 U496 ( .A(n382), .ZN(n394) );
  XOR2_X1 U497 ( .A(G134), .B(G131), .Z(n374) );
  INV_X1 U498 ( .A(G902), .ZN(n451) );
  AND2_X1 U499 ( .A1(n802), .A2(KEYINPUT2), .ZN(n375) );
  NOR2_X1 U500 ( .A1(n631), .A2(n630), .ZN(n376) );
  AND2_X1 U501 ( .A1(n383), .A2(n566), .ZN(n377) );
  INV_X1 U502 ( .A(KEYINPUT1), .ZN(n448) );
  XOR2_X1 U503 ( .A(KEYINPUT113), .B(KEYINPUT41), .Z(n378) );
  XNOR2_X2 U504 ( .A(n515), .B(KEYINPUT19), .ZN(n635) );
  AND2_X1 U505 ( .A1(n629), .A2(n376), .ZN(n408) );
  XNOR2_X1 U506 ( .A(n507), .B(n458), .ZN(n457) );
  NAND2_X1 U507 ( .A1(n446), .A2(n453), .ZN(n381) );
  NAND2_X1 U508 ( .A1(n446), .A2(n453), .ZN(n445) );
  NAND2_X1 U509 ( .A1(n447), .A2(n381), .ZN(n382) );
  XNOR2_X1 U510 ( .A(n641), .B(KEYINPUT47), .ZN(n417) );
  BUF_X1 U511 ( .A(n740), .Z(n383) );
  NAND2_X1 U512 ( .A1(n447), .A2(n445), .ZN(n739) );
  BUF_X1 U513 ( .A(n684), .Z(n384) );
  XNOR2_X1 U514 ( .A(n509), .B(n508), .ZN(n684) );
  OR2_X2 U515 ( .A1(n623), .A2(n631), .ZN(n611) );
  BUF_X1 U516 ( .A(n623), .Z(n737) );
  NOR2_X2 U517 ( .A1(n402), .A2(n631), .ZN(n515) );
  XNOR2_X2 U518 ( .A(n666), .B(KEYINPUT65), .ZN(n769) );
  XNOR2_X2 U519 ( .A(n369), .B(KEYINPUT65), .ZN(n385) );
  BUF_X1 U520 ( .A(n370), .Z(n386) );
  NAND2_X1 U521 ( .A1(n387), .A2(KEYINPUT44), .ZN(n594) );
  NAND2_X2 U522 ( .A1(n388), .A2(n629), .ZN(n505) );
  AND2_X1 U523 ( .A1(n388), .A2(n562), .ZN(n746) );
  XNOR2_X2 U524 ( .A(n490), .B(KEYINPUT77), .ZN(n388) );
  NOR2_X2 U525 ( .A1(n621), .A2(n477), .ZN(n478) );
  XNOR2_X2 U526 ( .A(n389), .B(n373), .ZN(n621) );
  NAND2_X1 U527 ( .A1(n390), .A2(n721), .ZN(n434) );
  NAND2_X1 U528 ( .A1(n390), .A2(n377), .ZN(n568) );
  NAND2_X1 U529 ( .A1(n436), .A2(n390), .ZN(n435) );
  AND2_X1 U530 ( .A1(n391), .A2(n394), .ZN(n588) );
  XNOR2_X2 U531 ( .A(n426), .B(G125), .ZN(n392) );
  XNOR2_X2 U532 ( .A(n393), .B(n374), .ZN(n439) );
  XNOR2_X1 U533 ( .A(n403), .B(n393), .ZN(n508) );
  XNOR2_X2 U534 ( .A(n551), .B(n427), .ZN(n393) );
  INV_X1 U535 ( .A(n728), .ZN(n398) );
  NAND2_X1 U536 ( .A1(n725), .A2(n378), .ZN(n400) );
  NAND2_X1 U537 ( .A1(n728), .A2(n378), .ZN(n401) );
  XNOR2_X2 U538 ( .A(n415), .B(KEYINPUT112), .ZN(n728) );
  XNOR2_X1 U539 ( .A(n370), .B(n614), .ZN(n723) );
  NOR2_X1 U540 ( .A1(n649), .A2(n386), .ZN(n632) );
  NOR2_X1 U541 ( .A1(n643), .A2(n386), .ZN(n644) );
  AND2_X1 U542 ( .A1(n386), .A2(n652), .ZN(n716) );
  XNOR2_X2 U543 ( .A(n479), .B(G128), .ZN(n551) );
  NAND2_X1 U544 ( .A1(n444), .A2(KEYINPUT1), .ZN(n443) );
  BUF_X1 U545 ( .A(n692), .Z(n405) );
  XNOR2_X1 U546 ( .A(n632), .B(n407), .ZN(n633) );
  XNOR2_X1 U547 ( .A(n438), .B(n555), .ZN(n591) );
  NOR2_X1 U548 ( .A1(n690), .A2(n575), .ZN(n576) );
  NAND2_X1 U549 ( .A1(n692), .A2(n711), .ZN(n574) );
  XNOR2_X2 U550 ( .A(n568), .B(n567), .ZN(n692) );
  NAND2_X1 U551 ( .A1(n409), .A2(n645), .ZN(n438) );
  NAND2_X1 U552 ( .A1(n433), .A2(n435), .ZN(n409) );
  XNOR2_X2 U553 ( .A(n499), .B(n488), .ZN(n765) );
  NAND2_X1 U554 ( .A1(n723), .A2(n722), .ZN(n415) );
  NAND2_X1 U555 ( .A1(n420), .A2(n416), .ZN(n648) );
  NAND2_X1 U556 ( .A1(n714), .A2(n419), .ZN(n418) );
  INV_X1 U557 ( .A(n704), .ZN(n419) );
  XNOR2_X1 U558 ( .A(n421), .B(n628), .ZN(n420) );
  NAND2_X1 U559 ( .A1(n803), .A2(n672), .ZN(n421) );
  XNOR2_X2 U560 ( .A(n627), .B(KEYINPUT42), .ZN(n803) );
  NAND2_X1 U561 ( .A1(n794), .A2(G224), .ZN(n423) );
  AND2_X1 U562 ( .A1(n428), .A2(n375), .ZN(n665) );
  XNOR2_X2 U563 ( .A(n429), .B(KEYINPUT0), .ZN(n563) );
  NOR2_X2 U564 ( .A1(n635), .A2(n524), .ZN(n429) );
  NAND2_X1 U565 ( .A1(n431), .A2(n662), .ZN(n430) );
  NAND2_X1 U566 ( .A1(n432), .A2(n793), .ZN(n431) );
  XNOR2_X2 U567 ( .A(n460), .B(KEYINPUT85), .ZN(n793) );
  XNOR2_X1 U568 ( .A(n459), .B(n600), .ZN(n432) );
  NAND2_X1 U569 ( .A1(n434), .A2(n525), .ZN(n433) );
  INV_X1 U570 ( .A(n525), .ZN(n437) );
  XNOR2_X2 U571 ( .A(n439), .B(n426), .ZN(n499) );
  OR2_X1 U572 ( .A1(n765), .A2(n450), .ZN(n449) );
  INV_X1 U573 ( .A(n444), .ZN(n453) );
  INV_X1 U574 ( .A(n440), .ZN(n447) );
  NAND2_X1 U575 ( .A1(n443), .A2(n441), .ZN(n440) );
  OR2_X1 U576 ( .A1(n765), .A2(n442), .ZN(n441) );
  NAND2_X1 U577 ( .A1(n453), .A2(n449), .ZN(n625) );
  INV_X1 U578 ( .A(n489), .ZN(n452) );
  NAND2_X1 U579 ( .A1(n765), .A2(n489), .ZN(n455) );
  XNOR2_X2 U580 ( .A(KEYINPUT3), .B(G119), .ZN(n492) );
  NAND2_X1 U581 ( .A1(n668), .A2(n451), .ZN(n501) );
  NOR2_X2 U582 ( .A1(n663), .A2(n660), .ZN(n459) );
  XNOR2_X2 U583 ( .A(n465), .B(G107), .ZN(n548) );
  XNOR2_X2 U584 ( .A(n493), .B(n492), .ZN(n783) );
  BUF_X1 U585 ( .A(n591), .Z(n689) );
  BUF_X1 U586 ( .A(n385), .Z(n773) );
  INV_X1 U587 ( .A(G137), .ZN(n495) );
  XNOR2_X1 U588 ( .A(n496), .B(n495), .ZN(n497) );
  INV_X1 U589 ( .A(KEYINPUT48), .ZN(n647) );
  INV_X1 U590 ( .A(KEYINPUT24), .ZN(n469) );
  XNOR2_X1 U591 ( .A(n530), .B(n529), .ZN(n531) );
  AND2_X1 U592 ( .A1(n618), .A2(n734), .ZN(n557) );
  XNOR2_X1 U593 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U594 ( .A(n551), .B(KEYINPUT9), .ZN(n552) );
  INV_X1 U595 ( .A(n777), .ZN(n671) );
  NAND2_X1 U596 ( .A1(G234), .A2(n794), .ZN(n468) );
  XOR2_X1 U597 ( .A(G110), .B(KEYINPUT23), .Z(n470) );
  XNOR2_X1 U598 ( .A(G140), .B(G137), .ZN(n484) );
  XNOR2_X2 U599 ( .A(G902), .B(KEYINPUT15), .ZN(n660) );
  NAND2_X1 U600 ( .A1(G234), .A2(n660), .ZN(n472) );
  XNOR2_X1 U601 ( .A(KEYINPUT20), .B(n472), .ZN(n475) );
  NAND2_X1 U602 ( .A1(n475), .A2(G217), .ZN(n474) );
  XOR2_X1 U603 ( .A(KEYINPUT98), .B(KEYINPUT25), .Z(n473) );
  NAND2_X1 U604 ( .A1(n475), .A2(G221), .ZN(n476) );
  XOR2_X1 U605 ( .A(KEYINPUT21), .B(n476), .Z(n734) );
  INV_X1 U606 ( .A(n734), .ZN(n477) );
  XNOR2_X1 U607 ( .A(n494), .B(n480), .ZN(n481) );
  XNOR2_X1 U608 ( .A(n506), .B(n481), .ZN(n487) );
  NAND2_X1 U609 ( .A1(n794), .A2(G227), .ZN(n482) );
  XNOR2_X1 U610 ( .A(n483), .B(n482), .ZN(n485) );
  XNOR2_X1 U611 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U612 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U613 ( .A(KEYINPUT72), .B(G469), .ZN(n489) );
  XOR2_X1 U614 ( .A(KEYINPUT79), .B(KEYINPUT5), .Z(n496) );
  NAND2_X1 U615 ( .A1(n526), .A2(G210), .ZN(n498) );
  INV_X1 U616 ( .A(G472), .ZN(n500) );
  XNOR2_X2 U617 ( .A(n501), .B(n500), .ZN(n623) );
  XNOR2_X1 U618 ( .A(n623), .B(KEYINPUT6), .ZN(n629) );
  INV_X1 U619 ( .A(n629), .ZN(n502) );
  INV_X1 U620 ( .A(KEYINPUT73), .ZN(n503) );
  XNOR2_X1 U621 ( .A(n503), .B(KEYINPUT33), .ZN(n504) );
  XNOR2_X2 U622 ( .A(n505), .B(n504), .ZN(n721) );
  NAND2_X1 U623 ( .A1(n684), .A2(n660), .ZN(n512) );
  XOR2_X1 U624 ( .A(KEYINPUT78), .B(n510), .Z(n513) );
  NAND2_X1 U625 ( .A1(n513), .A2(G210), .ZN(n511) );
  NAND2_X1 U626 ( .A1(n513), .A2(G214), .ZN(n514) );
  XOR2_X1 U627 ( .A(n514), .B(KEYINPUT93), .Z(n722) );
  INV_X1 U628 ( .A(n722), .ZN(n631) );
  OR2_X1 U629 ( .A1(G898), .A2(n602), .ZN(n516) );
  NAND2_X1 U630 ( .A1(n794), .A2(G952), .ZN(n601) );
  NAND2_X1 U631 ( .A1(n516), .A2(n601), .ZN(n518) );
  XNOR2_X1 U632 ( .A(KEYINPUT14), .B(n517), .ZN(n606) );
  NAND2_X1 U633 ( .A1(n518), .A2(n606), .ZN(n519) );
  NAND2_X1 U634 ( .A1(KEYINPUT94), .A2(n519), .ZN(n523) );
  INV_X1 U635 ( .A(n606), .ZN(n753) );
  NOR2_X1 U636 ( .A1(n753), .A2(n602), .ZN(n521) );
  NOR2_X1 U637 ( .A1(G898), .A2(KEYINPUT94), .ZN(n520) );
  NAND2_X1 U638 ( .A1(n521), .A2(n520), .ZN(n522) );
  NAND2_X1 U639 ( .A1(n523), .A2(n522), .ZN(n524) );
  XOR2_X1 U640 ( .A(KEYINPUT74), .B(KEYINPUT34), .Z(n525) );
  NAND2_X1 U641 ( .A1(G214), .A2(n526), .ZN(n527) );
  XNOR2_X1 U642 ( .A(n528), .B(n527), .ZN(n532) );
  XNOR2_X1 U643 ( .A(n532), .B(n531), .ZN(n538) );
  XNOR2_X1 U644 ( .A(n534), .B(n533), .ZN(n537) );
  INV_X1 U645 ( .A(n535), .ZN(n536) );
  NAND2_X1 U646 ( .A1(n674), .A2(n451), .ZN(n542) );
  XOR2_X1 U647 ( .A(KEYINPUT13), .B(KEYINPUT103), .Z(n540) );
  XNOR2_X1 U648 ( .A(KEYINPUT102), .B(G475), .ZN(n539) );
  XOR2_X1 U649 ( .A(n540), .B(n539), .Z(n541) );
  NAND2_X1 U650 ( .A1(G217), .A2(n543), .ZN(n547) );
  INV_X1 U651 ( .A(KEYINPUT105), .ZN(n544) );
  XNOR2_X1 U652 ( .A(n547), .B(n546), .ZN(n550) );
  XNOR2_X1 U653 ( .A(n548), .B(n361), .ZN(n549) );
  XNOR2_X1 U654 ( .A(n550), .B(n549), .ZN(n553) );
  NAND2_X1 U655 ( .A1(n771), .A2(n451), .ZN(n554) );
  AND2_X1 U656 ( .A1(n570), .A2(n572), .ZN(n645) );
  INV_X1 U657 ( .A(KEYINPUT35), .ZN(n555) );
  INV_X1 U658 ( .A(n591), .ZN(n556) );
  NAND2_X1 U659 ( .A1(n556), .A2(KEYINPUT44), .ZN(n577) );
  NOR2_X1 U660 ( .A1(n570), .A2(n572), .ZN(n618) );
  NAND2_X1 U661 ( .A1(n563), .A2(n557), .ZN(n558) );
  INV_X1 U662 ( .A(KEYINPUT87), .ZN(n559) );
  XNOR2_X1 U663 ( .A(n584), .B(n559), .ZN(n561) );
  BUF_X1 U664 ( .A(n621), .Z(n580) );
  INV_X1 U665 ( .A(n580), .ZN(n735) );
  NOR2_X1 U666 ( .A1(n580), .A2(n382), .ZN(n560) );
  INV_X1 U667 ( .A(n737), .ZN(n562) );
  NAND2_X1 U668 ( .A1(n746), .A2(n371), .ZN(n565) );
  XOR2_X1 U669 ( .A(KEYINPUT31), .B(KEYINPUT100), .Z(n564) );
  AND2_X1 U670 ( .A1(n737), .A2(n625), .ZN(n566) );
  INV_X1 U671 ( .A(KEYINPUT99), .ZN(n567) );
  INV_X1 U672 ( .A(KEYINPUT104), .ZN(n569) );
  XNOR2_X1 U673 ( .A(n570), .B(n569), .ZN(n571) );
  NAND2_X1 U674 ( .A1(n656), .A2(n708), .ZN(n573) );
  XNOR2_X1 U675 ( .A(n573), .B(KEYINPUT107), .ZN(n727) );
  INV_X1 U676 ( .A(n727), .ZN(n639) );
  AND2_X1 U677 ( .A1(n574), .A2(n639), .ZN(n575) );
  NAND2_X1 U678 ( .A1(n577), .A2(n576), .ZN(n579) );
  INV_X1 U679 ( .A(KEYINPUT88), .ZN(n578) );
  XNOR2_X1 U680 ( .A(n579), .B(n578), .ZN(n597) );
  NAND2_X1 U681 ( .A1(n580), .A2(n382), .ZN(n582) );
  INV_X1 U682 ( .A(KEYINPUT108), .ZN(n581) );
  XNOR2_X1 U683 ( .A(n582), .B(n581), .ZN(n583) );
  NAND2_X1 U684 ( .A1(n584), .A2(n583), .ZN(n586) );
  INV_X1 U685 ( .A(KEYINPUT32), .ZN(n585) );
  INV_X1 U686 ( .A(KEYINPUT109), .ZN(n587) );
  XNOR2_X1 U687 ( .A(n588), .B(n587), .ZN(n590) );
  AND2_X1 U688 ( .A1(n580), .A2(n737), .ZN(n589) );
  AND2_X1 U689 ( .A1(n590), .A2(n589), .ZN(n698) );
  INV_X1 U690 ( .A(KEYINPUT44), .ZN(n592) );
  NAND2_X1 U691 ( .A1(n595), .A2(n594), .ZN(n596) );
  NAND2_X1 U692 ( .A1(n597), .A2(n596), .ZN(n599) );
  INV_X1 U693 ( .A(KEYINPUT45), .ZN(n598) );
  XNOR2_X1 U694 ( .A(n599), .B(n598), .ZN(n663) );
  INV_X1 U695 ( .A(KEYINPUT83), .ZN(n600) );
  INV_X1 U696 ( .A(n601), .ZN(n604) );
  NOR2_X1 U697 ( .A1(G900), .A2(n602), .ZN(n603) );
  OR2_X1 U698 ( .A1(n604), .A2(n603), .ZN(n605) );
  NAND2_X1 U699 ( .A1(n606), .A2(n605), .ZN(n608) );
  INV_X1 U700 ( .A(KEYINPUT82), .ZN(n607) );
  XNOR2_X1 U701 ( .A(n608), .B(n607), .ZN(n619) );
  AND2_X1 U702 ( .A1(n625), .A2(n619), .ZN(n609) );
  AND2_X1 U703 ( .A1(n740), .A2(n609), .ZN(n613) );
  INV_X1 U704 ( .A(KEYINPUT30), .ZN(n610) );
  XNOR2_X1 U705 ( .A(n611), .B(n610), .ZN(n612) );
  XNOR2_X1 U706 ( .A(KEYINPUT76), .B(KEYINPUT38), .ZN(n614) );
  NAND2_X1 U707 ( .A1(n642), .A2(n723), .ZN(n615) );
  NAND2_X1 U708 ( .A1(n658), .A2(n705), .ZN(n617) );
  XOR2_X1 U709 ( .A(KEYINPUT111), .B(KEYINPUT40), .Z(n616) );
  INV_X1 U710 ( .A(n618), .ZN(n725) );
  NAND2_X1 U711 ( .A1(n619), .A2(n734), .ZN(n620) );
  XNOR2_X1 U712 ( .A(n620), .B(KEYINPUT71), .ZN(n622) );
  NAND2_X1 U713 ( .A1(n622), .A2(n621), .ZN(n630) );
  NOR2_X1 U714 ( .A1(n623), .A2(n630), .ZN(n624) );
  XNOR2_X1 U715 ( .A(n624), .B(KEYINPUT28), .ZN(n626) );
  AND2_X1 U716 ( .A1(n626), .A2(n625), .ZN(n634) );
  INV_X1 U717 ( .A(n634), .ZN(n637) );
  BUF_X1 U718 ( .A(n635), .Z(n636) );
  NOR2_X1 U719 ( .A1(n637), .A2(n636), .ZN(n706) );
  INV_X1 U720 ( .A(KEYINPUT69), .ZN(n638) );
  AND2_X1 U721 ( .A1(n706), .A2(n638), .ZN(n640) );
  NAND2_X1 U722 ( .A1(n640), .A2(n639), .ZN(n641) );
  INV_X1 U723 ( .A(n642), .ZN(n643) );
  XNOR2_X1 U724 ( .A(n644), .B(KEYINPUT110), .ZN(n646) );
  AND2_X1 U725 ( .A1(n646), .A2(n645), .ZN(n704) );
  XNOR2_X1 U726 ( .A(n648), .B(n647), .ZN(n654) );
  NOR2_X1 U727 ( .A1(n649), .A2(n382), .ZN(n651) );
  INV_X1 U728 ( .A(KEYINPUT43), .ZN(n650) );
  XNOR2_X1 U729 ( .A(n651), .B(n650), .ZN(n652) );
  INV_X1 U730 ( .A(n716), .ZN(n653) );
  NAND2_X1 U731 ( .A1(n654), .A2(n653), .ZN(n655) );
  INV_X1 U732 ( .A(n656), .ZN(n657) );
  NAND2_X1 U733 ( .A1(n658), .A2(n657), .ZN(n659) );
  XNOR2_X1 U734 ( .A(n659), .B(KEYINPUT114), .ZN(n802) );
  XOR2_X1 U735 ( .A(KEYINPUT84), .B(n660), .Z(n661) );
  NAND2_X1 U736 ( .A1(n661), .A2(KEYINPUT2), .ZN(n662) );
  BUF_X1 U737 ( .A(n663), .Z(n664) );
  INV_X1 U738 ( .A(n664), .ZN(n778) );
  NAND2_X1 U739 ( .A1(n778), .A2(n665), .ZN(n719) );
  NAND2_X1 U740 ( .A1(n385), .A2(G472), .ZN(n669) );
  XNOR2_X1 U741 ( .A(KEYINPUT115), .B(KEYINPUT62), .ZN(n667) );
  INV_X1 U742 ( .A(G952), .ZN(n670) );
  AND2_X1 U743 ( .A1(n670), .A2(G953), .ZN(n777) );
  XNOR2_X1 U744 ( .A(n672), .B(G131), .ZN(G33) );
  NAND2_X1 U745 ( .A1(n769), .A2(G475), .ZN(n676) );
  XOR2_X1 U746 ( .A(KEYINPUT91), .B(KEYINPUT59), .Z(n673) );
  XNOR2_X1 U747 ( .A(KEYINPUT126), .B(KEYINPUT60), .ZN(n678) );
  XNOR2_X1 U748 ( .A(n678), .B(KEYINPUT66), .ZN(n679) );
  XNOR2_X1 U749 ( .A(n680), .B(n679), .ZN(G60) );
  NAND2_X1 U750 ( .A1(n769), .A2(G210), .ZN(n686) );
  XOR2_X1 U751 ( .A(KEYINPUT89), .B(KEYINPUT90), .Z(n682) );
  XNOR2_X1 U752 ( .A(KEYINPUT55), .B(KEYINPUT54), .ZN(n681) );
  XNOR2_X1 U753 ( .A(n682), .B(n681), .ZN(n683) );
  XNOR2_X1 U754 ( .A(n384), .B(n683), .ZN(n685) );
  XNOR2_X1 U755 ( .A(n688), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U756 ( .A(n689), .B(G122), .ZN(G24) );
  XOR2_X1 U757 ( .A(G101), .B(n690), .Z(G3) );
  NOR2_X1 U758 ( .A1(n708), .A2(n405), .ZN(n691) );
  XOR2_X1 U759 ( .A(G104), .B(n691), .Z(G6) );
  NOR2_X1 U760 ( .A1(n710), .A2(n405), .ZN(n697) );
  XOR2_X1 U761 ( .A(KEYINPUT27), .B(KEYINPUT117), .Z(n694) );
  XNOR2_X1 U762 ( .A(G107), .B(KEYINPUT116), .ZN(n693) );
  XNOR2_X1 U763 ( .A(n694), .B(n693), .ZN(n695) );
  XNOR2_X1 U764 ( .A(KEYINPUT26), .B(n695), .ZN(n696) );
  XNOR2_X1 U765 ( .A(n697), .B(n696), .ZN(G9) );
  XOR2_X1 U766 ( .A(G110), .B(n698), .Z(n699) );
  XNOR2_X1 U767 ( .A(KEYINPUT118), .B(n699), .ZN(G12) );
  XOR2_X1 U768 ( .A(KEYINPUT119), .B(KEYINPUT29), .Z(n702) );
  NAND2_X1 U769 ( .A1(n706), .A2(n700), .ZN(n701) );
  XNOR2_X1 U770 ( .A(n702), .B(n701), .ZN(n703) );
  XOR2_X1 U771 ( .A(G128), .B(n703), .Z(G30) );
  XOR2_X1 U772 ( .A(G143), .B(n704), .Z(G45) );
  NAND2_X1 U773 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U774 ( .A(n707), .B(G146), .ZN(G48) );
  NOR2_X1 U775 ( .A1(n711), .A2(n708), .ZN(n709) );
  XOR2_X1 U776 ( .A(G113), .B(n709), .Z(G15) );
  NOR2_X1 U777 ( .A1(n711), .A2(n710), .ZN(n712) );
  XOR2_X1 U778 ( .A(KEYINPUT120), .B(n712), .Z(n713) );
  XNOR2_X1 U779 ( .A(n361), .B(n713), .ZN(G18) );
  XOR2_X1 U780 ( .A(n714), .B(G125), .Z(n715) );
  XNOR2_X1 U781 ( .A(n715), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U782 ( .A(G140), .B(n716), .Z(G42) );
  NAND2_X1 U783 ( .A1(n793), .A2(n778), .ZN(n718) );
  INV_X1 U784 ( .A(KEYINPUT2), .ZN(n717) );
  NAND2_X1 U785 ( .A1(n718), .A2(n717), .ZN(n720) );
  NAND2_X1 U786 ( .A1(n720), .A2(n719), .ZN(n761) );
  NOR2_X1 U787 ( .A1(n723), .A2(n722), .ZN(n724) );
  NOR2_X1 U788 ( .A1(n725), .A2(n724), .ZN(n726) );
  XOR2_X1 U789 ( .A(KEYINPUT122), .B(n726), .Z(n731) );
  NOR2_X1 U790 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U791 ( .A(KEYINPUT123), .B(n729), .ZN(n730) );
  NAND2_X1 U792 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U793 ( .A1(n757), .A2(n732), .ZN(n733) );
  XNOR2_X1 U794 ( .A(n733), .B(KEYINPUT124), .ZN(n750) );
  NOR2_X1 U795 ( .A1(n735), .A2(n734), .ZN(n736) );
  XNOR2_X1 U796 ( .A(n736), .B(KEYINPUT49), .ZN(n738) );
  NAND2_X1 U797 ( .A1(n738), .A2(n737), .ZN(n744) );
  NOR2_X1 U798 ( .A1(n383), .A2(n382), .ZN(n741) );
  XOR2_X1 U799 ( .A(KEYINPUT121), .B(n741), .Z(n742) );
  XNOR2_X1 U800 ( .A(n742), .B(KEYINPUT50), .ZN(n743) );
  NOR2_X1 U801 ( .A1(n744), .A2(n743), .ZN(n745) );
  NOR2_X1 U802 ( .A1(n746), .A2(n745), .ZN(n747) );
  XNOR2_X1 U803 ( .A(KEYINPUT51), .B(n747), .ZN(n748) );
  NAND2_X1 U804 ( .A1(n748), .A2(n756), .ZN(n749) );
  NAND2_X1 U805 ( .A1(n750), .A2(n749), .ZN(n751) );
  XOR2_X1 U806 ( .A(KEYINPUT52), .B(n751), .Z(n752) );
  NOR2_X1 U807 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U808 ( .A1(n754), .A2(G952), .ZN(n755) );
  NAND2_X1 U809 ( .A1(n755), .A2(n794), .ZN(n759) );
  AND2_X1 U810 ( .A1(n757), .A2(n756), .ZN(n758) );
  NOR2_X1 U811 ( .A1(n759), .A2(n758), .ZN(n760) );
  NAND2_X1 U812 ( .A1(n761), .A2(n760), .ZN(n762) );
  XOR2_X1 U813 ( .A(KEYINPUT53), .B(n762), .Z(G75) );
  NAND2_X1 U814 ( .A1(n773), .A2(G469), .ZN(n767) );
  XOR2_X1 U815 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n763) );
  XOR2_X1 U816 ( .A(n763), .B(KEYINPUT125), .Z(n764) );
  XNOR2_X1 U817 ( .A(n765), .B(n764), .ZN(n766) );
  XNOR2_X1 U818 ( .A(n767), .B(n766), .ZN(n768) );
  NOR2_X1 U819 ( .A1(n777), .A2(n768), .ZN(G54) );
  NAND2_X1 U820 ( .A1(n385), .A2(G478), .ZN(n770) );
  XOR2_X1 U821 ( .A(n771), .B(n770), .Z(n772) );
  NOR2_X1 U822 ( .A1(n777), .A2(n772), .ZN(G63) );
  NAND2_X1 U823 ( .A1(n773), .A2(G217), .ZN(n775) );
  XNOR2_X1 U824 ( .A(n774), .B(n775), .ZN(n776) );
  NOR2_X1 U825 ( .A1(n777), .A2(n776), .ZN(G66) );
  NAND2_X1 U826 ( .A1(n778), .A2(n794), .ZN(n782) );
  NAND2_X1 U827 ( .A1(G953), .A2(G224), .ZN(n779) );
  XNOR2_X1 U828 ( .A(KEYINPUT61), .B(n779), .ZN(n780) );
  NAND2_X1 U829 ( .A1(n780), .A2(G898), .ZN(n781) );
  NAND2_X1 U830 ( .A1(n782), .A2(n781), .ZN(n790) );
  OR2_X1 U831 ( .A1(G898), .A2(n794), .ZN(n787) );
  XOR2_X1 U832 ( .A(n783), .B(G101), .Z(n784) );
  XNOR2_X1 U833 ( .A(n785), .B(n784), .ZN(n786) );
  NAND2_X1 U834 ( .A1(n787), .A2(n786), .ZN(n788) );
  XNOR2_X1 U835 ( .A(n788), .B(KEYINPUT127), .ZN(n789) );
  XNOR2_X1 U836 ( .A(n790), .B(n789), .ZN(G69) );
  XNOR2_X1 U837 ( .A(n791), .B(KEYINPUT96), .ZN(n792) );
  XNOR2_X1 U838 ( .A(n793), .B(n796), .ZN(n795) );
  NAND2_X1 U839 ( .A1(n795), .A2(n794), .ZN(n800) );
  XOR2_X1 U840 ( .A(G227), .B(n796), .Z(n797) );
  NAND2_X1 U841 ( .A1(n797), .A2(G900), .ZN(n798) );
  NAND2_X1 U842 ( .A1(n798), .A2(G953), .ZN(n799) );
  NAND2_X1 U843 ( .A1(n800), .A2(n799), .ZN(G72) );
  XOR2_X1 U844 ( .A(G119), .B(n801), .Z(G21) );
  XNOR2_X1 U845 ( .A(G134), .B(n802), .ZN(G36) );
  XNOR2_X1 U846 ( .A(n803), .B(G137), .ZN(G39) );
endmodule

