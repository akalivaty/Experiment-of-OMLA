//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 0 1 1 1 1 1 1 1 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 0 1 0 1 1 0 0 0 0 1 0 0 1 0 1 0 1 0 0 1 0 1 1 0 0 1 0 1 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n718, new_n719, new_n720,
    new_n721, new_n723, new_n724, new_n725, new_n727, new_n728, new_n729,
    new_n731, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n855, new_n856,
    new_n857, new_n858, new_n860, new_n861, new_n862, new_n863, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n904, new_n905, new_n907, new_n908, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n924, new_n925, new_n926, new_n928,
    new_n929, new_n930, new_n931, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n947, new_n948, new_n949, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962;
  XNOR2_X1  g000(.A(G197gat), .B(G204gat), .ZN(new_n202));
  INV_X1    g001(.A(G211gat), .ZN(new_n203));
  INV_X1    g002(.A(G218gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n202), .B1(KEYINPUT22), .B2(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(G211gat), .B(G218gat), .ZN(new_n207));
  XNOR2_X1  g006(.A(new_n206), .B(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(G226gat), .A2(G233gat), .ZN(new_n210));
  XOR2_X1   g009(.A(new_n210), .B(KEYINPUT75), .Z(new_n211));
  INV_X1    g010(.A(KEYINPUT64), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT24), .ZN(new_n213));
  INV_X1    g012(.A(G183gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(G190gat), .ZN(new_n215));
  INV_X1    g014(.A(G190gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(G183gat), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n213), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n213), .A2(G183gat), .A3(G190gat), .ZN(new_n219));
  INV_X1    g018(.A(new_n219), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n212), .B1(new_n218), .B2(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(G183gat), .B(G190gat), .ZN(new_n222));
  OAI211_X1 g021(.A(KEYINPUT64), .B(new_n219), .C1(new_n222), .C2(new_n213), .ZN(new_n223));
  INV_X1    g022(.A(G169gat), .ZN(new_n224));
  INV_X1    g023(.A(G176gat), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n224), .A2(new_n225), .A3(KEYINPUT23), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT23), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n227), .B1(G169gat), .B2(G176gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(G169gat), .A2(G176gat), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n226), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n221), .A2(new_n223), .A3(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT65), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT25), .ZN(new_n234));
  AND3_X1   g033(.A1(new_n232), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n233), .B1(new_n232), .B2(new_n234), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n219), .B1(new_n222), .B2(new_n213), .ZN(new_n237));
  NOR3_X1   g036(.A1(new_n237), .A2(new_n230), .A3(new_n234), .ZN(new_n238));
  NOR3_X1   g037(.A1(new_n235), .A2(new_n236), .A3(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(KEYINPUT27), .B(G183gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(new_n216), .ZN(new_n241));
  XOR2_X1   g040(.A(KEYINPUT66), .B(KEYINPUT28), .Z(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(G183gat), .A2(G190gat), .ZN(new_n244));
  NOR2_X1   g043(.A1(KEYINPUT66), .A2(KEYINPUT28), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n240), .A2(new_n216), .A3(new_n245), .ZN(new_n246));
  OR3_X1    g045(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n247));
  OAI21_X1  g046(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n247), .A2(new_n248), .A3(new_n229), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n243), .A2(new_n244), .A3(new_n246), .A4(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n211), .B1(new_n239), .B2(new_n251), .ZN(new_n252));
  OAI21_X1  g051(.A(KEYINPUT76), .B1(new_n239), .B2(new_n251), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n232), .A2(new_n234), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n238), .B1(new_n254), .B2(KEYINPUT65), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n232), .A2(new_n233), .A3(new_n234), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n251), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT76), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  AOI21_X1  g058(.A(KEYINPUT29), .B1(new_n253), .B2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(new_n210), .ZN(new_n261));
  OAI211_X1 g060(.A(new_n209), .B(new_n252), .C1(new_n260), .C2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT77), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(G8gat), .B(G36gat), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n265), .B(G64gat), .ZN(new_n266));
  INV_X1    g065(.A(G92gat), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n266), .B(new_n267), .ZN(new_n268));
  AOI211_X1 g067(.A(KEYINPUT76), .B(new_n251), .C1(new_n255), .C2(new_n256), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n254), .A2(KEYINPUT65), .ZN(new_n270));
  INV_X1    g069(.A(new_n238), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n270), .A2(new_n256), .A3(new_n271), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n258), .B1(new_n272), .B2(new_n250), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n261), .B1(new_n269), .B2(new_n273), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n257), .A2(KEYINPUT29), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n274), .B1(new_n211), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(new_n208), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT29), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n278), .B1(new_n269), .B2(new_n273), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(new_n210), .ZN(new_n280));
  NAND4_X1  g079(.A1(new_n280), .A2(KEYINPUT77), .A3(new_n209), .A4(new_n252), .ZN(new_n281));
  NAND4_X1  g080(.A1(new_n264), .A2(new_n268), .A3(new_n277), .A4(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT30), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  AOI22_X1  g083(.A1(new_n262), .A2(new_n263), .B1(new_n276), .B2(new_n208), .ZN(new_n285));
  NAND4_X1  g084(.A1(new_n285), .A2(KEYINPUT30), .A3(new_n268), .A4(new_n281), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n264), .A2(new_n281), .A3(new_n277), .ZN(new_n287));
  INV_X1    g086(.A(new_n268), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n284), .A2(new_n286), .A3(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT39), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT4), .ZN(new_n292));
  INV_X1    g091(.A(G113gat), .ZN(new_n293));
  INV_X1    g092(.A(G120gat), .ZN(new_n294));
  AOI21_X1  g093(.A(KEYINPUT1), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(G113gat), .A2(G120gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT67), .ZN(new_n298));
  INV_X1    g097(.A(G127gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(G134gat), .ZN(new_n300));
  INV_X1    g099(.A(G134gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(G127gat), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n298), .B1(new_n300), .B2(new_n302), .ZN(new_n303));
  AOI21_X1  g102(.A(KEYINPUT67), .B1(new_n299), .B2(G134gat), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n297), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND4_X1  g104(.A1(new_n295), .A2(new_n296), .A3(new_n300), .A4(new_n302), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n305), .A2(KEYINPUT68), .A3(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  AOI21_X1  g107(.A(KEYINPUT68), .B1(new_n305), .B2(new_n306), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  AND2_X1   g109(.A1(G155gat), .A2(G162gat), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(G155gat), .ZN(new_n313));
  INV_X1    g112(.A(G162gat), .ZN(new_n314));
  AND3_X1   g113(.A1(new_n313), .A2(new_n314), .A3(KEYINPUT78), .ZN(new_n315));
  AOI21_X1  g114(.A(KEYINPUT78), .B1(new_n313), .B2(new_n314), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n312), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT79), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  OAI211_X1 g118(.A(KEYINPUT79), .B(new_n312), .C1(new_n315), .C2(new_n316), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n312), .A2(KEYINPUT2), .ZN(new_n321));
  INV_X1    g120(.A(G141gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(G148gat), .ZN(new_n323));
  INV_X1    g122(.A(G148gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(G141gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n321), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n319), .A2(new_n320), .A3(new_n327), .ZN(new_n328));
  NOR2_X1   g127(.A1(G155gat), .A2(G162gat), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n311), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT80), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(new_n324), .ZN(new_n332));
  NAND2_X1  g131(.A1(KEYINPUT80), .A2(G148gat), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n332), .A2(G141gat), .A3(new_n333), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n330), .B1(new_n334), .B2(new_n323), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT82), .ZN(new_n336));
  XNOR2_X1  g135(.A(KEYINPUT81), .B(G155gat), .ZN(new_n337));
  OAI21_X1  g136(.A(KEYINPUT2), .B1(new_n337), .B2(new_n314), .ZN(new_n338));
  AND3_X1   g137(.A1(new_n335), .A2(new_n336), .A3(new_n338), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n336), .B1(new_n335), .B2(new_n338), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n328), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n292), .B1(new_n310), .B2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n330), .ZN(new_n343));
  AND2_X1   g142(.A1(KEYINPUT80), .A2(G148gat), .ZN(new_n344));
  NOR2_X1   g143(.A1(KEYINPUT80), .A2(G148gat), .ZN(new_n345));
  NOR3_X1   g144(.A1(new_n344), .A2(new_n345), .A3(new_n322), .ZN(new_n346));
  INV_X1    g145(.A(new_n323), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n343), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT2), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n313), .A2(KEYINPUT81), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT81), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(G155gat), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n349), .B1(new_n353), .B2(G162gat), .ZN(new_n354));
  OAI21_X1  g153(.A(KEYINPUT82), .B1(new_n348), .B2(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n335), .A2(new_n336), .A3(new_n338), .ZN(new_n356));
  AOI22_X1  g155(.A1(new_n317), .A2(new_n318), .B1(new_n321), .B2(new_n326), .ZN(new_n357));
  AOI22_X1  g156(.A1(new_n355), .A2(new_n356), .B1(new_n320), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n305), .A2(new_n306), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n358), .A2(KEYINPUT4), .A3(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT3), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n359), .B1(new_n358), .B2(new_n362), .ZN(new_n363));
  OAI211_X1 g162(.A(new_n362), .B(new_n328), .C1(new_n339), .C2(new_n340), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  OAI211_X1 g164(.A(new_n342), .B(new_n361), .C1(new_n363), .C2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT85), .ZN(new_n367));
  NAND2_X1  g166(.A1(G225gat), .A2(G233gat), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  AND3_X1   g168(.A1(new_n366), .A2(new_n367), .A3(new_n369), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n367), .B1(new_n366), .B2(new_n369), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n291), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n366), .A2(new_n369), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(KEYINPUT85), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n366), .A2(new_n367), .A3(new_n369), .ZN(new_n375));
  XNOR2_X1  g174(.A(new_n341), .B(new_n360), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n291), .B1(new_n376), .B2(new_n368), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n374), .A2(new_n375), .A3(new_n377), .ZN(new_n378));
  XNOR2_X1  g177(.A(G1gat), .B(G29gat), .ZN(new_n379));
  XNOR2_X1  g178(.A(new_n379), .B(KEYINPUT0), .ZN(new_n380));
  XNOR2_X1  g179(.A(new_n380), .B(G57gat), .ZN(new_n381));
  INV_X1    g180(.A(G85gat), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n381), .B(new_n382), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n372), .A2(new_n378), .A3(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT40), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  OR2_X1    g185(.A1(new_n369), .A2(KEYINPUT5), .ZN(new_n387));
  OR2_X1    g186(.A1(new_n366), .A2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(new_n309), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(new_n307), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n390), .A2(new_n358), .A3(KEYINPUT4), .ZN(new_n391));
  OAI22_X1  g190(.A1(new_n341), .A2(new_n359), .B1(new_n292), .B2(new_n369), .ZN(new_n392));
  OAI211_X1 g191(.A(new_n391), .B(new_n392), .C1(new_n363), .C2(new_n365), .ZN(new_n393));
  OAI211_X1 g192(.A(new_n393), .B(KEYINPUT5), .C1(new_n368), .C2(new_n376), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n388), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n383), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n386), .A2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT87), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n384), .A2(KEYINPUT86), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT86), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n372), .A2(new_n378), .A3(new_n402), .A4(new_n383), .ZN(new_n403));
  AND4_X1   g202(.A1(new_n400), .A2(new_n401), .A3(new_n385), .A4(new_n403), .ZN(new_n404));
  AOI21_X1  g203(.A(KEYINPUT40), .B1(new_n384), .B2(KEYINPUT86), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n400), .B1(new_n405), .B2(new_n403), .ZN(new_n406));
  OAI211_X1 g205(.A(new_n290), .B(new_n399), .C1(new_n404), .C2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT37), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n264), .A2(new_n408), .A3(new_n277), .A4(new_n281), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(new_n288), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n408), .B1(new_n285), .B2(new_n281), .ZN(new_n411));
  OAI21_X1  g210(.A(KEYINPUT38), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n408), .B1(new_n276), .B2(new_n209), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n280), .A2(new_n208), .A3(new_n252), .ZN(new_n414));
  AOI21_X1  g213(.A(KEYINPUT38), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n409), .A2(new_n415), .A3(new_n288), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT6), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n417), .B1(new_n395), .B2(new_n396), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(new_n397), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n398), .A2(KEYINPUT6), .ZN(new_n421));
  AND3_X1   g220(.A1(new_n420), .A2(new_n282), .A3(new_n421), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n412), .A2(new_n416), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n209), .A2(new_n278), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n358), .B1(new_n424), .B2(new_n362), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n209), .B1(new_n364), .B2(new_n278), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(G228gat), .ZN(new_n428));
  INV_X1    g227(.A(G233gat), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n427), .A2(new_n430), .ZN(new_n431));
  NOR4_X1   g230(.A1(new_n425), .A2(new_n426), .A3(new_n428), .A4(new_n429), .ZN(new_n432));
  NOR3_X1   g231(.A1(new_n431), .A2(new_n432), .A3(G22gat), .ZN(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  OAI21_X1  g233(.A(G22gat), .B1(new_n431), .B2(new_n432), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  XNOR2_X1  g235(.A(G78gat), .B(G106gat), .ZN(new_n437));
  XNOR2_X1  g236(.A(KEYINPUT31), .B(G50gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n437), .B(new_n438), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n439), .B1(new_n433), .B2(KEYINPUT84), .ZN(new_n440));
  XNOR2_X1  g239(.A(new_n436), .B(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n407), .A2(new_n423), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n418), .A2(KEYINPUT83), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT83), .ZN(new_n444));
  OAI211_X1 g243(.A(new_n444), .B(new_n417), .C1(new_n395), .C2(new_n396), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n443), .A2(new_n397), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(new_n421), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n447), .A2(new_n286), .A3(new_n289), .A4(new_n284), .ZN(new_n448));
  INV_X1    g247(.A(new_n441), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  XNOR2_X1  g249(.A(G15gat), .B(G43gat), .ZN(new_n451));
  XNOR2_X1  g250(.A(G71gat), .B(G99gat), .ZN(new_n452));
  XNOR2_X1  g251(.A(new_n451), .B(new_n452), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n390), .B1(new_n239), .B2(new_n251), .ZN(new_n454));
  NAND2_X1  g253(.A1(G227gat), .A2(G233gat), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n272), .A2(new_n310), .A3(new_n250), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n454), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT33), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n453), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT69), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n458), .A2(new_n461), .A3(KEYINPUT32), .ZN(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n461), .B1(new_n458), .B2(KEYINPUT32), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n460), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n458), .A2(KEYINPUT32), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT70), .ZN(new_n467));
  OR2_X1    g266(.A1(new_n453), .A2(new_n467), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n459), .B1(new_n453), .B2(new_n467), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n466), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n465), .A2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT73), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT34), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n456), .B1(new_n454), .B2(new_n457), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT71), .ZN(new_n476));
  OAI211_X1 g275(.A(KEYINPUT72), .B(new_n474), .C1(new_n475), .C2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT72), .ZN(new_n478));
  AOI211_X1 g277(.A(new_n251), .B(new_n390), .C1(new_n255), .C2(new_n256), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n310), .B1(new_n272), .B2(new_n250), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n455), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n478), .B1(new_n481), .B2(KEYINPUT71), .ZN(new_n482));
  AOI21_X1  g281(.A(KEYINPUT34), .B1(new_n481), .B2(new_n478), .ZN(new_n483));
  OAI211_X1 g282(.A(new_n473), .B(new_n477), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(new_n484), .ZN(new_n485));
  OAI21_X1  g284(.A(KEYINPUT72), .B1(new_n475), .B2(new_n476), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n474), .B1(new_n475), .B2(KEYINPUT72), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n473), .B1(new_n488), .B2(new_n477), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n472), .B1(new_n485), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n466), .A2(KEYINPUT69), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(new_n462), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n470), .B1(new_n492), .B2(new_n460), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n477), .B1(new_n482), .B2(new_n483), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(KEYINPUT73), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n493), .A2(new_n495), .A3(new_n484), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n490), .A2(KEYINPUT74), .A3(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT36), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT74), .ZN(new_n499));
  NAND4_X1  g298(.A1(new_n493), .A2(new_n495), .A3(new_n499), .A4(new_n484), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n497), .A2(new_n498), .A3(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n490), .A2(KEYINPUT36), .A3(new_n496), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n442), .A2(new_n450), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n497), .A2(new_n500), .ZN(new_n505));
  INV_X1    g304(.A(new_n290), .ZN(new_n506));
  AOI21_X1  g305(.A(KEYINPUT35), .B1(new_n420), .B2(new_n421), .ZN(new_n507));
  AND2_X1   g306(.A1(new_n507), .A2(new_n441), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n505), .A2(new_n506), .A3(new_n508), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n441), .A2(new_n490), .A3(new_n496), .ZN(new_n510));
  OAI21_X1  g309(.A(KEYINPUT35), .B1(new_n448), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n504), .A2(new_n512), .ZN(new_n513));
  XNOR2_X1  g312(.A(G15gat), .B(G22gat), .ZN(new_n514));
  INV_X1    g313(.A(G1gat), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(KEYINPUT16), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n517), .B1(G1gat), .B2(new_n514), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n518), .B(G8gat), .ZN(new_n519));
  INV_X1    g318(.A(G64gat), .ZN(new_n520));
  AND2_X1   g319(.A1(new_n520), .A2(G57gat), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n520), .A2(G57gat), .ZN(new_n522));
  AND2_X1   g321(.A1(G71gat), .A2(G78gat), .ZN(new_n523));
  OAI22_X1  g322(.A1(new_n521), .A2(new_n522), .B1(KEYINPUT9), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g323(.A1(G71gat), .A2(G78gat), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n524), .B(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n519), .B1(KEYINPUT21), .B2(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n529), .B(G183gat), .ZN(new_n530));
  XNOR2_X1  g329(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n531));
  NAND2_X1  g330(.A1(G231gat), .A2(G233gat), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n531), .B(new_n532), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n530), .B(new_n533), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n528), .A2(KEYINPUT21), .ZN(new_n535));
  XNOR2_X1  g334(.A(G127gat), .B(G155gat), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n535), .B(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n537), .B(new_n203), .ZN(new_n538));
  OR2_X1    g337(.A1(new_n534), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n534), .A2(new_n538), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  XNOR2_X1  g341(.A(G190gat), .B(G218gat), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT15), .ZN(new_n545));
  INV_X1    g344(.A(G50gat), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(G43gat), .ZN(new_n547));
  INV_X1    g346(.A(G43gat), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(G50gat), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT88), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n545), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n552), .B1(new_n551), .B2(new_n550), .ZN(new_n553));
  OR3_X1    g352(.A1(KEYINPUT89), .A2(G29gat), .A3(G36gat), .ZN(new_n554));
  OAI21_X1  g353(.A(KEYINPUT89), .B1(G29gat), .B2(G36gat), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n554), .A2(KEYINPUT14), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(G29gat), .A2(G36gat), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT90), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n557), .B(new_n558), .ZN(new_n559));
  OAI211_X1 g358(.A(new_n556), .B(new_n559), .C1(KEYINPUT14), .C2(new_n555), .ZN(new_n560));
  OAI21_X1  g359(.A(KEYINPUT91), .B1(new_n546), .B2(G43gat), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT91), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n562), .A2(new_n548), .A3(G50gat), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n561), .A2(new_n563), .A3(new_n547), .ZN(new_n564));
  AND2_X1   g363(.A1(new_n564), .A2(new_n545), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n553), .B1(new_n560), .B2(new_n565), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n566), .B1(new_n553), .B2(new_n560), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(KEYINPUT17), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n568), .B(KEYINPUT93), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n567), .B(KEYINPUT92), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT17), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(G99gat), .A2(G106gat), .ZN(new_n573));
  AOI22_X1  g372(.A1(KEYINPUT8), .A2(new_n573), .B1(new_n382), .B2(new_n267), .ZN(new_n574));
  NAND2_X1  g373(.A1(G85gat), .A2(G92gat), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT97), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT7), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n575), .B(KEYINPUT97), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n580), .A2(KEYINPUT7), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n574), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  XOR2_X1   g381(.A(G99gat), .B(G106gat), .Z(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n583), .ZN(new_n585));
  OAI211_X1 g384(.A(new_n585), .B(new_n574), .C1(new_n579), .C2(new_n581), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n584), .A2(new_n586), .A3(KEYINPUT98), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT98), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n582), .A2(new_n588), .A3(new_n583), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n569), .A2(new_n572), .A3(new_n591), .ZN(new_n592));
  AND2_X1   g391(.A1(G232gat), .A2(G233gat), .ZN(new_n593));
  AOI22_X1  g392(.A1(new_n570), .A2(new_n590), .B1(KEYINPUT41), .B2(new_n593), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n544), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT99), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n592), .A2(new_n544), .A3(new_n594), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n593), .A2(KEYINPUT41), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(KEYINPUT96), .ZN(new_n600));
  XOR2_X1   g399(.A(G134gat), .B(G162gat), .Z(new_n601));
  XOR2_X1   g400(.A(new_n600), .B(new_n601), .Z(new_n602));
  NAND4_X1  g401(.A1(new_n596), .A2(new_n597), .A3(new_n598), .A4(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n592), .A2(new_n594), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n597), .B1(new_n604), .B2(new_n543), .ZN(new_n605));
  INV_X1    g404(.A(new_n602), .ZN(new_n606));
  INV_X1    g405(.A(new_n598), .ZN(new_n607));
  OAI22_X1  g406(.A1(new_n605), .A2(new_n606), .B1(new_n607), .B2(new_n595), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n542), .B1(new_n603), .B2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n519), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n569), .A2(new_n572), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(G229gat), .A2(G233gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(KEYINPUT94), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n570), .A2(new_n519), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n612), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT18), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  OR2_X1    g418(.A1(new_n567), .A2(KEYINPUT92), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n567), .A2(KEYINPUT92), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n620), .A2(new_n621), .A3(new_n611), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT95), .ZN(new_n623));
  OR2_X1    g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n622), .A2(new_n623), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n624), .A2(new_n616), .A3(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n614), .B(KEYINPUT13), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND4_X1  g427(.A1(new_n612), .A2(KEYINPUT18), .A3(new_n615), .A4(new_n616), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n619), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(G113gat), .B(G141gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n631), .B(KEYINPUT11), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(new_n224), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(G197gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(KEYINPUT12), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n630), .A2(new_n636), .ZN(new_n637));
  NAND4_X1  g436(.A1(new_n619), .A2(new_n628), .A3(new_n635), .A4(new_n629), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(G230gat), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n641), .A2(new_n429), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n587), .A2(new_n589), .A3(new_n527), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT10), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n527), .B1(new_n582), .B2(new_n583), .ZN(new_n645));
  AND3_X1   g444(.A1(new_n645), .A2(KEYINPUT100), .A3(new_n586), .ZN(new_n646));
  AOI21_X1  g445(.A(KEYINPUT100), .B1(new_n645), .B2(new_n586), .ZN(new_n647));
  OAI211_X1 g446(.A(new_n643), .B(new_n644), .C1(new_n646), .C2(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n590), .A2(KEYINPUT10), .A3(new_n528), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n642), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n643), .B1(new_n646), .B2(new_n647), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n652), .A2(new_n642), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(G120gat), .B(G148gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(G176gat), .ZN(new_n656));
  INV_X1    g455(.A(G204gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n656), .B(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n654), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n654), .A2(new_n659), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NOR3_X1   g462(.A1(new_n610), .A2(new_n640), .A3(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n513), .A2(new_n664), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n665), .A2(new_n447), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(new_n515), .ZN(G1324gat));
  INV_X1    g466(.A(KEYINPUT101), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n513), .A2(new_n290), .A3(new_n664), .ZN(new_n669));
  XNOR2_X1  g468(.A(KEYINPUT16), .B(G8gat), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n668), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  OR2_X1    g470(.A1(new_n671), .A2(KEYINPUT42), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(KEYINPUT42), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n669), .A2(G8gat), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n672), .A2(new_n673), .A3(new_n674), .ZN(G1325gat));
  OAI21_X1  g474(.A(G15gat), .B1(new_n665), .B2(new_n503), .ZN(new_n676));
  INV_X1    g475(.A(new_n505), .ZN(new_n677));
  OR2_X1    g476(.A1(new_n677), .A2(G15gat), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n676), .B1(new_n665), .B2(new_n678), .ZN(G1326gat));
  NOR2_X1   g478(.A1(new_n665), .A2(new_n441), .ZN(new_n680));
  XOR2_X1   g479(.A(KEYINPUT43), .B(G22gat), .Z(new_n681));
  XNOR2_X1  g480(.A(new_n680), .B(new_n681), .ZN(G1327gat));
  NAND2_X1  g481(.A1(new_n608), .A2(new_n603), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  NOR3_X1   g483(.A1(new_n640), .A2(new_n541), .A3(new_n663), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n513), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  NOR3_X1   g485(.A1(new_n686), .A2(G29gat), .A3(new_n447), .ZN(new_n687));
  XOR2_X1   g486(.A(new_n687), .B(KEYINPUT45), .Z(new_n688));
  AOI22_X1  g487(.A1(new_n501), .A2(new_n502), .B1(new_n449), .B2(new_n448), .ZN(new_n689));
  AOI22_X1  g488(.A1(new_n689), .A2(new_n442), .B1(new_n511), .B2(new_n509), .ZN(new_n690));
  OAI21_X1  g489(.A(KEYINPUT44), .B1(new_n690), .B2(new_n683), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT44), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n513), .A2(new_n692), .A3(new_n684), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  AND2_X1   g493(.A1(new_n694), .A2(new_n685), .ZN(new_n695));
  INV_X1    g494(.A(new_n447), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n697), .A2(G29gat), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n688), .A2(new_n698), .ZN(G1328gat));
  INV_X1    g498(.A(G36gat), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n695), .A2(new_n290), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n700), .B1(new_n701), .B2(KEYINPUT102), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n702), .B1(KEYINPUT102), .B2(new_n701), .ZN(new_n703));
  NOR3_X1   g502(.A1(new_n686), .A2(G36gat), .A3(new_n506), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n704), .B(KEYINPUT46), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n703), .A2(new_n705), .ZN(G1329gat));
  NOR3_X1   g505(.A1(new_n686), .A2(G43gat), .A3(new_n677), .ZN(new_n707));
  INV_X1    g506(.A(new_n503), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n695), .A2(new_n708), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n707), .B1(new_n709), .B2(G43gat), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(KEYINPUT47), .ZN(G1330gat));
  NOR3_X1   g510(.A1(new_n686), .A2(G50gat), .A3(new_n441), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n695), .A2(new_n449), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n712), .B1(new_n713), .B2(G50gat), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT48), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n715), .B1(new_n712), .B2(KEYINPUT103), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n714), .B(new_n716), .ZN(G1331gat));
  INV_X1    g516(.A(new_n663), .ZN(new_n718));
  NOR4_X1   g517(.A1(new_n690), .A2(new_n639), .A3(new_n610), .A4(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(new_n696), .ZN(new_n720));
  XOR2_X1   g519(.A(KEYINPUT104), .B(G57gat), .Z(new_n721));
  XNOR2_X1  g520(.A(new_n720), .B(new_n721), .ZN(G1332gat));
  NAND2_X1  g521(.A1(new_n719), .A2(new_n290), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n723), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n724));
  XOR2_X1   g523(.A(KEYINPUT49), .B(G64gat), .Z(new_n725));
  OAI21_X1  g524(.A(new_n724), .B1(new_n723), .B2(new_n725), .ZN(G1333gat));
  NAND2_X1  g525(.A1(new_n719), .A2(new_n708), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n677), .A2(G71gat), .ZN(new_n728));
  AOI22_X1  g527(.A1(new_n727), .A2(G71gat), .B1(new_n719), .B2(new_n728), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g529(.A1(new_n719), .A2(new_n449), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g531(.A1(new_n639), .A2(new_n541), .ZN(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n734), .A2(new_n718), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n692), .B1(new_n513), .B2(new_n684), .ZN(new_n736));
  AOI211_X1 g535(.A(KEYINPUT44), .B(new_n683), .C1(new_n504), .C2(new_n512), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n735), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT105), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n694), .A2(KEYINPUT105), .A3(new_n735), .ZN(new_n741));
  AND2_X1   g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n382), .B1(new_n742), .B2(new_n696), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n513), .A2(new_n684), .A3(new_n733), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n718), .B1(new_n744), .B2(KEYINPUT51), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT51), .ZN(new_n746));
  NAND4_X1  g545(.A1(new_n513), .A2(new_n746), .A3(new_n684), .A4(new_n733), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  NOR3_X1   g547(.A1(new_n748), .A2(G85gat), .A3(new_n447), .ZN(new_n749));
  OR3_X1    g548(.A1(new_n743), .A2(KEYINPUT106), .A3(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(KEYINPUT106), .B1(new_n743), .B2(new_n749), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(G1336gat));
  NAND2_X1  g551(.A1(new_n744), .A2(KEYINPUT51), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n506), .A2(G92gat), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n753), .A2(new_n663), .A3(new_n747), .A4(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT109), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND4_X1  g556(.A1(new_n745), .A2(KEYINPUT109), .A3(new_n747), .A4(new_n754), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  OAI211_X1 g558(.A(new_n290), .B(new_n735), .C1(new_n736), .C2(new_n737), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT110), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND4_X1  g561(.A1(new_n694), .A2(KEYINPUT110), .A3(new_n290), .A4(new_n735), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n762), .A2(G92gat), .A3(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT52), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n759), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT111), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n759), .A2(new_n764), .A3(KEYINPUT111), .A4(new_n765), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT108), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n740), .A2(new_n290), .A3(new_n741), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(G92gat), .ZN(new_n773));
  NOR3_X1   g572(.A1(new_n690), .A2(new_n683), .A3(new_n734), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n746), .B1(new_n774), .B2(KEYINPUT107), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT107), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n744), .A2(new_n776), .A3(KEYINPUT51), .ZN(new_n777));
  AND4_X1   g576(.A1(new_n663), .A2(new_n775), .A3(new_n754), .A4(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n773), .A2(new_n779), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n771), .B1(new_n780), .B2(KEYINPUT52), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n778), .B1(new_n772), .B2(G92gat), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n782), .A2(KEYINPUT108), .A3(new_n765), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n770), .B1(new_n781), .B2(new_n783), .ZN(G1337gat));
  NAND3_X1  g583(.A1(new_n742), .A2(G99gat), .A3(new_n708), .ZN(new_n785));
  INV_X1    g584(.A(G99gat), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n786), .B1(new_n748), .B2(new_n677), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(KEYINPUT112), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT112), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n785), .A2(new_n790), .A3(new_n787), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n789), .A2(new_n791), .ZN(G1338gat));
  OAI21_X1  g591(.A(G106gat), .B1(new_n738), .B2(new_n441), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT53), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n441), .A2(G106gat), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n745), .A2(new_n747), .A3(new_n795), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n793), .A2(new_n794), .A3(new_n796), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n740), .A2(new_n449), .A3(new_n741), .ZN(new_n798));
  AND2_X1   g597(.A1(new_n798), .A2(G106gat), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n775), .A2(new_n663), .A3(new_n777), .A4(new_n795), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT113), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  AND2_X1   g601(.A1(new_n800), .A2(new_n801), .ZN(new_n803));
  NOR3_X1   g602(.A1(new_n799), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n797), .B1(new_n804), .B2(new_n794), .ZN(G1339gat));
  NAND3_X1  g604(.A1(new_n609), .A2(new_n640), .A3(new_n718), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(KEYINPUT114), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT114), .ZN(new_n808));
  NAND4_X1  g607(.A1(new_n609), .A2(new_n640), .A3(new_n808), .A4(new_n718), .ZN(new_n809));
  AND2_X1   g608(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  AOI211_X1 g609(.A(KEYINPUT54), .B(new_n642), .C1(new_n648), .C2(new_n649), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT115), .ZN(new_n812));
  NOR3_X1   g611(.A1(new_n811), .A2(new_n812), .A3(new_n658), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT54), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n650), .A2(new_n814), .ZN(new_n815));
  AOI21_X1  g614(.A(KEYINPUT115), .B1(new_n815), .B2(new_n659), .ZN(new_n816));
  AND3_X1   g615(.A1(new_n648), .A2(new_n642), .A3(new_n649), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n651), .A2(KEYINPUT54), .ZN(new_n818));
  OAI22_X1  g617(.A1(new_n813), .A2(new_n816), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT116), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT55), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n819), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n817), .A2(new_n650), .A3(new_n814), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n812), .B1(new_n811), .B2(new_n658), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n815), .A2(KEYINPUT115), .A3(new_n659), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n823), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  OAI21_X1  g625(.A(KEYINPUT116), .B1(new_n826), .B2(KEYINPUT55), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n822), .A2(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n660), .B1(new_n826), .B2(KEYINPUT55), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n626), .A2(new_n627), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n615), .B1(new_n612), .B2(new_n616), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n634), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  AND4_X1   g631(.A1(new_n638), .A2(new_n608), .A3(new_n832), .A4(new_n603), .ZN(new_n833));
  AND3_X1   g632(.A1(new_n828), .A2(new_n829), .A3(new_n833), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n820), .B1(new_n819), .B2(new_n821), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n826), .A2(KEYINPUT116), .A3(KEYINPUT55), .ZN(new_n836));
  OAI211_X1 g635(.A(new_n639), .B(new_n829), .C1(new_n835), .C2(new_n836), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n832), .A2(new_n638), .A3(new_n663), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n834), .B1(new_n839), .B2(new_n683), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n810), .B1(new_n840), .B2(new_n541), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n290), .A2(new_n447), .ZN(new_n842));
  AND2_X1   g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(new_n510), .ZN(new_n844));
  AND2_X1   g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g644(.A(G113gat), .B1(new_n845), .B2(new_n639), .ZN(new_n846));
  INV_X1    g645(.A(new_n841), .ZN(new_n847));
  NOR3_X1   g646(.A1(new_n847), .A2(new_n449), .A3(new_n677), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n848), .A2(new_n842), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n640), .A2(new_n293), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n846), .B1(new_n849), .B2(new_n850), .ZN(G1340gat));
  AOI21_X1  g650(.A(G120gat), .B1(new_n845), .B2(new_n663), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n718), .A2(new_n294), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n852), .B1(new_n849), .B2(new_n853), .ZN(G1341gat));
  NAND3_X1  g653(.A1(new_n849), .A2(G127gat), .A3(new_n541), .ZN(new_n855));
  AND2_X1   g654(.A1(new_n855), .A2(KEYINPUT117), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n855), .A2(KEYINPUT117), .ZN(new_n857));
  AOI21_X1  g656(.A(G127gat), .B1(new_n845), .B2(new_n541), .ZN(new_n858));
  NOR3_X1   g657(.A1(new_n856), .A2(new_n857), .A3(new_n858), .ZN(G1342gat));
  NAND3_X1  g658(.A1(new_n845), .A2(new_n301), .A3(new_n684), .ZN(new_n860));
  AND2_X1   g659(.A1(new_n860), .A2(KEYINPUT56), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n301), .B1(new_n849), .B2(new_n684), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n863), .B1(KEYINPUT56), .B2(new_n860), .ZN(G1343gat));
  AND2_X1   g663(.A1(new_n503), .A2(new_n842), .ZN(new_n865));
  AOI21_X1  g664(.A(KEYINPUT57), .B1(new_n841), .B2(new_n449), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n449), .A2(KEYINPUT57), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n819), .A2(new_n821), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n639), .A2(new_n829), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n684), .B1(new_n869), .B2(new_n838), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n542), .B1(new_n834), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n867), .B1(new_n810), .B2(new_n871), .ZN(new_n872));
  OAI211_X1 g671(.A(new_n639), .B(new_n865), .C1(new_n866), .C2(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n322), .B1(new_n873), .B2(KEYINPUT120), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n874), .B1(KEYINPUT120), .B2(new_n873), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT58), .ZN(new_n876));
  AND3_X1   g675(.A1(new_n843), .A2(new_n449), .A3(new_n503), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n877), .A2(new_n322), .A3(new_n639), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n875), .A2(new_n876), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n873), .A2(G141gat), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(KEYINPUT118), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT118), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n873), .A2(new_n882), .A3(G141gat), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n881), .A2(new_n883), .A3(new_n878), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT119), .ZN(new_n885));
  AND3_X1   g684(.A1(new_n884), .A2(new_n885), .A3(KEYINPUT58), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n885), .B1(new_n884), .B2(KEYINPUT58), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n879), .B1(new_n886), .B2(new_n887), .ZN(G1344gat));
  NAND2_X1  g687(.A1(new_n332), .A2(new_n333), .ZN(new_n889));
  INV_X1    g688(.A(new_n889), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n877), .A2(new_n890), .A3(new_n663), .ZN(new_n891));
  XNOR2_X1  g690(.A(new_n891), .B(KEYINPUT121), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n865), .B1(new_n866), .B2(new_n872), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n893), .A2(new_n718), .ZN(new_n894));
  NOR3_X1   g693(.A1(new_n894), .A2(KEYINPUT59), .A3(new_n890), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT59), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n847), .A2(new_n867), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n871), .A2(new_n806), .ZN(new_n898));
  AOI21_X1  g697(.A(KEYINPUT57), .B1(new_n898), .B2(new_n449), .ZN(new_n899));
  OR2_X1    g698(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n900), .A2(new_n663), .A3(new_n865), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n896), .B1(new_n901), .B2(G148gat), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n892), .B1(new_n895), .B2(new_n902), .ZN(G1345gat));
  NAND3_X1  g702(.A1(new_n877), .A2(new_n337), .A3(new_n541), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n353), .B1(new_n893), .B2(new_n542), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(G1346gat));
  NAND3_X1  g705(.A1(new_n877), .A2(new_n314), .A3(new_n684), .ZN(new_n907));
  OAI21_X1  g706(.A(G162gat), .B1(new_n893), .B2(new_n683), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(G1347gat));
  NOR2_X1   g708(.A1(new_n506), .A2(new_n696), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n841), .A2(new_n844), .A3(new_n910), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n911), .A2(G169gat), .A3(new_n640), .ZN(new_n912));
  XNOR2_X1  g711(.A(new_n912), .B(KEYINPUT122), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n848), .A2(new_n910), .ZN(new_n914));
  OAI21_X1  g713(.A(G169gat), .B1(new_n914), .B2(new_n640), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n913), .A2(new_n915), .ZN(G1348gat));
  NAND4_X1  g715(.A1(new_n848), .A2(G176gat), .A3(new_n663), .A4(new_n910), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT123), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n917), .A2(new_n918), .ZN(new_n920));
  INV_X1    g719(.A(new_n911), .ZN(new_n921));
  AOI21_X1  g720(.A(G176gat), .B1(new_n921), .B2(new_n663), .ZN(new_n922));
  NOR3_X1   g721(.A1(new_n919), .A2(new_n920), .A3(new_n922), .ZN(G1349gat));
  OAI21_X1  g722(.A(G183gat), .B1(new_n914), .B2(new_n542), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n921), .A2(new_n240), .A3(new_n541), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  XNOR2_X1  g725(.A(new_n926), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g726(.A1(new_n921), .A2(new_n216), .A3(new_n684), .ZN(new_n928));
  OAI21_X1  g727(.A(G190gat), .B1(new_n914), .B2(new_n683), .ZN(new_n929));
  AND2_X1   g728(.A1(new_n929), .A2(KEYINPUT61), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n929), .A2(KEYINPUT61), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n928), .B1(new_n930), .B2(new_n931), .ZN(G1351gat));
  INV_X1    g731(.A(G197gat), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n847), .A2(new_n441), .ZN(new_n934));
  AND2_X1   g733(.A1(new_n503), .A2(new_n910), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n933), .B1(new_n936), .B2(new_n640), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n900), .A2(KEYINPUT124), .ZN(new_n938));
  OR3_X1    g737(.A1(new_n897), .A2(KEYINPUT124), .A3(new_n899), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n938), .A2(new_n935), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n639), .A2(G197gat), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n937), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT125), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  OAI211_X1 g743(.A(KEYINPUT125), .B(new_n937), .C1(new_n940), .C2(new_n941), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(G1352gat));
  OAI21_X1  g745(.A(G204gat), .B1(new_n940), .B2(new_n718), .ZN(new_n947));
  NOR3_X1   g746(.A1(new_n936), .A2(G204gat), .A3(new_n718), .ZN(new_n948));
  XNOR2_X1  g747(.A(new_n948), .B(KEYINPUT62), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n947), .A2(new_n949), .ZN(G1353gat));
  OAI211_X1 g749(.A(new_n541), .B(new_n935), .C1(new_n897), .C2(new_n899), .ZN(new_n951));
  AND3_X1   g750(.A1(new_n951), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n952));
  AOI21_X1  g751(.A(KEYINPUT63), .B1(new_n951), .B2(G211gat), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n541), .A2(new_n203), .ZN(new_n954));
  OAI22_X1  g753(.A1(new_n952), .A2(new_n953), .B1(new_n936), .B2(new_n954), .ZN(new_n955));
  XNOR2_X1  g754(.A(new_n955), .B(KEYINPUT126), .ZN(G1354gat));
  OAI21_X1  g755(.A(new_n204), .B1(new_n936), .B2(new_n683), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n684), .A2(G218gat), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n957), .B1(new_n940), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n959), .A2(KEYINPUT127), .ZN(new_n960));
  INV_X1    g759(.A(KEYINPUT127), .ZN(new_n961));
  OAI211_X1 g760(.A(new_n961), .B(new_n957), .C1(new_n940), .C2(new_n958), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n960), .A2(new_n962), .ZN(G1355gat));
endmodule


