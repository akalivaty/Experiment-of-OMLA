

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U546 ( .A(KEYINPUT17), .ZN(n515) );
  XNOR2_X1 U547 ( .A(n739), .B(n738), .ZN(n753) );
  INV_X1 U548 ( .A(KEYINPUT96), .ZN(n738) );
  NAND2_X1 U549 ( .A1(n867), .A2(G138), .ZN(n536) );
  AND2_X1 U550 ( .A1(n512), .A2(n977), .ZN(n511) );
  OR2_X1 U551 ( .A1(n757), .A2(n748), .ZN(n512) );
  NOR2_X1 U552 ( .A1(n736), .A2(n735), .ZN(n513) );
  OR2_X1 U553 ( .A1(KEYINPUT33), .A2(n746), .ZN(n514) );
  NOR2_X1 U554 ( .A1(G299), .A2(n711), .ZN(n708) );
  NOR2_X1 U555 ( .A1(n715), .A2(n714), .ZN(n716) );
  INV_X1 U556 ( .A(KEYINPUT31), .ZN(n689) );
  XNOR2_X1 U557 ( .A(KEYINPUT98), .B(KEYINPUT32), .ZN(n732) );
  XNOR2_X1 U558 ( .A(n733), .B(n732), .ZN(n752) );
  NOR2_X1 U559 ( .A1(G2104), .A2(n521), .ZN(n871) );
  NOR2_X1 U560 ( .A1(G651), .A2(n640), .ZN(n642) );
  NOR2_X1 U561 ( .A1(G651), .A2(G543), .ZN(n637) );
  AND2_X1 U562 ( .A1(n526), .A2(n525), .ZN(G160) );
  NOR2_X1 U563 ( .A1(G2104), .A2(G2105), .ZN(n516) );
  XNOR2_X2 U564 ( .A(n516), .B(n515), .ZN(n867) );
  NAND2_X1 U565 ( .A1(n867), .A2(G137), .ZN(n518) );
  AND2_X1 U566 ( .A1(G2104), .A2(G2105), .ZN(n874) );
  NAND2_X1 U567 ( .A1(n874), .A2(G113), .ZN(n517) );
  AND2_X1 U568 ( .A1(n518), .A2(n517), .ZN(n526) );
  XOR2_X1 U569 ( .A(KEYINPUT64), .B(KEYINPUT23), .Z(n520) );
  INV_X1 U570 ( .A(G2105), .ZN(n521) );
  AND2_X1 U571 ( .A1(n521), .A2(G2104), .ZN(n866) );
  NAND2_X1 U572 ( .A1(G101), .A2(n866), .ZN(n519) );
  XNOR2_X1 U573 ( .A(n520), .B(n519), .ZN(n523) );
  NAND2_X1 U574 ( .A1(n871), .A2(G125), .ZN(n522) );
  NAND2_X1 U575 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U576 ( .A(KEYINPUT65), .B(n524), .ZN(n525) );
  XOR2_X1 U577 ( .A(KEYINPUT0), .B(G543), .Z(n640) );
  INV_X1 U578 ( .A(G651), .ZN(n530) );
  NOR2_X1 U579 ( .A1(n640), .A2(n530), .ZN(n633) );
  NAND2_X1 U580 ( .A1(G78), .A2(n633), .ZN(n528) );
  NAND2_X1 U581 ( .A1(G91), .A2(n637), .ZN(n527) );
  NAND2_X1 U582 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U583 ( .A(KEYINPUT69), .B(n529), .ZN(n535) );
  NOR2_X1 U584 ( .A1(G543), .A2(n530), .ZN(n531) );
  XOR2_X1 U585 ( .A(KEYINPUT1), .B(n531), .Z(n646) );
  NAND2_X1 U586 ( .A1(G65), .A2(n646), .ZN(n533) );
  NAND2_X1 U587 ( .A1(G53), .A2(n642), .ZN(n532) );
  AND2_X1 U588 ( .A1(n533), .A2(n532), .ZN(n534) );
  NAND2_X1 U589 ( .A1(n535), .A2(n534), .ZN(G299) );
  INV_X1 U590 ( .A(KEYINPUT83), .ZN(n539) );
  NAND2_X1 U591 ( .A1(G102), .A2(n866), .ZN(n537) );
  NAND2_X1 U592 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U593 ( .A(n539), .B(n538), .ZN(n544) );
  NAND2_X1 U594 ( .A1(G126), .A2(n871), .ZN(n541) );
  NAND2_X1 U595 ( .A1(G114), .A2(n874), .ZN(n540) );
  NAND2_X1 U596 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U597 ( .A(KEYINPUT82), .B(n542), .ZN(n543) );
  NOR2_X1 U598 ( .A1(n544), .A2(n543), .ZN(G164) );
  NAND2_X1 U599 ( .A1(G64), .A2(n646), .ZN(n546) );
  NAND2_X1 U600 ( .A1(G52), .A2(n642), .ZN(n545) );
  NAND2_X1 U601 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U602 ( .A(KEYINPUT68), .B(n547), .ZN(n552) );
  NAND2_X1 U603 ( .A1(G77), .A2(n633), .ZN(n549) );
  NAND2_X1 U604 ( .A1(G90), .A2(n637), .ZN(n548) );
  NAND2_X1 U605 ( .A1(n549), .A2(n548), .ZN(n550) );
  XOR2_X1 U606 ( .A(KEYINPUT9), .B(n550), .Z(n551) );
  NOR2_X1 U607 ( .A1(n552), .A2(n551), .ZN(G171) );
  AND2_X1 U608 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U609 ( .A(G132), .ZN(G219) );
  INV_X1 U610 ( .A(G82), .ZN(G220) );
  INV_X1 U611 ( .A(G120), .ZN(G236) );
  INV_X1 U612 ( .A(G57), .ZN(G237) );
  NAND2_X1 U613 ( .A1(G75), .A2(n633), .ZN(n554) );
  NAND2_X1 U614 ( .A1(G88), .A2(n637), .ZN(n553) );
  NAND2_X1 U615 ( .A1(n554), .A2(n553), .ZN(n558) );
  NAND2_X1 U616 ( .A1(G62), .A2(n646), .ZN(n556) );
  NAND2_X1 U617 ( .A1(G50), .A2(n642), .ZN(n555) );
  NAND2_X1 U618 ( .A1(n556), .A2(n555), .ZN(n557) );
  NOR2_X1 U619 ( .A1(n558), .A2(n557), .ZN(G166) );
  NAND2_X1 U620 ( .A1(n637), .A2(G89), .ZN(n559) );
  XNOR2_X1 U621 ( .A(n559), .B(KEYINPUT4), .ZN(n561) );
  NAND2_X1 U622 ( .A1(G76), .A2(n633), .ZN(n560) );
  NAND2_X1 U623 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U624 ( .A(n562), .B(KEYINPUT5), .ZN(n568) );
  XNOR2_X1 U625 ( .A(KEYINPUT6), .B(KEYINPUT73), .ZN(n566) );
  NAND2_X1 U626 ( .A1(G63), .A2(n646), .ZN(n564) );
  NAND2_X1 U627 ( .A1(G51), .A2(n642), .ZN(n563) );
  NAND2_X1 U628 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U629 ( .A(n566), .B(n565), .ZN(n567) );
  NAND2_X1 U630 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U631 ( .A(KEYINPUT7), .B(n569), .ZN(G168) );
  XOR2_X1 U632 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U633 ( .A1(G7), .A2(G661), .ZN(n570) );
  XNOR2_X1 U634 ( .A(n570), .B(KEYINPUT10), .ZN(n571) );
  XNOR2_X1 U635 ( .A(KEYINPUT70), .B(n571), .ZN(G223) );
  INV_X1 U636 ( .A(G223), .ZN(n815) );
  NAND2_X1 U637 ( .A1(n815), .A2(G567), .ZN(n572) );
  XOR2_X1 U638 ( .A(KEYINPUT11), .B(n572), .Z(G234) );
  NAND2_X1 U639 ( .A1(n646), .A2(G56), .ZN(n573) );
  XOR2_X1 U640 ( .A(KEYINPUT14), .B(n573), .Z(n580) );
  NAND2_X1 U641 ( .A1(n633), .A2(G68), .ZN(n574) );
  XNOR2_X1 U642 ( .A(KEYINPUT71), .B(n574), .ZN(n577) );
  NAND2_X1 U643 ( .A1(n637), .A2(G81), .ZN(n575) );
  XOR2_X1 U644 ( .A(KEYINPUT12), .B(n575), .Z(n576) );
  NOR2_X1 U645 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U646 ( .A(n578), .B(KEYINPUT13), .ZN(n579) );
  NOR2_X1 U647 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U648 ( .A(n581), .B(KEYINPUT72), .ZN(n583) );
  NAND2_X1 U649 ( .A1(G43), .A2(n642), .ZN(n582) );
  NAND2_X1 U650 ( .A1(n583), .A2(n582), .ZN(n983) );
  INV_X1 U651 ( .A(n983), .ZN(n584) );
  NAND2_X1 U652 ( .A1(n584), .A2(G860), .ZN(G153) );
  INV_X1 U653 ( .A(G171), .ZN(G301) );
  NAND2_X1 U654 ( .A1(G868), .A2(G301), .ZN(n593) );
  NAND2_X1 U655 ( .A1(G79), .A2(n633), .ZN(n586) );
  NAND2_X1 U656 ( .A1(G92), .A2(n637), .ZN(n585) );
  NAND2_X1 U657 ( .A1(n586), .A2(n585), .ZN(n590) );
  NAND2_X1 U658 ( .A1(G66), .A2(n646), .ZN(n588) );
  NAND2_X1 U659 ( .A1(G54), .A2(n642), .ZN(n587) );
  NAND2_X1 U660 ( .A1(n588), .A2(n587), .ZN(n589) );
  NOR2_X1 U661 ( .A1(n590), .A2(n589), .ZN(n591) );
  XOR2_X1 U662 ( .A(KEYINPUT15), .B(n591), .Z(n968) );
  INV_X1 U663 ( .A(n968), .ZN(n599) );
  INV_X1 U664 ( .A(G868), .ZN(n657) );
  NAND2_X1 U665 ( .A1(n599), .A2(n657), .ZN(n592) );
  NAND2_X1 U666 ( .A1(n593), .A2(n592), .ZN(G284) );
  NOR2_X1 U667 ( .A1(G868), .A2(G299), .ZN(n595) );
  NOR2_X1 U668 ( .A1(G286), .A2(n657), .ZN(n594) );
  NOR2_X1 U669 ( .A1(n595), .A2(n594), .ZN(G297) );
  INV_X1 U670 ( .A(G559), .ZN(n596) );
  NOR2_X1 U671 ( .A1(G860), .A2(n596), .ZN(n597) );
  XNOR2_X1 U672 ( .A(n597), .B(KEYINPUT74), .ZN(n598) );
  NOR2_X1 U673 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U674 ( .A(n600), .B(KEYINPUT16), .ZN(n601) );
  XNOR2_X1 U675 ( .A(n601), .B(KEYINPUT75), .ZN(G148) );
  NOR2_X1 U676 ( .A1(G868), .A2(n983), .ZN(n604) );
  NAND2_X1 U677 ( .A1(G868), .A2(n968), .ZN(n602) );
  NOR2_X1 U678 ( .A1(G559), .A2(n602), .ZN(n603) );
  NOR2_X1 U679 ( .A1(n604), .A2(n603), .ZN(G282) );
  NAND2_X1 U680 ( .A1(G123), .A2(n871), .ZN(n605) );
  XNOR2_X1 U681 ( .A(n605), .B(KEYINPUT18), .ZN(n612) );
  NAND2_X1 U682 ( .A1(G99), .A2(n866), .ZN(n607) );
  NAND2_X1 U683 ( .A1(G135), .A2(n867), .ZN(n606) );
  NAND2_X1 U684 ( .A1(n607), .A2(n606), .ZN(n610) );
  NAND2_X1 U685 ( .A1(n874), .A2(G111), .ZN(n608) );
  XOR2_X1 U686 ( .A(KEYINPUT76), .B(n608), .Z(n609) );
  NOR2_X1 U687 ( .A1(n610), .A2(n609), .ZN(n611) );
  NAND2_X1 U688 ( .A1(n612), .A2(n611), .ZN(n906) );
  XOR2_X1 U689 ( .A(n906), .B(G2096), .Z(n614) );
  XNOR2_X1 U690 ( .A(G2100), .B(KEYINPUT77), .ZN(n613) );
  NAND2_X1 U691 ( .A1(n614), .A2(n613), .ZN(G156) );
  NAND2_X1 U692 ( .A1(G559), .A2(n968), .ZN(n615) );
  XNOR2_X1 U693 ( .A(n615), .B(n983), .ZN(n655) );
  NOR2_X1 U694 ( .A1(n655), .A2(G860), .ZN(n622) );
  NAND2_X1 U695 ( .A1(G67), .A2(n646), .ZN(n617) );
  NAND2_X1 U696 ( .A1(G55), .A2(n642), .ZN(n616) );
  NAND2_X1 U697 ( .A1(n617), .A2(n616), .ZN(n621) );
  NAND2_X1 U698 ( .A1(G80), .A2(n633), .ZN(n619) );
  NAND2_X1 U699 ( .A1(G93), .A2(n637), .ZN(n618) );
  NAND2_X1 U700 ( .A1(n619), .A2(n618), .ZN(n620) );
  OR2_X1 U701 ( .A1(n621), .A2(n620), .ZN(n658) );
  XOR2_X1 U702 ( .A(n622), .B(n658), .Z(G145) );
  NAND2_X1 U703 ( .A1(n646), .A2(G60), .ZN(n629) );
  NAND2_X1 U704 ( .A1(G72), .A2(n633), .ZN(n624) );
  NAND2_X1 U705 ( .A1(G85), .A2(n637), .ZN(n623) );
  NAND2_X1 U706 ( .A1(n624), .A2(n623), .ZN(n627) );
  NAND2_X1 U707 ( .A1(n642), .A2(G47), .ZN(n625) );
  XOR2_X1 U708 ( .A(KEYINPUT66), .B(n625), .Z(n626) );
  NOR2_X1 U709 ( .A1(n627), .A2(n626), .ZN(n628) );
  NAND2_X1 U710 ( .A1(n629), .A2(n628), .ZN(n630) );
  XOR2_X1 U711 ( .A(KEYINPUT67), .B(n630), .Z(G290) );
  NAND2_X1 U712 ( .A1(G61), .A2(n646), .ZN(n632) );
  NAND2_X1 U713 ( .A1(G48), .A2(n642), .ZN(n631) );
  NAND2_X1 U714 ( .A1(n632), .A2(n631), .ZN(n636) );
  NAND2_X1 U715 ( .A1(G73), .A2(n633), .ZN(n634) );
  XOR2_X1 U716 ( .A(KEYINPUT2), .B(n634), .Z(n635) );
  NOR2_X1 U717 ( .A1(n636), .A2(n635), .ZN(n639) );
  NAND2_X1 U718 ( .A1(n637), .A2(G86), .ZN(n638) );
  NAND2_X1 U719 ( .A1(n639), .A2(n638), .ZN(G305) );
  NAND2_X1 U720 ( .A1(G87), .A2(n640), .ZN(n641) );
  XNOR2_X1 U721 ( .A(n641), .B(KEYINPUT78), .ZN(n648) );
  NAND2_X1 U722 ( .A1(G49), .A2(n642), .ZN(n644) );
  NAND2_X1 U723 ( .A1(G74), .A2(G651), .ZN(n643) );
  NAND2_X1 U724 ( .A1(n644), .A2(n643), .ZN(n645) );
  NOR2_X1 U725 ( .A1(n646), .A2(n645), .ZN(n647) );
  NAND2_X1 U726 ( .A1(n648), .A2(n647), .ZN(G288) );
  XNOR2_X1 U727 ( .A(KEYINPUT19), .B(KEYINPUT79), .ZN(n650) );
  XNOR2_X1 U728 ( .A(G305), .B(G166), .ZN(n649) );
  XNOR2_X1 U729 ( .A(n650), .B(n649), .ZN(n651) );
  XOR2_X1 U730 ( .A(n658), .B(n651), .Z(n652) );
  XNOR2_X1 U731 ( .A(n652), .B(G288), .ZN(n653) );
  XNOR2_X1 U732 ( .A(G290), .B(n653), .ZN(n654) );
  XNOR2_X1 U733 ( .A(G299), .B(n654), .ZN(n897) );
  XNOR2_X1 U734 ( .A(n655), .B(n897), .ZN(n656) );
  NAND2_X1 U735 ( .A1(n656), .A2(G868), .ZN(n660) );
  NAND2_X1 U736 ( .A1(n658), .A2(n657), .ZN(n659) );
  NAND2_X1 U737 ( .A1(n660), .A2(n659), .ZN(G295) );
  NAND2_X1 U738 ( .A1(G2078), .A2(G2084), .ZN(n661) );
  XOR2_X1 U739 ( .A(KEYINPUT20), .B(n661), .Z(n662) );
  NAND2_X1 U740 ( .A1(G2090), .A2(n662), .ZN(n663) );
  XNOR2_X1 U741 ( .A(KEYINPUT21), .B(n663), .ZN(n664) );
  NAND2_X1 U742 ( .A1(n664), .A2(G2072), .ZN(n665) );
  XNOR2_X1 U743 ( .A(KEYINPUT80), .B(n665), .ZN(G158) );
  XNOR2_X1 U744 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U745 ( .A1(G237), .A2(G236), .ZN(n666) );
  NAND2_X1 U746 ( .A1(G69), .A2(n666), .ZN(n667) );
  XNOR2_X1 U747 ( .A(KEYINPUT81), .B(n667), .ZN(n668) );
  NAND2_X1 U748 ( .A1(n668), .A2(G108), .ZN(n819) );
  NAND2_X1 U749 ( .A1(G567), .A2(n819), .ZN(n673) );
  NOR2_X1 U750 ( .A1(G220), .A2(G219), .ZN(n669) );
  XOR2_X1 U751 ( .A(KEYINPUT22), .B(n669), .Z(n670) );
  NOR2_X1 U752 ( .A1(G218), .A2(n670), .ZN(n671) );
  NAND2_X1 U753 ( .A1(G96), .A2(n671), .ZN(n820) );
  NAND2_X1 U754 ( .A1(G2106), .A2(n820), .ZN(n672) );
  NAND2_X1 U755 ( .A1(n673), .A2(n672), .ZN(n831) );
  NAND2_X1 U756 ( .A1(G483), .A2(G661), .ZN(n674) );
  NOR2_X1 U757 ( .A1(n831), .A2(n674), .ZN(n818) );
  NAND2_X1 U758 ( .A1(n818), .A2(G36), .ZN(G176) );
  INV_X1 U759 ( .A(G166), .ZN(G303) );
  XOR2_X1 U760 ( .A(KEYINPUT94), .B(KEYINPUT95), .Z(n681) );
  NAND2_X1 U761 ( .A1(G160), .A2(G40), .ZN(n779) );
  INV_X1 U762 ( .A(n779), .ZN(n675) );
  NOR2_X1 U763 ( .A1(G164), .A2(G1384), .ZN(n780) );
  NAND2_X1 U764 ( .A1(n675), .A2(n780), .ZN(n723) );
  NAND2_X1 U765 ( .A1(G8), .A2(n723), .ZN(n757) );
  NOR2_X1 U766 ( .A1(G1966), .A2(n757), .ZN(n736) );
  NOR2_X1 U767 ( .A1(n779), .A2(G2084), .ZN(n676) );
  AND2_X1 U768 ( .A1(n780), .A2(n676), .ZN(n734) );
  NOR2_X1 U769 ( .A1(n736), .A2(n734), .ZN(n678) );
  INV_X1 U770 ( .A(KEYINPUT93), .ZN(n677) );
  XNOR2_X1 U771 ( .A(n678), .B(n677), .ZN(n679) );
  NAND2_X1 U772 ( .A1(n679), .A2(G8), .ZN(n680) );
  XNOR2_X1 U773 ( .A(n681), .B(n680), .ZN(n682) );
  XNOR2_X1 U774 ( .A(n682), .B(KEYINPUT30), .ZN(n683) );
  NOR2_X1 U775 ( .A1(n683), .A2(G168), .ZN(n688) );
  INV_X1 U776 ( .A(n723), .ZN(n703) );
  NOR2_X1 U777 ( .A1(n703), .A2(G1961), .ZN(n684) );
  XNOR2_X1 U778 ( .A(n684), .B(KEYINPUT89), .ZN(n686) );
  XNOR2_X1 U779 ( .A(KEYINPUT25), .B(G2078), .ZN(n993) );
  NAND2_X1 U780 ( .A1(n703), .A2(n993), .ZN(n685) );
  NAND2_X1 U781 ( .A1(n686), .A2(n685), .ZN(n717) );
  NOR2_X1 U782 ( .A1(G171), .A2(n717), .ZN(n687) );
  NOR2_X1 U783 ( .A1(n688), .A2(n687), .ZN(n690) );
  XNOR2_X1 U784 ( .A(n690), .B(n689), .ZN(n721) );
  AND2_X1 U785 ( .A1(n703), .A2(G2067), .ZN(n692) );
  INV_X1 U786 ( .A(G1348), .ZN(n934) );
  NOR2_X1 U787 ( .A1(n703), .A2(n934), .ZN(n691) );
  NOR2_X1 U788 ( .A1(n692), .A2(n691), .ZN(n698) );
  NOR2_X1 U789 ( .A1(n968), .A2(n698), .ZN(n702) );
  NAND2_X1 U790 ( .A1(n703), .A2(G1996), .ZN(n694) );
  INV_X1 U791 ( .A(KEYINPUT26), .ZN(n693) );
  XOR2_X1 U792 ( .A(n694), .B(n693), .Z(n696) );
  NAND2_X1 U793 ( .A1(n723), .A2(G1341), .ZN(n695) );
  NAND2_X1 U794 ( .A1(n696), .A2(n695), .ZN(n697) );
  NOR2_X1 U795 ( .A1(n983), .A2(n697), .ZN(n700) );
  AND2_X1 U796 ( .A1(n698), .A2(n968), .ZN(n699) );
  NOR2_X1 U797 ( .A1(n700), .A2(n699), .ZN(n701) );
  NOR2_X1 U798 ( .A1(n702), .A2(n701), .ZN(n710) );
  AND2_X1 U799 ( .A1(n703), .A2(G2072), .ZN(n705) );
  XNOR2_X1 U800 ( .A(KEYINPUT90), .B(KEYINPUT27), .ZN(n704) );
  XNOR2_X1 U801 ( .A(n705), .B(n704), .ZN(n707) );
  NAND2_X1 U802 ( .A1(n723), .A2(G1956), .ZN(n706) );
  NAND2_X1 U803 ( .A1(n707), .A2(n706), .ZN(n711) );
  XNOR2_X1 U804 ( .A(n708), .B(KEYINPUT92), .ZN(n709) );
  NOR2_X1 U805 ( .A1(n710), .A2(n709), .ZN(n715) );
  NAND2_X1 U806 ( .A1(n711), .A2(G299), .ZN(n712) );
  XNOR2_X1 U807 ( .A(n712), .B(KEYINPUT91), .ZN(n713) );
  XNOR2_X1 U808 ( .A(n713), .B(KEYINPUT28), .ZN(n714) );
  XNOR2_X1 U809 ( .A(n716), .B(KEYINPUT29), .ZN(n719) );
  NAND2_X1 U810 ( .A1(G171), .A2(n717), .ZN(n718) );
  NAND2_X1 U811 ( .A1(n719), .A2(n718), .ZN(n720) );
  NAND2_X1 U812 ( .A1(n721), .A2(n720), .ZN(n737) );
  AND2_X1 U813 ( .A1(G286), .A2(G8), .ZN(n722) );
  NAND2_X1 U814 ( .A1(n737), .A2(n722), .ZN(n731) );
  INV_X1 U815 ( .A(G8), .ZN(n729) );
  NOR2_X1 U816 ( .A1(G2090), .A2(n723), .ZN(n724) );
  XNOR2_X1 U817 ( .A(KEYINPUT97), .B(n724), .ZN(n727) );
  NOR2_X1 U818 ( .A1(G1971), .A2(n757), .ZN(n725) );
  NOR2_X1 U819 ( .A1(G166), .A2(n725), .ZN(n726) );
  NAND2_X1 U820 ( .A1(n727), .A2(n726), .ZN(n728) );
  OR2_X1 U821 ( .A1(n729), .A2(n728), .ZN(n730) );
  AND2_X1 U822 ( .A1(n731), .A2(n730), .ZN(n733) );
  AND2_X1 U823 ( .A1(G8), .A2(n734), .ZN(n735) );
  AND2_X1 U824 ( .A1(n737), .A2(n513), .ZN(n739) );
  NAND2_X1 U825 ( .A1(G1976), .A2(G288), .ZN(n962) );
  AND2_X1 U826 ( .A1(n753), .A2(n962), .ZN(n740) );
  NAND2_X1 U827 ( .A1(n752), .A2(n740), .ZN(n744) );
  INV_X1 U828 ( .A(n962), .ZN(n742) );
  NOR2_X1 U829 ( .A1(G1976), .A2(G288), .ZN(n747) );
  NOR2_X1 U830 ( .A1(G1971), .A2(G303), .ZN(n741) );
  NOR2_X1 U831 ( .A1(n747), .A2(n741), .ZN(n963) );
  OR2_X1 U832 ( .A1(n742), .A2(n963), .ZN(n743) );
  AND2_X1 U833 ( .A1(n744), .A2(n743), .ZN(n745) );
  NOR2_X1 U834 ( .A1(n745), .A2(n757), .ZN(n746) );
  NAND2_X1 U835 ( .A1(n747), .A2(KEYINPUT33), .ZN(n748) );
  XOR2_X1 U836 ( .A(G1981), .B(G305), .Z(n977) );
  NAND2_X1 U837 ( .A1(n514), .A2(n511), .ZN(n749) );
  XNOR2_X1 U838 ( .A(n749), .B(KEYINPUT99), .ZN(n805) );
  NOR2_X1 U839 ( .A1(G1981), .A2(G305), .ZN(n750) );
  XOR2_X1 U840 ( .A(n750), .B(KEYINPUT24), .Z(n751) );
  OR2_X1 U841 ( .A1(n757), .A2(n751), .ZN(n761) );
  NAND2_X1 U842 ( .A1(n753), .A2(n752), .ZN(n756) );
  NOR2_X1 U843 ( .A1(G2090), .A2(G303), .ZN(n754) );
  NAND2_X1 U844 ( .A1(G8), .A2(n754), .ZN(n755) );
  NAND2_X1 U845 ( .A1(n756), .A2(n755), .ZN(n758) );
  NAND2_X1 U846 ( .A1(n758), .A2(n757), .ZN(n759) );
  XNOR2_X1 U847 ( .A(n759), .B(KEYINPUT100), .ZN(n760) );
  NAND2_X1 U848 ( .A1(n761), .A2(n760), .ZN(n803) );
  XOR2_X1 U849 ( .A(KEYINPUT86), .B(KEYINPUT38), .Z(n763) );
  NAND2_X1 U850 ( .A1(G105), .A2(n866), .ZN(n762) );
  XNOR2_X1 U851 ( .A(n763), .B(n762), .ZN(n767) );
  NAND2_X1 U852 ( .A1(G117), .A2(n874), .ZN(n765) );
  NAND2_X1 U853 ( .A1(G141), .A2(n867), .ZN(n764) );
  NAND2_X1 U854 ( .A1(n765), .A2(n764), .ZN(n766) );
  NOR2_X1 U855 ( .A1(n767), .A2(n766), .ZN(n769) );
  NAND2_X1 U856 ( .A1(n871), .A2(G129), .ZN(n768) );
  NAND2_X1 U857 ( .A1(n769), .A2(n768), .ZN(n882) );
  NOR2_X1 U858 ( .A1(G1996), .A2(n882), .ZN(n922) );
  NAND2_X1 U859 ( .A1(G1996), .A2(n882), .ZN(n770) );
  XNOR2_X1 U860 ( .A(n770), .B(KEYINPUT87), .ZN(n778) );
  INV_X1 U861 ( .A(G1991), .ZN(n991) );
  NAND2_X1 U862 ( .A1(G95), .A2(n866), .ZN(n772) );
  NAND2_X1 U863 ( .A1(G107), .A2(n874), .ZN(n771) );
  NAND2_X1 U864 ( .A1(n772), .A2(n771), .ZN(n776) );
  NAND2_X1 U865 ( .A1(G119), .A2(n871), .ZN(n774) );
  NAND2_X1 U866 ( .A1(G131), .A2(n867), .ZN(n773) );
  NAND2_X1 U867 ( .A1(n774), .A2(n773), .ZN(n775) );
  NOR2_X1 U868 ( .A1(n776), .A2(n775), .ZN(n888) );
  NOR2_X1 U869 ( .A1(n991), .A2(n888), .ZN(n777) );
  NOR2_X1 U870 ( .A1(n778), .A2(n777), .ZN(n924) );
  NOR2_X1 U871 ( .A1(n780), .A2(n779), .ZN(n806) );
  XOR2_X1 U872 ( .A(KEYINPUT88), .B(n806), .Z(n781) );
  NOR2_X1 U873 ( .A1(n924), .A2(n781), .ZN(n808) );
  AND2_X1 U874 ( .A1(n991), .A2(n888), .ZN(n909) );
  NOR2_X1 U875 ( .A1(G1986), .A2(G290), .ZN(n782) );
  XOR2_X1 U876 ( .A(n782), .B(KEYINPUT101), .Z(n783) );
  NOR2_X1 U877 ( .A1(n909), .A2(n783), .ZN(n784) );
  NOR2_X1 U878 ( .A1(n808), .A2(n784), .ZN(n785) );
  NOR2_X1 U879 ( .A1(n922), .A2(n785), .ZN(n786) );
  XNOR2_X1 U880 ( .A(n786), .B(KEYINPUT39), .ZN(n798) );
  XNOR2_X1 U881 ( .A(G2067), .B(KEYINPUT37), .ZN(n799) );
  NAND2_X1 U882 ( .A1(G104), .A2(n866), .ZN(n788) );
  NAND2_X1 U883 ( .A1(G140), .A2(n867), .ZN(n787) );
  NAND2_X1 U884 ( .A1(n788), .A2(n787), .ZN(n789) );
  XNOR2_X1 U885 ( .A(KEYINPUT34), .B(n789), .ZN(n795) );
  NAND2_X1 U886 ( .A1(n871), .A2(G128), .ZN(n790) );
  XNOR2_X1 U887 ( .A(n790), .B(KEYINPUT84), .ZN(n792) );
  NAND2_X1 U888 ( .A1(G116), .A2(n874), .ZN(n791) );
  NAND2_X1 U889 ( .A1(n792), .A2(n791), .ZN(n793) );
  XOR2_X1 U890 ( .A(n793), .B(KEYINPUT35), .Z(n794) );
  NOR2_X1 U891 ( .A1(n795), .A2(n794), .ZN(n796) );
  XOR2_X1 U892 ( .A(KEYINPUT36), .B(n796), .Z(n797) );
  XNOR2_X1 U893 ( .A(KEYINPUT85), .B(n797), .ZN(n887) );
  OR2_X1 U894 ( .A1(n799), .A2(n887), .ZN(n910) );
  NAND2_X1 U895 ( .A1(n798), .A2(n910), .ZN(n800) );
  NAND2_X1 U896 ( .A1(n799), .A2(n887), .ZN(n919) );
  NAND2_X1 U897 ( .A1(n800), .A2(n919), .ZN(n801) );
  NAND2_X1 U898 ( .A1(n801), .A2(n806), .ZN(n811) );
  INV_X1 U899 ( .A(n811), .ZN(n802) );
  OR2_X1 U900 ( .A1(n803), .A2(n802), .ZN(n804) );
  NOR2_X1 U901 ( .A1(n805), .A2(n804), .ZN(n813) );
  XOR2_X1 U902 ( .A(G1986), .B(G290), .Z(n972) );
  NAND2_X1 U903 ( .A1(n972), .A2(n910), .ZN(n807) );
  AND2_X1 U904 ( .A1(n807), .A2(n806), .ZN(n809) );
  OR2_X1 U905 ( .A1(n809), .A2(n808), .ZN(n810) );
  AND2_X1 U906 ( .A1(n811), .A2(n810), .ZN(n812) );
  NOR2_X1 U907 ( .A1(n813), .A2(n812), .ZN(n814) );
  XNOR2_X1 U908 ( .A(n814), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U909 ( .A1(G2106), .A2(n815), .ZN(G217) );
  AND2_X1 U910 ( .A1(G15), .A2(G2), .ZN(n816) );
  NAND2_X1 U911 ( .A1(G661), .A2(n816), .ZN(G259) );
  NAND2_X1 U912 ( .A1(G3), .A2(G1), .ZN(n817) );
  NAND2_X1 U913 ( .A1(n818), .A2(n817), .ZN(G188) );
  XNOR2_X1 U914 ( .A(G69), .B(KEYINPUT103), .ZN(G235) );
  INV_X1 U916 ( .A(G108), .ZN(G238) );
  INV_X1 U917 ( .A(G96), .ZN(G221) );
  NOR2_X1 U918 ( .A1(n820), .A2(n819), .ZN(G325) );
  INV_X1 U919 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U920 ( .A(G1348), .B(G2454), .ZN(n821) );
  XNOR2_X1 U921 ( .A(n821), .B(G2430), .ZN(n822) );
  XNOR2_X1 U922 ( .A(n822), .B(G1341), .ZN(n828) );
  XOR2_X1 U923 ( .A(G2443), .B(G2427), .Z(n824) );
  XNOR2_X1 U924 ( .A(G2438), .B(G2446), .ZN(n823) );
  XNOR2_X1 U925 ( .A(n824), .B(n823), .ZN(n826) );
  XOR2_X1 U926 ( .A(G2451), .B(G2435), .Z(n825) );
  XNOR2_X1 U927 ( .A(n826), .B(n825), .ZN(n827) );
  XNOR2_X1 U928 ( .A(n828), .B(n827), .ZN(n829) );
  NAND2_X1 U929 ( .A1(n829), .A2(G14), .ZN(n830) );
  XOR2_X1 U930 ( .A(KEYINPUT102), .B(n830), .Z(G401) );
  XOR2_X1 U931 ( .A(KEYINPUT104), .B(n831), .Z(G319) );
  XOR2_X1 U932 ( .A(G1986), .B(G1966), .Z(n833) );
  XNOR2_X1 U933 ( .A(G1961), .B(G1956), .ZN(n832) );
  XNOR2_X1 U934 ( .A(n833), .B(n832), .ZN(n834) );
  XOR2_X1 U935 ( .A(n834), .B(G2474), .Z(n836) );
  XNOR2_X1 U936 ( .A(G1971), .B(G1976), .ZN(n835) );
  XNOR2_X1 U937 ( .A(n836), .B(n835), .ZN(n840) );
  XOR2_X1 U938 ( .A(KEYINPUT41), .B(G1991), .Z(n838) );
  XNOR2_X1 U939 ( .A(G1981), .B(G1996), .ZN(n837) );
  XNOR2_X1 U940 ( .A(n838), .B(n837), .ZN(n839) );
  XNOR2_X1 U941 ( .A(n840), .B(n839), .ZN(G229) );
  XOR2_X1 U942 ( .A(KEYINPUT105), .B(G2084), .Z(n842) );
  XNOR2_X1 U943 ( .A(G2090), .B(G2078), .ZN(n841) );
  XNOR2_X1 U944 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U945 ( .A(n843), .B(G2100), .Z(n845) );
  XNOR2_X1 U946 ( .A(G2067), .B(G2072), .ZN(n844) );
  XNOR2_X1 U947 ( .A(n845), .B(n844), .ZN(n849) );
  XOR2_X1 U948 ( .A(G2096), .B(G2678), .Z(n847) );
  XNOR2_X1 U949 ( .A(KEYINPUT42), .B(KEYINPUT43), .ZN(n846) );
  XNOR2_X1 U950 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U951 ( .A(n849), .B(n848), .Z(G227) );
  NAND2_X1 U952 ( .A1(G124), .A2(n871), .ZN(n850) );
  XNOR2_X1 U953 ( .A(n850), .B(KEYINPUT106), .ZN(n851) );
  XNOR2_X1 U954 ( .A(n851), .B(KEYINPUT44), .ZN(n853) );
  NAND2_X1 U955 ( .A1(G112), .A2(n874), .ZN(n852) );
  NAND2_X1 U956 ( .A1(n853), .A2(n852), .ZN(n857) );
  NAND2_X1 U957 ( .A1(G100), .A2(n866), .ZN(n855) );
  NAND2_X1 U958 ( .A1(G136), .A2(n867), .ZN(n854) );
  NAND2_X1 U959 ( .A1(n855), .A2(n854), .ZN(n856) );
  NOR2_X1 U960 ( .A1(n857), .A2(n856), .ZN(G162) );
  NAND2_X1 U961 ( .A1(G127), .A2(n871), .ZN(n859) );
  NAND2_X1 U962 ( .A1(G115), .A2(n874), .ZN(n858) );
  NAND2_X1 U963 ( .A1(n859), .A2(n858), .ZN(n860) );
  XNOR2_X1 U964 ( .A(n860), .B(KEYINPUT47), .ZN(n862) );
  NAND2_X1 U965 ( .A1(G139), .A2(n867), .ZN(n861) );
  NAND2_X1 U966 ( .A1(n862), .A2(n861), .ZN(n865) );
  NAND2_X1 U967 ( .A1(n866), .A2(G103), .ZN(n863) );
  XOR2_X1 U968 ( .A(KEYINPUT108), .B(n863), .Z(n864) );
  NOR2_X1 U969 ( .A1(n865), .A2(n864), .ZN(n912) );
  XNOR2_X1 U970 ( .A(n912), .B(G162), .ZN(n879) );
  NAND2_X1 U971 ( .A1(G106), .A2(n866), .ZN(n869) );
  NAND2_X1 U972 ( .A1(G142), .A2(n867), .ZN(n868) );
  NAND2_X1 U973 ( .A1(n869), .A2(n868), .ZN(n870) );
  XNOR2_X1 U974 ( .A(n870), .B(KEYINPUT45), .ZN(n873) );
  NAND2_X1 U975 ( .A1(G130), .A2(n871), .ZN(n872) );
  NAND2_X1 U976 ( .A1(n873), .A2(n872), .ZN(n877) );
  NAND2_X1 U977 ( .A1(G118), .A2(n874), .ZN(n875) );
  XNOR2_X1 U978 ( .A(KEYINPUT107), .B(n875), .ZN(n876) );
  NOR2_X1 U979 ( .A1(n877), .A2(n876), .ZN(n878) );
  XNOR2_X1 U980 ( .A(n879), .B(n878), .ZN(n886) );
  XOR2_X1 U981 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n881) );
  XNOR2_X1 U982 ( .A(KEYINPUT110), .B(KEYINPUT109), .ZN(n880) );
  XNOR2_X1 U983 ( .A(n881), .B(n880), .ZN(n883) );
  XNOR2_X1 U984 ( .A(n883), .B(n882), .ZN(n884) );
  XNOR2_X1 U985 ( .A(n884), .B(n906), .ZN(n885) );
  XOR2_X1 U986 ( .A(n886), .B(n885), .Z(n890) );
  XOR2_X1 U987 ( .A(n888), .B(n887), .Z(n889) );
  XNOR2_X1 U988 ( .A(n890), .B(n889), .ZN(n892) );
  XNOR2_X1 U989 ( .A(G160), .B(G164), .ZN(n891) );
  XNOR2_X1 U990 ( .A(n892), .B(n891), .ZN(n893) );
  NOR2_X1 U991 ( .A1(G37), .A2(n893), .ZN(G395) );
  XNOR2_X1 U992 ( .A(n983), .B(n968), .ZN(n895) );
  XNOR2_X1 U993 ( .A(G286), .B(G171), .ZN(n894) );
  XNOR2_X1 U994 ( .A(n895), .B(n894), .ZN(n896) );
  XOR2_X1 U995 ( .A(n897), .B(n896), .Z(n898) );
  NOR2_X1 U996 ( .A1(G37), .A2(n898), .ZN(n899) );
  XOR2_X1 U997 ( .A(KEYINPUT111), .B(n899), .Z(G397) );
  NOR2_X1 U998 ( .A1(G229), .A2(G227), .ZN(n900) );
  XOR2_X1 U999 ( .A(KEYINPUT49), .B(n900), .Z(n901) );
  NAND2_X1 U1000 ( .A1(G319), .A2(n901), .ZN(n902) );
  NOR2_X1 U1001 ( .A1(G401), .A2(n902), .ZN(n905) );
  NOR2_X1 U1002 ( .A1(G395), .A2(G397), .ZN(n903) );
  XNOR2_X1 U1003 ( .A(n903), .B(KEYINPUT112), .ZN(n904) );
  NAND2_X1 U1004 ( .A1(n905), .A2(n904), .ZN(G225) );
  INV_X1 U1005 ( .A(G225), .ZN(G308) );
  INV_X1 U1006 ( .A(KEYINPUT55), .ZN(n931) );
  XNOR2_X1 U1007 ( .A(KEYINPUT52), .B(KEYINPUT114), .ZN(n929) );
  XNOR2_X1 U1008 ( .A(G160), .B(G2084), .ZN(n907) );
  NAND2_X1 U1009 ( .A1(n907), .A2(n906), .ZN(n908) );
  NOR2_X1 U1010 ( .A1(n909), .A2(n908), .ZN(n911) );
  NAND2_X1 U1011 ( .A1(n911), .A2(n910), .ZN(n918) );
  XNOR2_X1 U1012 ( .A(G2072), .B(n912), .ZN(n914) );
  XNOR2_X1 U1013 ( .A(G164), .B(G2078), .ZN(n913) );
  NAND2_X1 U1014 ( .A1(n914), .A2(n913), .ZN(n915) );
  XOR2_X1 U1015 ( .A(KEYINPUT113), .B(n915), .Z(n916) );
  XNOR2_X1 U1016 ( .A(KEYINPUT50), .B(n916), .ZN(n917) );
  NOR2_X1 U1017 ( .A1(n918), .A2(n917), .ZN(n920) );
  NAND2_X1 U1018 ( .A1(n920), .A2(n919), .ZN(n927) );
  XOR2_X1 U1019 ( .A(G2090), .B(G162), .Z(n921) );
  NOR2_X1 U1020 ( .A1(n922), .A2(n921), .ZN(n923) );
  XOR2_X1 U1021 ( .A(KEYINPUT51), .B(n923), .Z(n925) );
  NAND2_X1 U1022 ( .A1(n925), .A2(n924), .ZN(n926) );
  NOR2_X1 U1023 ( .A1(n927), .A2(n926), .ZN(n928) );
  XNOR2_X1 U1024 ( .A(n929), .B(n928), .ZN(n930) );
  NAND2_X1 U1025 ( .A1(n931), .A2(n930), .ZN(n932) );
  NAND2_X1 U1026 ( .A1(n932), .A2(G29), .ZN(n933) );
  XNOR2_X1 U1027 ( .A(n933), .B(KEYINPUT115), .ZN(n960) );
  XOR2_X1 U1028 ( .A(G16), .B(KEYINPUT124), .Z(n957) );
  XNOR2_X1 U1029 ( .A(KEYINPUT59), .B(G4), .ZN(n935) );
  XNOR2_X1 U1030 ( .A(n935), .B(n934), .ZN(n937) );
  XNOR2_X1 U1031 ( .A(G6), .B(G1981), .ZN(n936) );
  NOR2_X1 U1032 ( .A1(n937), .A2(n936), .ZN(n941) );
  XNOR2_X1 U1033 ( .A(G1341), .B(G19), .ZN(n939) );
  XNOR2_X1 U1034 ( .A(G1956), .B(G20), .ZN(n938) );
  NOR2_X1 U1035 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1036 ( .A1(n941), .A2(n940), .ZN(n942) );
  XNOR2_X1 U1037 ( .A(n942), .B(KEYINPUT125), .ZN(n943) );
  XNOR2_X1 U1038 ( .A(KEYINPUT60), .B(n943), .ZN(n947) );
  XNOR2_X1 U1039 ( .A(G1961), .B(G5), .ZN(n945) );
  XNOR2_X1 U1040 ( .A(G1966), .B(G21), .ZN(n944) );
  NOR2_X1 U1041 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1042 ( .A1(n947), .A2(n946), .ZN(n954) );
  XNOR2_X1 U1043 ( .A(G1971), .B(G22), .ZN(n949) );
  XNOR2_X1 U1044 ( .A(G23), .B(G1976), .ZN(n948) );
  NOR2_X1 U1045 ( .A1(n949), .A2(n948), .ZN(n951) );
  XOR2_X1 U1046 ( .A(G1986), .B(G24), .Z(n950) );
  NAND2_X1 U1047 ( .A1(n951), .A2(n950), .ZN(n952) );
  XNOR2_X1 U1048 ( .A(KEYINPUT58), .B(n952), .ZN(n953) );
  NOR2_X1 U1049 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1050 ( .A(n955), .B(KEYINPUT61), .ZN(n956) );
  NAND2_X1 U1051 ( .A1(n957), .A2(n956), .ZN(n958) );
  NAND2_X1 U1052 ( .A1(G11), .A2(n958), .ZN(n959) );
  NOR2_X1 U1053 ( .A1(n960), .A2(n959), .ZN(n1015) );
  XOR2_X1 U1054 ( .A(G16), .B(KEYINPUT56), .Z(n988) );
  INV_X1 U1055 ( .A(G1971), .ZN(n961) );
  NOR2_X1 U1056 ( .A1(G166), .A2(n961), .ZN(n965) );
  NAND2_X1 U1057 ( .A1(n963), .A2(n962), .ZN(n964) );
  NOR2_X1 U1058 ( .A1(n965), .A2(n964), .ZN(n967) );
  XOR2_X1 U1059 ( .A(G1956), .B(G299), .Z(n966) );
  NAND2_X1 U1060 ( .A1(n967), .A2(n966), .ZN(n975) );
  XNOR2_X1 U1061 ( .A(n968), .B(G1348), .ZN(n970) );
  XNOR2_X1 U1062 ( .A(G171), .B(G1961), .ZN(n969) );
  NAND2_X1 U1063 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1064 ( .A(KEYINPUT121), .B(n971), .ZN(n973) );
  NAND2_X1 U1065 ( .A1(n973), .A2(n972), .ZN(n974) );
  NOR2_X1 U1066 ( .A1(n975), .A2(n974), .ZN(n976) );
  XNOR2_X1 U1067 ( .A(KEYINPUT122), .B(n976), .ZN(n982) );
  XNOR2_X1 U1068 ( .A(G168), .B(G1966), .ZN(n978) );
  NAND2_X1 U1069 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1070 ( .A(n979), .B(KEYINPUT120), .ZN(n980) );
  XNOR2_X1 U1071 ( .A(KEYINPUT57), .B(n980), .ZN(n981) );
  NAND2_X1 U1072 ( .A1(n982), .A2(n981), .ZN(n985) );
  XNOR2_X1 U1073 ( .A(G1341), .B(n983), .ZN(n984) );
  NOR2_X1 U1074 ( .A1(n985), .A2(n984), .ZN(n986) );
  XOR2_X1 U1075 ( .A(KEYINPUT123), .B(n986), .Z(n987) );
  NOR2_X1 U1076 ( .A1(n988), .A2(n987), .ZN(n1013) );
  XNOR2_X1 U1077 ( .A(G2067), .B(G26), .ZN(n990) );
  XNOR2_X1 U1078 ( .A(G33), .B(G2072), .ZN(n989) );
  NOR2_X1 U1079 ( .A1(n990), .A2(n989), .ZN(n1001) );
  XNOR2_X1 U1080 ( .A(G25), .B(n991), .ZN(n992) );
  NAND2_X1 U1081 ( .A1(n992), .A2(G28), .ZN(n999) );
  XNOR2_X1 U1082 ( .A(n993), .B(G27), .ZN(n996) );
  XNOR2_X1 U1083 ( .A(G1996), .B(G32), .ZN(n994) );
  XNOR2_X1 U1084 ( .A(n994), .B(KEYINPUT117), .ZN(n995) );
  NAND2_X1 U1085 ( .A1(n996), .A2(n995), .ZN(n997) );
  XNOR2_X1 U1086 ( .A(n997), .B(KEYINPUT118), .ZN(n998) );
  NOR2_X1 U1087 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1088 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1089 ( .A(KEYINPUT119), .B(n1002), .ZN(n1003) );
  XOR2_X1 U1090 ( .A(KEYINPUT53), .B(n1003), .Z(n1006) );
  XOR2_X1 U1091 ( .A(KEYINPUT54), .B(G34), .Z(n1004) );
  XNOR2_X1 U1092 ( .A(G2084), .B(n1004), .ZN(n1005) );
  NAND2_X1 U1093 ( .A1(n1006), .A2(n1005), .ZN(n1009) );
  XNOR2_X1 U1094 ( .A(KEYINPUT116), .B(G2090), .ZN(n1007) );
  XNOR2_X1 U1095 ( .A(G35), .B(n1007), .ZN(n1008) );
  NOR2_X1 U1096 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XOR2_X1 U1097 ( .A(KEYINPUT55), .B(n1010), .Z(n1011) );
  NOR2_X1 U1098 ( .A1(G29), .A2(n1011), .ZN(n1012) );
  NOR2_X1 U1099 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1100 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1101 ( .A(KEYINPUT62), .B(n1016), .ZN(n1017) );
  XNOR2_X1 U1102 ( .A(KEYINPUT126), .B(n1017), .ZN(G150) );
  INV_X1 U1103 ( .A(G150), .ZN(G311) );
endmodule

