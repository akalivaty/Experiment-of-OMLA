//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 1 0 0 0 0 1 1 0 1 0 0 1 1 1 0 0 0 0 1 1 1 0 1 1 1 1 0 0 1 0 0 0 0 1 1 1 1 1 1 0 1 0 1 1 0 1 1 0 0 1 0 0 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:50 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1260, new_n1261, new_n1262, new_n1263;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(G13), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XOR2_X1   g0009(.A(new_n209), .B(KEYINPUT0), .Z(new_n210));
  AOI22_X1  g0010(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G87), .A2(G250), .ZN(new_n212));
  INV_X1    g0012(.A(G97), .ZN(new_n213));
  INV_X1    g0013(.A(G257), .ZN(new_n214));
  OAI211_X1 g0014(.A(new_n211), .B(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(KEYINPUT64), .ZN(new_n216));
  AOI21_X1  g0016(.A(new_n216), .B1(G50), .B2(G226), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n215), .A2(KEYINPUT64), .ZN(new_n218));
  INV_X1    g0018(.A(G68), .ZN(new_n219));
  INV_X1    g0019(.A(G238), .ZN(new_n220));
  OAI211_X1 g0020(.A(new_n217), .B(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  AOI21_X1  g0021(.A(new_n221), .B1(G116), .B2(G270), .ZN(new_n222));
  INV_X1    g0022(.A(G77), .ZN(new_n223));
  INV_X1    g0023(.A(G244), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n222), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n225), .B1(new_n203), .B2(new_n204), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT1), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n228), .A2(new_n204), .ZN(new_n229));
  OAI21_X1  g0029(.A(G50), .B1(G58), .B2(G68), .ZN(new_n230));
  INV_X1    g0030(.A(new_n230), .ZN(new_n231));
  AOI211_X1 g0031(.A(new_n210), .B(new_n227), .C1(new_n229), .C2(new_n231), .ZN(G361));
  XNOR2_X1  g0032(.A(KEYINPUT2), .B(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT65), .B(G250), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n236), .B(new_n240), .ZN(G358));
  XOR2_X1   g0041(.A(G68), .B(G77), .Z(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G58), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G87), .B(G97), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n244), .B(new_n247), .Z(G351));
  XNOR2_X1  g0048(.A(KEYINPUT3), .B(G33), .ZN(new_n249));
  INV_X1    g0049(.A(G1698), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(G222), .ZN(new_n251));
  INV_X1    g0051(.A(G223), .ZN(new_n252));
  OAI211_X1 g0052(.A(new_n249), .B(new_n251), .C1(new_n252), .C2(new_n250), .ZN(new_n253));
  INV_X1    g0053(.A(G33), .ZN(new_n254));
  INV_X1    g0054(.A(G41), .ZN(new_n255));
  OAI211_X1 g0055(.A(G1), .B(G13), .C1(new_n254), .C2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  OAI211_X1 g0057(.A(new_n253), .B(new_n257), .C1(G77), .C2(new_n249), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n203), .B1(G41), .B2(G45), .ZN(new_n259));
  INV_X1    g0059(.A(G274), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G226), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n256), .A2(new_n259), .ZN(new_n264));
  OAI211_X1 g0064(.A(new_n258), .B(new_n262), .C1(new_n263), .C2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G190), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n267), .B1(G200), .B2(new_n265), .ZN(new_n268));
  NAND3_X1  g0068(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(new_n228), .ZN(new_n270));
  INV_X1    g0070(.A(G150), .ZN(new_n271));
  NOR2_X1   g0071(.A1(G20), .A2(G33), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  NOR3_X1   g0073(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n274));
  OAI22_X1  g0074(.A1(new_n271), .A2(new_n273), .B1(new_n274), .B2(new_n204), .ZN(new_n275));
  XNOR2_X1  g0075(.A(KEYINPUT8), .B(G58), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n204), .A2(G33), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n270), .B1(new_n275), .B2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT66), .ZN(new_n280));
  XNOR2_X1  g0080(.A(new_n279), .B(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n203), .A2(G13), .A3(G20), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n282), .A2(G50), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n203), .A2(G20), .ZN(new_n284));
  INV_X1    g0084(.A(new_n270), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n284), .B1(new_n285), .B2(KEYINPUT67), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n286), .B1(KEYINPUT67), .B2(new_n285), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n283), .B1(new_n287), .B2(G50), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n281), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT9), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n281), .A2(KEYINPUT9), .A3(new_n288), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n268), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT10), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n265), .A2(G200), .ZN(new_n295));
  OAI211_X1 g0095(.A(new_n295), .B(KEYINPUT68), .C1(new_n266), .C2(new_n265), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n293), .A2(new_n294), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(new_n294), .ZN(new_n298));
  NAND4_X1  g0098(.A1(new_n298), .A2(new_n268), .A3(new_n291), .A4(new_n292), .ZN(new_n299));
  INV_X1    g0099(.A(G169), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n265), .A2(new_n300), .ZN(new_n301));
  OAI211_X1 g0101(.A(new_n289), .B(new_n301), .C1(G179), .C2(new_n265), .ZN(new_n302));
  AND3_X1   g0102(.A1(new_n297), .A2(new_n299), .A3(new_n302), .ZN(new_n303));
  NOR2_X1   g0103(.A1(G226), .A2(G1698), .ZN(new_n304));
  INV_X1    g0104(.A(G232), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n304), .B1(new_n305), .B2(G1698), .ZN(new_n306));
  AND2_X1   g0106(.A1(new_n306), .A2(new_n249), .ZN(new_n307));
  NAND2_X1  g0107(.A1(G33), .A2(G97), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(KEYINPUT69), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT69), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n310), .A2(G33), .A3(G97), .ZN(new_n311));
  AND2_X1   g0111(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n257), .B1(new_n307), .B2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT13), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n256), .A2(G238), .A3(new_n259), .ZN(new_n315));
  NAND4_X1  g0115(.A1(new_n313), .A2(new_n314), .A3(new_n262), .A4(new_n315), .ZN(new_n316));
  AOI22_X1  g0116(.A1(new_n306), .A2(new_n249), .B1(new_n311), .B2(new_n309), .ZN(new_n317));
  OAI211_X1 g0117(.A(new_n262), .B(new_n315), .C1(new_n317), .C2(new_n256), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(KEYINPUT13), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT70), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n316), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  OR3_X1    g0121(.A1(new_n318), .A2(new_n320), .A3(KEYINPUT13), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n321), .A2(new_n322), .A3(G169), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(KEYINPUT14), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT14), .ZN(new_n325));
  NAND4_X1  g0125(.A1(new_n321), .A2(new_n322), .A3(new_n325), .A4(G169), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n316), .A2(new_n319), .A3(G179), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n324), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n219), .A2(G20), .ZN(new_n329));
  INV_X1    g0129(.A(G50), .ZN(new_n330));
  OAI221_X1 g0130(.A(new_n329), .B1(new_n277), .B2(new_n223), .C1(new_n273), .C2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(new_n270), .ZN(new_n332));
  XNOR2_X1  g0132(.A(new_n332), .B(KEYINPUT11), .ZN(new_n333));
  NOR3_X1   g0133(.A1(new_n329), .A2(G1), .A3(new_n206), .ZN(new_n334));
  XNOR2_X1  g0134(.A(new_n334), .B(KEYINPUT12), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n285), .A2(new_n284), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n335), .B1(G68), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n333), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n328), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n321), .A2(new_n322), .A3(G200), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n316), .A2(new_n319), .A3(G190), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n341), .A2(new_n338), .A3(new_n333), .A4(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(G238), .A2(G1698), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n249), .B(new_n344), .C1(new_n305), .C2(G1698), .ZN(new_n345));
  OAI211_X1 g0145(.A(new_n345), .B(new_n257), .C1(G107), .C2(new_n249), .ZN(new_n346));
  OAI211_X1 g0146(.A(new_n346), .B(new_n262), .C1(new_n224), .C2(new_n264), .ZN(new_n347));
  OR2_X1    g0147(.A1(new_n347), .A2(G179), .ZN(new_n348));
  INV_X1    g0148(.A(new_n276), .ZN(new_n349));
  AOI22_X1  g0149(.A1(new_n349), .A2(new_n272), .B1(G20), .B2(G77), .ZN(new_n350));
  XOR2_X1   g0150(.A(KEYINPUT15), .B(G87), .Z(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n350), .B1(new_n277), .B2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n282), .ZN(new_n354));
  AOI22_X1  g0154(.A1(new_n353), .A2(new_n270), .B1(new_n223), .B2(new_n354), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n355), .B1(new_n223), .B2(new_n336), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n347), .A2(new_n300), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n348), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  AND4_X1   g0158(.A1(new_n303), .A2(new_n340), .A3(new_n343), .A4(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT16), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT7), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n361), .B1(new_n249), .B2(G20), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n254), .A2(KEYINPUT3), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT3), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(G33), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n366), .A2(KEYINPUT7), .A3(new_n204), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n219), .B1(new_n362), .B2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(G58), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n369), .A2(new_n219), .ZN(new_n370));
  NOR2_X1   g0170(.A1(G58), .A2(G68), .ZN(new_n371));
  OAI21_X1  g0171(.A(G20), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n272), .A2(G159), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n360), .B1(new_n368), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(KEYINPUT71), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n362), .A2(new_n367), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n374), .B1(new_n377), .B2(G68), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n285), .B1(new_n378), .B2(KEYINPUT16), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT71), .ZN(new_n380));
  OAI211_X1 g0180(.A(new_n380), .B(new_n360), .C1(new_n368), .C2(new_n374), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n376), .A2(new_n379), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(KEYINPUT72), .ZN(new_n383));
  INV_X1    g0183(.A(G200), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n252), .A2(new_n250), .ZN(new_n385));
  OAI211_X1 g0185(.A(new_n249), .B(new_n385), .C1(G226), .C2(new_n250), .ZN(new_n386));
  NAND2_X1  g0186(.A1(G33), .A2(G87), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(new_n257), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n262), .B1(new_n264), .B2(new_n305), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(KEYINPUT73), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n256), .B1(new_n386), .B2(new_n387), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT73), .ZN(new_n394));
  NOR3_X1   g0194(.A1(new_n393), .A2(new_n394), .A3(new_n390), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n384), .B1(new_n392), .B2(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n389), .A2(new_n266), .A3(new_n391), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n349), .A2(new_n282), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n399), .B1(new_n287), .B2(new_n349), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT72), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n376), .A2(new_n379), .A3(new_n401), .A4(new_n381), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n383), .A2(new_n398), .A3(new_n400), .A4(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT74), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT17), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n403), .A2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  NOR2_X1   g0208(.A1(KEYINPUT74), .A2(KEYINPUT17), .ZN(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n406), .B1(new_n403), .B2(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n383), .A2(new_n400), .A3(new_n402), .ZN(new_n412));
  INV_X1    g0212(.A(new_n395), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n394), .B1(new_n393), .B2(new_n390), .ZN(new_n414));
  AOI21_X1  g0214(.A(G169), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NOR3_X1   g0215(.A1(new_n393), .A2(G179), .A3(new_n390), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  AND3_X1   g0217(.A1(new_n412), .A2(KEYINPUT18), .A3(new_n417), .ZN(new_n418));
  AOI21_X1  g0218(.A(KEYINPUT18), .B1(new_n412), .B2(new_n417), .ZN(new_n419));
  OAI22_X1  g0219(.A1(new_n408), .A2(new_n411), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(new_n420), .ZN(new_n421));
  AND2_X1   g0221(.A1(new_n347), .A2(G200), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n347), .A2(new_n266), .ZN(new_n423));
  OR3_X1    g0223(.A1(new_n356), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n359), .A2(new_n421), .A3(new_n424), .ZN(new_n425));
  OAI211_X1 g0225(.A(new_n203), .B(G45), .C1(new_n255), .C2(KEYINPUT5), .ZN(new_n426));
  XNOR2_X1  g0226(.A(new_n426), .B(KEYINPUT76), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n255), .A2(KEYINPUT5), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n427), .A2(G274), .A3(new_n256), .A4(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(G264), .A2(G1698), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n249), .B(new_n430), .C1(new_n214), .C2(G1698), .ZN(new_n431));
  OAI211_X1 g0231(.A(new_n431), .B(new_n257), .C1(G303), .C2(new_n249), .ZN(new_n432));
  INV_X1    g0232(.A(G45), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n433), .A2(G1), .ZN(new_n434));
  OAI211_X1 g0234(.A(new_n434), .B(KEYINPUT76), .C1(KEYINPUT5), .C2(new_n255), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT76), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n426), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n435), .A2(new_n437), .A3(new_n428), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n438), .A2(G270), .A3(new_n256), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n429), .A2(new_n432), .A3(new_n439), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n206), .A2(G1), .ZN(new_n441));
  INV_X1    g0241(.A(G116), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n441), .A2(G20), .A3(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT78), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n441), .A2(KEYINPUT78), .A3(G20), .A4(new_n442), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n203), .A2(G33), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n285), .A2(G116), .A3(new_n282), .A4(new_n448), .ZN(new_n449));
  AOI22_X1  g0249(.A1(new_n269), .A2(new_n228), .B1(G20), .B2(new_n442), .ZN(new_n450));
  NAND2_X1  g0250(.A1(G33), .A2(G283), .ZN(new_n451));
  OAI211_X1 g0251(.A(new_n451), .B(new_n204), .C1(G33), .C2(new_n213), .ZN(new_n452));
  AND3_X1   g0252(.A1(new_n450), .A2(KEYINPUT20), .A3(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(KEYINPUT20), .B1(new_n450), .B2(new_n452), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n447), .B(new_n449), .C1(new_n453), .C2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT21), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(KEYINPUT80), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n440), .A2(G169), .A3(new_n455), .A4(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n440), .A2(G169), .A3(new_n455), .ZN(new_n459));
  XOR2_X1   g0259(.A(KEYINPUT80), .B(KEYINPUT21), .Z(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n429), .A2(G179), .A3(new_n432), .A4(new_n439), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  AOI21_X1  g0263(.A(KEYINPUT79), .B1(new_n463), .B2(new_n455), .ZN(new_n464));
  INV_X1    g0264(.A(new_n455), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT79), .ZN(new_n466));
  NOR3_X1   g0266(.A1(new_n462), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n458), .B(new_n461), .C1(new_n464), .C2(new_n467), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n363), .A2(new_n365), .A3(new_n204), .A4(G87), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(KEYINPUT22), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT22), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n249), .A2(new_n471), .A3(new_n204), .A4(G87), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n254), .A2(new_n442), .ZN(new_n473));
  AOI22_X1  g0273(.A1(new_n470), .A2(new_n472), .B1(new_n204), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n204), .A2(G107), .ZN(new_n475));
  XNOR2_X1  g0275(.A(new_n475), .B(KEYINPUT23), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT24), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n474), .A2(KEYINPUT24), .A3(new_n476), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n479), .A2(new_n270), .A3(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(G107), .ZN(new_n482));
  OR2_X1    g0282(.A1(KEYINPUT81), .A2(KEYINPUT25), .ZN(new_n483));
  NAND2_X1  g0283(.A1(KEYINPUT81), .A2(KEYINPUT25), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n354), .A2(new_n482), .A3(new_n483), .A4(new_n484), .ZN(new_n485));
  OAI211_X1 g0285(.A(KEYINPUT81), .B(KEYINPUT25), .C1(new_n282), .C2(G107), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n285), .A2(new_n282), .A3(new_n448), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n487), .A2(new_n482), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n481), .A2(new_n485), .A3(new_n486), .A4(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(G250), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(new_n250), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n214), .A2(G1698), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n249), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(G33), .A2(G294), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n496), .A2(KEYINPUT82), .A3(new_n257), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n438), .A2(G264), .A3(new_n256), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n496), .A2(new_n257), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n435), .A2(new_n437), .A3(G274), .A4(new_n428), .ZN(new_n501));
  OAI21_X1  g0301(.A(KEYINPUT82), .B1(new_n501), .B2(new_n257), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n499), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  OAI21_X1  g0303(.A(KEYINPUT83), .B1(new_n503), .B2(new_n300), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n429), .A2(new_n498), .A3(new_n500), .ZN(new_n505));
  INV_X1    g0305(.A(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(G179), .ZN(new_n507));
  AND2_X1   g0307(.A1(new_n497), .A2(new_n498), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n502), .A2(new_n500), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT83), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n510), .A2(new_n511), .A3(G169), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n504), .A2(new_n507), .A3(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n468), .B1(new_n490), .B2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT4), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n515), .B1(new_n366), .B2(new_n224), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n249), .A2(KEYINPUT4), .A3(G244), .A4(new_n250), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n516), .A2(new_n517), .A3(new_n451), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n249), .A2(G250), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n250), .B1(new_n519), .B2(KEYINPUT4), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n257), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n438), .A2(G257), .A3(new_n256), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n521), .A2(new_n429), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(G200), .ZN(new_n524));
  INV_X1    g0324(.A(new_n487), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(G97), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n282), .A2(G97), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n377), .A2(G107), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT75), .ZN(new_n529));
  NAND2_X1  g0329(.A1(KEYINPUT6), .A2(G97), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n529), .B1(new_n530), .B2(G107), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n482), .A2(KEYINPUT75), .A3(KEYINPUT6), .A4(G97), .ZN(new_n532));
  AND2_X1   g0332(.A1(G97), .A2(G107), .ZN(new_n533));
  NOR2_X1   g0333(.A1(G97), .A2(G107), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n531), .B(new_n532), .C1(new_n535), .C2(KEYINPUT6), .ZN(new_n536));
  AOI22_X1  g0336(.A1(new_n536), .A2(G20), .B1(G77), .B2(new_n272), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n528), .A2(new_n537), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n527), .B1(new_n538), .B2(new_n270), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n521), .A2(G190), .A3(new_n429), .A4(new_n522), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n524), .A2(new_n526), .A3(new_n539), .A4(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n523), .A2(new_n300), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n536), .A2(G20), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n272), .A2(G77), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n482), .B1(new_n362), .B2(new_n367), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n270), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(new_n527), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n547), .A2(new_n526), .A3(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(G179), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n521), .A2(new_n550), .A3(new_n429), .A4(new_n522), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n542), .A2(new_n549), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n525), .A2(new_n351), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n352), .A2(new_n354), .ZN(new_n554));
  NOR3_X1   g0354(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n309), .A2(new_n311), .A3(KEYINPUT19), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n555), .B1(new_n556), .B2(new_n204), .ZN(new_n557));
  NOR3_X1   g0357(.A1(new_n366), .A2(G20), .A3(new_n219), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n277), .A2(new_n213), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n559), .A2(KEYINPUT19), .ZN(new_n560));
  NOR3_X1   g0360(.A1(new_n557), .A2(new_n558), .A3(new_n560), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n553), .B(new_n554), .C1(new_n561), .C2(new_n285), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n434), .A2(new_n260), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n491), .B1(new_n433), .B2(G1), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n563), .A2(new_n256), .A3(new_n564), .ZN(new_n565));
  NOR2_X1   g0365(.A1(G238), .A2(G1698), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n566), .B1(new_n224), .B2(G1698), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n473), .B1(new_n567), .B2(new_n249), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n565), .B1(new_n568), .B2(new_n256), .ZN(new_n569));
  INV_X1    g0369(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n550), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n569), .A2(new_n300), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n562), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n525), .A2(G87), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n574), .B(new_n554), .C1(new_n561), .C2(new_n285), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n570), .A2(new_n384), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  OAI211_X1 g0377(.A(G190), .B(new_n565), .C1(new_n568), .C2(new_n256), .ZN(new_n578));
  XNOR2_X1  g0378(.A(new_n578), .B(KEYINPUT77), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n541), .A2(new_n552), .A3(new_n573), .A4(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n508), .A2(new_n509), .A3(new_n266), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n505), .A2(new_n384), .ZN(new_n583));
  AND2_X1   g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n490), .A2(new_n584), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n581), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n440), .A2(G200), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n587), .B(new_n465), .C1(new_n266), .C2(new_n440), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n514), .A2(new_n586), .A3(new_n588), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n425), .A2(new_n589), .ZN(G372));
  OR2_X1    g0390(.A1(new_n418), .A2(new_n419), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n408), .A2(new_n411), .ZN(new_n592));
  INV_X1    g0392(.A(new_n358), .ZN(new_n593));
  AOI22_X1  g0393(.A1(new_n328), .A2(new_n339), .B1(new_n343), .B2(new_n593), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n591), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n595), .A2(new_n299), .A3(new_n297), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(new_n302), .ZN(new_n597));
  INV_X1    g0397(.A(new_n597), .ZN(new_n598));
  AND2_X1   g0398(.A1(new_n562), .A2(new_n572), .ZN(new_n599));
  AOI22_X1  g0399(.A1(new_n599), .A2(new_n571), .B1(new_n577), .B2(new_n579), .ZN(new_n600));
  INV_X1    g0400(.A(new_n552), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(KEYINPUT26), .ZN(new_n603));
  XOR2_X1   g0403(.A(new_n573), .B(KEYINPUT84), .Z(new_n604));
  AND3_X1   g0404(.A1(new_n474), .A2(KEYINPUT24), .A3(new_n476), .ZN(new_n605));
  AOI21_X1  g0405(.A(KEYINPUT24), .B1(new_n474), .B2(new_n476), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n488), .B1(new_n607), .B2(new_n270), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n582), .A2(new_n583), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n608), .A2(new_n485), .A3(new_n609), .A4(new_n486), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n610), .A2(new_n600), .A3(new_n552), .A4(new_n541), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n603), .B(new_n604), .C1(new_n514), .C2(new_n611), .ZN(new_n612));
  XOR2_X1   g0412(.A(KEYINPUT85), .B(KEYINPUT26), .Z(new_n613));
  NOR2_X1   g0413(.A1(new_n602), .A2(new_n613), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n598), .B1(new_n425), .B2(new_n615), .ZN(G369));
  NAND2_X1  g0416(.A1(new_n513), .A2(new_n490), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n441), .A2(new_n204), .ZN(new_n618));
  OR2_X1    g0418(.A1(new_n618), .A2(KEYINPUT27), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(KEYINPUT27), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n619), .A2(new_n620), .A3(G213), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(G343), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n490), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n617), .A2(new_n610), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n468), .A2(new_n623), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n513), .A2(new_n490), .A3(new_n624), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n626), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n468), .B1(new_n465), .B2(new_n623), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n462), .A2(new_n465), .ZN(new_n631));
  XNOR2_X1  g0431(.A(new_n631), .B(KEYINPUT79), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n623), .A2(new_n465), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n632), .A2(new_n458), .A3(new_n461), .A4(new_n633), .ZN(new_n634));
  AND3_X1   g0434(.A1(new_n630), .A2(new_n634), .A3(new_n588), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n629), .A2(new_n635), .A3(G330), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n585), .B1(new_n490), .B2(new_n513), .ZN(new_n637));
  INV_X1    g0437(.A(new_n627), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n513), .A2(new_n490), .ZN(new_n639));
  AOI22_X1  g0439(.A1(new_n637), .A2(new_n638), .B1(new_n639), .B2(new_n623), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n636), .A2(new_n640), .ZN(G399));
  NOR2_X1   g0441(.A1(new_n207), .A2(G41), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  AND2_X1   g0443(.A1(new_n555), .A2(new_n442), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n643), .A2(G1), .A3(new_n644), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n645), .B1(new_n230), .B2(new_n643), .ZN(new_n646));
  XNOR2_X1  g0446(.A(new_n646), .B(KEYINPUT28), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n523), .A2(new_n569), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n498), .A2(new_n500), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n462), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT30), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n523), .A2(new_n550), .A3(new_n440), .A4(new_n569), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n653), .B1(new_n506), .B2(new_n654), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n651), .A2(new_n652), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n624), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n514), .A2(new_n586), .A3(new_n588), .A4(new_n623), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n658), .B1(new_n659), .B2(KEYINPUT31), .ZN(new_n660));
  XOR2_X1   g0460(.A(KEYINPUT86), .B(KEYINPUT31), .Z(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n654), .A2(new_n506), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n663), .B1(new_n652), .B2(new_n651), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT87), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n656), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n655), .A2(KEYINPUT87), .ZN(new_n667));
  AOI211_X1 g0467(.A(new_n623), .B(new_n662), .C1(new_n666), .C2(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(G330), .B1(new_n660), .B2(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n604), .B1(new_n514), .B2(new_n611), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n602), .A2(new_n613), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n671), .B1(KEYINPUT26), .B2(new_n602), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n623), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(KEYINPUT29), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT29), .ZN(new_n675));
  OAI211_X1 g0475(.A(new_n675), .B(new_n623), .C1(new_n612), .C2(new_n614), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n669), .A2(new_n674), .A3(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n647), .B1(new_n678), .B2(G1), .ZN(G364));
  NAND3_X1  g0479(.A1(new_n630), .A2(new_n634), .A3(new_n588), .ZN(new_n680));
  INV_X1    g0480(.A(G330), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g0482(.A(new_n682), .B(KEYINPUT88), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n630), .A2(new_n634), .A3(G330), .A4(new_n588), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n206), .A2(G20), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(G45), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n643), .A2(G1), .A3(new_n686), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n683), .A2(new_n684), .A3(new_n687), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n228), .B1(G20), .B2(new_n300), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n384), .A2(G179), .ZN(new_n691));
  XNOR2_X1  g0491(.A(new_n691), .B(KEYINPUT91), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n204), .A2(new_n266), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(G87), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(new_n249), .ZN(new_n697));
  XNOR2_X1  g0497(.A(new_n697), .B(KEYINPUT92), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n204), .A2(G190), .ZN(new_n699));
  NOR2_X1   g0499(.A1(G179), .A2(G200), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(G159), .ZN(new_n703));
  XNOR2_X1  g0503(.A(new_n703), .B(KEYINPUT32), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n692), .A2(new_n699), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n550), .A2(G200), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(new_n699), .ZN(new_n707));
  OAI22_X1  g0507(.A1(new_n705), .A2(new_n482), .B1(new_n223), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n700), .A2(G190), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(G20), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NAND3_X1  g0511(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n712), .A2(new_n266), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  OAI22_X1  g0514(.A1(new_n711), .A2(new_n213), .B1(new_n330), .B2(new_n714), .ZN(new_n715));
  NOR4_X1   g0515(.A1(new_n698), .A2(new_n704), .A3(new_n708), .A4(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n693), .A2(new_n706), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n712), .A2(G190), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  OAI221_X1 g0519(.A(new_n716), .B1(new_n369), .B2(new_n717), .C1(new_n219), .C2(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(KEYINPUT33), .A2(G317), .ZN(new_n721));
  AND2_X1   g0521(.A1(KEYINPUT33), .A2(G317), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n718), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(G311), .ZN(new_n724));
  INV_X1    g0524(.A(G329), .ZN(new_n725));
  OAI221_X1 g0525(.A(new_n723), .B1(new_n724), .B2(new_n707), .C1(new_n725), .C2(new_n701), .ZN(new_n726));
  INV_X1    g0526(.A(G283), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n705), .A2(new_n727), .ZN(new_n728));
  AOI211_X1 g0528(.A(new_n726), .B(new_n728), .C1(G303), .C2(new_n695), .ZN(new_n729));
  INV_X1    g0529(.A(new_n717), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(G322), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n710), .A2(G294), .ZN(new_n732));
  XNOR2_X1  g0532(.A(KEYINPUT93), .B(G326), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n249), .B1(new_n713), .B2(new_n733), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n729), .A2(new_n731), .A3(new_n732), .A4(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n690), .B1(new_n720), .B2(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(G13), .A2(G33), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n738), .A2(G20), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n680), .A2(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n739), .A2(new_n689), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n208), .A2(new_n366), .ZN(new_n742));
  XNOR2_X1  g0542(.A(new_n742), .B(KEYINPUT90), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n743), .B1(G45), .B2(new_n230), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n244), .A2(new_n433), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n208), .A2(new_n249), .ZN(new_n746));
  XOR2_X1   g0546(.A(G355), .B(KEYINPUT89), .Z(new_n747));
  OAI22_X1  g0547(.A1(new_n744), .A2(new_n745), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n208), .A2(G116), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n741), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n687), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n740), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n688), .B1(new_n736), .B2(new_n752), .ZN(G396));
  NAND2_X1  g0553(.A1(new_n356), .A2(new_n624), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n424), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(new_n358), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n593), .A2(new_n623), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n758), .B1(new_n615), .B2(new_n624), .ZN(new_n759));
  INV_X1    g0559(.A(new_n758), .ZN(new_n760));
  OAI211_X1 g0560(.A(new_n760), .B(new_n623), .C1(new_n612), .C2(new_n614), .ZN(new_n761));
  AND2_X1   g0561(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g0562(.A(new_n762), .B(new_n669), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(new_n687), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n758), .A2(new_n737), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n689), .A2(new_n737), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(new_n223), .ZN(new_n767));
  OAI22_X1  g0567(.A1(new_n711), .A2(new_n213), .B1(new_n727), .B2(new_n719), .ZN(new_n768));
  INV_X1    g0568(.A(new_n707), .ZN(new_n769));
  AOI211_X1 g0569(.A(new_n249), .B(new_n768), .C1(G116), .C2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n705), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(G87), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n713), .A2(G303), .ZN(new_n773));
  INV_X1    g0573(.A(G294), .ZN(new_n774));
  OAI22_X1  g0574(.A1(new_n717), .A2(new_n774), .B1(new_n701), .B2(new_n724), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n775), .B1(new_n695), .B2(G107), .ZN(new_n776));
  NAND4_X1  g0576(.A1(new_n770), .A2(new_n772), .A3(new_n773), .A4(new_n776), .ZN(new_n777));
  AOI22_X1  g0577(.A1(new_n730), .A2(G143), .B1(G150), .B2(new_n718), .ZN(new_n778));
  INV_X1    g0578(.A(G137), .ZN(new_n779));
  INV_X1    g0579(.A(G159), .ZN(new_n780));
  OAI221_X1 g0580(.A(new_n778), .B1(new_n779), .B2(new_n714), .C1(new_n780), .C2(new_n707), .ZN(new_n781));
  INV_X1    g0581(.A(KEYINPUT34), .ZN(new_n782));
  OR2_X1    g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  AOI22_X1  g0583(.A1(new_n781), .A2(new_n782), .B1(G50), .B2(new_n695), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n771), .A2(G68), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n702), .A2(G132), .ZN(new_n786));
  NAND4_X1  g0586(.A1(new_n783), .A2(new_n784), .A3(new_n785), .A4(new_n786), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n249), .B1(new_n711), .B2(new_n369), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n777), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(new_n689), .ZN(new_n790));
  NAND4_X1  g0590(.A1(new_n765), .A2(new_n751), .A3(new_n767), .A4(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n764), .A2(new_n791), .ZN(G384));
  NAND2_X1  g0592(.A1(new_n339), .A2(new_n624), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n340), .A2(new_n343), .A3(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(KEYINPUT94), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n328), .A2(new_n339), .A3(new_n624), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n794), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n795), .B1(new_n794), .B2(new_n796), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n659), .A2(new_n657), .A3(new_n661), .ZN(new_n801));
  OR2_X1    g0601(.A1(new_n657), .A2(KEYINPUT31), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n801), .A2(new_n760), .A3(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n800), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n379), .A2(new_n375), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n805), .A2(new_n400), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n420), .A2(new_n622), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n412), .A2(new_n417), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n412), .A2(new_n622), .ZN(new_n809));
  INV_X1    g0609(.A(KEYINPUT37), .ZN(new_n810));
  NAND4_X1  g0610(.A1(new_n808), .A2(new_n809), .A3(new_n810), .A4(new_n403), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n621), .B1(new_n415), .B2(new_n416), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(new_n806), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(new_n403), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n814), .A2(KEYINPUT37), .ZN(new_n815));
  AOI21_X1  g0615(.A(KEYINPUT95), .B1(new_n811), .B2(new_n815), .ZN(new_n816));
  AND3_X1   g0616(.A1(new_n811), .A2(KEYINPUT95), .A3(new_n815), .ZN(new_n817));
  OAI211_X1 g0617(.A(new_n807), .B(KEYINPUT38), .C1(new_n816), .C2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n811), .A2(new_n815), .ZN(new_n820));
  INV_X1    g0620(.A(KEYINPUT95), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n811), .A2(KEYINPUT95), .A3(new_n815), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  AOI21_X1  g0624(.A(KEYINPUT38), .B1(new_n824), .B2(new_n807), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n804), .B1(new_n819), .B2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(KEYINPUT40), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n827), .A2(KEYINPUT98), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n827), .A2(KEYINPUT98), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n826), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n809), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n808), .A2(new_n809), .A3(new_n403), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(KEYINPUT37), .ZN(new_n834));
  AOI22_X1  g0634(.A1(new_n420), .A2(new_n832), .B1(new_n834), .B2(new_n811), .ZN(new_n835));
  OAI211_X1 g0635(.A(new_n818), .B(KEYINPUT97), .C1(KEYINPUT38), .C2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT97), .ZN(new_n837));
  NAND4_X1  g0637(.A1(new_n824), .A2(new_n837), .A3(KEYINPUT38), .A4(new_n807), .ZN(new_n838));
  NAND4_X1  g0638(.A1(new_n836), .A2(KEYINPUT40), .A3(new_n804), .A4(new_n838), .ZN(new_n839));
  AND2_X1   g0639(.A1(new_n831), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n801), .A2(new_n802), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n425), .A2(new_n841), .ZN(new_n842));
  XOR2_X1   g0642(.A(new_n842), .B(KEYINPUT99), .Z(new_n843));
  OAI21_X1  g0643(.A(G330), .B1(new_n840), .B2(new_n843), .ZN(new_n844));
  XNOR2_X1  g0644(.A(new_n844), .B(KEYINPUT100), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n840), .A2(new_n843), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT96), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n761), .A2(new_n757), .ZN(new_n849));
  INV_X1    g0649(.A(new_n799), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(new_n797), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT38), .ZN(new_n853));
  INV_X1    g0653(.A(new_n807), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n817), .A2(new_n816), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n853), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n852), .B1(new_n818), .B2(new_n856), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n591), .A2(new_n622), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n848), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n858), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n819), .A2(new_n825), .ZN(new_n861));
  OAI211_X1 g0661(.A(KEYINPUT96), .B(new_n860), .C1(new_n861), .C2(new_n852), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT39), .ZN(new_n863));
  OAI21_X1  g0663(.A(KEYINPUT97), .B1(new_n835), .B2(KEYINPUT38), .ZN(new_n864));
  OAI211_X1 g0664(.A(new_n863), .B(new_n838), .C1(new_n819), .C2(new_n864), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n340), .A2(new_n624), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n856), .A2(KEYINPUT39), .A3(new_n818), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n859), .A2(new_n862), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n674), .A2(new_n676), .ZN(new_n870));
  NAND4_X1  g0670(.A1(new_n870), .A2(new_n359), .A3(new_n421), .A4(new_n424), .ZN(new_n871));
  INV_X1    g0671(.A(new_n871), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n872), .A2(new_n597), .ZN(new_n873));
  XNOR2_X1  g0673(.A(new_n869), .B(new_n873), .ZN(new_n874));
  XNOR2_X1  g0674(.A(new_n847), .B(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n875), .B1(new_n203), .B2(new_n685), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n442), .B1(new_n536), .B2(KEYINPUT35), .ZN(new_n877));
  OAI211_X1 g0677(.A(new_n877), .B(new_n229), .C1(KEYINPUT35), .C2(new_n536), .ZN(new_n878));
  XNOR2_X1  g0678(.A(new_n878), .B(KEYINPUT36), .ZN(new_n879));
  OAI21_X1  g0679(.A(G77), .B1(new_n369), .B2(new_n219), .ZN(new_n880));
  OAI22_X1  g0680(.A1(new_n880), .A2(new_n230), .B1(G50), .B2(new_n219), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n881), .A2(G1), .A3(new_n206), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n876), .A2(new_n879), .A3(new_n882), .ZN(new_n883));
  XOR2_X1   g0683(.A(new_n883), .B(KEYINPUT101), .Z(G367));
  INV_X1    g0684(.A(KEYINPUT107), .ZN(new_n885));
  NAND4_X1  g0685(.A1(new_n684), .A2(new_n627), .A3(new_n626), .A4(new_n628), .ZN(new_n886));
  NAND4_X1  g0686(.A1(new_n617), .A2(new_n468), .A3(new_n610), .A4(new_n623), .ZN(new_n887));
  AND3_X1   g0687(.A1(new_n636), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  AND4_X1   g0688(.A1(new_n674), .A2(new_n669), .A3(new_n888), .A4(new_n676), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT105), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n549), .A2(new_n624), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n541), .A2(new_n552), .A3(new_n891), .ZN(new_n892));
  NAND4_X1  g0692(.A1(new_n542), .A2(new_n549), .A3(new_n551), .A4(new_n624), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(KEYINPUT102), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT102), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n892), .A2(new_n896), .A3(new_n893), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  OAI21_X1  g0698(.A(KEYINPUT44), .B1(new_n640), .B2(new_n898), .ZN(new_n899));
  XOR2_X1   g0699(.A(KEYINPUT104), .B(KEYINPUT45), .Z(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n513), .A2(new_n490), .A3(new_n623), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n887), .A2(new_n902), .ZN(new_n903));
  AND3_X1   g0703(.A1(new_n892), .A2(new_n896), .A3(new_n893), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n896), .B1(new_n892), .B2(new_n893), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n901), .B1(new_n903), .B2(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n640), .A2(new_n898), .A3(new_n900), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT44), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n903), .A2(new_n906), .A3(new_n909), .ZN(new_n910));
  AND4_X1   g0710(.A1(new_n899), .A2(new_n907), .A3(new_n908), .A4(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n890), .B1(new_n911), .B2(new_n636), .ZN(new_n912));
  NAND4_X1  g0712(.A1(new_n899), .A2(new_n907), .A3(new_n908), .A4(new_n910), .ZN(new_n913));
  INV_X1    g0713(.A(new_n636), .ZN(new_n914));
  NOR3_X1   g0714(.A1(new_n913), .A2(KEYINPUT105), .A3(new_n914), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n889), .B1(new_n912), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(KEYINPUT106), .ZN(new_n917));
  AND2_X1   g0717(.A1(new_n899), .A2(new_n910), .ZN(new_n918));
  AND2_X1   g0718(.A1(new_n907), .A2(new_n908), .ZN(new_n919));
  NAND4_X1  g0719(.A1(new_n918), .A2(new_n919), .A3(new_n890), .A4(new_n636), .ZN(new_n920));
  OAI21_X1  g0720(.A(KEYINPUT105), .B1(new_n913), .B2(new_n914), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT106), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n922), .A2(new_n923), .A3(new_n889), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n677), .B1(new_n917), .B2(new_n924), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n642), .B(KEYINPUT41), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n885), .B1(new_n925), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n686), .A2(G1), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  AND3_X1   g0730(.A1(new_n922), .A2(new_n923), .A3(new_n889), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n923), .B1(new_n922), .B2(new_n889), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n678), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n933), .A2(KEYINPUT107), .A3(new_n926), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n928), .A2(new_n930), .A3(new_n934), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n906), .A2(new_n887), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n936), .B(KEYINPUT42), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n601), .B1(new_n898), .B2(new_n639), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n937), .B1(new_n624), .B2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT43), .ZN(new_n940));
  INV_X1    g0740(.A(new_n575), .ZN(new_n941));
  OR3_X1    g0741(.A1(new_n604), .A2(new_n941), .A3(new_n623), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n600), .B1(new_n941), .B2(new_n623), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n939), .B1(new_n940), .B2(new_n945), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n944), .A2(KEYINPUT43), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n946), .B(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT103), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n636), .A2(new_n906), .ZN(new_n951));
  NOR3_X1   g0751(.A1(new_n949), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n946), .B(new_n947), .ZN(new_n953));
  INV_X1    g0753(.A(new_n951), .ZN(new_n954));
  AOI21_X1  g0754(.A(KEYINPUT103), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n952), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n949), .A2(new_n951), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n935), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n945), .A2(new_n739), .ZN(new_n959));
  AOI22_X1  g0759(.A1(new_n695), .A2(G58), .B1(G150), .B2(new_n730), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n702), .A2(G137), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n366), .B1(new_n713), .B2(G143), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n710), .A2(G68), .ZN(new_n963));
  NAND4_X1  g0763(.A1(new_n960), .A2(new_n961), .A3(new_n962), .A4(new_n963), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n705), .A2(new_n223), .ZN(new_n965));
  AOI22_X1  g0765(.A1(new_n769), .A2(G50), .B1(G159), .B2(new_n718), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT108), .ZN(new_n967));
  NOR3_X1   g0767(.A1(new_n964), .A2(new_n965), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n771), .A2(G97), .ZN(new_n969));
  INV_X1    g0769(.A(G317), .ZN(new_n970));
  OAI221_X1 g0770(.A(new_n969), .B1(new_n724), .B2(new_n714), .C1(new_n970), .C2(new_n701), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n694), .A2(new_n442), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(KEYINPUT46), .ZN(new_n973));
  AOI22_X1  g0773(.A1(new_n730), .A2(G303), .B1(new_n710), .B2(G107), .ZN(new_n974));
  OAI211_X1 g0774(.A(new_n974), .B(new_n366), .C1(new_n774), .C2(new_n719), .ZN(new_n975));
  NOR3_X1   g0775(.A1(new_n971), .A2(new_n973), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n769), .A2(G283), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n968), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  XOR2_X1   g0778(.A(new_n978), .B(KEYINPUT47), .Z(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(new_n689), .ZN(new_n980));
  INV_X1    g0780(.A(new_n743), .ZN(new_n981));
  OAI221_X1 g0781(.A(new_n741), .B1(new_n208), .B2(new_n352), .C1(new_n981), .C2(new_n240), .ZN(new_n982));
  NAND4_X1  g0782(.A1(new_n959), .A2(new_n751), .A3(new_n980), .A4(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n958), .A2(new_n983), .ZN(G387));
  NOR2_X1   g0784(.A1(new_n678), .A2(new_n888), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n643), .B1(new_n985), .B2(KEYINPUT111), .ZN(new_n986));
  INV_X1    g0786(.A(new_n889), .ZN(new_n987));
  OAI211_X1 g0787(.A(new_n986), .B(new_n987), .C1(KEYINPUT111), .C2(new_n985), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n888), .A2(new_n929), .ZN(new_n989));
  AOI22_X1  g0789(.A1(new_n769), .A2(G303), .B1(G311), .B2(new_n718), .ZN(new_n990));
  XOR2_X1   g0790(.A(KEYINPUT109), .B(G322), .Z(new_n991));
  OAI221_X1 g0791(.A(new_n990), .B1(new_n970), .B2(new_n717), .C1(new_n714), .C2(new_n991), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT48), .ZN(new_n993));
  OAI221_X1 g0793(.A(new_n993), .B1(new_n727), .B2(new_n711), .C1(new_n774), .C2(new_n694), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n994), .B(KEYINPUT49), .Z(new_n995));
  AOI21_X1  g0795(.A(new_n249), .B1(new_n702), .B2(new_n733), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n996), .B1(new_n705), .B2(new_n442), .ZN(new_n997));
  OAI22_X1  g0797(.A1(new_n780), .A2(new_n714), .B1(new_n719), .B2(new_n276), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n969), .B1(new_n330), .B2(new_n717), .ZN(new_n999));
  AOI211_X1 g0799(.A(new_n998), .B(new_n999), .C1(G77), .C2(new_n695), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n710), .A2(new_n351), .ZN(new_n1001));
  OAI211_X1 g0801(.A(new_n1000), .B(new_n1001), .C1(new_n271), .C2(new_n701), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n249), .B1(new_n707), .B2(new_n219), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n995), .A2(new_n997), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  XOR2_X1   g0804(.A(new_n1004), .B(KEYINPUT110), .Z(new_n1005));
  OAI21_X1  g0805(.A(new_n743), .B1(new_n236), .B2(new_n433), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1006), .B1(new_n644), .B2(new_n746), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n276), .A2(G50), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT50), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(G68), .A2(G77), .ZN(new_n1010));
  NAND4_X1  g0810(.A1(new_n1009), .A2(new_n433), .A3(new_n1010), .A4(new_n644), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1007), .A2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(G107), .B2(new_n208), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n1005), .A2(new_n689), .B1(new_n741), .B2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n626), .A2(new_n628), .A3(new_n739), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1014), .A2(new_n751), .A3(new_n1015), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n988), .A2(new_n989), .A3(new_n1016), .ZN(G393));
  NAND2_X1  g0817(.A1(new_n913), .A2(new_n914), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT112), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1019), .A2(new_n922), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1020), .A2(new_n987), .ZN(new_n1021));
  OAI211_X1 g0821(.A(new_n1021), .B(new_n642), .C1(new_n931), .C2(new_n932), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n1020), .A2(new_n930), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n743), .A2(new_n247), .ZN(new_n1024));
  OAI211_X1 g0824(.A(new_n1024), .B(new_n741), .C1(new_n213), .C2(new_n208), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n714), .A2(new_n970), .B1(new_n717), .B2(new_n724), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT52), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n1027), .B1(new_n482), .B2(new_n705), .C1(new_n727), .C2(new_n694), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n711), .A2(new_n442), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n991), .A2(new_n701), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n366), .B1(new_n707), .B2(new_n774), .ZN(new_n1031));
  NOR4_X1   g0831(.A1(new_n1028), .A2(new_n1029), .A3(new_n1030), .A4(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n718), .A2(G303), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n730), .A2(G159), .B1(G150), .B2(new_n713), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1034), .A2(KEYINPUT51), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n702), .A2(G143), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n772), .B(new_n1036), .C1(new_n276), .C2(new_n707), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n694), .A2(new_n219), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n366), .B1(new_n718), .B2(G50), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n710), .A2(G77), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n1039), .B(new_n1040), .C1(new_n1034), .C2(KEYINPUT51), .ZN(new_n1041));
  NOR3_X1   g0841(.A1(new_n1037), .A2(new_n1038), .A3(new_n1041), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n1032), .A2(new_n1033), .B1(new_n1035), .B2(new_n1042), .ZN(new_n1043));
  OAI211_X1 g0843(.A(new_n751), .B(new_n1025), .C1(new_n1043), .C2(new_n690), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1044), .B1(new_n739), .B2(new_n906), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n1023), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1022), .A2(new_n1046), .ZN(G390));
  NOR3_X1   g0847(.A1(new_n425), .A2(new_n681), .A3(new_n841), .ZN(new_n1048));
  NOR3_X1   g0848(.A1(new_n872), .A2(new_n1048), .A3(new_n597), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n756), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n673), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n757), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NAND4_X1  g0853(.A1(new_n801), .A2(G330), .A3(new_n760), .A4(new_n802), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1054), .A2(new_n800), .ZN(new_n1055));
  OAI211_X1 g0855(.A(G330), .B(new_n760), .C1(new_n660), .C2(new_n668), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n1053), .B(new_n1055), .C1(new_n800), .C2(new_n1056), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n1057), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n1054), .A2(new_n800), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1056), .A2(new_n800), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n1060), .A2(new_n1061), .B1(new_n757), .B2(new_n761), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1049), .B1(new_n1058), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1063), .A2(KEYINPUT114), .ZN(new_n1064));
  INV_X1    g0864(.A(KEYINPUT114), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n1049), .B(new_n1065), .C1(new_n1058), .C2(new_n1062), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1064), .A2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n865), .A2(new_n867), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n866), .B1(new_n849), .B2(new_n851), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1068), .A2(new_n1070), .ZN(new_n1071));
  OR2_X1    g0871(.A1(new_n1056), .A2(new_n800), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n851), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n866), .B(KEYINPUT113), .ZN(new_n1074));
  NAND4_X1  g0874(.A1(new_n836), .A2(new_n838), .A3(new_n1073), .A4(new_n1074), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1071), .A2(new_n1072), .A3(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1069), .B1(new_n865), .B2(new_n867), .ZN(new_n1077));
  AND4_X1   g0877(.A1(new_n836), .A2(new_n838), .A3(new_n1073), .A4(new_n1074), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1059), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1076), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1067), .A2(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n1048), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1082), .A2(new_n598), .A3(new_n871), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1062), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1083), .B1(new_n1084), .B2(new_n1057), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1076), .A2(new_n1079), .A3(new_n1085), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1081), .A2(new_n642), .A3(new_n1086), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1076), .A2(new_n929), .A3(new_n1079), .ZN(new_n1088));
  INV_X1    g0888(.A(KEYINPUT116), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n694), .A2(new_n271), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(new_n1090), .B(new_n1091), .ZN(new_n1092));
  XOR2_X1   g0892(.A(KEYINPUT54), .B(G143), .Z(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1092), .B1(new_n707), .B2(new_n1094), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n719), .A2(new_n779), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n705), .A2(new_n330), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n730), .A2(G132), .B1(new_n710), .B2(G159), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n366), .B1(new_n713), .B2(G128), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n702), .A2(G125), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1098), .A2(new_n1099), .A3(new_n1100), .ZN(new_n1101));
  NOR4_X1   g0901(.A1(new_n1095), .A2(new_n1096), .A3(new_n1097), .A4(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n713), .A2(G283), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n696), .A2(new_n785), .A3(new_n1040), .A4(new_n1103), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n707), .A2(new_n213), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n717), .A2(new_n442), .ZN(new_n1106));
  OAI221_X1 g0906(.A(new_n366), .B1(new_n701), .B2(new_n774), .C1(new_n719), .C2(new_n482), .ZN(new_n1107));
  NOR4_X1   g0907(.A1(new_n1104), .A2(new_n1105), .A3(new_n1106), .A4(new_n1107), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n689), .B1(new_n1102), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n766), .A2(new_n276), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1109), .A2(new_n751), .A3(new_n1110), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n1068), .A2(new_n737), .B1(new_n1089), .B2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1112), .B1(new_n1089), .B2(new_n1111), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1087), .A2(new_n1088), .A3(new_n1113), .ZN(G378));
  AND3_X1   g0914(.A1(new_n831), .A2(G330), .A3(new_n839), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1115), .A2(new_n869), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n831), .A2(G330), .A3(new_n839), .ZN(new_n1117));
  NAND4_X1  g0917(.A1(new_n1117), .A2(new_n862), .A3(new_n868), .A4(new_n859), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1119));
  XOR2_X1   g0919(.A(new_n303), .B(KEYINPUT55), .Z(new_n1120));
  NAND2_X1  g0920(.A1(new_n289), .A2(new_n622), .ZN(new_n1121));
  XNOR2_X1  g0921(.A(new_n1120), .B(new_n1121), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(KEYINPUT123), .B(KEYINPUT56), .ZN(new_n1123));
  OR2_X1    g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1119), .A2(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1126), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1116), .A2(new_n1118), .A3(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1127), .A2(new_n929), .A3(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1126), .A2(new_n737), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n771), .A2(G58), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(new_n1132), .B(KEYINPUT118), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n694), .A2(new_n223), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n769), .A2(new_n351), .B1(new_n710), .B2(G68), .ZN(new_n1136));
  OAI221_X1 g0936(.A(new_n1136), .B1(new_n482), .B2(new_n717), .C1(new_n719), .C2(new_n213), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n249), .A2(G41), .ZN(new_n1138));
  OAI221_X1 g0938(.A(new_n1138), .B1(new_n727), .B2(new_n701), .C1(new_n442), .C2(new_n714), .ZN(new_n1139));
  NOR4_X1   g0939(.A1(new_n1134), .A2(new_n1135), .A3(new_n1137), .A4(new_n1139), .ZN(new_n1140));
  XOR2_X1   g0940(.A(new_n1140), .B(KEYINPUT58), .Z(new_n1141));
  NAND2_X1  g0941(.A1(new_n254), .A2(new_n255), .ZN(new_n1142));
  XNOR2_X1  g0942(.A(new_n1142), .B(KEYINPUT117), .ZN(new_n1143));
  OR3_X1    g0943(.A1(new_n1143), .A2(new_n1138), .A3(G50), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n707), .A2(new_n779), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n718), .A2(G132), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1146), .B1(new_n711), .B2(new_n271), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n695), .A2(new_n1093), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1147), .B1(new_n1148), .B2(KEYINPUT119), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n730), .A2(G128), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n1149), .B(new_n1150), .C1(KEYINPUT119), .C2(new_n1148), .ZN(new_n1151));
  AOI211_X1 g0951(.A(new_n1145), .B(new_n1151), .C1(G125), .C2(new_n713), .ZN(new_n1152));
  XOR2_X1   g0952(.A(new_n1152), .B(KEYINPUT59), .Z(new_n1153));
  OR2_X1    g0953(.A1(KEYINPUT120), .A2(G124), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(KEYINPUT120), .A2(G124), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n702), .A2(new_n1154), .A3(new_n1155), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n1143), .B(new_n1156), .C1(new_n705), .C2(new_n780), .ZN(new_n1157));
  XOR2_X1   g0957(.A(new_n1157), .B(KEYINPUT121), .Z(new_n1158));
  OAI211_X1 g0958(.A(new_n1141), .B(new_n1144), .C1(new_n1153), .C2(new_n1158), .ZN(new_n1159));
  XOR2_X1   g0959(.A(new_n1159), .B(KEYINPUT122), .Z(new_n1160));
  NAND2_X1  g0960(.A1(new_n1160), .A2(new_n689), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n766), .A2(new_n330), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n1131), .A2(new_n751), .A3(new_n1161), .A4(new_n1162), .ZN(new_n1163));
  AND2_X1   g0963(.A1(new_n1130), .A2(new_n1163), .ZN(new_n1164));
  AND3_X1   g0964(.A1(new_n1116), .A2(new_n1118), .A3(new_n1128), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1128), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1086), .A2(new_n1049), .ZN(new_n1168));
  AOI21_X1  g0968(.A(KEYINPUT57), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  NAND4_X1  g0969(.A1(new_n1127), .A2(KEYINPUT57), .A3(new_n1129), .A4(new_n1168), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1170), .A2(new_n642), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1164), .B1(new_n1169), .B2(new_n1171), .ZN(G375));
  NOR2_X1   g0972(.A1(new_n1062), .A2(new_n1058), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(new_n1083), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1067), .A2(new_n926), .A3(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1173), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n766), .A2(new_n219), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n851), .A2(new_n738), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1134), .B1(G137), .B2(new_n730), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n769), .A2(G150), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n713), .A2(G132), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(new_n702), .A2(G128), .B1(new_n710), .B2(G50), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1182), .B1(new_n719), .B2(new_n1094), .ZN(new_n1183));
  AOI211_X1 g0983(.A(new_n366), .B(new_n1183), .C1(G159), .C2(new_n695), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n1179), .A2(new_n1180), .A3(new_n1181), .A4(new_n1184), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1001), .B1(new_n482), .B2(new_n707), .ZN(new_n1186));
  AOI211_X1 g0986(.A(new_n249), .B(new_n1186), .C1(G294), .C2(new_n713), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n730), .A2(G283), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n965), .B1(G303), .B2(new_n702), .ZN(new_n1189));
  AND3_X1   g0989(.A1(new_n1187), .A2(new_n1188), .A3(new_n1189), .ZN(new_n1190));
  OAI221_X1 g0990(.A(new_n1190), .B1(new_n213), .B2(new_n694), .C1(new_n442), .C2(new_n719), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n690), .B1(new_n1185), .B2(new_n1191), .ZN(new_n1192));
  NOR3_X1   g0992(.A1(new_n1178), .A2(new_n687), .A3(new_n1192), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n1176), .A2(new_n929), .B1(new_n1177), .B2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1175), .A2(new_n1194), .ZN(G381));
  NAND3_X1  g0995(.A1(new_n1127), .A2(new_n1129), .A3(new_n1168), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT57), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1198), .A2(new_n642), .A3(new_n1170), .ZN(new_n1199));
  AND3_X1   g0999(.A1(new_n1087), .A2(new_n1088), .A3(new_n1113), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1199), .A2(new_n1200), .A3(new_n1164), .ZN(new_n1201));
  NOR3_X1   g1001(.A1(new_n1201), .A2(G396), .A3(G393), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(G381), .A2(G384), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(G387), .A2(G390), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1202), .A2(new_n1203), .A3(new_n1204), .ZN(G407));
  OAI211_X1 g1005(.A(G407), .B(G213), .C1(G343), .C2(new_n1201), .ZN(G409));
  INV_X1    g1006(.A(G390), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(G387), .A2(new_n1207), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n958), .A2(G390), .A3(new_n983), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1208), .A2(KEYINPUT125), .A3(new_n1209), .ZN(new_n1210));
  XOR2_X1   g1010(.A(G393), .B(G396), .Z(new_n1211));
  INV_X1    g1011(.A(KEYINPUT125), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n958), .A2(G390), .A3(new_n1212), .A4(new_n983), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1210), .A2(new_n1211), .A3(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT126), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1210), .A2(new_n1211), .A3(KEYINPUT126), .A4(new_n1213), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1209), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n1219), .A2(new_n1211), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1220), .A2(new_n1208), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1218), .A2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(G375), .A2(G378), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT60), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n643), .B1(new_n1174), .B2(new_n1224), .ZN(new_n1225));
  OAI211_X1 g1025(.A(new_n1225), .B(new_n1063), .C1(new_n1224), .C2(new_n1174), .ZN(new_n1226));
  AND3_X1   g1026(.A1(new_n1226), .A2(G384), .A3(new_n1194), .ZN(new_n1227));
  AOI21_X1  g1027(.A(G384), .B1(new_n1226), .B2(new_n1194), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(G213), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1230), .A2(G343), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  OAI211_X1 g1032(.A(new_n1130), .B(new_n1163), .C1(new_n1196), .C2(new_n927), .ZN(new_n1233));
  OR2_X1    g1033(.A1(new_n1233), .A2(G378), .ZN(new_n1234));
  NAND4_X1  g1034(.A1(new_n1223), .A2(new_n1229), .A3(new_n1232), .A4(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT124), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1235), .B1(new_n1236), .B2(KEYINPUT63), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1200), .B1(new_n1199), .B2(new_n1164), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1233), .A2(G378), .ZN(new_n1239));
  NOR3_X1   g1039(.A1(new_n1238), .A2(new_n1231), .A3(new_n1239), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1236), .A2(KEYINPUT63), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1240), .A2(new_n1229), .A3(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1237), .A2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT61), .ZN(new_n1244));
  INV_X1    g1044(.A(G2897), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1229), .B1(new_n1245), .B2(new_n1232), .ZN(new_n1246));
  OAI211_X1 g1046(.A(G2897), .B(new_n1231), .C1(new_n1227), .C2(new_n1228), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1244), .B1(new_n1240), .B2(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1222), .A2(new_n1243), .A3(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1231), .B1(G375), .B2(G378), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1252), .A2(KEYINPUT124), .A3(new_n1234), .A4(new_n1229), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT127), .ZN(new_n1254));
  AOI21_X1  g1054(.A(KEYINPUT62), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1236), .B1(new_n1254), .B2(KEYINPUT62), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1256), .B1(new_n1240), .B2(new_n1229), .ZN(new_n1257));
  NOR3_X1   g1057(.A1(new_n1255), .A2(new_n1249), .A3(new_n1257), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1251), .B1(new_n1258), .B2(new_n1222), .ZN(G405));
  NAND2_X1  g1059(.A1(new_n1223), .A2(new_n1201), .ZN(new_n1260));
  OR2_X1    g1060(.A1(new_n1260), .A2(new_n1229), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1260), .A2(new_n1229), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  XNOR2_X1  g1063(.A(new_n1222), .B(new_n1263), .ZN(G402));
endmodule


