//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 1 0 0 1 1 1 0 1 1 1 0 1 1 0 0 0 0 1 1 0 0 1 0 1 0 0 1 1 1 0 1 1 0 0 0 1 1 0 1 0 0 1 0 1 0 1 0 0 1 1 1 0 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:39 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1233, new_n1234, new_n1235, new_n1236, new_n1237,
    new_n1238, new_n1239, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  AOI211_X1 g0005(.A(G50), .B(G77), .C1(new_n203), .C2(new_n205), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  AOI22_X1  g0007(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n211));
  NAND4_X1  g0011(.A1(new_n208), .A2(new_n209), .A3(new_n210), .A4(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(G1), .ZN(new_n213));
  INV_X1    g0013(.A(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n212), .A2(new_n216), .ZN(new_n217));
  OR2_X1    g0017(.A1(new_n217), .A2(KEYINPUT1), .ZN(new_n218));
  XNOR2_X1  g0018(.A(new_n218), .B(KEYINPUT65), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n216), .A2(G13), .ZN(new_n220));
  OAI211_X1 g0020(.A(new_n220), .B(G250), .C1(G257), .C2(G264), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(KEYINPUT0), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G13), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n223), .A2(new_n214), .ZN(new_n224));
  INV_X1    g0024(.A(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n203), .A2(new_n205), .ZN(new_n226));
  INV_X1    g0026(.A(G50), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n222), .B1(new_n225), .B2(new_n229), .ZN(new_n230));
  AOI211_X1 g0030(.A(new_n219), .B(new_n230), .C1(KEYINPUT1), .C2(new_n217), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XNOR2_X1  g0039(.A(G87), .B(G97), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT66), .ZN(new_n241));
  XOR2_X1   g0041(.A(G107), .B(G116), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n243), .B(KEYINPUT67), .Z(new_n244));
  NAND2_X1  g0044(.A1(new_n227), .A2(G68), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n202), .A2(G50), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G58), .B(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n244), .B(new_n249), .ZN(G351));
  INV_X1    g0050(.A(G41), .ZN(new_n251));
  INV_X1    g0051(.A(G45), .ZN(new_n252));
  AOI21_X1  g0052(.A(G1), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(G33), .A2(G41), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n254), .A2(G1), .A3(G13), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n253), .A2(new_n255), .A3(G274), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n223), .B1(G33), .B2(G41), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n257), .A2(new_n253), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G226), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n256), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT3), .ZN(new_n263));
  INV_X1    g0063(.A(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(KEYINPUT3), .A2(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G1698), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n267), .A2(G222), .A3(new_n268), .ZN(new_n269));
  XNOR2_X1  g0069(.A(new_n269), .B(KEYINPUT68), .ZN(new_n270));
  AND2_X1   g0070(.A1(KEYINPUT3), .A2(G33), .ZN(new_n271));
  NOR2_X1   g0071(.A1(KEYINPUT3), .A2(G33), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n273), .A2(new_n268), .ZN(new_n274));
  AOI22_X1  g0074(.A1(new_n274), .A2(G223), .B1(G77), .B2(new_n273), .ZN(new_n275));
  AND2_X1   g0075(.A1(new_n270), .A2(new_n275), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n262), .B1(new_n276), .B2(new_n255), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G179), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT70), .ZN(new_n281));
  NAND4_X1  g0081(.A1(KEYINPUT69), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n282));
  AND2_X1   g0082(.A1(new_n282), .A2(new_n223), .ZN(new_n283));
  NAND3_X1  g0083(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT69), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n281), .B1(new_n283), .B2(new_n286), .ZN(new_n287));
  NAND4_X1  g0087(.A1(new_n286), .A2(new_n281), .A3(new_n223), .A4(new_n282), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G13), .ZN(new_n291));
  NOR3_X1   g0091(.A1(new_n291), .A2(new_n214), .A3(G1), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT71), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n294), .B1(new_n214), .B2(G1), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n213), .A2(KEYINPUT71), .A3(G20), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n293), .A2(G50), .A3(new_n297), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n214), .B1(new_n226), .B2(new_n227), .ZN(new_n299));
  XNOR2_X1  g0099(.A(KEYINPUT8), .B(G58), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n264), .A2(G20), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G150), .ZN(new_n303));
  NOR2_X1   g0103(.A1(G20), .A2(G33), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  OAI22_X1  g0105(.A1(new_n300), .A2(new_n302), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  OR2_X1    g0106(.A1(new_n299), .A2(new_n306), .ZN(new_n307));
  AOI22_X1  g0107(.A1(new_n307), .A2(new_n290), .B1(new_n227), .B2(new_n292), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n298), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(G169), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n277), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n280), .A2(new_n309), .A3(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  OR2_X1    g0113(.A1(new_n309), .A2(KEYINPUT9), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n309), .A2(KEYINPUT9), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n278), .A2(G190), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n277), .A2(G200), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  OAI21_X1  g0120(.A(KEYINPUT10), .B1(new_n317), .B2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT10), .ZN(new_n322));
  NAND4_X1  g0122(.A1(new_n316), .A2(new_n322), .A3(new_n319), .A4(new_n318), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n313), .B1(new_n321), .B2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(G77), .ZN(new_n325));
  OAI22_X1  g0125(.A1(new_n302), .A2(new_n325), .B1(new_n214), .B2(G68), .ZN(new_n326));
  OAI22_X1  g0126(.A1(new_n326), .A2(KEYINPUT74), .B1(new_n227), .B2(new_n305), .ZN(new_n327));
  AND2_X1   g0127(.A1(new_n326), .A2(KEYINPUT74), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n290), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT11), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  OAI211_X1 g0131(.A(KEYINPUT11), .B(new_n290), .C1(new_n327), .C2(new_n328), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n292), .A2(new_n202), .ZN(new_n333));
  XNOR2_X1  g0133(.A(new_n333), .B(KEYINPUT12), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n286), .A2(new_n223), .A3(new_n282), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(KEYINPUT70), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(new_n288), .ZN(new_n337));
  INV_X1    g0137(.A(new_n292), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n337), .A2(G68), .A3(new_n338), .A4(new_n297), .ZN(new_n339));
  NAND4_X1  g0139(.A1(new_n331), .A2(new_n332), .A3(new_n334), .A4(new_n339), .ZN(new_n340));
  AND3_X1   g0140(.A1(new_n253), .A2(new_n255), .A3(G274), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n341), .B1(G238), .B2(new_n258), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT72), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n260), .A2(new_n268), .ZN(new_n344));
  INV_X1    g0144(.A(G232), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(G1698), .ZN(new_n346));
  OAI211_X1 g0146(.A(new_n344), .B(new_n346), .C1(new_n271), .C2(new_n272), .ZN(new_n347));
  NAND2_X1  g0147(.A1(G33), .A2(G97), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n343), .B1(new_n349), .B2(new_n257), .ZN(new_n350));
  AOI211_X1 g0150(.A(KEYINPUT72), .B(new_n255), .C1(new_n347), .C2(new_n348), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n342), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(KEYINPUT13), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT13), .ZN(new_n354));
  OAI211_X1 g0154(.A(new_n354), .B(new_n342), .C1(new_n350), .C2(new_n351), .ZN(new_n355));
  AND2_X1   g0155(.A1(new_n355), .A2(G190), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n340), .B1(new_n353), .B2(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n353), .A2(KEYINPUT73), .A3(new_n355), .ZN(new_n358));
  OR2_X1    g0158(.A1(new_n350), .A2(new_n351), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT73), .ZN(new_n360));
  NAND4_X1  g0160(.A1(new_n359), .A2(new_n360), .A3(new_n354), .A4(new_n342), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n358), .A2(G200), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n357), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n353), .A2(G179), .A3(new_n355), .ZN(new_n365));
  INV_X1    g0165(.A(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n358), .A2(G169), .A3(new_n361), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n366), .B1(new_n367), .B2(KEYINPUT14), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT14), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n358), .A2(new_n361), .A3(new_n369), .A4(G169), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT75), .ZN(new_n371));
  AND2_X1   g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n370), .A2(new_n371), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n368), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n364), .B1(new_n374), .B2(new_n340), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n300), .B1(new_n295), .B2(new_n296), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n337), .A2(new_n338), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n300), .A2(new_n292), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n265), .A2(new_n214), .A3(new_n266), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT7), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n273), .A2(KEYINPUT7), .A3(new_n214), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n202), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(G58), .A2(G68), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n203), .A2(new_n205), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(G20), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n304), .A2(G159), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  OAI21_X1  g0189(.A(KEYINPUT16), .B1(new_n384), .B2(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(KEYINPUT7), .B1(new_n273), .B2(new_n214), .ZN(new_n391));
  NOR4_X1   g0191(.A1(new_n271), .A2(new_n272), .A3(new_n381), .A4(G20), .ZN(new_n392));
  OAI21_X1  g0192(.A(G68), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT16), .ZN(new_n394));
  AOI22_X1  g0194(.A1(new_n386), .A2(G20), .B1(G159), .B2(new_n304), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n393), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n390), .A2(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n379), .B1(new_n397), .B2(new_n290), .ZN(new_n398));
  INV_X1    g0198(.A(G87), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n264), .A2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n260), .A2(G1698), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n402), .B1(G223), .B2(G1698), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n401), .B1(new_n403), .B2(new_n273), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n341), .B1(new_n404), .B2(new_n257), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n213), .B1(G41), .B2(G45), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n255), .A2(G232), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(KEYINPUT76), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT76), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n255), .A2(new_n406), .A3(new_n409), .A4(G232), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  AND3_X1   g0211(.A1(new_n405), .A2(G190), .A3(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(G200), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n413), .B1(new_n405), .B2(new_n411), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT77), .ZN(new_n415));
  NOR3_X1   g0215(.A1(new_n412), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(new_n411), .ZN(new_n417));
  NOR2_X1   g0217(.A1(G223), .A2(G1698), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n418), .B1(new_n260), .B2(G1698), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n400), .B1(new_n419), .B2(new_n267), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n256), .B1(new_n420), .B2(new_n255), .ZN(new_n421));
  OAI21_X1  g0221(.A(G200), .B1(new_n417), .B2(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n405), .A2(G190), .A3(new_n411), .ZN(new_n423));
  AOI21_X1  g0223(.A(KEYINPUT77), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n398), .B1(new_n416), .B2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT17), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n398), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT18), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n405), .A2(new_n411), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(new_n310), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n405), .A2(new_n279), .A3(new_n411), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n428), .A2(new_n429), .A3(new_n431), .A4(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n337), .B1(new_n390), .B2(new_n396), .ZN(new_n434));
  OAI211_X1 g0234(.A(new_n431), .B(new_n432), .C1(new_n434), .C2(new_n379), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(KEYINPUT18), .ZN(new_n436));
  OAI211_X1 g0236(.A(new_n398), .B(KEYINPUT17), .C1(new_n416), .C2(new_n424), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n427), .A2(new_n433), .A3(new_n436), .A4(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n345), .A2(new_n268), .ZN(new_n440));
  OR2_X1    g0240(.A1(new_n268), .A2(G238), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n273), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(G107), .ZN(new_n443));
  AOI211_X1 g0243(.A(new_n255), .B(new_n442), .C1(new_n443), .C2(new_n273), .ZN(new_n444));
  INV_X1    g0244(.A(G244), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n256), .B1(new_n259), .B2(new_n445), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(G190), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n448), .B1(new_n413), .B2(new_n447), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n293), .A2(G77), .A3(new_n297), .ZN(new_n450));
  INV_X1    g0250(.A(new_n300), .ZN(new_n451));
  AOI22_X1  g0251(.A1(new_n451), .A2(new_n304), .B1(G20), .B2(G77), .ZN(new_n452));
  XNOR2_X1  g0252(.A(KEYINPUT15), .B(G87), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n452), .B1(new_n302), .B2(new_n453), .ZN(new_n454));
  AOI22_X1  g0254(.A1(new_n454), .A2(new_n290), .B1(new_n325), .B2(new_n292), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n450), .A2(new_n455), .ZN(new_n456));
  OR2_X1    g0256(.A1(new_n449), .A2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n447), .A2(new_n279), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n310), .B1(new_n444), .B2(new_n446), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n459), .A2(new_n456), .A3(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n458), .A2(new_n462), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n324), .A2(new_n375), .A3(new_n439), .A4(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT4), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n268), .A2(G244), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n467), .B1(new_n265), .B2(new_n266), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n466), .B1(new_n468), .B2(KEYINPUT78), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n445), .A2(G1698), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n470), .B(KEYINPUT78), .C1(new_n272), .C2(new_n271), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  OAI21_X1  g0272(.A(KEYINPUT79), .B1(new_n469), .B2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT78), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n474), .B1(new_n273), .B2(new_n467), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT79), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n475), .A2(new_n476), .A3(new_n466), .A4(new_n471), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n267), .A2(KEYINPUT4), .A3(new_n470), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n267), .A2(G250), .A3(G1698), .ZN(new_n479));
  NAND2_X1  g0279(.A1(G33), .A2(G283), .ZN(new_n480));
  AND3_X1   g0280(.A1(new_n478), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n473), .A2(new_n477), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(new_n257), .ZN(new_n483));
  AND2_X1   g0283(.A1(KEYINPUT5), .A2(G41), .ZN(new_n484));
  NOR2_X1   g0284(.A1(KEYINPUT5), .A2(G41), .ZN(new_n485));
  OR2_X1    g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n252), .A2(G1), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n486), .A2(G274), .A3(new_n255), .A4(new_n487), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n487), .B1(new_n484), .B2(new_n485), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(new_n255), .ZN(new_n490));
  INV_X1    g0290(.A(G257), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n488), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n310), .B1(new_n483), .B2(new_n493), .ZN(new_n494));
  AOI211_X1 g0294(.A(new_n279), .B(new_n492), .C1(new_n482), .C2(new_n257), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT80), .ZN(new_n496));
  OAI21_X1  g0296(.A(G107), .B1(new_n391), .B2(new_n392), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT6), .ZN(new_n498));
  AND2_X1   g0298(.A1(G97), .A2(G107), .ZN(new_n499));
  NOR2_X1   g0299(.A1(G97), .A2(G107), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n443), .A2(KEYINPUT6), .A3(G97), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AOI22_X1  g0303(.A1(new_n503), .A2(G20), .B1(G77), .B2(new_n304), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n497), .A2(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(G97), .ZN(new_n506));
  AOI22_X1  g0306(.A1(new_n505), .A2(new_n290), .B1(new_n506), .B2(new_n292), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n213), .A2(G33), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n337), .A2(G97), .A3(new_n338), .A4(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n496), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n304), .A2(G77), .ZN(new_n511));
  INV_X1    g0311(.A(new_n502), .ZN(new_n512));
  XNOR2_X1  g0312(.A(G97), .B(G107), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n512), .B1(new_n498), .B2(new_n513), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n511), .B1(new_n514), .B2(new_n214), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n443), .B1(new_n382), .B2(new_n383), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n290), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n292), .A2(new_n506), .ZN(new_n518));
  AND4_X1   g0318(.A1(new_n496), .A2(new_n517), .A3(new_n509), .A4(new_n518), .ZN(new_n519));
  OAI22_X1  g0319(.A1(new_n494), .A2(new_n495), .B1(new_n510), .B2(new_n519), .ZN(new_n520));
  AND2_X1   g0320(.A1(new_n507), .A2(new_n509), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n483), .A2(G190), .A3(new_n493), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n492), .B1(new_n482), .B2(new_n257), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n521), .B(new_n522), .C1(new_n523), .C2(new_n413), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n255), .A2(G274), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n213), .A2(G45), .ZN(new_n527));
  AND2_X1   g0327(.A1(new_n527), .A2(G250), .ZN(new_n528));
  AOI22_X1  g0328(.A1(new_n526), .A2(new_n487), .B1(new_n255), .B2(new_n528), .ZN(new_n529));
  NOR2_X1   g0329(.A1(G238), .A2(G1698), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n530), .B1(new_n445), .B2(G1698), .ZN(new_n531));
  AOI22_X1  g0331(.A1(new_n531), .A2(new_n267), .B1(G33), .B2(G116), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n529), .B1(new_n255), .B2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(G190), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n535), .B1(G200), .B2(new_n533), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT19), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n301), .A2(new_n537), .A3(G97), .ZN(new_n538));
  AOI22_X1  g0338(.A1(new_n500), .A2(new_n399), .B1(new_n348), .B2(new_n214), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n538), .B1(new_n539), .B2(new_n537), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n267), .A2(new_n214), .A3(G68), .ZN(new_n541));
  INV_X1    g0341(.A(new_n541), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n540), .B1(new_n542), .B2(KEYINPUT81), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT81), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n541), .A2(new_n544), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n290), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n453), .A2(new_n292), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n337), .A2(G87), .A3(new_n338), .A4(new_n508), .ZN(new_n548));
  AND3_X1   g0348(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(new_n453), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n337), .A2(new_n338), .A3(new_n508), .A4(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n546), .A2(new_n547), .A3(new_n551), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n532), .A2(new_n255), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n528), .A2(new_n255), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n554), .B1(new_n527), .B2(new_n525), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n310), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n529), .B(new_n279), .C1(new_n255), .C2(new_n532), .ZN(new_n557));
  AND2_X1   g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  AOI22_X1  g0358(.A1(new_n536), .A2(new_n549), .B1(new_n552), .B2(new_n558), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n520), .A2(new_n524), .A3(new_n559), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n337), .A2(G107), .A3(new_n338), .A4(new_n508), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n292), .A2(new_n443), .ZN(new_n562));
  XOR2_X1   g0362(.A(new_n562), .B(KEYINPUT25), .Z(new_n563));
  NAND2_X1  g0363(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n489), .A2(G264), .A3(new_n255), .ZN(new_n566));
  NOR2_X1   g0366(.A1(G250), .A2(G1698), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n567), .B1(new_n491), .B2(G1698), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n568), .A2(new_n267), .B1(G33), .B2(G294), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n488), .B(new_n566), .C1(new_n569), .C2(new_n255), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n413), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n491), .A2(G1698), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n572), .B1(G250), .B2(G1698), .ZN(new_n573));
  INV_X1    g0373(.A(G294), .ZN(new_n574));
  OAI22_X1  g0374(.A1(new_n573), .A2(new_n273), .B1(new_n264), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n257), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n576), .A2(new_n534), .A3(new_n488), .A4(new_n566), .ZN(new_n577));
  AND2_X1   g0377(.A1(new_n571), .A2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n214), .B(G87), .C1(new_n271), .C2(new_n272), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(KEYINPUT22), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT22), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n267), .A2(new_n582), .A3(new_n214), .A4(G87), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT82), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n585), .B1(new_n214), .B2(G107), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(KEYINPUT23), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT23), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n585), .B(new_n588), .C1(new_n214), .C2(G107), .ZN(new_n589));
  AOI22_X1  g0389(.A1(new_n587), .A2(new_n589), .B1(G116), .B2(new_n301), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n584), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(KEYINPUT24), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT24), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n584), .A2(new_n593), .A3(new_n590), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  AOI21_X1  g0395(.A(KEYINPUT83), .B1(new_n595), .B2(new_n290), .ZN(new_n596));
  AND3_X1   g0396(.A1(new_n584), .A2(new_n593), .A3(new_n590), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n593), .B1(new_n584), .B2(new_n590), .ZN(new_n598));
  OAI211_X1 g0398(.A(KEYINPUT83), .B(new_n290), .C1(new_n597), .C2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(new_n599), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n565), .B(new_n579), .C1(new_n596), .C2(new_n600), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n290), .B1(new_n597), .B2(new_n598), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT83), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n564), .B1(new_n604), .B2(new_n599), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n570), .A2(new_n310), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n606), .B1(G179), .B2(new_n570), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n601), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n525), .A2(new_n489), .ZN(new_n609));
  INV_X1    g0409(.A(new_n490), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n609), .B1(new_n610), .B2(G270), .ZN(new_n611));
  NOR2_X1   g0411(.A1(G257), .A2(G1698), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n268), .A2(G264), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n267), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n614), .B(new_n257), .C1(G303), .C2(new_n267), .ZN(new_n615));
  AND2_X1   g0415(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n616), .A2(new_n413), .ZN(new_n617));
  AOI21_X1  g0417(.A(G20), .B1(G33), .B2(G283), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n264), .A2(G97), .ZN(new_n619));
  INV_X1    g0419(.A(G116), .ZN(new_n620));
  AOI22_X1  g0420(.A1(new_n618), .A2(new_n619), .B1(G20), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n335), .A2(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT20), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n335), .A2(new_n621), .A3(KEYINPUT20), .ZN(new_n625));
  AOI22_X1  g0425(.A1(new_n624), .A2(new_n625), .B1(new_n620), .B2(new_n292), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n337), .A2(G116), .A3(new_n338), .A4(new_n508), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n611), .A2(new_n615), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n629), .A2(new_n534), .ZN(new_n630));
  OR3_X1    g0430(.A1(new_n617), .A2(new_n628), .A3(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT21), .ZN(new_n632));
  INV_X1    g0432(.A(new_n628), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n629), .A2(G169), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n632), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n628), .A2(new_n616), .A3(G179), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n628), .A2(KEYINPUT21), .A3(G169), .A4(new_n629), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n631), .A2(new_n635), .A3(new_n636), .A4(new_n637), .ZN(new_n638));
  NOR3_X1   g0438(.A1(new_n560), .A2(new_n608), .A3(new_n638), .ZN(new_n639));
  AND2_X1   g0439(.A1(new_n465), .A2(new_n639), .ZN(G372));
  AND2_X1   g0440(.A1(new_n552), .A2(new_n558), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n520), .A2(new_n601), .A3(new_n524), .A4(new_n559), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n604), .A2(new_n599), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n607), .B1(new_n644), .B2(new_n565), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n635), .A2(new_n636), .A3(new_n637), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n642), .B1(new_n643), .B2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n559), .ZN(new_n649));
  OAI21_X1  g0449(.A(KEYINPUT26), .B1(new_n649), .B2(new_n520), .ZN(new_n650));
  OR2_X1    g0450(.A1(new_n494), .A2(new_n495), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT26), .ZN(new_n652));
  INV_X1    g0452(.A(new_n521), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n651), .A2(new_n652), .A3(new_n559), .A4(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n650), .A2(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n465), .B1(new_n648), .B2(new_n655), .ZN(new_n656));
  XNOR2_X1  g0456(.A(new_n656), .B(KEYINPUT84), .ZN(new_n657));
  XNOR2_X1  g0457(.A(new_n435), .B(new_n429), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n367), .A2(KEYINPUT14), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(new_n365), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n370), .A2(new_n371), .ZN(new_n662));
  OR2_X1    g0462(.A1(new_n370), .A2(new_n371), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n661), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n340), .ZN(new_n665));
  OAI22_X1  g0465(.A1(new_n664), .A2(new_n665), .B1(new_n364), .B2(new_n461), .ZN(new_n666));
  INV_X1    g0466(.A(new_n437), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n415), .B1(new_n412), .B2(new_n414), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n422), .A2(KEYINPUT77), .A3(new_n423), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  AOI21_X1  g0470(.A(KEYINPUT17), .B1(new_n670), .B2(new_n398), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n667), .A2(new_n671), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n659), .B1(new_n666), .B2(new_n672), .ZN(new_n673));
  AND2_X1   g0473(.A1(new_n321), .A2(new_n323), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n312), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  OR2_X1    g0475(.A1(new_n657), .A2(new_n675), .ZN(G369));
  AOI211_X1 g0476(.A(new_n564), .B(new_n578), .C1(new_n604), .C2(new_n599), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n645), .A2(new_n677), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n213), .A2(new_n214), .A3(G13), .ZN(new_n679));
  XNOR2_X1  g0479(.A(new_n679), .B(KEYINPUT85), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT27), .ZN(new_n681));
  OR2_X1    g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n680), .A2(new_n681), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n682), .A2(new_n683), .A3(G213), .ZN(new_n684));
  INV_X1    g0484(.A(G343), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n678), .B1(new_n605), .B2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n645), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n688), .B1(new_n689), .B2(new_n687), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n687), .A2(new_n633), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n646), .A2(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n692), .B1(new_n638), .B2(new_n691), .ZN(new_n693));
  AND2_X1   g0493(.A1(new_n693), .A2(G330), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n690), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n646), .A2(new_n687), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n608), .A2(new_n696), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n697), .B1(new_n645), .B2(new_n687), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n695), .A2(new_n698), .ZN(G399));
  INV_X1    g0499(.A(new_n220), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n700), .A2(G41), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n500), .A2(new_n399), .A3(new_n620), .ZN(new_n702));
  NOR3_X1   g0502(.A1(new_n701), .A2(new_n702), .A3(new_n213), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n703), .B1(new_n228), .B2(new_n701), .ZN(new_n704));
  XOR2_X1   g0504(.A(new_n704), .B(KEYINPUT28), .Z(new_n705));
  NAND3_X1  g0505(.A1(new_n651), .A2(new_n653), .A3(new_n559), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(KEYINPUT26), .ZN(new_n707));
  OR2_X1    g0507(.A1(new_n510), .A2(new_n519), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n651), .A2(new_n708), .A3(new_n559), .A4(new_n652), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  OAI211_X1 g0510(.A(KEYINPUT29), .B(new_n687), .C1(new_n710), .C2(new_n648), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n687), .B1(new_n648), .B2(new_n655), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  OAI211_X1 g0513(.A(KEYINPUT87), .B(new_n711), .C1(new_n713), .C2(KEYINPUT29), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n483), .A2(new_n493), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n553), .A2(new_n555), .ZN(new_n716));
  AND2_X1   g0516(.A1(new_n576), .A2(new_n566), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n616), .A2(G179), .A3(new_n716), .A4(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n715), .A2(new_n718), .ZN(new_n719));
  AND2_X1   g0519(.A1(new_n719), .A2(KEYINPUT30), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n716), .A2(G179), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n715), .A2(new_n629), .A3(new_n570), .A4(new_n721), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n722), .B1(new_n719), .B2(KEYINPUT30), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n686), .B1(new_n720), .B2(new_n723), .ZN(new_n724));
  XNOR2_X1  g0524(.A(new_n724), .B(KEYINPUT31), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT86), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n726), .B1(new_n639), .B2(new_n687), .ZN(new_n727));
  AND3_X1   g0527(.A1(new_n520), .A2(new_n524), .A3(new_n559), .ZN(new_n728));
  NOR3_X1   g0528(.A1(new_n617), .A2(new_n628), .A3(new_n630), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n646), .A2(new_n729), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n728), .A2(new_n678), .A3(new_n730), .A4(new_n687), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(KEYINPUT86), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n725), .B1(new_n727), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(G330), .ZN(new_n734));
  OR2_X1    g0534(.A1(new_n711), .A2(KEYINPUT87), .ZN(new_n735));
  AND3_X1   g0535(.A1(new_n714), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n705), .B1(new_n736), .B2(G1), .ZN(G364));
  INV_X1    g0537(.A(KEYINPUT88), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n291), .A2(G20), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n213), .B1(new_n739), .B2(G45), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n738), .B1(new_n701), .B2(new_n741), .ZN(new_n742));
  OAI211_X1 g0542(.A(KEYINPUT88), .B(new_n740), .C1(new_n700), .C2(G41), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n694), .A2(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n746), .B1(G330), .B2(new_n693), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n700), .A2(new_n273), .ZN(new_n748));
  OR2_X1    g0548(.A1(G355), .A2(KEYINPUT89), .ZN(new_n749));
  NAND2_X1  g0549(.A1(G355), .A2(KEYINPUT89), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n748), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n700), .A2(new_n267), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n752), .B1(new_n229), .B2(G45), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n249), .A2(new_n252), .ZN(new_n754));
  OAI221_X1 g0554(.A(new_n751), .B1(G116), .B2(new_n220), .C1(new_n753), .C2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(G13), .A2(G33), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(G20), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n223), .B1(G20), .B2(new_n310), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n744), .B1(new_n755), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n413), .A2(G190), .ZN(new_n762));
  NOR3_X1   g0562(.A1(new_n762), .A2(new_n214), .A3(new_n279), .ZN(new_n763));
  XOR2_X1   g0563(.A(new_n763), .B(KEYINPUT90), .Z(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(new_n201), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n214), .A2(new_n279), .ZN(new_n766));
  NOR2_X1   g0566(.A1(G190), .A2(G200), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n766), .A2(G200), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(new_n534), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  OAI221_X1 g0571(.A(new_n267), .B1(new_n325), .B2(new_n768), .C1(new_n771), .C2(new_n227), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n769), .A2(G190), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n214), .A2(G179), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n775), .A2(G190), .A3(G200), .ZN(new_n776));
  OAI22_X1  g0576(.A1(new_n774), .A2(new_n202), .B1(new_n776), .B2(new_n399), .ZN(new_n777));
  NOR3_X1   g0577(.A1(new_n765), .A2(new_n772), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n775), .A2(new_n767), .ZN(new_n779));
  INV_X1    g0579(.A(G159), .ZN(new_n780));
  NOR3_X1   g0580(.A1(new_n779), .A2(KEYINPUT32), .A3(new_n780), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n775), .A2(new_n534), .A3(G200), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(G107), .ZN(new_n784));
  OAI21_X1  g0584(.A(KEYINPUT32), .B1(new_n779), .B2(new_n780), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  OAI21_X1  g0586(.A(G20), .B1(new_n762), .B2(G179), .ZN(new_n787));
  INV_X1    g0587(.A(KEYINPUT91), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n787), .A2(new_n788), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  AOI211_X1 g0593(.A(new_n781), .B(new_n786), .C1(new_n793), .C2(G97), .ZN(new_n794));
  INV_X1    g0594(.A(new_n779), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n267), .B1(new_n795), .B2(G329), .ZN(new_n796));
  INV_X1    g0596(.A(G311), .ZN(new_n797));
  INV_X1    g0597(.A(G322), .ZN(new_n798));
  INV_X1    g0598(.A(new_n763), .ZN(new_n799));
  OAI221_X1 g0599(.A(new_n796), .B1(new_n797), .B2(new_n768), .C1(new_n798), .C2(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n770), .A2(G326), .ZN(new_n801));
  INV_X1    g0601(.A(G303), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n801), .B1(new_n802), .B2(new_n776), .ZN(new_n803));
  XOR2_X1   g0603(.A(KEYINPUT33), .B(G317), .Z(new_n804));
  INV_X1    g0604(.A(G283), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n774), .A2(new_n804), .B1(new_n782), .B2(new_n805), .ZN(new_n806));
  NOR3_X1   g0606(.A1(new_n800), .A2(new_n803), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n793), .A2(G294), .ZN(new_n808));
  AOI22_X1  g0608(.A1(new_n778), .A2(new_n794), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n759), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n761), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  XOR2_X1   g0611(.A(new_n811), .B(KEYINPUT92), .Z(new_n812));
  INV_X1    g0612(.A(new_n758), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n812), .B1(new_n693), .B2(new_n813), .ZN(new_n814));
  AND2_X1   g0614(.A1(new_n747), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(G396));
  NAND2_X1  g0616(.A1(new_n810), .A2(new_n757), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n745), .B1(G77), .B2(new_n817), .ZN(new_n818));
  OAI221_X1 g0618(.A(new_n273), .B1(new_n779), .B2(new_n797), .C1(new_n799), .C2(new_n574), .ZN(new_n819));
  OAI22_X1  g0619(.A1(new_n771), .A2(new_n802), .B1(new_n782), .B2(new_n399), .ZN(new_n820));
  INV_X1    g0620(.A(new_n776), .ZN(new_n821));
  AOI211_X1 g0621(.A(new_n819), .B(new_n820), .C1(G107), .C2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n768), .ZN(new_n823));
  AOI22_X1  g0623(.A1(new_n773), .A2(G283), .B1(new_n823), .B2(G116), .ZN(new_n824));
  AOI22_X1  g0624(.A1(new_n793), .A2(G97), .B1(KEYINPUT93), .B2(new_n824), .ZN(new_n825));
  OAI211_X1 g0625(.A(new_n822), .B(new_n825), .C1(KEYINPUT93), .C2(new_n824), .ZN(new_n826));
  XOR2_X1   g0626(.A(new_n826), .B(KEYINPUT94), .Z(new_n827));
  AOI22_X1  g0627(.A1(new_n770), .A2(G137), .B1(new_n823), .B2(G159), .ZN(new_n828));
  INV_X1    g0628(.A(G143), .ZN(new_n829));
  OAI221_X1 g0629(.A(new_n828), .B1(new_n303), .B2(new_n774), .C1(new_n764), .C2(new_n829), .ZN(new_n830));
  XOR2_X1   g0630(.A(new_n830), .B(KEYINPUT34), .Z(new_n831));
  NOR2_X1   g0631(.A1(new_n782), .A2(new_n202), .ZN(new_n832));
  INV_X1    g0632(.A(G132), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n267), .B1(new_n779), .B2(new_n833), .ZN(new_n834));
  AOI211_X1 g0634(.A(new_n832), .B(new_n834), .C1(G50), .C2(new_n821), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n835), .B1(new_n201), .B2(new_n792), .ZN(new_n836));
  XNOR2_X1  g0636(.A(new_n836), .B(KEYINPUT95), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n827), .B1(new_n831), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n818), .B1(new_n838), .B2(new_n759), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n456), .A2(new_n686), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n462), .B1(new_n457), .B2(new_n840), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n461), .A2(new_n686), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n839), .B1(new_n757), .B2(new_n843), .ZN(new_n844));
  XOR2_X1   g0644(.A(new_n844), .B(KEYINPUT96), .Z(new_n845));
  XNOR2_X1  g0645(.A(new_n712), .B(new_n843), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n847), .A2(new_n734), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n745), .B1(new_n847), .B2(new_n734), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n845), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(G384));
  OAI211_X1 g0652(.A(new_n368), .B(new_n363), .C1(new_n372), .C2(new_n373), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n665), .A2(new_n687), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(KEYINPUT98), .ZN(new_n856));
  INV_X1    g0656(.A(new_n854), .ZN(new_n857));
  OAI211_X1 g0657(.A(new_n363), .B(new_n857), .C1(new_n664), .C2(new_n665), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT98), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n853), .A2(new_n859), .A3(new_n854), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n856), .A2(new_n858), .A3(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n684), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n862), .B1(new_n434), .B2(new_n379), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n863), .B1(new_n672), .B2(new_n658), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n425), .A2(new_n435), .A3(new_n863), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT37), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND4_X1  g0667(.A1(new_n425), .A2(KEYINPUT37), .A3(new_n435), .A4(new_n863), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NOR3_X1   g0669(.A1(new_n864), .A2(KEYINPUT38), .A3(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT38), .ZN(new_n871));
  AND2_X1   g0671(.A1(new_n867), .A2(new_n868), .ZN(new_n872));
  INV_X1    g0672(.A(new_n863), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n438), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n871), .B1(new_n872), .B2(new_n874), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n870), .A2(new_n875), .ZN(new_n876));
  NAND4_X1  g0676(.A1(new_n733), .A2(new_n861), .A3(new_n843), .A4(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT40), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT101), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n877), .A2(KEYINPUT101), .A3(new_n878), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  AND3_X1   g0683(.A1(new_n733), .A2(new_n861), .A3(new_n843), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n864), .A2(new_n869), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT100), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n871), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n872), .A2(new_n874), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n888), .A2(KEYINPUT100), .A3(KEYINPUT38), .ZN(new_n889));
  AND3_X1   g0689(.A1(new_n887), .A2(KEYINPUT40), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n884), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n883), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n465), .A2(new_n733), .ZN(new_n893));
  OR2_X1    g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n892), .A2(new_n893), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n894), .A2(G330), .A3(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT39), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n887), .A2(new_n897), .A3(new_n889), .ZN(new_n898));
  OAI21_X1  g0698(.A(KEYINPUT39), .B1(new_n870), .B2(new_n875), .ZN(new_n899));
  AND2_X1   g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n374), .A2(new_n340), .A3(new_n687), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT99), .ZN(new_n902));
  OR2_X1    g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n901), .A2(new_n902), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n900), .A2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(new_n842), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n907), .B1(new_n712), .B2(new_n841), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n908), .A2(new_n861), .A3(new_n876), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n659), .A2(new_n684), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n906), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n464), .B1(new_n714), .B2(new_n735), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n912), .A2(new_n675), .ZN(new_n913));
  XOR2_X1   g0713(.A(new_n911), .B(new_n913), .Z(new_n914));
  NAND2_X1  g0714(.A1(new_n896), .A2(new_n914), .ZN(new_n915));
  OR2_X1    g0715(.A1(new_n915), .A2(KEYINPUT102), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(KEYINPUT102), .ZN(new_n917));
  OR2_X1    g0717(.A1(new_n896), .A2(new_n914), .ZN(new_n918));
  OAI21_X1  g0718(.A(G1), .B1(new_n291), .B2(G20), .ZN(new_n919));
  NAND4_X1  g0719(.A1(new_n916), .A2(new_n917), .A3(new_n918), .A4(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n385), .A2(G77), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n245), .B1(new_n229), .B2(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n922), .A2(G1), .A3(new_n291), .ZN(new_n923));
  AOI211_X1 g0723(.A(new_n620), .B(new_n225), .C1(new_n503), .C2(KEYINPUT35), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n924), .B1(KEYINPUT35), .B2(new_n503), .ZN(new_n925));
  XNOR2_X1  g0725(.A(KEYINPUT97), .B(KEYINPUT36), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n925), .B(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n920), .A2(new_n923), .A3(new_n927), .ZN(G367));
  INV_X1    g0728(.A(new_n752), .ZN(new_n929));
  OAI221_X1 g0729(.A(new_n760), .B1(new_n220), .B2(new_n453), .C1(new_n929), .C2(new_n238), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n745), .A2(new_n930), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n931), .B(KEYINPUT107), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n793), .A2(G68), .ZN(new_n933));
  INV_X1    g0733(.A(G137), .ZN(new_n934));
  OAI22_X1  g0734(.A1(new_n768), .A2(new_n227), .B1(new_n779), .B2(new_n934), .ZN(new_n935));
  AOI211_X1 g0735(.A(new_n273), .B(new_n935), .C1(G150), .C2(new_n763), .ZN(new_n936));
  AOI22_X1  g0736(.A1(G143), .A2(new_n770), .B1(new_n773), .B2(G159), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n782), .A2(new_n325), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n938), .B1(G58), .B2(new_n821), .ZN(new_n939));
  NAND4_X1  g0739(.A1(new_n933), .A2(new_n936), .A3(new_n937), .A4(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(G317), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n273), .B1(new_n779), .B2(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n942), .B1(G97), .B2(new_n783), .ZN(new_n943));
  AOI22_X1  g0743(.A1(new_n793), .A2(G107), .B1(KEYINPUT108), .B2(new_n943), .ZN(new_n944));
  OAI22_X1  g0744(.A1(new_n774), .A2(new_n574), .B1(new_n768), .B2(new_n805), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n945), .B1(G311), .B2(new_n770), .ZN(new_n946));
  OAI211_X1 g0746(.A(new_n944), .B(new_n946), .C1(KEYINPUT108), .C2(new_n943), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n821), .A2(KEYINPUT46), .A3(G116), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT46), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n949), .B1(new_n776), .B2(new_n620), .ZN(new_n950));
  OAI211_X1 g0750(.A(new_n948), .B(new_n950), .C1(new_n764), .C2(new_n802), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n940), .B1(new_n947), .B2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT47), .ZN(new_n953));
  OR2_X1    g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n810), .B1(new_n952), .B2(new_n953), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n932), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  OR3_X1    g0756(.A1(new_n642), .A2(new_n549), .A3(new_n687), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT103), .ZN(new_n958));
  OR2_X1    g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n559), .B1(new_n549), .B2(new_n687), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n957), .A2(new_n958), .A3(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n956), .B1(new_n963), .B2(new_n813), .ZN(new_n964));
  OAI211_X1 g0764(.A(new_n520), .B(new_n524), .C1(new_n521), .C2(new_n687), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n651), .A2(new_n653), .A3(new_n686), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  AOI22_X1  g0767(.A1(new_n967), .A2(new_n645), .B1(new_n651), .B2(new_n708), .ZN(new_n968));
  AOI21_X1  g0768(.A(KEYINPUT42), .B1(new_n967), .B2(new_n697), .ZN(new_n969));
  AND3_X1   g0769(.A1(new_n967), .A2(KEYINPUT42), .A3(new_n697), .ZN(new_n970));
  OAI22_X1  g0770(.A1(new_n968), .A2(new_n686), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  OR3_X1    g0771(.A1(new_n971), .A2(KEYINPUT43), .A3(new_n963), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n962), .B(KEYINPUT43), .ZN(new_n973));
  AND2_X1   g0773(.A1(new_n973), .A2(new_n971), .ZN(new_n974));
  OR2_X1    g0774(.A1(new_n974), .A2(KEYINPUT104), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(KEYINPUT104), .ZN(new_n976));
  INV_X1    g0776(.A(new_n695), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n977), .A2(new_n967), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT105), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND4_X1  g0780(.A1(new_n972), .A2(new_n975), .A3(new_n976), .A4(new_n980), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n978), .A2(new_n979), .ZN(new_n982));
  INV_X1    g0782(.A(new_n982), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n981), .B(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n698), .A2(new_n967), .ZN(new_n985));
  XOR2_X1   g0785(.A(new_n985), .B(KEYINPUT45), .Z(new_n986));
  NOR2_X1   g0786(.A1(new_n698), .A2(new_n967), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT44), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(new_n977), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n986), .A2(new_n695), .A3(new_n988), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(new_n697), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT106), .ZN(new_n994));
  INV_X1    g0794(.A(new_n696), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n993), .B1(new_n694), .B2(new_n994), .C1(new_n690), .C2(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n694), .A2(new_n994), .ZN(new_n997));
  XOR2_X1   g0797(.A(new_n996), .B(new_n997), .Z(new_n998));
  NAND2_X1  g0798(.A1(new_n998), .A2(new_n736), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n736), .B1(new_n992), .B2(new_n999), .ZN(new_n1000));
  XOR2_X1   g0800(.A(new_n701), .B(KEYINPUT41), .Z(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n741), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n964), .B1(new_n984), .B2(new_n1003), .ZN(G387));
  NAND2_X1  g0804(.A1(new_n998), .A2(new_n741), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n764), .A2(new_n941), .B1(new_n802), .B2(new_n768), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1006), .ZN(new_n1007));
  OR2_X1    g0807(.A1(new_n1007), .A2(KEYINPUT111), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1007), .A2(KEYINPUT111), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(G311), .A2(new_n773), .B1(new_n770), .B2(G322), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1008), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT48), .ZN(new_n1012));
  OR2_X1    g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(new_n793), .A2(G283), .B1(G294), .B2(new_n821), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1013), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  XOR2_X1   g0816(.A(new_n1016), .B(KEYINPUT49), .Z(new_n1017));
  OR2_X1    g0817(.A1(new_n1017), .A2(KEYINPUT112), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1017), .A2(KEYINPUT112), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n782), .A2(new_n620), .ZN(new_n1020));
  AOI211_X1 g0820(.A(new_n267), .B(new_n1020), .C1(G326), .C2(new_n795), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1018), .A2(new_n1019), .A3(new_n1021), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n792), .A2(new_n453), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n823), .A2(G68), .B1(new_n763), .B2(G50), .ZN(new_n1024));
  OAI211_X1 g0824(.A(new_n1024), .B(new_n267), .C1(new_n303), .C2(new_n779), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n771), .A2(new_n780), .B1(new_n782), .B2(new_n506), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n774), .A2(new_n300), .B1(new_n325), .B2(new_n776), .ZN(new_n1027));
  NOR4_X1   g0827(.A1(new_n1023), .A2(new_n1025), .A3(new_n1026), .A4(new_n1027), .ZN(new_n1028));
  XOR2_X1   g0828(.A(new_n1028), .B(KEYINPUT110), .Z(new_n1029));
  AOI21_X1  g0829(.A(new_n810), .B1(new_n1022), .B2(new_n1029), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n748), .A2(new_n702), .B1(new_n443), .B2(new_n700), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n235), .A2(new_n252), .ZN(new_n1032));
  AOI211_X1 g0832(.A(G45), .B(new_n702), .C1(G68), .C2(G77), .ZN(new_n1033));
  XOR2_X1   g0833(.A(KEYINPUT109), .B(KEYINPUT50), .Z(new_n1034));
  OR3_X1    g0834(.A1(new_n1034), .A2(G50), .A3(new_n300), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1034), .B1(G50), .B2(new_n300), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1033), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1037), .A2(new_n752), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1031), .B1(new_n1032), .B2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n744), .B1(new_n1039), .B2(new_n760), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1040), .B1(new_n690), .B2(new_n813), .ZN(new_n1041));
  XOR2_X1   g0841(.A(new_n701), .B(KEYINPUT113), .Z(new_n1042));
  NAND2_X1  g0842(.A1(new_n999), .A2(new_n1042), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n998), .A2(new_n736), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n1005), .B1(new_n1030), .B2(new_n1041), .C1(new_n1043), .C2(new_n1044), .ZN(G393));
  NOR2_X1   g0845(.A1(new_n243), .A2(new_n929), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n760), .B1(new_n506), .B2(new_n220), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n745), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n774), .A2(new_n227), .B1(new_n300), .B2(new_n768), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1049), .B1(new_n793), .B2(G77), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1050), .B(KEYINPUT114), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n770), .A2(G150), .B1(G159), .B2(new_n763), .ZN(new_n1052));
  XOR2_X1   g0852(.A(new_n1052), .B(KEYINPUT51), .Z(new_n1053));
  OAI221_X1 g0853(.A(new_n267), .B1(new_n779), .B2(new_n829), .C1(new_n399), .C2(new_n782), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(G68), .B2(new_n821), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1051), .A2(new_n1053), .A3(new_n1055), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n774), .A2(new_n802), .B1(new_n768), .B2(new_n574), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1057), .B1(new_n793), .B2(G116), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT115), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n770), .A2(G317), .B1(G311), .B2(new_n763), .ZN(new_n1060));
  XOR2_X1   g0860(.A(new_n1060), .B(KEYINPUT52), .Z(new_n1061));
  OAI211_X1 g0861(.A(new_n784), .B(new_n273), .C1(new_n798), .C2(new_n779), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1062), .B1(G283), .B2(new_n821), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1056), .B1(new_n1059), .B2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1048), .B1(new_n1065), .B2(new_n759), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1066), .B1(new_n967), .B2(new_n813), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1067), .B1(new_n992), .B2(new_n740), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n992), .A2(new_n999), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n1042), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n992), .A2(new_n999), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1068), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1073), .ZN(G390));
  OAI21_X1  g0874(.A(new_n687), .B1(new_n710), .B2(new_n648), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n907), .B1(new_n1075), .B2(new_n841), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1076), .A2(new_n861), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n905), .ZN(new_n1078));
  NAND4_X1  g0878(.A1(new_n1077), .A2(new_n1078), .A3(new_n887), .A4(new_n889), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n843), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n731), .A2(KEYINPUT86), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n560), .A2(new_n608), .ZN(new_n1082));
  NAND4_X1  g0882(.A1(new_n1082), .A2(new_n726), .A3(new_n730), .A4(new_n687), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1080), .B1(new_n1084), .B2(new_n725), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1085), .A2(G330), .A3(new_n861), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n905), .B1(new_n908), .B2(new_n861), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n1079), .B(new_n1086), .C1(new_n1087), .C2(new_n900), .ZN(new_n1088));
  AND4_X1   g0888(.A1(G330), .A2(new_n733), .A3(new_n843), .A4(new_n861), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n908), .A2(new_n861), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(new_n1090), .A2(new_n1078), .B1(new_n898), .B2(new_n899), .ZN(new_n1091));
  NAND4_X1  g0891(.A1(new_n887), .A2(new_n903), .A3(new_n904), .A4(new_n889), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(new_n861), .B2(new_n1076), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1089), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1088), .A2(new_n1094), .A3(new_n741), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n817), .A2(new_n451), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n744), .A2(new_n1096), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(KEYINPUT54), .B(G143), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n774), .A2(new_n934), .B1(new_n768), .B2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1099), .B1(new_n793), .B2(G159), .ZN(new_n1100));
  XOR2_X1   g0900(.A(new_n1100), .B(KEYINPUT116), .Z(new_n1101));
  OAI21_X1  g0901(.A(new_n267), .B1(new_n782), .B2(new_n227), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(new_n1102), .B(KEYINPUT117), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n795), .A2(G125), .B1(new_n763), .B2(G132), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n770), .A2(G128), .ZN(new_n1105));
  OAI21_X1  g0905(.A(KEYINPUT53), .B1(new_n776), .B2(new_n303), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1104), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  NOR3_X1   g0907(.A1(new_n776), .A2(KEYINPUT53), .A3(new_n303), .ZN(new_n1108));
  NOR3_X1   g0908(.A1(new_n1103), .A2(new_n1107), .A3(new_n1108), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n792), .A2(new_n325), .B1(new_n620), .B2(new_n799), .ZN(new_n1110));
  XOR2_X1   g0910(.A(new_n1110), .B(KEYINPUT119), .Z(new_n1111));
  OAI22_X1  g0911(.A1(new_n782), .A2(new_n202), .B1(new_n779), .B2(new_n574), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(new_n1112), .B(KEYINPUT118), .ZN(new_n1113));
  OAI22_X1  g0913(.A1(new_n443), .A2(new_n774), .B1(new_n771), .B2(new_n805), .ZN(new_n1114));
  OAI221_X1 g0914(.A(new_n273), .B1(new_n768), .B2(new_n506), .C1(new_n399), .C2(new_n776), .ZN(new_n1115));
  NOR3_X1   g0915(.A1(new_n1113), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n1101), .A2(new_n1109), .B1(new_n1111), .B2(new_n1116), .ZN(new_n1117));
  OAI221_X1 g0917(.A(new_n1097), .B1(new_n810), .B2(new_n1117), .C1(new_n900), .C2(new_n757), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1095), .A2(new_n1118), .ZN(new_n1119));
  XOR2_X1   g0919(.A(new_n1119), .B(KEYINPUT120), .Z(new_n1120));
  AOI21_X1  g0920(.A(new_n861), .B1(new_n1085), .B2(G330), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n908), .B1(new_n1089), .B2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n733), .A2(G330), .A3(new_n843), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n861), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1076), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1125), .A2(new_n1126), .A3(new_n1086), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1122), .A2(new_n1127), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n734), .A2(new_n464), .ZN(new_n1129));
  NOR3_X1   g0929(.A1(new_n912), .A2(new_n1129), .A3(new_n675), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1088), .A2(new_n1094), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NAND4_X1  g0933(.A1(new_n1128), .A2(new_n1094), .A3(new_n1088), .A4(new_n1130), .ZN(new_n1134));
  AND3_X1   g0934(.A1(new_n1133), .A2(new_n1042), .A3(new_n1134), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1120), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(G378));
  INV_X1    g0937(.A(new_n911), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n309), .A2(new_n862), .ZN(new_n1139));
  OR2_X1    g0939(.A1(new_n324), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n324), .A2(new_n1139), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1142));
  AND3_X1   g0942(.A1(new_n1140), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1142), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(G330), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1146), .B1(new_n884), .B2(new_n890), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1145), .B1(new_n883), .B2(new_n1147), .ZN(new_n1148));
  AND3_X1   g0948(.A1(new_n877), .A2(KEYINPUT101), .A3(new_n878), .ZN(new_n1149));
  AOI21_X1  g0949(.A(KEYINPUT101), .B1(new_n877), .B2(new_n878), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n1145), .B(new_n1147), .C1(new_n1149), .C2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1138), .B1(new_n1148), .B2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1147), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1145), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1156), .A2(new_n911), .A3(new_n1151), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1153), .A2(KEYINPUT123), .A3(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n911), .B1(new_n1156), .B2(new_n1151), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT123), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1158), .A2(new_n741), .A3(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1145), .A2(new_n756), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n745), .B1(G50), .B2(new_n817), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n506), .A2(new_n774), .B1(new_n771), .B2(new_n620), .ZN(new_n1165));
  OAI22_X1  g0965(.A1(new_n201), .A2(new_n782), .B1(new_n776), .B2(new_n325), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n273), .A2(new_n251), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1168), .B1(G283), .B2(new_n795), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(new_n823), .A2(new_n550), .B1(new_n763), .B2(G107), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n1167), .A2(new_n933), .A3(new_n1169), .A4(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT58), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n1168), .B(new_n227), .C1(G33), .C2(G41), .ZN(new_n1174));
  AND2_X1   g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n770), .A2(G125), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1176), .B1(new_n776), .B2(new_n1098), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n823), .A2(G137), .B1(new_n763), .B2(G128), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1178), .B1(new_n833), .B2(new_n774), .ZN(new_n1179));
  AOI211_X1 g0979(.A(new_n1177), .B(new_n1179), .C1(G150), .C2(new_n793), .ZN(new_n1180));
  XNOR2_X1  g0980(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n1181));
  XOR2_X1   g0981(.A(new_n1180), .B(new_n1181), .Z(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1183), .A2(KEYINPUT122), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n783), .A2(G159), .ZN(new_n1185));
  AOI211_X1 g0985(.A(G33), .B(G41), .C1(new_n795), .C2(G124), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1184), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n1183), .A2(KEYINPUT122), .ZN(new_n1188));
  OAI221_X1 g0988(.A(new_n1175), .B1(new_n1172), .B2(new_n1171), .C1(new_n1187), .C2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1164), .B1(new_n1189), .B2(new_n759), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1163), .A2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1162), .A2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1134), .A2(new_n1130), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1158), .A2(new_n1193), .A3(new_n1161), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT57), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1195), .B1(new_n1134), .B2(new_n1130), .ZN(new_n1197));
  AND3_X1   g0997(.A1(new_n1156), .A2(new_n911), .A3(new_n1151), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1197), .B1(new_n1198), .B2(new_n1159), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1199), .A2(new_n1042), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1192), .B1(new_n1196), .B2(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(G375));
  NAND2_X1  g1003(.A1(new_n1128), .A2(new_n741), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n745), .B1(G68), .B2(new_n817), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n201), .A2(new_n782), .B1(new_n776), .B2(new_n780), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n764), .A2(new_n934), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n833), .A2(new_n771), .B1(new_n774), .B2(new_n1098), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n273), .B1(new_n795), .B2(G128), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1209), .B1(new_n303), .B2(new_n768), .ZN(new_n1210));
  OR4_X1    g1010(.A1(new_n1206), .A2(new_n1207), .A3(new_n1208), .A4(new_n1210), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n792), .A2(new_n227), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n799), .A2(new_n805), .B1(new_n768), .B2(new_n443), .ZN(new_n1213));
  AOI211_X1 g1013(.A(new_n267), .B(new_n1213), .C1(G303), .C2(new_n795), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n938), .B1(G116), .B2(new_n773), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n770), .A2(G294), .B1(new_n821), .B2(G97), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1214), .A2(new_n1215), .A3(new_n1216), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n1211), .A2(new_n1212), .B1(new_n1217), .B2(new_n1023), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1205), .B1(new_n1218), .B2(new_n759), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1219), .B1(new_n861), .B2(new_n757), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1204), .A2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1131), .A2(new_n1002), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1222), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  XOR2_X1   g1025(.A(new_n1225), .B(KEYINPUT124), .Z(G381));
  INV_X1    g1026(.A(G387), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(G393), .A2(G396), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1227), .A2(new_n851), .A3(new_n1073), .A4(new_n1228), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1135), .A2(new_n1119), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1230), .ZN(new_n1231));
  OR4_X1    g1031(.A1(G375), .A2(new_n1229), .A3(G381), .A4(new_n1231), .ZN(G407));
  NAND2_X1  g1032(.A1(new_n685), .A2(G213), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1233), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1202), .A2(new_n1230), .A3(new_n1234), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(G407), .A2(G213), .A3(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT125), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(G407), .A2(KEYINPUT125), .A3(G213), .A4(new_n1235), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1238), .A2(new_n1239), .ZN(G409));
  NAND2_X1  g1040(.A1(new_n1131), .A2(KEYINPUT60), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1241), .B1(new_n1130), .B2(new_n1128), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1223), .A2(KEYINPUT60), .A3(new_n1131), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1242), .A2(new_n1042), .A3(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1244), .A2(new_n1222), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1245), .A2(new_n851), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1244), .A2(G384), .A3(new_n1222), .ZN(new_n1247));
  AND2_X1   g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1200), .B1(new_n1195), .B2(new_n1194), .ZN(new_n1249));
  NOR3_X1   g1049(.A1(new_n1249), .A2(new_n1136), .A3(new_n1192), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n740), .B1(new_n1153), .B2(new_n1157), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1251), .B1(new_n1163), .B2(new_n1190), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1158), .A2(new_n1193), .A3(new_n1002), .A4(new_n1161), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1231), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1254));
  OAI211_X1 g1054(.A(new_n1233), .B(new_n1248), .C1(new_n1250), .C2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1255), .A2(KEYINPUT62), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT61), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1234), .A2(G2897), .ZN(new_n1258));
  AND3_X1   g1058(.A1(new_n1246), .A2(new_n1247), .A3(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1258), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1254), .B1(new_n1202), .B2(G378), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1261), .B1(new_n1262), .B2(new_n1234), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1196), .A2(new_n1201), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1192), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1264), .A2(G378), .A3(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1254), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT62), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1268), .A2(new_n1269), .A3(new_n1233), .A4(new_n1248), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1256), .A2(new_n1257), .A3(new_n1263), .A4(new_n1270), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(G387), .A2(new_n1073), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(new_n1273));
  XNOR2_X1  g1073(.A(G393), .B(new_n815), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(G387), .A2(new_n1073), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT126), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1273), .A2(new_n1275), .A3(new_n1276), .A4(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1276), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1277), .B1(G387), .B2(new_n1073), .ZN(new_n1280));
  OAI22_X1  g1080(.A1(new_n1279), .A2(new_n1272), .B1(new_n1280), .B2(new_n1274), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1278), .A2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1271), .A2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT63), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1283), .B1(new_n1255), .B2(new_n1285), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1268), .A2(KEYINPUT63), .A3(new_n1233), .A4(new_n1248), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1286), .A2(new_n1257), .A3(new_n1287), .A4(new_n1263), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1284), .A2(new_n1288), .ZN(G405));
  NAND2_X1  g1089(.A1(new_n1248), .A2(KEYINPUT127), .ZN(new_n1290));
  XNOR2_X1  g1090(.A(new_n1282), .B(new_n1290), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1248), .A2(KEYINPUT127), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(G375), .A2(new_n1230), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1292), .B1(new_n1293), .B2(new_n1266), .ZN(new_n1294));
  XNOR2_X1  g1094(.A(new_n1291), .B(new_n1294), .ZN(G402));
endmodule


