

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749;

  AND2_X1 U377 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U378 ( .A(n521), .B(n520), .ZN(n676) );
  INV_X1 U379 ( .A(n454), .ZN(n357) );
  INV_X1 U380 ( .A(n509), .ZN(n627) );
  XNOR2_X1 U381 ( .A(n596), .B(n504), .ZN(n509) );
  NOR2_X1 U382 ( .A1(n706), .A2(G902), .ZN(n503) );
  XNOR2_X1 U383 ( .A(n359), .B(n433), .ZN(n467) );
  XNOR2_X1 U384 ( .A(n441), .B(n410), .ZN(n472) );
  XOR2_X1 U385 ( .A(G101), .B(G119), .Z(n359) );
  XNOR2_X1 U386 ( .A(KEYINPUT3), .B(KEYINPUT90), .ZN(n433) );
  INV_X2 U387 ( .A(G953), .ZN(n736) );
  NAND2_X1 U388 ( .A1(n649), .A2(n735), .ZN(n373) );
  XNOR2_X2 U389 ( .A(n547), .B(KEYINPUT45), .ZN(n649) );
  OR2_X2 U390 ( .A1(n559), .A2(n538), .ZN(n517) );
  XNOR2_X2 U391 ( .A(n358), .B(n357), .ZN(n534) );
  NAND2_X1 U392 ( .A1(n590), .A2(n453), .ZN(n358) );
  XNOR2_X2 U393 ( .A(n513), .B(KEYINPUT70), .ZN(n533) );
  XNOR2_X2 U394 ( .A(G143), .B(G128), .ZN(n441) );
  NAND2_X2 U395 ( .A1(n528), .A2(n505), .ZN(n506) );
  NOR2_X2 U396 ( .A1(n373), .A2(n656), .ZN(n372) );
  NOR2_X2 U397 ( .A1(n531), .A2(n530), .ZN(n693) );
  NOR2_X2 U398 ( .A1(n583), .A2(n585), .ZN(n597) );
  XNOR2_X1 U399 ( .A(n470), .B(n471), .ZN(n392) );
  INV_X1 U400 ( .A(G469), .ZN(n388) );
  NAND2_X1 U401 ( .A1(n746), .A2(n687), .ZN(n525) );
  XNOR2_X1 U402 ( .A(n517), .B(n516), .ZN(n519) );
  NAND2_X1 U403 ( .A1(n385), .A2(n384), .ZN(n559) );
  XNOR2_X1 U404 ( .A(n459), .B(n458), .ZN(n507) );
  AND2_X1 U405 ( .A1(n383), .A2(n386), .ZN(n385) );
  XNOR2_X1 U406 ( .A(n395), .B(KEYINPUT39), .ZN(n634) );
  OR2_X1 U407 ( .A1(n533), .A2(n360), .ZN(n384) );
  NOR2_X1 U408 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U409 ( .A(n413), .B(n412), .ZN(n531) );
  NOR2_X1 U410 ( .A1(G953), .A2(G237), .ZN(n466) );
  OR2_X1 U411 ( .A1(n676), .A2(n525), .ZN(n526) );
  INV_X1 U412 ( .A(G134), .ZN(n410) );
  NOR2_X1 U413 ( .A1(n531), .A2(n529), .ZN(n561) );
  XNOR2_X1 U414 ( .A(G113), .B(G104), .ZN(n419) );
  XOR2_X1 U415 ( .A(G116), .B(G107), .Z(n432) );
  XNOR2_X1 U416 ( .A(n730), .B(n445), .ZN(n672) );
  AND2_X1 U417 ( .A1(n747), .A2(n748), .ZN(n625) );
  XNOR2_X1 U418 ( .A(n744), .B(n375), .ZN(n374) );
  AND2_X1 U419 ( .A1(n619), .A2(n377), .ZN(n376) );
  INV_X1 U420 ( .A(KEYINPUT86), .ZN(n375) );
  XNOR2_X1 U421 ( .A(G113), .B(KEYINPUT5), .ZN(n460) );
  XOR2_X1 U422 ( .A(KEYINPUT98), .B(KEYINPUT99), .Z(n461) );
  XNOR2_X1 U423 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U424 ( .A(G137), .B(G116), .ZN(n463) );
  NOR2_X1 U425 ( .A1(n584), .A2(n585), .ZN(n608) );
  XNOR2_X1 U426 ( .A(n508), .B(n478), .ZN(n609) );
  XNOR2_X1 U427 ( .A(n382), .B(n381), .ZN(n486) );
  INV_X1 U428 ( .A(KEYINPUT8), .ZN(n381) );
  NAND2_X1 U429 ( .A1(n736), .A2(G234), .ZN(n382) );
  XNOR2_X1 U430 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U431 ( .A(G140), .B(G137), .ZN(n495) );
  INV_X1 U432 ( .A(G110), .ZN(n497) );
  XNOR2_X1 U433 ( .A(G104), .B(G101), .ZN(n498) );
  NAND2_X1 U434 ( .A1(n672), .A2(n656), .ZN(n368) );
  NAND2_X1 U435 ( .A1(n714), .A2(n474), .ZN(n413) );
  XNOR2_X1 U436 ( .A(n424), .B(n423), .ZN(n710) );
  XNOR2_X1 U437 ( .A(n422), .B(n421), .ZN(n423) );
  NAND2_X2 U438 ( .A1(n371), .A2(n661), .ZN(n716) );
  INV_X1 U439 ( .A(KEYINPUT48), .ZN(n389) );
  XNOR2_X1 U440 ( .A(n414), .B(G125), .ZN(n438) );
  INV_X1 U441 ( .A(G146), .ZN(n414) );
  NAND2_X1 U442 ( .A1(n597), .A2(n627), .ZN(n513) );
  NAND2_X1 U443 ( .A1(G234), .A2(G237), .ZN(n450) );
  XNOR2_X1 U444 ( .A(n428), .B(n427), .ZN(n529) );
  XNOR2_X1 U445 ( .A(n426), .B(n425), .ZN(n427) );
  NOR2_X1 U446 ( .A1(G902), .A2(n710), .ZN(n428) );
  XNOR2_X1 U447 ( .A(n465), .B(n464), .ZN(n469) );
  XOR2_X1 U448 ( .A(KEYINPUT67), .B(KEYINPUT24), .Z(n481) );
  XNOR2_X1 U449 ( .A(n438), .B(n415), .ZN(n479) );
  INV_X1 U450 ( .A(KEYINPUT10), .ZN(n415) );
  XOR2_X1 U451 ( .A(G140), .B(KEYINPUT12), .Z(n418) );
  BUF_X1 U452 ( .A(n649), .Z(n721) );
  INV_X1 U453 ( .A(n660), .ZN(n369) );
  XNOR2_X1 U454 ( .A(n396), .B(KEYINPUT107), .ZN(n629) );
  AND2_X1 U455 ( .A1(n693), .A2(n609), .ZN(n397) );
  NOR2_X1 U456 ( .A1(n620), .A2(n394), .ZN(n393) );
  XNOR2_X1 U457 ( .A(n457), .B(KEYINPUT69), .ZN(n458) );
  XNOR2_X1 U458 ( .A(n492), .B(n493), .ZN(n398) );
  OR2_X1 U459 ( .A1(n717), .A2(G902), .ZN(n399) );
  XNOR2_X1 U460 ( .A(n434), .B(n435), .ZN(n730) );
  XNOR2_X1 U461 ( .A(n380), .B(n379), .ZN(n714) );
  XNOR2_X1 U462 ( .A(n411), .B(n406), .ZN(n379) );
  XNOR2_X1 U463 ( .A(n409), .B(n405), .ZN(n380) );
  XNOR2_X1 U464 ( .A(n370), .B(n502), .ZN(n706) );
  AND2_X1 U465 ( .A1(n367), .A2(n365), .ZN(n712) );
  AND2_X1 U466 ( .A1(n366), .A2(n365), .ZN(n675) );
  OR2_X1 U467 ( .A1(n514), .A2(n387), .ZN(n360) );
  AND2_X1 U468 ( .A1(n600), .A2(n601), .ZN(n361) );
  AND2_X1 U469 ( .A1(n376), .A2(n374), .ZN(n362) );
  XNOR2_X1 U470 ( .A(n710), .B(KEYINPUT59), .ZN(n363) );
  XOR2_X1 U471 ( .A(n672), .B(n671), .Z(n364) );
  AND2_X1 U472 ( .A1(n666), .A2(G953), .ZN(n720) );
  INV_X1 U473 ( .A(n720), .ZN(n365) );
  XNOR2_X1 U474 ( .A(n673), .B(n364), .ZN(n366) );
  XNOR2_X1 U475 ( .A(n711), .B(n363), .ZN(n367) );
  XNOR2_X2 U476 ( .A(n368), .B(n446), .ZN(n632) );
  NOR2_X1 U477 ( .A1(n369), .A2(n373), .ZN(n655) );
  NAND2_X1 U478 ( .A1(n649), .A2(n645), .ZN(n660) );
  XNOR2_X1 U479 ( .A(n370), .B(n473), .ZN(n663) );
  XNOR2_X2 U480 ( .A(n734), .B(G146), .ZN(n370) );
  NAND2_X1 U481 ( .A1(n372), .A2(n660), .ZN(n371) );
  XNOR2_X2 U482 ( .A(n615), .B(n614), .ZN(n744) );
  NAND2_X1 U483 ( .A1(n378), .A2(n562), .ZN(n377) );
  OR2_X1 U484 ( .A1(n617), .A2(KEYINPUT81), .ZN(n378) );
  XNOR2_X2 U485 ( .A(KEYINPUT40), .B(n621), .ZN(n747) );
  NAND2_X1 U486 ( .A1(n533), .A2(n387), .ZN(n383) );
  NAND2_X1 U487 ( .A1(n514), .A2(n387), .ZN(n386) );
  INV_X1 U488 ( .A(KEYINPUT33), .ZN(n387) );
  XNOR2_X2 U489 ( .A(n503), .B(n388), .ZN(n596) );
  NAND2_X2 U490 ( .A1(n647), .A2(n646), .ZN(n648) );
  XNOR2_X2 U491 ( .A(n390), .B(n389), .ZN(n647) );
  NAND2_X1 U492 ( .A1(n391), .A2(n362), .ZN(n390) );
  XNOR2_X1 U493 ( .A(n625), .B(KEYINPUT46), .ZN(n391) );
  XNOR2_X2 U494 ( .A(n472), .B(n392), .ZN(n734) );
  XNOR2_X2 U495 ( .A(KEYINPUT66), .B(G131), .ZN(n471) );
  XNOR2_X2 U496 ( .A(KEYINPUT64), .B(KEYINPUT4), .ZN(n470) );
  NAND2_X1 U497 ( .A1(n600), .A2(n393), .ZN(n395) );
  INV_X1 U498 ( .A(n601), .ZN(n394) );
  NAND2_X1 U499 ( .A1(n634), .A2(n693), .ZN(n621) );
  NAND2_X1 U500 ( .A1(n608), .A2(n397), .ZN(n396) );
  XNOR2_X2 U501 ( .A(n399), .B(n398), .ZN(n583) );
  XNOR2_X1 U502 ( .A(n488), .B(n487), .ZN(n489) );
  AND2_X1 U503 ( .A1(n466), .A2(G210), .ZN(n400) );
  XNOR2_X1 U504 ( .A(G110), .B(KEYINPUT16), .ZN(n401) );
  XNOR2_X1 U505 ( .A(n525), .B(KEYINPUT87), .ZN(n523) );
  INV_X1 U506 ( .A(KEYINPUT71), .ZN(n462) );
  XNOR2_X1 U507 ( .A(n467), .B(n400), .ZN(n468) );
  INV_X1 U508 ( .A(KEYINPUT30), .ZN(n594) );
  INV_X1 U509 ( .A(G475), .ZN(n425) );
  XNOR2_X1 U510 ( .A(n469), .B(n468), .ZN(n473) );
  INV_X1 U511 ( .A(KEYINPUT100), .ZN(n407) );
  XNOR2_X1 U512 ( .A(n595), .B(n594), .ZN(n599) );
  INV_X1 U513 ( .A(KEYINPUT22), .ZN(n457) );
  XNOR2_X1 U514 ( .A(n654), .B(n653), .ZN(G75) );
  XNOR2_X1 U515 ( .A(G902), .B(KEYINPUT15), .ZN(n656) );
  NAND2_X1 U516 ( .A1(G234), .A2(n656), .ZN(n402) );
  XNOR2_X1 U517 ( .A(KEYINPUT20), .B(n402), .ZN(n491) );
  NAND2_X1 U518 ( .A1(n491), .A2(G221), .ZN(n403) );
  XOR2_X1 U519 ( .A(KEYINPUT21), .B(n403), .Z(n404) );
  XNOR2_X1 U520 ( .A(n404), .B(KEYINPUT97), .ZN(n585) );
  XOR2_X1 U521 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n406) );
  NAND2_X1 U522 ( .A1(G217), .A2(n486), .ZN(n405) );
  XNOR2_X1 U523 ( .A(n432), .B(G122), .ZN(n408) );
  INV_X1 U524 ( .A(n472), .ZN(n411) );
  INV_X1 U525 ( .A(G902), .ZN(n474) );
  XOR2_X1 U526 ( .A(KEYINPUT101), .B(G478), .Z(n412) );
  INV_X1 U527 ( .A(n479), .ZN(n416) );
  XNOR2_X1 U528 ( .A(KEYINPUT11), .B(n416), .ZN(n424) );
  NAND2_X1 U529 ( .A1(G214), .A2(n466), .ZN(n417) );
  XNOR2_X1 U530 ( .A(n418), .B(n417), .ZN(n420) );
  XNOR2_X1 U531 ( .A(n419), .B(G122), .ZN(n431) );
  XNOR2_X1 U532 ( .A(n420), .B(n431), .ZN(n422) );
  XOR2_X1 U533 ( .A(n471), .B(G143), .Z(n421) );
  INV_X1 U534 ( .A(KEYINPUT13), .ZN(n426) );
  INV_X1 U535 ( .A(n561), .ZN(n429) );
  NOR2_X1 U536 ( .A1(n585), .A2(n429), .ZN(n430) );
  XNOR2_X1 U537 ( .A(n430), .B(KEYINPUT104), .ZN(n456) );
  XNOR2_X1 U538 ( .A(n432), .B(n431), .ZN(n435) );
  XNOR2_X1 U539 ( .A(n467), .B(n401), .ZN(n434) );
  NAND2_X1 U540 ( .A1(G224), .A2(n736), .ZN(n436) );
  XNOR2_X1 U541 ( .A(n470), .B(n436), .ZN(n437) );
  XNOR2_X1 U542 ( .A(n438), .B(n437), .ZN(n444) );
  XOR2_X1 U543 ( .A(KEYINPUT18), .B(KEYINPUT91), .Z(n440) );
  XNOR2_X1 U544 ( .A(KEYINPUT74), .B(KEYINPUT17), .ZN(n439) );
  XNOR2_X1 U545 ( .A(n440), .B(n439), .ZN(n442) );
  XNOR2_X1 U546 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U547 ( .A(n444), .B(n443), .ZN(n445) );
  OR2_X1 U548 ( .A1(G237), .A2(G902), .ZN(n447) );
  NAND2_X1 U549 ( .A1(n447), .A2(G210), .ZN(n446) );
  NAND2_X1 U550 ( .A1(n447), .A2(G214), .ZN(n448) );
  XOR2_X1 U551 ( .A(KEYINPUT92), .B(n448), .Z(n626) );
  NOR2_X2 U552 ( .A1(n632), .A2(n626), .ZN(n610) );
  INV_X1 U553 ( .A(KEYINPUT19), .ZN(n449) );
  XNOR2_X1 U554 ( .A(n610), .B(n449), .ZN(n590) );
  XOR2_X1 U555 ( .A(n450), .B(KEYINPUT14), .Z(n579) );
  NOR2_X1 U556 ( .A1(G898), .A2(n736), .ZN(n729) );
  NAND2_X1 U557 ( .A1(n729), .A2(G902), .ZN(n451) );
  NAND2_X1 U558 ( .A1(G952), .A2(n736), .ZN(n577) );
  AND2_X1 U559 ( .A1(n451), .A2(n577), .ZN(n452) );
  NOR2_X1 U560 ( .A1(n579), .A2(n452), .ZN(n453) );
  XNOR2_X1 U561 ( .A(KEYINPUT88), .B(KEYINPUT0), .ZN(n454) );
  NAND2_X1 U562 ( .A1(n456), .A2(n534), .ZN(n459) );
  XNOR2_X1 U563 ( .A(n461), .B(n460), .ZN(n465) );
  NAND2_X1 U564 ( .A1(n663), .A2(n474), .ZN(n476) );
  INV_X1 U565 ( .A(G472), .ZN(n475) );
  XNOR2_X2 U566 ( .A(n476), .B(n475), .ZN(n508) );
  INV_X1 U567 ( .A(KEYINPUT103), .ZN(n477) );
  XNOR2_X1 U568 ( .A(n477), .B(KEYINPUT6), .ZN(n478) );
  NOR2_X2 U569 ( .A1(n507), .A2(n609), .ZN(n528) );
  XNOR2_X1 U570 ( .A(n479), .B(n495), .ZN(n733) );
  XNOR2_X1 U571 ( .A(G128), .B(KEYINPUT94), .ZN(n480) );
  XNOR2_X1 U572 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U573 ( .A(n733), .B(n482), .ZN(n490) );
  XOR2_X1 U574 ( .A(KEYINPUT72), .B(KEYINPUT23), .Z(n484) );
  XNOR2_X1 U575 ( .A(G119), .B(G110), .ZN(n483) );
  XNOR2_X1 U576 ( .A(n484), .B(n483), .ZN(n485) );
  XOR2_X1 U577 ( .A(n485), .B(KEYINPUT95), .Z(n488) );
  AND2_X1 U578 ( .A1(n486), .A2(G221), .ZN(n487) );
  XNOR2_X1 U579 ( .A(n490), .B(n489), .ZN(n717) );
  NAND2_X1 U580 ( .A1(G217), .A2(n491), .ZN(n492) );
  XNOR2_X1 U581 ( .A(KEYINPUT96), .B(KEYINPUT25), .ZN(n493) );
  NAND2_X1 U582 ( .A1(n736), .A2(G227), .ZN(n494) );
  XNOR2_X1 U583 ( .A(n494), .B(KEYINPUT73), .ZN(n496) );
  XNOR2_X1 U584 ( .A(n496), .B(n495), .ZN(n501) );
  XNOR2_X1 U585 ( .A(n497), .B(G107), .ZN(n499) );
  XNOR2_X1 U586 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U587 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U588 ( .A(KEYINPUT65), .B(KEYINPUT1), .ZN(n504) );
  AND2_X1 U589 ( .A1(n583), .A2(n627), .ZN(n505) );
  XNOR2_X2 U590 ( .A(n506), .B(KEYINPUT32), .ZN(n746) );
  INV_X1 U591 ( .A(n507), .ZN(n512) );
  XNOR2_X1 U592 ( .A(n508), .B(KEYINPUT106), .ZN(n593) );
  AND2_X1 U593 ( .A1(n583), .A2(n509), .ZN(n510) );
  AND2_X1 U594 ( .A1(n593), .A2(n510), .ZN(n511) );
  NAND2_X1 U595 ( .A1(n512), .A2(n511), .ZN(n687) );
  XNOR2_X1 U596 ( .A(n534), .B(KEYINPUT93), .ZN(n538) );
  INV_X1 U597 ( .A(n609), .ZN(n514) );
  INV_X1 U598 ( .A(KEYINPUT76), .ZN(n515) );
  XNOR2_X1 U599 ( .A(n515), .B(KEYINPUT34), .ZN(n516) );
  NAND2_X1 U600 ( .A1(n529), .A2(n531), .ZN(n602) );
  XNOR2_X1 U601 ( .A(n602), .B(KEYINPUT75), .ZN(n518) );
  NAND2_X1 U602 ( .A1(n519), .A2(n518), .ZN(n521) );
  XNOR2_X1 U603 ( .A(KEYINPUT84), .B(KEYINPUT35), .ZN(n520) );
  NOR2_X1 U604 ( .A1(n676), .A2(KEYINPUT44), .ZN(n522) );
  NAND2_X1 U605 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U606 ( .A(n524), .B(KEYINPUT68), .ZN(n546) );
  NAND2_X1 U607 ( .A1(n526), .A2(KEYINPUT44), .ZN(n544) );
  NOR2_X1 U608 ( .A1(n583), .A2(n627), .ZN(n527) );
  AND2_X1 U609 ( .A1(n528), .A2(n527), .ZN(n677) );
  INV_X1 U610 ( .A(n529), .ZN(n530) );
  NAND2_X1 U611 ( .A1(n531), .A2(n530), .ZN(n532) );
  XOR2_X1 U612 ( .A(n532), .B(KEYINPUT102), .Z(n698) );
  NOR2_X1 U613 ( .A1(n693), .A2(n698), .ZN(n618) );
  NOR2_X1 U614 ( .A1(n533), .A2(n508), .ZN(n554) );
  NAND2_X1 U615 ( .A1(n534), .A2(n554), .ZN(n535) );
  XNOR2_X1 U616 ( .A(n535), .B(KEYINPUT31), .ZN(n697) );
  AND2_X1 U617 ( .A1(n508), .A2(n596), .ZN(n536) );
  NAND2_X1 U618 ( .A1(n597), .A2(n536), .ZN(n537) );
  NOR2_X1 U619 ( .A1(n538), .A2(n537), .ZN(n682) );
  NOR2_X1 U620 ( .A1(n697), .A2(n682), .ZN(n539) );
  NOR2_X1 U621 ( .A1(n618), .A2(n539), .ZN(n540) );
  NOR2_X1 U622 ( .A1(n677), .A2(n540), .ZN(n542) );
  INV_X1 U623 ( .A(KEYINPUT105), .ZN(n541) );
  XNOR2_X1 U624 ( .A(n542), .B(n541), .ZN(n543) );
  NAND2_X1 U625 ( .A1(n546), .A2(n545), .ZN(n547) );
  XOR2_X1 U626 ( .A(KEYINPUT38), .B(n632), .Z(n620) );
  NOR2_X1 U627 ( .A1(n620), .A2(n626), .ZN(n563) );
  NAND2_X1 U628 ( .A1(n561), .A2(n563), .ZN(n548) );
  XNOR2_X1 U629 ( .A(n548), .B(KEYINPUT41), .ZN(n623) );
  NAND2_X1 U630 ( .A1(n583), .A2(n585), .ZN(n549) );
  XNOR2_X1 U631 ( .A(n549), .B(KEYINPUT49), .ZN(n553) );
  NOR2_X1 U632 ( .A1(n597), .A2(n627), .ZN(n550) );
  XOR2_X1 U633 ( .A(KEYINPUT50), .B(n550), .Z(n551) );
  NAND2_X1 U634 ( .A1(n508), .A2(n551), .ZN(n552) );
  NOR2_X1 U635 ( .A1(n553), .A2(n552), .ZN(n555) );
  NOR2_X1 U636 ( .A1(n555), .A2(n554), .ZN(n557) );
  XOR2_X1 U637 ( .A(KEYINPUT51), .B(KEYINPUT119), .Z(n556) );
  XNOR2_X1 U638 ( .A(n557), .B(n556), .ZN(n558) );
  NAND2_X1 U639 ( .A1(n623), .A2(n558), .ZN(n568) );
  INV_X1 U640 ( .A(n559), .ZN(n573) );
  NAND2_X1 U641 ( .A1(n620), .A2(n626), .ZN(n560) );
  NAND2_X1 U642 ( .A1(n561), .A2(n560), .ZN(n565) );
  INV_X1 U643 ( .A(n618), .ZN(n562) );
  NAND2_X1 U644 ( .A1(n563), .A2(n562), .ZN(n564) );
  NAND2_X1 U645 ( .A1(n565), .A2(n564), .ZN(n566) );
  NAND2_X1 U646 ( .A1(n573), .A2(n566), .ZN(n567) );
  NAND2_X1 U647 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U648 ( .A(KEYINPUT52), .B(n569), .Z(n570) );
  NOR2_X1 U649 ( .A1(n579), .A2(n570), .ZN(n571) );
  NAND2_X1 U650 ( .A1(G952), .A2(n571), .ZN(n572) );
  XNOR2_X1 U651 ( .A(n572), .B(KEYINPUT120), .ZN(n575) );
  NAND2_X1 U652 ( .A1(n573), .A2(n623), .ZN(n574) );
  AND2_X1 U653 ( .A1(n575), .A2(n574), .ZN(n640) );
  INV_X1 U654 ( .A(KEYINPUT81), .ZN(n605) );
  NAND2_X1 U655 ( .A1(n605), .A2(n618), .ZN(n591) );
  NOR2_X1 U656 ( .A1(G900), .A2(n736), .ZN(n576) );
  NAND2_X1 U657 ( .A1(n576), .A2(G902), .ZN(n578) );
  NAND2_X1 U658 ( .A1(n578), .A2(n577), .ZN(n581) );
  INV_X1 U659 ( .A(n579), .ZN(n580) );
  NAND2_X1 U660 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U661 ( .A(KEYINPUT77), .B(n582), .ZN(n601) );
  NAND2_X1 U662 ( .A1(n601), .A2(n583), .ZN(n584) );
  INV_X1 U663 ( .A(n593), .ZN(n586) );
  NAND2_X1 U664 ( .A1(n608), .A2(n586), .ZN(n588) );
  XNOR2_X1 U665 ( .A(KEYINPUT28), .B(KEYINPUT109), .ZN(n587) );
  XNOR2_X1 U666 ( .A(n588), .B(n587), .ZN(n589) );
  AND2_X1 U667 ( .A1(n589), .A2(n596), .ZN(n622) );
  AND2_X1 U668 ( .A1(n590), .A2(n622), .ZN(n691) );
  NAND2_X1 U669 ( .A1(n591), .A2(n691), .ZN(n592) );
  NAND2_X1 U670 ( .A1(n592), .A2(KEYINPUT47), .ZN(n604) );
  NOR2_X1 U671 ( .A1(n593), .A2(n626), .ZN(n595) );
  NAND2_X1 U672 ( .A1(n597), .A2(n596), .ZN(n598) );
  NOR2_X1 U673 ( .A1(n632), .A2(n602), .ZN(n603) );
  NAND2_X1 U674 ( .A1(n361), .A2(n603), .ZN(n690) );
  NAND2_X1 U675 ( .A1(n604), .A2(n690), .ZN(n607) );
  NOR2_X1 U676 ( .A1(KEYINPUT47), .A2(n605), .ZN(n606) );
  NOR2_X1 U677 ( .A1(n607), .A2(n606), .ZN(n619) );
  NAND2_X1 U678 ( .A1(n629), .A2(n610), .ZN(n612) );
  INV_X1 U679 ( .A(KEYINPUT36), .ZN(n611) );
  XNOR2_X1 U680 ( .A(n612), .B(n611), .ZN(n613) );
  NAND2_X1 U681 ( .A1(n613), .A2(n627), .ZN(n615) );
  INV_X1 U682 ( .A(KEYINPUT110), .ZN(n614) );
  INV_X1 U683 ( .A(n691), .ZN(n616) );
  NOR2_X1 U684 ( .A1(KEYINPUT47), .A2(n616), .ZN(n617) );
  NAND2_X1 U685 ( .A1(n623), .A2(n622), .ZN(n624) );
  XNOR2_X1 U686 ( .A(n624), .B(KEYINPUT42), .ZN(n748) );
  INV_X1 U687 ( .A(n647), .ZN(n638) );
  NOR2_X1 U688 ( .A1(n627), .A2(n626), .ZN(n628) );
  NAND2_X1 U689 ( .A1(n629), .A2(n628), .ZN(n630) );
  XNOR2_X1 U690 ( .A(KEYINPUT43), .B(n630), .ZN(n631) );
  XNOR2_X1 U691 ( .A(n631), .B(KEYINPUT108), .ZN(n633) );
  NAND2_X1 U692 ( .A1(n633), .A2(n632), .ZN(n703) );
  NAND2_X1 U693 ( .A1(n698), .A2(n634), .ZN(n701) );
  NAND2_X1 U694 ( .A1(KEYINPUT2), .A2(n701), .ZN(n635) );
  XOR2_X1 U695 ( .A(KEYINPUT78), .B(n635), .Z(n636) );
  NAND2_X1 U696 ( .A1(n703), .A2(n636), .ZN(n637) );
  NOR2_X1 U697 ( .A1(n638), .A2(n637), .ZN(n645) );
  AND2_X1 U698 ( .A1(n640), .A2(n645), .ZN(n639) );
  NAND2_X1 U699 ( .A1(n721), .A2(n639), .ZN(n644) );
  INV_X1 U700 ( .A(n640), .ZN(n642) );
  XNOR2_X1 U701 ( .A(KEYINPUT80), .B(KEYINPUT2), .ZN(n641) );
  OR2_X1 U702 ( .A1(n642), .A2(n641), .ZN(n643) );
  AND2_X1 U703 ( .A1(n644), .A2(n643), .ZN(n650) );
  AND2_X1 U704 ( .A1(n703), .A2(n701), .ZN(n646) );
  XNOR2_X2 U705 ( .A(n648), .B(KEYINPUT83), .ZN(n735) );
  NOR2_X1 U706 ( .A1(n650), .A2(n655), .ZN(n651) );
  XNOR2_X1 U707 ( .A(n651), .B(KEYINPUT121), .ZN(n652) );
  NOR2_X1 U708 ( .A1(G953), .A2(n652), .ZN(n654) );
  XNOR2_X1 U709 ( .A(KEYINPUT122), .B(KEYINPUT53), .ZN(n653) );
  XNOR2_X1 U710 ( .A(n656), .B(KEYINPUT82), .ZN(n658) );
  INV_X1 U711 ( .A(KEYINPUT2), .ZN(n657) );
  NOR2_X1 U712 ( .A1(n658), .A2(n657), .ZN(n659) );
  NAND2_X1 U713 ( .A1(n660), .A2(n659), .ZN(n661) );
  NAND2_X1 U714 ( .A1(n716), .A2(G472), .ZN(n665) );
  XNOR2_X1 U715 ( .A(KEYINPUT111), .B(KEYINPUT62), .ZN(n662) );
  XNOR2_X1 U716 ( .A(n663), .B(n662), .ZN(n664) );
  XNOR2_X1 U717 ( .A(n665), .B(n664), .ZN(n667) );
  INV_X1 U718 ( .A(G952), .ZN(n666) );
  NOR2_X2 U719 ( .A1(n667), .A2(n720), .ZN(n669) );
  XNOR2_X1 U720 ( .A(KEYINPUT89), .B(KEYINPUT63), .ZN(n668) );
  XNOR2_X1 U721 ( .A(n669), .B(n668), .ZN(G57) );
  NAND2_X1 U722 ( .A1(n716), .A2(G210), .ZN(n673) );
  XOR2_X1 U723 ( .A(KEYINPUT79), .B(KEYINPUT54), .Z(n670) );
  XNOR2_X1 U724 ( .A(n670), .B(KEYINPUT55), .ZN(n671) );
  XOR2_X1 U725 ( .A(KEYINPUT85), .B(KEYINPUT56), .Z(n674) );
  XNOR2_X1 U726 ( .A(n675), .B(n674), .ZN(G51) );
  XOR2_X1 U727 ( .A(G122), .B(n676), .Z(G24) );
  XOR2_X1 U728 ( .A(G101), .B(n677), .Z(n678) );
  XNOR2_X1 U729 ( .A(KEYINPUT112), .B(n678), .ZN(G3) );
  NAND2_X1 U730 ( .A1(n682), .A2(n693), .ZN(n679) );
  XNOR2_X1 U731 ( .A(n679), .B(G104), .ZN(G6) );
  XOR2_X1 U732 ( .A(KEYINPUT115), .B(KEYINPUT27), .Z(n681) );
  XNOR2_X1 U733 ( .A(KEYINPUT113), .B(KEYINPUT114), .ZN(n680) );
  XNOR2_X1 U734 ( .A(n681), .B(n680), .ZN(n686) );
  XNOR2_X1 U735 ( .A(G107), .B(KEYINPUT26), .ZN(n684) );
  NAND2_X1 U736 ( .A1(n682), .A2(n698), .ZN(n683) );
  XNOR2_X1 U737 ( .A(n684), .B(n683), .ZN(n685) );
  XNOR2_X1 U738 ( .A(n686), .B(n685), .ZN(G9) );
  XNOR2_X1 U739 ( .A(G110), .B(n687), .ZN(G12) );
  XOR2_X1 U740 ( .A(G128), .B(KEYINPUT29), .Z(n689) );
  NAND2_X1 U741 ( .A1(n691), .A2(n698), .ZN(n688) );
  XNOR2_X1 U742 ( .A(n689), .B(n688), .ZN(G30) );
  XNOR2_X1 U743 ( .A(G143), .B(n690), .ZN(G45) );
  NAND2_X1 U744 ( .A1(n691), .A2(n693), .ZN(n692) );
  XNOR2_X1 U745 ( .A(n692), .B(G146), .ZN(G48) );
  XOR2_X1 U746 ( .A(KEYINPUT116), .B(KEYINPUT117), .Z(n695) );
  NAND2_X1 U747 ( .A1(n697), .A2(n693), .ZN(n694) );
  XNOR2_X1 U748 ( .A(n695), .B(n694), .ZN(n696) );
  XNOR2_X1 U749 ( .A(G113), .B(n696), .ZN(G15) );
  NAND2_X1 U750 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U751 ( .A(n699), .B(KEYINPUT118), .ZN(n700) );
  XNOR2_X1 U752 ( .A(G116), .B(n700), .ZN(G18) );
  INV_X1 U753 ( .A(n701), .ZN(n702) );
  XOR2_X1 U754 ( .A(G134), .B(n702), .Z(G36) );
  XNOR2_X1 U755 ( .A(G140), .B(n703), .ZN(G42) );
  NAND2_X1 U756 ( .A1(n716), .A2(G469), .ZN(n708) );
  XOR2_X1 U757 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n704) );
  XOR2_X1 U758 ( .A(n704), .B(KEYINPUT123), .Z(n705) );
  XNOR2_X1 U759 ( .A(n706), .B(n705), .ZN(n707) );
  XNOR2_X1 U760 ( .A(n708), .B(n707), .ZN(n709) );
  NOR2_X1 U761 ( .A1(n720), .A2(n709), .ZN(G54) );
  NAND2_X1 U762 ( .A1(n716), .A2(G475), .ZN(n711) );
  XNOR2_X1 U763 ( .A(n712), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U764 ( .A1(n716), .A2(G478), .ZN(n713) );
  XOR2_X1 U765 ( .A(n714), .B(n713), .Z(n715) );
  NOR2_X1 U766 ( .A1(n720), .A2(n715), .ZN(G63) );
  NAND2_X1 U767 ( .A1(n716), .A2(G217), .ZN(n718) );
  XNOR2_X1 U768 ( .A(n718), .B(n717), .ZN(n719) );
  NOR2_X1 U769 ( .A1(n720), .A2(n719), .ZN(G66) );
  INV_X1 U770 ( .A(n721), .ZN(n722) );
  NOR2_X1 U771 ( .A1(n722), .A2(G953), .ZN(n728) );
  NAND2_X1 U772 ( .A1(G224), .A2(G953), .ZN(n723) );
  XNOR2_X1 U773 ( .A(n723), .B(KEYINPUT124), .ZN(n724) );
  XNOR2_X1 U774 ( .A(KEYINPUT61), .B(n724), .ZN(n725) );
  NAND2_X1 U775 ( .A1(n725), .A2(G898), .ZN(n726) );
  XNOR2_X1 U776 ( .A(n726), .B(KEYINPUT125), .ZN(n727) );
  NOR2_X1 U777 ( .A1(n728), .A2(n727), .ZN(n732) );
  NOR2_X1 U778 ( .A1(n730), .A2(n729), .ZN(n731) );
  XOR2_X1 U779 ( .A(n732), .B(n731), .Z(G69) );
  XOR2_X1 U780 ( .A(n734), .B(n733), .Z(n738) );
  XNOR2_X1 U781 ( .A(n735), .B(n738), .ZN(n737) );
  NAND2_X1 U782 ( .A1(n737), .A2(n736), .ZN(n743) );
  XOR2_X1 U783 ( .A(n738), .B(G227), .Z(n739) );
  XNOR2_X1 U784 ( .A(n739), .B(KEYINPUT126), .ZN(n740) );
  NAND2_X1 U785 ( .A1(n740), .A2(G900), .ZN(n741) );
  NAND2_X1 U786 ( .A1(G953), .A2(n741), .ZN(n742) );
  NAND2_X1 U787 ( .A1(n743), .A2(n742), .ZN(G72) );
  XNOR2_X1 U788 ( .A(G125), .B(KEYINPUT37), .ZN(n745) );
  XNOR2_X1 U789 ( .A(n745), .B(n744), .ZN(G27) );
  XNOR2_X1 U790 ( .A(n746), .B(G119), .ZN(G21) );
  XNOR2_X1 U791 ( .A(G131), .B(n747), .ZN(G33) );
  XOR2_X1 U792 ( .A(G137), .B(n748), .Z(n749) );
  XNOR2_X1 U793 ( .A(KEYINPUT127), .B(n749), .ZN(G39) );
endmodule

