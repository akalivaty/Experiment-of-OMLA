//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 1 0 1 0 1 0 0 0 0 1 1 1 0 0 1 1 0 0 1 0 1 1 1 1 0 0 1 0 0 1 1 1 1 0 0 1 0 1 0 0 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n715, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n736, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n759, new_n760, new_n761, new_n763, new_n764,
    new_n765, new_n766, new_n768, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n863,
    new_n864, new_n866, new_n867, new_n868, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n922, new_n923, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n938, new_n939, new_n940, new_n942,
    new_n943, new_n944, new_n945, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n967, new_n968, new_n969, new_n970, new_n972, new_n973, new_n974,
    new_n975, new_n976;
  XNOR2_X1  g000(.A(KEYINPUT84), .B(KEYINPUT31), .ZN(new_n202));
  NAND2_X1  g001(.A1(G228gat), .A2(G233gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(G211gat), .B(G218gat), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT22), .ZN(new_n205));
  INV_X1    g004(.A(G211gat), .ZN(new_n206));
  INV_X1    g005(.A(G218gat), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n205), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(G197gat), .B(G204gat), .ZN(new_n209));
  AOI21_X1  g008(.A(new_n204), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n204), .A2(new_n209), .A3(new_n208), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(G155gat), .B(G162gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT2), .ZN(new_n215));
  INV_X1    g014(.A(G141gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(G148gat), .ZN(new_n217));
  INV_X1    g016(.A(G148gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(G141gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n214), .B1(new_n215), .B2(new_n220), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n217), .A2(new_n219), .A3(KEYINPUT79), .ZN(new_n222));
  INV_X1    g021(.A(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT79), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n224), .A2(new_n216), .A3(G148gat), .ZN(new_n225));
  NOR3_X1   g024(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n226));
  AND2_X1   g025(.A1(G155gat), .A2(G162gat), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n225), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  OAI21_X1  g027(.A(KEYINPUT80), .B1(new_n223), .B2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(new_n227), .ZN(new_n230));
  INV_X1    g029(.A(G155gat), .ZN(new_n231));
  INV_X1    g030(.A(G162gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n230), .B1(KEYINPUT2), .B2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT80), .ZN(new_n235));
  NAND4_X1  g034(.A1(new_n234), .A2(new_n235), .A3(new_n222), .A4(new_n225), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n221), .B1(new_n229), .B2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT29), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n213), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(new_n213), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n238), .B1(new_n243), .B2(KEYINPUT29), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n229), .A2(new_n236), .ZN(new_n245));
  INV_X1    g044(.A(new_n221), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(KEYINPUT81), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT81), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n237), .A2(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n244), .A2(new_n248), .A3(new_n250), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n203), .B1(new_n242), .B2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT85), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n211), .A2(new_n253), .A3(new_n212), .ZN(new_n254));
  AOI21_X1  g053(.A(KEYINPUT29), .B1(new_n210), .B2(KEYINPUT85), .ZN(new_n255));
  AOI21_X1  g054(.A(KEYINPUT3), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n203), .B1(new_n256), .B2(new_n237), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n257), .A2(new_n241), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n202), .B1(new_n252), .B2(new_n258), .ZN(new_n259));
  OR2_X1    g058(.A1(new_n257), .A2(new_n241), .ZN(new_n260));
  INV_X1    g059(.A(new_n202), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n237), .A2(new_n249), .ZN(new_n262));
  AOI211_X1 g061(.A(KEYINPUT81), .B(new_n221), .C1(new_n229), .C2(new_n236), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n241), .B1(new_n264), .B2(new_n244), .ZN(new_n265));
  OAI211_X1 g064(.A(new_n260), .B(new_n261), .C1(new_n265), .C2(new_n203), .ZN(new_n266));
  XNOR2_X1  g065(.A(G78gat), .B(G106gat), .ZN(new_n267));
  INV_X1    g066(.A(G50gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n267), .B(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n269), .B(G22gat), .ZN(new_n270));
  AND3_X1   g069(.A1(new_n259), .A2(new_n266), .A3(new_n270), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n270), .B1(new_n259), .B2(new_n266), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(G227gat), .A2(G233gat), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT25), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT23), .ZN(new_n277));
  AOI22_X1  g076(.A1(new_n277), .A2(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT65), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(KEYINPUT23), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(G169gat), .ZN(new_n282));
  INV_X1    g081(.A(G176gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n281), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT24), .ZN(new_n286));
  INV_X1    g085(.A(G183gat), .ZN(new_n287));
  INV_X1    g086(.A(G190gat), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n286), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NAND3_X1  g088(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n290));
  OAI211_X1 g089(.A(new_n289), .B(new_n290), .C1(G183gat), .C2(G190gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n285), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n282), .A2(new_n283), .A3(KEYINPUT23), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n293), .B(KEYINPUT64), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n276), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n293), .A2(KEYINPUT25), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n296), .B1(new_n281), .B2(new_n284), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n287), .A2(KEYINPUT67), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT67), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(G183gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n288), .A2(KEYINPUT68), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT68), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(G190gat), .ZN(new_n303));
  NAND4_X1  g102(.A1(new_n298), .A2(new_n300), .A3(new_n301), .A4(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n290), .A2(KEYINPUT66), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT66), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n306), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n304), .A2(new_n308), .A3(new_n289), .ZN(new_n309));
  AND3_X1   g108(.A1(new_n297), .A2(new_n309), .A3(KEYINPUT69), .ZN(new_n310));
  AOI21_X1  g109(.A(KEYINPUT69), .B1(new_n297), .B2(new_n309), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n295), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  XOR2_X1   g111(.A(G113gat), .B(G120gat), .Z(new_n313));
  INV_X1    g112(.A(KEYINPUT1), .ZN(new_n314));
  XNOR2_X1  g113(.A(G127gat), .B(G134gat), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT73), .ZN(new_n316));
  OAI211_X1 g115(.A(new_n313), .B(new_n314), .C1(new_n315), .C2(new_n316), .ZN(new_n317));
  XOR2_X1   g116(.A(G127gat), .B(G134gat), .Z(new_n318));
  NAND2_X1  g117(.A1(new_n316), .A2(new_n314), .ZN(new_n319));
  XNOR2_X1  g118(.A(G113gat), .B(G120gat), .ZN(new_n320));
  OAI211_X1 g119(.A(new_n318), .B(new_n319), .C1(new_n320), .C2(KEYINPUT1), .ZN(new_n321));
  AND2_X1   g120(.A1(new_n317), .A2(new_n321), .ZN(new_n322));
  OR3_X1    g121(.A1(new_n284), .A2(KEYINPUT72), .A3(KEYINPUT26), .ZN(new_n323));
  OAI21_X1  g122(.A(KEYINPUT72), .B1(new_n284), .B2(KEYINPUT26), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n282), .A2(new_n283), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n326), .B1(KEYINPUT26), .B2(new_n284), .ZN(new_n327));
  AOI22_X1  g126(.A1(new_n325), .A2(new_n327), .B1(G183gat), .B2(G190gat), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT28), .ZN(new_n329));
  XNOR2_X1  g128(.A(KEYINPUT68), .B(G190gat), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT27), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n331), .B1(new_n298), .B2(new_n300), .ZN(new_n332));
  NOR2_X1   g131(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n330), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n301), .A2(new_n303), .A3(KEYINPUT28), .ZN(new_n335));
  AND2_X1   g134(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n336), .A2(new_n333), .ZN(new_n337));
  OAI21_X1  g136(.A(KEYINPUT70), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(KEYINPUT27), .B(G183gat), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT70), .ZN(new_n340));
  NAND4_X1  g139(.A1(new_n330), .A2(new_n339), .A3(new_n340), .A4(KEYINPUT28), .ZN(new_n341));
  AOI22_X1  g140(.A1(new_n329), .A2(new_n334), .B1(new_n338), .B2(new_n341), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n328), .B1(new_n342), .B2(KEYINPUT71), .ZN(new_n343));
  AND2_X1   g142(.A1(new_n338), .A2(new_n341), .ZN(new_n344));
  INV_X1    g143(.A(new_n333), .ZN(new_n345));
  XNOR2_X1  g144(.A(KEYINPUT67), .B(G183gat), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n345), .B1(new_n346), .B2(new_n331), .ZN(new_n347));
  AOI21_X1  g146(.A(KEYINPUT28), .B1(new_n347), .B2(new_n330), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT71), .ZN(new_n349));
  NOR3_X1   g148(.A1(new_n344), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  OAI211_X1 g149(.A(new_n312), .B(new_n322), .C1(new_n343), .C2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n349), .B1(new_n344), .B2(new_n348), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n342), .A2(KEYINPUT71), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n353), .A2(new_n354), .A3(new_n328), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n322), .B1(new_n355), .B2(new_n312), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n275), .B1(new_n352), .B2(new_n356), .ZN(new_n357));
  XNOR2_X1  g156(.A(G15gat), .B(G43gat), .ZN(new_n358));
  XNOR2_X1  g157(.A(G71gat), .B(G99gat), .ZN(new_n359));
  XNOR2_X1  g158(.A(new_n358), .B(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT33), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n357), .A2(KEYINPUT32), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(KEYINPUT74), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT32), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n312), .B1(new_n343), .B2(new_n350), .ZN(new_n367));
  INV_X1    g166(.A(new_n322), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(new_n351), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n366), .B1(new_n370), .B2(new_n275), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT74), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n371), .A2(new_n372), .A3(new_n363), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n365), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n360), .B1(new_n357), .B2(KEYINPUT32), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n357), .A2(new_n361), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n374), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n369), .A2(new_n274), .A3(new_n351), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT34), .ZN(new_n380));
  XNOR2_X1  g179(.A(new_n379), .B(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n273), .B1(new_n378), .B2(new_n382), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n372), .B1(new_n371), .B2(new_n363), .ZN(new_n384));
  AND4_X1   g183(.A1(new_n372), .A2(new_n357), .A3(KEYINPUT32), .A4(new_n363), .ZN(new_n385));
  OAI211_X1 g184(.A(new_n381), .B(new_n377), .C1(new_n384), .C2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT75), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  AOI22_X1  g187(.A1(new_n365), .A2(new_n373), .B1(new_n376), .B2(new_n375), .ZN(new_n389));
  AOI21_X1  g188(.A(KEYINPUT75), .B1(new_n389), .B2(new_n381), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n383), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  AND3_X1   g190(.A1(new_n237), .A2(KEYINPUT4), .A3(new_n322), .ZN(new_n392));
  AOI21_X1  g191(.A(KEYINPUT4), .B1(new_n237), .B2(new_n322), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(G225gat), .A2(G233gat), .ZN(new_n395));
  XOR2_X1   g194(.A(new_n395), .B(KEYINPUT82), .Z(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  NOR3_X1   g196(.A1(new_n262), .A2(new_n263), .A3(new_n238), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n239), .A2(new_n368), .ZN(new_n399));
  OAI211_X1 g198(.A(new_n394), .B(new_n397), .C1(new_n398), .C2(new_n399), .ZN(new_n400));
  NOR3_X1   g199(.A1(new_n262), .A2(new_n263), .A3(new_n322), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n247), .A2(new_n368), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n396), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n400), .A2(KEYINPUT5), .A3(new_n403), .ZN(new_n404));
  XNOR2_X1  g203(.A(G1gat), .B(G29gat), .ZN(new_n405));
  XNOR2_X1  g204(.A(new_n405), .B(KEYINPUT0), .ZN(new_n406));
  XNOR2_X1  g205(.A(G57gat), .B(G85gat), .ZN(new_n407));
  XOR2_X1   g206(.A(new_n406), .B(new_n407), .Z(new_n408));
  NAND3_X1  g207(.A1(new_n248), .A2(KEYINPUT3), .A3(new_n250), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n409), .A2(new_n368), .A3(new_n239), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT5), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n410), .A2(new_n411), .A3(new_n397), .A4(new_n394), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n404), .A2(new_n408), .A3(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT6), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n408), .B1(new_n404), .B2(new_n412), .ZN(new_n416));
  OAI21_X1  g215(.A(KEYINPUT83), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n416), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT83), .ZN(new_n419));
  NAND4_X1  g218(.A1(new_n418), .A2(new_n419), .A3(new_n414), .A4(new_n413), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n416), .A2(KEYINPUT6), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n417), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(G226gat), .A2(G233gat), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n424), .B1(new_n367), .B2(new_n240), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n423), .B1(new_n355), .B2(new_n312), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n243), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n367), .A2(new_n424), .ZN(new_n428));
  AOI21_X1  g227(.A(KEYINPUT29), .B1(new_n355), .B2(new_n312), .ZN(new_n429));
  OAI211_X1 g228(.A(new_n428), .B(new_n213), .C1(new_n429), .C2(new_n424), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n427), .A2(new_n430), .ZN(new_n431));
  XNOR2_X1  g230(.A(G8gat), .B(G36gat), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n432), .B(KEYINPUT76), .ZN(new_n433));
  XOR2_X1   g232(.A(G64gat), .B(G92gat), .Z(new_n434));
  XNOR2_X1  g233(.A(new_n433), .B(new_n434), .ZN(new_n435));
  XNOR2_X1  g234(.A(new_n435), .B(KEYINPUT77), .ZN(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n431), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT30), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n427), .A2(new_n430), .A3(new_n435), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n438), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT78), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n442), .B1(new_n440), .B2(new_n439), .ZN(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n440), .A2(new_n442), .A3(new_n439), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n441), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n422), .A2(new_n446), .ZN(new_n447));
  OAI21_X1  g246(.A(KEYINPUT35), .B1(new_n391), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(KEYINPUT90), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT90), .ZN(new_n450));
  OAI211_X1 g249(.A(new_n450), .B(KEYINPUT35), .C1(new_n391), .C2(new_n447), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n404), .A2(new_n412), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT87), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n404), .A2(KEYINPUT87), .A3(new_n412), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n408), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n421), .B1(new_n456), .B2(new_n415), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT35), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  AND3_X1   g258(.A1(new_n427), .A2(new_n430), .A3(new_n435), .ZN(new_n460));
  AOI22_X1  g259(.A1(new_n460), .A2(KEYINPUT30), .B1(new_n431), .B2(new_n437), .ZN(new_n461));
  INV_X1    g260(.A(new_n445), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n461), .B1(new_n462), .B2(new_n443), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT86), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  OAI211_X1 g264(.A(new_n461), .B(KEYINPUT86), .C1(new_n462), .C2(new_n443), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n459), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(new_n391), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n449), .A2(new_n451), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n386), .A2(new_n387), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n389), .A2(KEYINPUT75), .A3(new_n381), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT36), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n378), .A2(new_n382), .ZN(new_n475));
  AND3_X1   g274(.A1(new_n473), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n474), .B1(new_n473), .B2(new_n475), .ZN(new_n477));
  INV_X1    g276(.A(new_n273), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n478), .B1(new_n422), .B2(new_n446), .ZN(new_n479));
  NOR3_X1   g278(.A1(new_n476), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT40), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n397), .B1(new_n410), .B2(new_n394), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT39), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(new_n408), .ZN(new_n485));
  OR3_X1    g284(.A1(new_n401), .A2(new_n396), .A3(new_n402), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(KEYINPUT39), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n487), .A2(new_n482), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n481), .B1(new_n485), .B2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(new_n408), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n490), .B1(new_n482), .B2(new_n483), .ZN(new_n491));
  OAI211_X1 g290(.A(new_n491), .B(KEYINPUT40), .C1(new_n482), .C2(new_n487), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n493), .A2(new_n456), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n465), .A2(new_n466), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(KEYINPUT88), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT88), .ZN(new_n497));
  NAND4_X1  g296(.A1(new_n465), .A2(new_n494), .A3(new_n497), .A4(new_n466), .ZN(new_n498));
  XOR2_X1   g297(.A(KEYINPUT89), .B(KEYINPUT37), .Z(new_n499));
  OR2_X1    g298(.A1(new_n431), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n431), .A2(KEYINPUT37), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n436), .A2(KEYINPUT38), .ZN(new_n502));
  AND3_X1   g301(.A1(new_n500), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT38), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n435), .B1(new_n431), .B2(KEYINPUT37), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n504), .B1(new_n500), .B2(new_n505), .ZN(new_n506));
  NOR3_X1   g305(.A1(new_n503), .A2(new_n506), .A3(new_n460), .ZN(new_n507));
  INV_X1    g306(.A(new_n457), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n273), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n496), .A2(new_n498), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n480), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n470), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(G71gat), .A2(G78gat), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT9), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(G57gat), .ZN(new_n516));
  AND2_X1   g315(.A1(new_n516), .A2(G64gat), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n516), .A2(G64gat), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n515), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(G71gat), .B(G78gat), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n520), .A2(KEYINPUT99), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT99), .ZN(new_n522));
  OR2_X1    g321(.A1(G71gat), .A2(G78gat), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n522), .B1(new_n523), .B2(new_n513), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n519), .B1(new_n521), .B2(new_n524), .ZN(new_n525));
  OR2_X1    g324(.A1(KEYINPUT100), .A2(G57gat), .ZN(new_n526));
  NAND2_X1  g325(.A1(KEYINPUT100), .A2(G57gat), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n526), .A2(KEYINPUT101), .A3(G64gat), .A4(new_n527), .ZN(new_n528));
  AND3_X1   g327(.A1(new_n526), .A2(G64gat), .A3(new_n527), .ZN(new_n529));
  OR2_X1    g328(.A1(new_n518), .A2(KEYINPUT101), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT102), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n520), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n523), .A2(KEYINPUT102), .A3(new_n513), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n533), .A2(new_n515), .A3(new_n534), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n525), .B1(new_n531), .B2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT21), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(G231gat), .A2(G233gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n538), .B(new_n539), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n540), .B(G127gat), .ZN(new_n541));
  XNOR2_X1  g340(.A(G15gat), .B(G22gat), .ZN(new_n542));
  INV_X1    g341(.A(G1gat), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(KEYINPUT16), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n542), .A2(G1gat), .ZN(new_n547));
  NOR3_X1   g346(.A1(new_n546), .A2(new_n547), .A3(G8gat), .ZN(new_n548));
  INV_X1    g347(.A(G8gat), .ZN(new_n549));
  OR2_X1    g348(.A1(new_n542), .A2(G1gat), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n549), .B1(new_n550), .B2(new_n545), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT103), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n536), .B(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n553), .B1(new_n555), .B2(KEYINPUT21), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n541), .B(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n558), .B(new_n231), .ZN(new_n559));
  XOR2_X1   g358(.A(G183gat), .B(G211gat), .Z(new_n560));
  XNOR2_X1  g359(.A(new_n559), .B(new_n560), .ZN(new_n561));
  XOR2_X1   g360(.A(new_n557), .B(new_n561), .Z(new_n562));
  AND2_X1   g361(.A1(G232gat), .A2(G233gat), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n563), .A2(KEYINPUT41), .ZN(new_n564));
  XNOR2_X1  g363(.A(G134gat), .B(G162gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n564), .B(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT106), .ZN(new_n568));
  NAND2_X1  g367(.A1(G99gat), .A2(G106gat), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n569), .A2(KEYINPUT8), .ZN(new_n570));
  NAND2_X1  g369(.A1(G85gat), .A2(G92gat), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT7), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  OR2_X1    g372(.A1(G85gat), .A2(G92gat), .ZN(new_n574));
  NAND3_X1  g373(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n575));
  AND4_X1   g374(.A1(new_n570), .A2(new_n573), .A3(new_n574), .A4(new_n575), .ZN(new_n576));
  AND2_X1   g375(.A1(G99gat), .A2(G106gat), .ZN(new_n577));
  NOR2_X1   g376(.A1(G99gat), .A2(G106gat), .ZN(new_n578));
  OAI21_X1  g377(.A(KEYINPUT104), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(G99gat), .ZN(new_n580));
  INV_X1    g379(.A(G106gat), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT104), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n582), .A2(new_n583), .A3(new_n569), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n579), .A2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT105), .ZN(new_n586));
  AND3_X1   g385(.A1(new_n576), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n586), .B1(new_n576), .B2(new_n585), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n568), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  AND2_X1   g388(.A1(new_n579), .A2(new_n584), .ZN(new_n590));
  NAND4_X1  g389(.A1(new_n570), .A2(new_n573), .A3(new_n574), .A4(new_n575), .ZN(new_n591));
  OAI21_X1  g390(.A(KEYINPUT105), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n576), .A2(new_n585), .A3(new_n586), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n592), .A2(KEYINPUT106), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n589), .A2(new_n594), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n576), .A2(new_n585), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(G43gat), .B(G50gat), .ZN(new_n599));
  OR3_X1    g398(.A1(new_n599), .A2(KEYINPUT94), .A3(KEYINPUT15), .ZN(new_n600));
  OAI21_X1  g399(.A(KEYINPUT15), .B1(new_n599), .B2(KEYINPUT94), .ZN(new_n601));
  NAND2_X1  g400(.A1(G29gat), .A2(G36gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(KEYINPUT92), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT14), .ZN(new_n604));
  INV_X1    g403(.A(G29gat), .ZN(new_n605));
  INV_X1    g404(.A(G36gat), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  OAI21_X1  g406(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND4_X1  g408(.A1(new_n600), .A2(new_n601), .A3(new_n603), .A4(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n599), .A2(KEYINPUT15), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT91), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n607), .A2(new_n612), .ZN(new_n613));
  NAND4_X1  g412(.A1(new_n604), .A2(new_n605), .A3(new_n606), .A4(KEYINPUT91), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n613), .A2(new_n608), .A3(new_n614), .ZN(new_n615));
  AOI211_X1 g414(.A(KEYINPUT93), .B(new_n611), .C1(new_n615), .C2(new_n603), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT93), .ZN(new_n617));
  NOR3_X1   g416(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n608), .B1(new_n618), .B2(KEYINPUT91), .ZN(new_n619));
  INV_X1    g418(.A(new_n614), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n603), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n611), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n617), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  OAI211_X1 g422(.A(KEYINPUT17), .B(new_n610), .C1(new_n616), .C2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n610), .ZN(new_n625));
  INV_X1    g424(.A(new_n623), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n621), .A2(new_n617), .A3(new_n622), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n625), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  XOR2_X1   g427(.A(KEYINPUT95), .B(KEYINPUT17), .Z(new_n629));
  OAI211_X1 g428(.A(new_n598), .B(new_n624), .C1(new_n628), .C2(new_n629), .ZN(new_n630));
  XOR2_X1   g429(.A(G190gat), .B(G218gat), .Z(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n596), .B1(new_n589), .B2(new_n594), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n610), .B1(new_n616), .B2(new_n623), .ZN(new_n634));
  AOI22_X1  g433(.A1(new_n633), .A2(new_n634), .B1(KEYINPUT41), .B2(new_n563), .ZN(new_n635));
  AND3_X1   g434(.A1(new_n630), .A2(new_n632), .A3(new_n635), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n632), .B1(new_n630), .B2(new_n635), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n567), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n630), .A2(new_n635), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n639), .A2(new_n631), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n630), .A2(new_n632), .A3(new_n635), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n640), .A2(new_n566), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n638), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(G230gat), .A2(G233gat), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n598), .A2(new_n536), .ZN(new_n646));
  INV_X1    g445(.A(new_n536), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n592), .A2(new_n593), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n647), .A2(new_n597), .A3(new_n648), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n645), .B1(new_n646), .B2(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(G120gat), .B(G148gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(G176gat), .B(G204gat), .ZN(new_n652));
  XOR2_X1   g451(.A(new_n651), .B(new_n652), .Z(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n650), .A2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT10), .ZN(new_n656));
  OAI211_X1 g455(.A(new_n656), .B(new_n649), .C1(new_n633), .C2(new_n647), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n555), .A2(KEYINPUT10), .A3(new_n633), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(new_n645), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n655), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n645), .B(KEYINPUT107), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n662), .B1(new_n657), .B2(new_n658), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n654), .B1(new_n663), .B2(new_n650), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  NOR3_X1   g464(.A1(new_n562), .A2(new_n644), .A3(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n634), .A2(new_n553), .ZN(new_n667));
  OAI211_X1 g466(.A(new_n552), .B(new_n610), .C1(new_n623), .C2(new_n616), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n667), .A2(KEYINPUT96), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(G229gat), .A2(G233gat), .ZN(new_n670));
  XOR2_X1   g469(.A(new_n670), .B(KEYINPUT13), .Z(new_n671));
  INV_X1    g470(.A(KEYINPUT96), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n634), .A2(new_n553), .A3(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n669), .A2(new_n671), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n674), .A2(KEYINPUT97), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT97), .ZN(new_n676));
  NAND4_X1  g475(.A1(new_n669), .A2(new_n676), .A3(new_n671), .A4(new_n673), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g477(.A(G113gat), .B(G141gat), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(G197gat), .ZN(new_n680));
  XNOR2_X1  g479(.A(KEYINPUT11), .B(G169gat), .ZN(new_n681));
  XOR2_X1   g480(.A(new_n680), .B(new_n681), .Z(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(KEYINPUT12), .ZN(new_n683));
  OAI211_X1 g482(.A(new_n624), .B(new_n552), .C1(new_n628), .C2(new_n629), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n684), .A2(new_n670), .A3(new_n667), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT18), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND4_X1  g486(.A1(new_n684), .A2(KEYINPUT18), .A3(new_n670), .A4(new_n667), .ZN(new_n688));
  NAND4_X1  g487(.A1(new_n678), .A2(new_n683), .A3(new_n687), .A4(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT98), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  AND2_X1   g490(.A1(new_n687), .A2(new_n688), .ZN(new_n692));
  NAND4_X1  g491(.A1(new_n692), .A2(new_n678), .A3(KEYINPUT98), .A4(new_n683), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n692), .A2(new_n678), .ZN(new_n695));
  INV_X1    g494(.A(new_n683), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n694), .A2(new_n697), .ZN(new_n698));
  AND2_X1   g497(.A1(new_n666), .A2(new_n698), .ZN(new_n699));
  AND2_X1   g498(.A1(new_n512), .A2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n422), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(G1gat), .ZN(G1324gat));
  INV_X1    g502(.A(new_n700), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n465), .A2(new_n466), .ZN(new_n705));
  XNOR2_X1  g504(.A(KEYINPUT16), .B(G8gat), .ZN(new_n706));
  NOR3_X1   g505(.A1(new_n704), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(new_n705), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n549), .B1(new_n700), .B2(new_n708), .ZN(new_n709));
  OAI21_X1  g508(.A(KEYINPUT42), .B1(new_n707), .B2(new_n709), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n710), .B1(KEYINPUT42), .B2(new_n707), .ZN(G1325gat));
  NAND2_X1  g510(.A1(new_n473), .A2(new_n475), .ZN(new_n712));
  OR3_X1    g511(.A1(new_n704), .A2(G15gat), .A3(new_n712), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n476), .A2(new_n477), .ZN(new_n714));
  OAI21_X1  g513(.A(G15gat), .B1(new_n704), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n713), .A2(new_n715), .ZN(G1326gat));
  NAND2_X1  g515(.A1(new_n700), .A2(new_n273), .ZN(new_n717));
  XNOR2_X1  g516(.A(KEYINPUT43), .B(G22gat), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n717), .B(new_n718), .ZN(G1327gat));
  AOI21_X1  g518(.A(new_n643), .B1(new_n470), .B2(new_n511), .ZN(new_n720));
  INV_X1    g519(.A(new_n562), .ZN(new_n721));
  INV_X1    g520(.A(new_n698), .ZN(new_n722));
  NOR3_X1   g521(.A1(new_n721), .A2(new_n722), .A3(new_n665), .ZN(new_n723));
  AND2_X1   g522(.A1(new_n720), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n724), .A2(new_n605), .A3(new_n701), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(KEYINPUT45), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT44), .ZN(new_n727));
  AOI22_X1  g526(.A1(new_n448), .A2(KEYINPUT90), .B1(new_n467), .B2(new_n468), .ZN(new_n728));
  AOI22_X1  g527(.A1(new_n728), .A2(new_n451), .B1(new_n480), .B2(new_n510), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n727), .B1(new_n729), .B2(new_n643), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n512), .A2(KEYINPUT44), .A3(new_n644), .ZN(new_n731));
  AND2_X1   g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(new_n723), .ZN(new_n733));
  OAI21_X1  g532(.A(G29gat), .B1(new_n733), .B2(new_n422), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n726), .A2(new_n734), .ZN(G1328gat));
  NAND3_X1  g534(.A1(new_n724), .A2(new_n606), .A3(new_n708), .ZN(new_n736));
  XOR2_X1   g535(.A(new_n736), .B(KEYINPUT46), .Z(new_n737));
  OAI21_X1  g536(.A(G36gat), .B1(new_n733), .B2(new_n705), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(G1329gat));
  INV_X1    g538(.A(new_n714), .ZN(new_n740));
  NAND4_X1  g539(.A1(new_n730), .A2(new_n731), .A3(new_n740), .A4(new_n723), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(G43gat), .ZN(new_n742));
  INV_X1    g541(.A(G43gat), .ZN(new_n743));
  INV_X1    g542(.A(new_n712), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n724), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n742), .A2(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT47), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n746), .B(new_n747), .ZN(G1330gat));
  NOR2_X1   g547(.A1(new_n478), .A2(new_n268), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n730), .A2(new_n731), .A3(new_n723), .A4(new_n749), .ZN(new_n750));
  AND2_X1   g549(.A1(new_n724), .A2(new_n273), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n750), .B1(new_n751), .B2(G50gat), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(KEYINPUT48), .ZN(G1331gat));
  NAND3_X1  g552(.A1(new_n721), .A2(new_n643), .A3(new_n665), .ZN(new_n754));
  NOR3_X1   g553(.A1(new_n729), .A2(new_n698), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(new_n701), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n526), .A2(new_n527), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n756), .B(new_n757), .ZN(G1332gat));
  NAND2_X1  g557(.A1(new_n755), .A2(new_n708), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n759), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n760));
  XOR2_X1   g559(.A(KEYINPUT49), .B(G64gat), .Z(new_n761));
  OAI21_X1  g560(.A(new_n760), .B1(new_n759), .B2(new_n761), .ZN(G1333gat));
  NAND2_X1  g561(.A1(new_n755), .A2(new_n740), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n712), .A2(G71gat), .ZN(new_n764));
  AOI22_X1  g563(.A1(new_n763), .A2(G71gat), .B1(new_n755), .B2(new_n764), .ZN(new_n765));
  XNOR2_X1  g564(.A(KEYINPUT108), .B(KEYINPUT50), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n765), .B(new_n766), .ZN(G1334gat));
  NAND2_X1  g566(.A1(new_n755), .A2(new_n273), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g568(.A1(new_n721), .A2(new_n698), .ZN(new_n770));
  INV_X1    g569(.A(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(new_n665), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n732), .A2(new_n701), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(G85gat), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n512), .A2(new_n644), .A3(new_n770), .ZN(new_n776));
  OR2_X1    g575(.A1(new_n776), .A2(KEYINPUT51), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(KEYINPUT51), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  OR3_X1    g578(.A1(new_n422), .A2(G85gat), .A3(new_n772), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n775), .B1(new_n779), .B2(new_n780), .ZN(G1336gat));
  NAND4_X1  g580(.A1(new_n730), .A2(new_n731), .A3(new_n708), .A4(new_n773), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT109), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n782), .A2(new_n783), .A3(G92gat), .ZN(new_n784));
  NOR3_X1   g583(.A1(new_n705), .A2(G92gat), .A3(new_n772), .ZN(new_n785));
  NOR2_X1   g584(.A1(KEYINPUT110), .A2(KEYINPUT51), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n776), .A2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(new_n786), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n788), .B1(new_n720), .B2(new_n770), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n785), .B1(new_n787), .B2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n784), .A2(new_n790), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n783), .B1(new_n782), .B2(G92gat), .ZN(new_n792));
  OAI21_X1  g591(.A(KEYINPUT52), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n782), .A2(G92gat), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT52), .ZN(new_n795));
  INV_X1    g594(.A(new_n785), .ZN(new_n796));
  OAI211_X1 g595(.A(new_n794), .B(new_n795), .C1(new_n779), .C2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n793), .A2(new_n797), .ZN(G1337gat));
  NAND4_X1  g597(.A1(new_n730), .A2(new_n731), .A3(new_n740), .A4(new_n773), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT111), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n580), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n801), .B1(new_n800), .B2(new_n799), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n744), .A2(new_n580), .A3(new_n665), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n802), .B1(new_n779), .B2(new_n803), .ZN(G1338gat));
  NOR3_X1   g603(.A1(new_n478), .A2(G106gat), .A3(new_n772), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n777), .A2(new_n778), .A3(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT53), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n730), .A2(new_n731), .A3(new_n273), .A4(new_n773), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(G106gat), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n806), .A2(new_n807), .A3(new_n809), .ZN(new_n810));
  OR2_X1    g609(.A1(new_n787), .A2(new_n789), .ZN(new_n811));
  AOI22_X1  g610(.A1(new_n811), .A2(new_n805), .B1(G106gat), .B2(new_n808), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n810), .B1(new_n812), .B2(new_n807), .ZN(G1339gat));
  INV_X1    g612(.A(KEYINPUT114), .ZN(new_n814));
  XOR2_X1   g613(.A(KEYINPUT113), .B(KEYINPUT54), .Z(new_n815));
  AOI21_X1  g614(.A(new_n653), .B1(new_n663), .B2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT112), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n657), .A2(new_n658), .A3(new_n662), .ZN(new_n818));
  AND4_X1   g617(.A1(new_n817), .A2(new_n660), .A3(KEYINPUT54), .A4(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT54), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n820), .B1(new_n659), .B2(new_n645), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n817), .B1(new_n821), .B2(new_n818), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n816), .B1(new_n819), .B2(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT55), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  OAI211_X1 g624(.A(KEYINPUT55), .B(new_n816), .C1(new_n819), .C2(new_n822), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n825), .A2(new_n661), .A3(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(new_n682), .ZN(new_n828));
  AND2_X1   g627(.A1(new_n669), .A2(new_n673), .ZN(new_n829));
  OR2_X1    g628(.A1(new_n829), .A2(new_n671), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n684), .A2(new_n667), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n831), .A2(G229gat), .A3(G233gat), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n828), .B1(new_n830), .B2(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n694), .A2(new_n644), .A3(new_n834), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n814), .B1(new_n827), .B2(new_n835), .ZN(new_n836));
  AOI211_X1 g635(.A(new_n833), .B(new_n643), .C1(new_n691), .C2(new_n693), .ZN(new_n837));
  INV_X1    g636(.A(new_n661), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n838), .B1(new_n823), .B2(new_n824), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n837), .A2(KEYINPUT114), .A3(new_n826), .A4(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n836), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n698), .A2(new_n826), .A3(new_n839), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n694), .A2(new_n665), .A3(new_n834), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n644), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n562), .B1(new_n841), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n666), .A2(new_n722), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n391), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n708), .A2(new_n422), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(new_n698), .ZN(new_n850));
  XNOR2_X1  g649(.A(new_n850), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g650(.A1(new_n849), .A2(new_n665), .ZN(new_n852));
  INV_X1    g651(.A(G120gat), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(KEYINPUT115), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(KEYINPUT116), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n853), .A2(KEYINPUT115), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT116), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n852), .A2(new_n858), .A3(new_n854), .ZN(new_n859));
  AND3_X1   g658(.A1(new_n856), .A2(new_n857), .A3(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n857), .B1(new_n856), .B2(new_n859), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n860), .A2(new_n861), .ZN(G1341gat));
  NAND2_X1  g661(.A1(new_n849), .A2(new_n721), .ZN(new_n863));
  XNOR2_X1  g662(.A(KEYINPUT117), .B(G127gat), .ZN(new_n864));
  XNOR2_X1  g663(.A(new_n863), .B(new_n864), .ZN(G1342gat));
  AOI21_X1  g664(.A(new_n643), .B1(KEYINPUT56), .B2(G134gat), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n849), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g666(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n868));
  XOR2_X1   g667(.A(new_n867), .B(new_n868), .Z(G1343gat));
  NAND2_X1  g668(.A1(new_n714), .A2(new_n848), .ZN(new_n870));
  INV_X1    g669(.A(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT57), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n478), .A2(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(new_n846), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n875), .B1(new_n845), .B2(KEYINPUT118), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT118), .ZN(new_n877));
  OAI211_X1 g676(.A(new_n877), .B(new_n562), .C1(new_n841), .C2(new_n844), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n874), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n845), .A2(new_n846), .ZN(new_n880));
  AOI21_X1  g679(.A(KEYINPUT57), .B1(new_n880), .B2(new_n273), .ZN(new_n881));
  OAI211_X1 g680(.A(new_n698), .B(new_n871), .C1(new_n879), .C2(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(G141gat), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(KEYINPUT120), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n880), .A2(new_n701), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(KEYINPUT119), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT119), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n880), .A2(new_n887), .A3(new_n701), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n714), .A2(new_n273), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n889), .A2(new_n708), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n722), .A2(G141gat), .ZN(new_n891));
  NAND4_X1  g690(.A1(new_n886), .A2(new_n888), .A3(new_n890), .A4(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n883), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n884), .A2(new_n893), .A3(KEYINPUT58), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT58), .ZN(new_n895));
  OAI211_X1 g694(.A(new_n883), .B(new_n892), .C1(KEYINPUT120), .C2(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n894), .A2(new_n896), .ZN(G1344gat));
  NOR2_X1   g696(.A1(new_n772), .A2(G148gat), .ZN(new_n898));
  NAND4_X1  g697(.A1(new_n886), .A2(new_n888), .A3(new_n890), .A4(new_n898), .ZN(new_n899));
  XOR2_X1   g698(.A(new_n899), .B(KEYINPUT121), .Z(new_n900));
  XOR2_X1   g699(.A(KEYINPUT122), .B(KEYINPUT59), .Z(new_n901));
  NOR2_X1   g700(.A1(new_n827), .A2(new_n835), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n562), .B1(new_n844), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(new_n846), .ZN(new_n904));
  AOI21_X1  g703(.A(KEYINPUT57), .B1(new_n904), .B2(new_n273), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n874), .B1(new_n845), .B2(new_n846), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n907), .A2(new_n772), .A3(new_n870), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n901), .B1(new_n908), .B2(new_n218), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n218), .A2(KEYINPUT59), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n871), .B1(new_n879), .B2(new_n881), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n910), .B1(new_n911), .B2(new_n772), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n909), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n900), .A2(new_n913), .ZN(G1345gat));
  AND4_X1   g713(.A1(new_n721), .A2(new_n886), .A3(new_n888), .A4(new_n890), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT123), .ZN(new_n916));
  OR2_X1    g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g716(.A(G155gat), .B1(new_n915), .B2(new_n916), .ZN(new_n918));
  INV_X1    g717(.A(new_n911), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n562), .A2(new_n231), .ZN(new_n920));
  AOI22_X1  g719(.A1(new_n917), .A2(new_n918), .B1(new_n919), .B2(new_n920), .ZN(G1346gat));
  NOR2_X1   g720(.A1(new_n643), .A2(new_n232), .ZN(new_n922));
  NAND4_X1  g721(.A1(new_n886), .A2(new_n644), .A3(new_n888), .A4(new_n890), .ZN(new_n923));
  AOI22_X1  g722(.A1(new_n919), .A2(new_n922), .B1(new_n923), .B2(new_n232), .ZN(G1347gat));
  NOR2_X1   g723(.A1(new_n705), .A2(new_n701), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n847), .A2(new_n925), .ZN(new_n926));
  NOR3_X1   g725(.A1(new_n926), .A2(new_n282), .A3(new_n722), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n880), .A2(new_n422), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT124), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n705), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n880), .A2(KEYINPUT124), .A3(new_n422), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n930), .A2(new_n468), .A3(new_n931), .ZN(new_n932));
  OR2_X1    g731(.A1(new_n932), .A2(new_n722), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n927), .B1(new_n933), .B2(new_n282), .ZN(G1348gat));
  OAI21_X1  g733(.A(G176gat), .B1(new_n926), .B2(new_n772), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n665), .A2(new_n283), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n935), .B1(new_n932), .B2(new_n936), .ZN(G1349gat));
  NAND2_X1  g736(.A1(new_n721), .A2(new_n339), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n926), .A2(new_n562), .ZN(new_n939));
  OAI22_X1  g738(.A1(new_n932), .A2(new_n938), .B1(new_n346), .B2(new_n939), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n940), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g740(.A(G190gat), .B1(new_n926), .B2(new_n643), .ZN(new_n942));
  AND2_X1   g741(.A1(new_n942), .A2(KEYINPUT61), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n942), .A2(KEYINPUT61), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n644), .A2(new_n330), .ZN(new_n945));
  OAI22_X1  g744(.A1(new_n943), .A2(new_n944), .B1(new_n932), .B2(new_n945), .ZN(G1351gat));
  NAND2_X1  g745(.A1(new_n928), .A2(new_n929), .ZN(new_n947));
  INV_X1    g746(.A(new_n889), .ZN(new_n948));
  NAND4_X1  g747(.A1(new_n947), .A2(new_n708), .A3(new_n948), .A4(new_n931), .ZN(new_n949));
  INV_X1    g748(.A(new_n949), .ZN(new_n950));
  AOI21_X1  g749(.A(G197gat), .B1(new_n950), .B2(new_n698), .ZN(new_n951));
  INV_X1    g750(.A(new_n907), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n714), .A2(new_n925), .ZN(new_n953));
  XOR2_X1   g752(.A(new_n953), .B(KEYINPUT125), .Z(new_n954));
  NAND2_X1  g753(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  INV_X1    g754(.A(new_n955), .ZN(new_n956));
  AND2_X1   g755(.A1(new_n698), .A2(G197gat), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n951), .B1(new_n956), .B2(new_n957), .ZN(G1352gat));
  OR2_X1    g757(.A1(new_n772), .A2(G204gat), .ZN(new_n959));
  OAI21_X1  g758(.A(KEYINPUT62), .B1(new_n949), .B2(new_n959), .ZN(new_n960));
  OAI21_X1  g759(.A(G204gat), .B1(new_n955), .B2(new_n772), .ZN(new_n961));
  NOR3_X1   g760(.A1(new_n949), .A2(KEYINPUT62), .A3(new_n959), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n962), .A2(KEYINPUT126), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT126), .ZN(new_n964));
  NOR4_X1   g763(.A1(new_n949), .A2(new_n964), .A3(KEYINPUT62), .A4(new_n959), .ZN(new_n965));
  OAI211_X1 g764(.A(new_n960), .B(new_n961), .C1(new_n963), .C2(new_n965), .ZN(G1353gat));
  NAND3_X1  g765(.A1(new_n950), .A2(new_n206), .A3(new_n721), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n952), .A2(new_n721), .A3(new_n954), .ZN(new_n968));
  AND3_X1   g767(.A1(new_n968), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n969));
  AOI21_X1  g768(.A(KEYINPUT63), .B1(new_n968), .B2(G211gat), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n967), .B1(new_n969), .B2(new_n970), .ZN(G1354gat));
  OAI21_X1  g770(.A(new_n207), .B1(new_n949), .B2(new_n643), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n972), .A2(KEYINPUT127), .ZN(new_n973));
  INV_X1    g772(.A(KEYINPUT127), .ZN(new_n974));
  OAI211_X1 g773(.A(new_n974), .B(new_n207), .C1(new_n949), .C2(new_n643), .ZN(new_n975));
  NOR2_X1   g774(.A1(new_n643), .A2(new_n207), .ZN(new_n976));
  AOI22_X1  g775(.A1(new_n973), .A2(new_n975), .B1(new_n956), .B2(new_n976), .ZN(G1355gat));
endmodule


