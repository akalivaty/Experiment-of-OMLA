//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 1 1 1 1 0 0 0 0 0 0 0 1 1 1 0 1 0 0 0 1 1 0 1 1 0 1 0 1 1 1 1 0 0 0 0 0 0 1 0 0 0 0 0 0 0 1 0 0 1 0 0 1 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:37 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n545, new_n546, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n561, new_n562,
    new_n563, new_n565, new_n566, new_n567, new_n568, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n593, new_n596, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT65), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  INV_X1    g022(.A(G567), .ZN(new_n448));
  NOR2_X1   g023(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT66), .Z(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT67), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(G2106), .ZN(new_n458));
  OAI22_X1  g033(.A1(new_n453), .A2(new_n458), .B1(new_n448), .B2(new_n454), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  NAND2_X1  g035(.A1(G113), .A2(G2104), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G125), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n461), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n462), .A2(KEYINPUT68), .A3(KEYINPUT3), .ZN(new_n470));
  AND2_X1   g045(.A1(new_n470), .A2(new_n465), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT68), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n473), .B1(new_n464), .B2(G2104), .ZN(new_n474));
  NAND4_X1  g049(.A1(new_n471), .A2(G137), .A3(new_n472), .A4(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n462), .A2(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G101), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n469), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G160));
  NAND3_X1  g054(.A1(new_n471), .A2(G2105), .A3(new_n474), .ZN(new_n480));
  INV_X1    g055(.A(G124), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n472), .A2(G112), .ZN(new_n482));
  OAI21_X1  g057(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n483));
  OAI22_X1  g058(.A1(new_n480), .A2(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND4_X1  g059(.A1(new_n474), .A2(new_n470), .A3(new_n472), .A4(new_n465), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n484), .B1(G136), .B2(new_n486), .ZN(G162));
  AND2_X1   g062(.A1(KEYINPUT4), .A2(G138), .ZN(new_n488));
  NAND4_X1  g063(.A1(new_n474), .A2(new_n470), .A3(new_n465), .A4(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(G102), .A2(G2104), .ZN(new_n490));
  AOI21_X1  g065(.A(G2105), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n474), .A2(new_n470), .A3(G126), .A4(new_n465), .ZN(new_n492));
  NAND2_X1  g067(.A1(G114), .A2(G2104), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n472), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  XNOR2_X1  g069(.A(KEYINPUT3), .B(G2104), .ZN(new_n495));
  AND2_X1   g070(.A1(new_n472), .A2(G138), .ZN(new_n496));
  AOI21_X1  g071(.A(KEYINPUT4), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NOR3_X1   g072(.A1(new_n491), .A2(new_n494), .A3(new_n497), .ZN(G164));
  INV_X1    g073(.A(G543), .ZN(new_n499));
  OR2_X1    g074(.A1(KEYINPUT6), .A2(G651), .ZN(new_n500));
  NAND2_X1  g075(.A1(KEYINPUT6), .A2(G651), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G50), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n500), .A2(new_n501), .ZN(new_n504));
  XNOR2_X1  g079(.A(KEYINPUT5), .B(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  XOR2_X1   g081(.A(KEYINPUT69), .B(G88), .Z(new_n507));
  OAI21_X1  g082(.A(new_n503), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n505), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n509));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n508), .A2(new_n511), .ZN(G166));
  NAND3_X1  g087(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n513));
  XNOR2_X1  g088(.A(new_n513), .B(KEYINPUT7), .ZN(new_n514));
  INV_X1    g089(.A(new_n502), .ZN(new_n515));
  XOR2_X1   g090(.A(KEYINPUT70), .B(G51), .Z(new_n516));
  OAI21_X1  g091(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  AND2_X1   g092(.A1(KEYINPUT5), .A2(G543), .ZN(new_n518));
  NOR2_X1   g093(.A1(KEYINPUT5), .A2(G543), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n504), .A2(G89), .ZN(new_n521));
  NAND2_X1  g096(.A1(G63), .A2(G651), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n517), .A2(new_n523), .ZN(G168));
  NAND2_X1  g099(.A1(new_n502), .A2(G52), .ZN(new_n525));
  INV_X1    g100(.A(G90), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n525), .B1(new_n526), .B2(new_n506), .ZN(new_n527));
  AOI22_X1  g102(.A1(new_n505), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n528), .A2(new_n510), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n527), .A2(new_n529), .ZN(G171));
  NAND2_X1  g105(.A1(G68), .A2(G543), .ZN(new_n531));
  INV_X1    g106(.A(G56), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n531), .B1(new_n520), .B2(new_n532), .ZN(new_n533));
  AOI21_X1  g108(.A(KEYINPUT71), .B1(new_n533), .B2(G651), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n502), .A2(G43), .ZN(new_n535));
  INV_X1    g110(.A(G81), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n535), .B1(new_n536), .B2(new_n506), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n534), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n533), .A2(KEYINPUT71), .A3(G651), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G860), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n542), .B(KEYINPUT72), .ZN(G153));
  NAND4_X1  g118(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g119(.A1(G1), .A2(G3), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT8), .ZN(new_n546));
  NAND4_X1  g121(.A1(G319), .A2(G483), .A3(G661), .A4(new_n546), .ZN(G188));
  NAND2_X1  g122(.A1(new_n502), .A2(G53), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT9), .ZN(new_n549));
  INV_X1    g124(.A(KEYINPUT73), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n506), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n504), .A2(new_n505), .A3(KEYINPUT73), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n551), .A2(G91), .A3(new_n552), .ZN(new_n553));
  XNOR2_X1  g128(.A(KEYINPUT74), .B(G65), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n520), .A2(new_n554), .ZN(new_n555));
  AOI21_X1  g130(.A(new_n555), .B1(G78), .B2(G543), .ZN(new_n556));
  OAI211_X1 g131(.A(new_n549), .B(new_n553), .C1(new_n510), .C2(new_n556), .ZN(G299));
  INV_X1    g132(.A(G171), .ZN(G301));
  INV_X1    g133(.A(G168), .ZN(G286));
  INV_X1    g134(.A(G166), .ZN(G303));
  NAND3_X1  g135(.A1(new_n551), .A2(G87), .A3(new_n552), .ZN(new_n561));
  OR2_X1    g136(.A1(new_n505), .A2(G74), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n562), .A2(G651), .B1(new_n502), .B2(G49), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n561), .A2(new_n563), .ZN(G288));
  AOI22_X1  g139(.A1(new_n505), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n565));
  INV_X1    g140(.A(new_n565), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n566), .A2(G651), .B1(G48), .B2(new_n502), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n551), .A2(G86), .A3(new_n552), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n567), .A2(new_n568), .ZN(G305));
  NAND2_X1  g144(.A1(new_n502), .A2(G47), .ZN(new_n570));
  INV_X1    g145(.A(G85), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n570), .B1(new_n571), .B2(new_n506), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n505), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n573));
  NOR2_X1   g148(.A1(new_n573), .A2(new_n510), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT75), .ZN(new_n575));
  OR3_X1    g150(.A1(new_n572), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n572), .B2(new_n574), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(G290));
  INV_X1    g153(.A(G868), .ZN(new_n579));
  NOR2_X1   g154(.A1(G171), .A2(new_n579), .ZN(new_n580));
  XNOR2_X1  g155(.A(new_n580), .B(KEYINPUT76), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n502), .A2(G54), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n505), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n582), .B1(new_n583), .B2(new_n510), .ZN(new_n584));
  AND2_X1   g159(.A1(new_n551), .A2(new_n552), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n585), .A2(G92), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT10), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n585), .A2(KEYINPUT10), .A3(G92), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n584), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n581), .B1(G868), .B2(new_n590), .ZN(G284));
  OAI21_X1  g166(.A(new_n581), .B1(G868), .B2(new_n590), .ZN(G321));
  NAND2_X1  g167(.A1(G299), .A2(new_n579), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n593), .B1(new_n579), .B2(G168), .ZN(G297));
  OAI21_X1  g169(.A(new_n593), .B1(new_n579), .B2(G168), .ZN(G280));
  INV_X1    g170(.A(G559), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n590), .B1(new_n596), .B2(G860), .ZN(G148));
  NAND2_X1  g172(.A1(new_n540), .A2(new_n579), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n588), .A2(new_n589), .ZN(new_n599));
  INV_X1    g174(.A(new_n584), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n601), .A2(G559), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n598), .B1(new_n602), .B2(new_n579), .ZN(G323));
  XNOR2_X1  g178(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g179(.A1(new_n495), .A2(new_n476), .ZN(new_n605));
  XOR2_X1   g180(.A(new_n605), .B(KEYINPUT12), .Z(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(KEYINPUT13), .ZN(new_n607));
  XOR2_X1   g182(.A(new_n607), .B(G2100), .Z(new_n608));
  INV_X1    g183(.A(G123), .ZN(new_n609));
  NOR2_X1   g184(.A1(new_n472), .A2(G111), .ZN(new_n610));
  OAI21_X1  g185(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n611));
  OAI22_X1  g186(.A1(new_n480), .A2(new_n609), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  AND2_X1   g187(.A1(new_n486), .A2(G135), .ZN(new_n613));
  NOR2_X1   g188(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(new_n614), .ZN(new_n615));
  OR2_X1    g190(.A1(new_n615), .A2(G2096), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n615), .A2(G2096), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n608), .A2(new_n616), .A3(new_n617), .ZN(G156));
  XNOR2_X1  g193(.A(KEYINPUT15), .B(G2435), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(G2438), .ZN(new_n620));
  XNOR2_X1  g195(.A(G2427), .B(G2430), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n622), .A2(KEYINPUT14), .ZN(new_n623));
  AND2_X1   g198(.A1(new_n623), .A2(KEYINPUT77), .ZN(new_n624));
  NOR2_X1   g199(.A1(new_n623), .A2(KEYINPUT77), .ZN(new_n625));
  OAI22_X1  g200(.A1(new_n624), .A2(new_n625), .B1(new_n620), .B2(new_n621), .ZN(new_n626));
  XOR2_X1   g201(.A(G2443), .B(G2446), .Z(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(G2451), .B(G2454), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT16), .ZN(new_n630));
  INV_X1    g205(.A(new_n630), .ZN(new_n631));
  OR2_X1    g206(.A1(new_n628), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n628), .A2(new_n631), .ZN(new_n633));
  XNOR2_X1  g208(.A(G1341), .B(G1348), .ZN(new_n634));
  INV_X1    g209(.A(new_n634), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n632), .A2(new_n633), .A3(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT78), .ZN(new_n637));
  INV_X1    g212(.A(G14), .ZN(new_n638));
  AOI21_X1  g213(.A(new_n635), .B1(new_n632), .B2(new_n633), .ZN(new_n639));
  NOR3_X1   g214(.A1(new_n637), .A2(new_n638), .A3(new_n639), .ZN(G401));
  XOR2_X1   g215(.A(G2072), .B(G2078), .Z(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2067), .B(G2678), .ZN(new_n643));
  XOR2_X1   g218(.A(G2084), .B(G2090), .Z(new_n644));
  NAND3_X1  g219(.A1(new_n642), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n645), .B(KEYINPUT18), .Z(new_n646));
  INV_X1    g221(.A(new_n643), .ZN(new_n647));
  AOI21_X1  g222(.A(new_n644), .B1(new_n647), .B2(new_n641), .ZN(new_n648));
  XOR2_X1   g223(.A(KEYINPUT79), .B(KEYINPUT17), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n641), .B(new_n649), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n648), .B1(new_n650), .B2(new_n647), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n650), .A2(new_n647), .A3(new_n644), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n646), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(G2096), .B(G2100), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(G227));
  XNOR2_X1  g230(.A(G1991), .B(G1996), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G1971), .B(G1976), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT19), .ZN(new_n659));
  XOR2_X1   g234(.A(G1956), .B(G2474), .Z(new_n660));
  XOR2_X1   g235(.A(G1961), .B(G1966), .Z(new_n661));
  AND2_X1   g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT20), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n660), .A2(new_n661), .ZN(new_n665));
  NOR3_X1   g240(.A1(new_n659), .A2(new_n662), .A3(new_n665), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n666), .B1(new_n659), .B2(new_n665), .ZN(new_n667));
  AND2_X1   g242(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(G1981), .ZN(new_n669));
  INV_X1    g244(.A(G1986), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT80), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n671), .A2(new_n673), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n657), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  OR2_X1    g252(.A1(new_n671), .A2(new_n673), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n678), .A2(new_n656), .A3(new_n674), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n677), .A2(new_n679), .ZN(G229));
  INV_X1    g255(.A(G29), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n681), .A2(G35), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n682), .B1(G162), .B2(new_n681), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n683), .B(KEYINPUT29), .Z(new_n684));
  INV_X1    g259(.A(G2090), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT98), .ZN(new_n687));
  NAND2_X1  g262(.A1(G299), .A2(G16), .ZN(new_n688));
  INV_X1    g263(.A(G16), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n689), .A2(G20), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT99), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT23), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n688), .A2(new_n692), .ZN(new_n693));
  XOR2_X1   g268(.A(new_n693), .B(KEYINPUT100), .Z(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(G1956), .ZN(new_n695));
  OR2_X1    g270(.A1(new_n684), .A2(new_n685), .ZN(new_n696));
  OR2_X1    g271(.A1(new_n694), .A2(G1956), .ZN(new_n697));
  NAND4_X1  g272(.A1(new_n687), .A2(new_n695), .A3(new_n696), .A4(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(G168), .A2(G16), .ZN(new_n699));
  OAI211_X1 g274(.A(new_n699), .B(KEYINPUT91), .C1(G16), .C2(G21), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n700), .B1(KEYINPUT91), .B2(new_n699), .ZN(new_n701));
  XOR2_X1   g276(.A(KEYINPUT92), .B(G1966), .Z(new_n702));
  XOR2_X1   g277(.A(new_n701), .B(new_n702), .Z(new_n703));
  NAND2_X1  g278(.A1(new_n689), .A2(G19), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(new_n541), .B2(new_n689), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(G1341), .ZN(new_n706));
  NOR2_X1   g281(.A1(G171), .A2(new_n689), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n707), .B1(G5), .B2(new_n689), .ZN(new_n708));
  INV_X1    g283(.A(G1961), .ZN(new_n709));
  INV_X1    g284(.A(G2084), .ZN(new_n710));
  INV_X1    g285(.A(KEYINPUT24), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n681), .B1(new_n711), .B2(G34), .ZN(new_n712));
  OR2_X1    g287(.A1(new_n712), .A2(KEYINPUT89), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n712), .A2(KEYINPUT89), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n711), .A2(G34), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n713), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(new_n478), .B2(new_n681), .ZN(new_n717));
  OAI22_X1  g292(.A1(new_n708), .A2(new_n709), .B1(new_n710), .B2(new_n717), .ZN(new_n718));
  NOR3_X1   g293(.A1(new_n703), .A2(new_n706), .A3(new_n718), .ZN(new_n719));
  XOR2_X1   g294(.A(KEYINPUT31), .B(G11), .Z(new_n720));
  INV_X1    g295(.A(KEYINPUT30), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n681), .B1(new_n721), .B2(G28), .ZN(new_n722));
  INV_X1    g297(.A(KEYINPUT93), .ZN(new_n723));
  OR2_X1    g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  AOI22_X1  g299(.A1(new_n722), .A2(new_n723), .B1(new_n721), .B2(G28), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n720), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(new_n615), .B2(new_n681), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(KEYINPUT94), .Z(new_n728));
  XOR2_X1   g303(.A(KEYINPUT97), .B(G2078), .Z(new_n729));
  NAND2_X1  g304(.A1(new_n681), .A2(G27), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(KEYINPUT96), .Z(new_n731));
  NAND2_X1  g306(.A1(new_n489), .A2(new_n490), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n732), .A2(new_n472), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n492), .A2(new_n493), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(G2105), .ZN(new_n735));
  INV_X1    g310(.A(new_n497), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n733), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n731), .B1(new_n737), .B2(G29), .ZN(new_n738));
  OAI211_X1 g313(.A(new_n719), .B(new_n728), .C1(new_n729), .C2(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n681), .A2(G26), .ZN(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(KEYINPUT28), .Z(new_n741));
  NAND2_X1  g316(.A1(new_n486), .A2(G140), .ZN(new_n742));
  INV_X1    g317(.A(G128), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n472), .A2(G116), .ZN(new_n744));
  OAI21_X1  g319(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n745));
  OAI221_X1 g320(.A(new_n742), .B1(new_n480), .B2(new_n743), .C1(new_n744), .C2(new_n745), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT84), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n741), .B1(new_n747), .B2(G29), .ZN(new_n748));
  INV_X1    g323(.A(G2067), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  NOR2_X1   g325(.A1(G4), .A2(G16), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(new_n590), .B2(G16), .ZN(new_n752));
  OR2_X1    g327(.A1(new_n752), .A2(G1348), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n738), .A2(new_n729), .ZN(new_n754));
  INV_X1    g329(.A(KEYINPUT90), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(G29), .B2(G32), .ZN(new_n756));
  NAND3_X1  g331(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT26), .ZN(new_n758));
  OR2_X1    g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n757), .A2(new_n758), .ZN(new_n760));
  AOI22_X1  g335(.A1(new_n759), .A2(new_n760), .B1(G105), .B2(new_n476), .ZN(new_n761));
  INV_X1    g336(.A(G129), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n761), .B1(new_n480), .B2(new_n762), .ZN(new_n763));
  AND2_X1   g338(.A1(new_n486), .A2(G141), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n765), .A2(G29), .ZN(new_n766));
  MUX2_X1   g341(.A(new_n755), .B(new_n756), .S(new_n766), .Z(new_n767));
  XNOR2_X1  g342(.A(KEYINPUT27), .B(G1996), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n752), .A2(G1348), .ZN(new_n770));
  NAND4_X1  g345(.A1(new_n753), .A2(new_n754), .A3(new_n769), .A4(new_n770), .ZN(new_n771));
  NOR4_X1   g346(.A1(new_n698), .A2(new_n739), .A3(new_n750), .A4(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n689), .A2(G6), .ZN(new_n773));
  INV_X1    g348(.A(G305), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n773), .B1(new_n774), .B2(new_n689), .ZN(new_n775));
  XOR2_X1   g350(.A(KEYINPUT32), .B(G1981), .Z(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  NOR2_X1   g352(.A1(G16), .A2(G23), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT83), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G288), .B2(new_n689), .ZN(new_n780));
  XNOR2_X1  g355(.A(KEYINPUT33), .B(G1976), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  OR2_X1    g357(.A1(new_n780), .A2(new_n781), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n689), .A2(G22), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(G166), .B2(new_n689), .ZN(new_n785));
  INV_X1    g360(.A(G1971), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NAND4_X1  g362(.A1(new_n777), .A2(new_n782), .A3(new_n783), .A4(new_n787), .ZN(new_n788));
  OR2_X1    g363(.A1(new_n788), .A2(KEYINPUT34), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n788), .A2(KEYINPUT34), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n689), .A2(G24), .ZN(new_n791));
  INV_X1    g366(.A(G290), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n791), .B1(new_n792), .B2(new_n689), .ZN(new_n793));
  XOR2_X1   g368(.A(KEYINPUT82), .B(G1986), .Z(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n681), .A2(G25), .ZN(new_n796));
  INV_X1    g371(.A(G119), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n480), .A2(new_n797), .ZN(new_n798));
  XOR2_X1   g373(.A(new_n798), .B(KEYINPUT81), .Z(new_n799));
  OAI21_X1  g374(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n800));
  INV_X1    g375(.A(G107), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n800), .B1(new_n801), .B2(G2105), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(new_n486), .B2(G131), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n799), .A2(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(new_n804), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n796), .B1(new_n805), .B2(new_n681), .ZN(new_n806));
  XOR2_X1   g381(.A(KEYINPUT35), .B(G1991), .Z(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  NAND4_X1  g383(.A1(new_n789), .A2(new_n790), .A3(new_n795), .A4(new_n808), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT36), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n681), .A2(G33), .ZN(new_n811));
  NAND3_X1  g386(.A1(new_n472), .A2(G103), .A3(G2104), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT86), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  OR2_X1    g389(.A1(new_n814), .A2(KEYINPUT85), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n814), .A2(KEYINPUT85), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT25), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(G139), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n485), .A2(new_n820), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT87), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n815), .A2(KEYINPUT25), .A3(new_n816), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n819), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT88), .ZN(new_n825));
  AOI22_X1  g400(.A1(new_n495), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n826), .A2(new_n472), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n811), .B1(new_n828), .B2(new_n681), .ZN(new_n829));
  OR2_X1    g404(.A1(new_n829), .A2(G2072), .ZN(new_n830));
  AOI22_X1  g405(.A1(new_n708), .A2(new_n709), .B1(new_n710), .B2(new_n717), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n831), .B1(new_n767), .B2(new_n768), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT95), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n829), .A2(G2072), .ZN(new_n834));
  AND3_X1   g409(.A1(new_n830), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n772), .A2(new_n810), .A3(new_n835), .ZN(G150));
  INV_X1    g411(.A(G150), .ZN(G311));
  NAND2_X1  g412(.A1(new_n590), .A2(G559), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(KEYINPUT38), .Z(new_n839));
  NAND2_X1  g414(.A1(G80), .A2(G543), .ZN(new_n840));
  INV_X1    g415(.A(G67), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n840), .B1(new_n520), .B2(new_n841), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n510), .B1(new_n842), .B2(KEYINPUT101), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n843), .B1(KEYINPUT101), .B2(new_n842), .ZN(new_n844));
  AND2_X1   g419(.A1(new_n504), .A2(new_n505), .ZN(new_n845));
  AOI22_X1  g420(.A1(new_n845), .A2(G93), .B1(G55), .B2(new_n502), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  OR2_X1    g422(.A1(new_n847), .A2(new_n540), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n847), .A2(new_n540), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n839), .B(new_n850), .ZN(new_n851));
  AND2_X1   g426(.A1(new_n851), .A2(KEYINPUT39), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n851), .A2(KEYINPUT39), .ZN(new_n853));
  NOR3_X1   g428(.A1(new_n852), .A2(new_n853), .A3(G860), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n847), .A2(G860), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(KEYINPUT37), .ZN(new_n856));
  OR2_X1    g431(.A1(new_n854), .A2(new_n856), .ZN(G145));
  XNOR2_X1  g432(.A(new_n614), .B(new_n478), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(G162), .ZN(new_n859));
  OR2_X1    g434(.A1(G106), .A2(G2105), .ZN(new_n860));
  OAI211_X1 g435(.A(new_n860), .B(G2104), .C1(G118), .C2(new_n472), .ZN(new_n861));
  INV_X1    g436(.A(G130), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n861), .B1(new_n480), .B2(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n863), .B1(G142), .B2(new_n486), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n805), .A2(KEYINPUT102), .ZN(new_n866));
  INV_X1    g441(.A(new_n606), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT102), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n804), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n866), .A2(new_n867), .A3(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n867), .B1(new_n866), .B2(new_n869), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n865), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n872), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n874), .A2(new_n864), .A3(new_n870), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT103), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n747), .B(new_n737), .ZN(new_n880));
  AND2_X1   g455(.A1(new_n828), .A2(new_n880), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n828), .A2(new_n880), .ZN(new_n882));
  INV_X1    g457(.A(new_n765), .ZN(new_n883));
  OR3_X1    g458(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n883), .B1(new_n881), .B2(new_n882), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n859), .B1(new_n879), .B2(new_n886), .ZN(new_n887));
  NAND4_X1  g462(.A1(new_n877), .A2(new_n884), .A3(new_n878), .A4(new_n885), .ZN(new_n888));
  AOI21_X1  g463(.A(G37), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n886), .A2(new_n876), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n877), .B1(new_n884), .B2(new_n885), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n859), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  AND3_X1   g467(.A1(new_n889), .A2(new_n892), .A3(KEYINPUT40), .ZN(new_n893));
  AOI21_X1  g468(.A(KEYINPUT40), .B1(new_n889), .B2(new_n892), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n893), .A2(new_n894), .ZN(G395));
  NAND2_X1  g470(.A1(new_n847), .A2(new_n579), .ZN(new_n896));
  OR2_X1    g471(.A1(new_n601), .A2(G299), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n601), .A2(G299), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT41), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n897), .A2(KEYINPUT41), .A3(new_n898), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n602), .B(new_n850), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n899), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n905), .B1(new_n906), .B2(new_n904), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n907), .B(KEYINPUT42), .ZN(new_n908));
  XNOR2_X1  g483(.A(G290), .B(G305), .ZN(new_n909));
  XNOR2_X1  g484(.A(G288), .B(G166), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n909), .B(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n912), .A2(KEYINPUT104), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n908), .B(new_n913), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n896), .B1(new_n914), .B2(new_n579), .ZN(G295));
  OAI21_X1  g490(.A(new_n896), .B1(new_n914), .B2(new_n579), .ZN(G331));
  INV_X1    g491(.A(KEYINPUT44), .ZN(new_n917));
  XNOR2_X1  g492(.A(G171), .B(KEYINPUT106), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n918), .B1(new_n848), .B2(new_n849), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n848), .A2(new_n849), .A3(new_n918), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n920), .A2(G168), .A3(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n921), .ZN(new_n923));
  OAI21_X1  g498(.A(G286), .B1(new_n923), .B2(new_n919), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n906), .A2(new_n922), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n922), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  OAI211_X1 g502(.A(new_n912), .B(new_n925), .C1(new_n927), .C2(new_n903), .ZN(new_n928));
  INV_X1    g503(.A(G37), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n925), .B1(new_n927), .B2(new_n903), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n912), .B1(new_n931), .B2(KEYINPUT107), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT107), .ZN(new_n933));
  OAI211_X1 g508(.A(new_n933), .B(new_n925), .C1(new_n927), .C2(new_n903), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n930), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  XNOR2_X1  g510(.A(KEYINPUT105), .B(KEYINPUT43), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n917), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  AND2_X1   g512(.A1(new_n901), .A2(new_n902), .ZN(new_n938));
  AOI22_X1  g513(.A1(new_n938), .A2(new_n926), .B1(new_n925), .B2(KEYINPUT108), .ZN(new_n939));
  OR2_X1    g514(.A1(new_n925), .A2(KEYINPUT108), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n912), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  OAI21_X1  g516(.A(KEYINPUT43), .B1(new_n941), .B2(new_n930), .ZN(new_n942));
  AOI21_X1  g517(.A(KEYINPUT109), .B1(new_n937), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n931), .A2(KEYINPUT107), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n944), .A2(new_n911), .A3(new_n934), .ZN(new_n945));
  INV_X1    g520(.A(new_n930), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n945), .A2(new_n936), .A3(new_n946), .ZN(new_n947));
  AND4_X1   g522(.A1(KEYINPUT109), .A2(new_n947), .A3(new_n942), .A4(KEYINPUT44), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n935), .A2(new_n936), .ZN(new_n949));
  INV_X1    g524(.A(new_n936), .ZN(new_n950));
  NOR3_X1   g525(.A1(new_n941), .A2(new_n950), .A3(new_n930), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  OAI22_X1  g527(.A1(new_n943), .A2(new_n948), .B1(new_n952), .B2(KEYINPUT44), .ZN(G397));
  NAND2_X1  g528(.A1(new_n792), .A2(new_n670), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT45), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n955), .B1(G164), .B2(G1384), .ZN(new_n956));
  INV_X1    g531(.A(new_n956), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n469), .A2(G40), .A3(new_n475), .A4(new_n477), .ZN(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n954), .A2(new_n960), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n961), .B(KEYINPUT127), .ZN(new_n962));
  XOR2_X1   g537(.A(new_n962), .B(KEYINPUT48), .Z(new_n963));
  NOR2_X1   g538(.A1(new_n960), .A2(G1996), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n964), .B(KEYINPUT110), .ZN(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(new_n960), .ZN(new_n967));
  XNOR2_X1  g542(.A(new_n747), .B(new_n749), .ZN(new_n968));
  INV_X1    g543(.A(G1996), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n968), .B1(new_n969), .B2(new_n765), .ZN(new_n970));
  AOI22_X1  g545(.A1(new_n966), .A2(new_n765), .B1(new_n967), .B2(new_n970), .ZN(new_n971));
  AND2_X1   g546(.A1(new_n805), .A2(new_n807), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n805), .A2(new_n807), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n967), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n971), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT126), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n963), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n977), .B1(new_n976), .B2(new_n975), .ZN(new_n978));
  AND2_X1   g553(.A1(new_n971), .A2(new_n972), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n747), .A2(G2067), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n981), .A2(new_n960), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n960), .B1(new_n968), .B2(new_n765), .ZN(new_n983));
  OR2_X1    g558(.A1(new_n965), .A2(KEYINPUT46), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n965), .A2(KEYINPUT46), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n983), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  XNOR2_X1  g561(.A(new_n986), .B(KEYINPUT47), .ZN(new_n987));
  NOR3_X1   g562(.A1(new_n978), .A2(new_n982), .A3(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(G290), .A2(G1986), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n960), .B1(new_n954), .B2(new_n989), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n975), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(G8), .ZN(new_n992));
  NOR2_X1   g567(.A1(G168), .A2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(new_n993), .ZN(new_n994));
  OAI21_X1  g569(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n995));
  NOR2_X1   g570(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n958), .B1(new_n737), .B2(new_n996), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n995), .A2(new_n997), .A3(new_n710), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(KEYINPUT118), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT118), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n995), .A2(new_n997), .A3(new_n1000), .A4(new_n710), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n497), .B1(new_n734), .B2(G2105), .ZN(new_n1002));
  AOI21_X1  g577(.A(G1384), .B1(new_n1002), .B2(new_n733), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n959), .B1(new_n1003), .B2(KEYINPUT45), .ZN(new_n1004));
  NOR3_X1   g579(.A1(G164), .A2(new_n955), .A3(G1384), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n702), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n999), .A2(new_n1001), .A3(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(KEYINPUT122), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT122), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n999), .A2(new_n1009), .A3(new_n1006), .A4(new_n1001), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n994), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1008), .A2(G168), .A3(new_n1010), .ZN(new_n1012));
  AND2_X1   g587(.A1(KEYINPUT51), .A2(G8), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1007), .A2(G8), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n993), .A2(KEYINPUT51), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1011), .B1(new_n1014), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT62), .ZN(new_n1019));
  OAI21_X1  g594(.A(KEYINPUT124), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n992), .B1(new_n1003), .B2(new_n959), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n502), .A2(G48), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n504), .A2(new_n505), .A3(G86), .ZN(new_n1024));
  OAI211_X1 g599(.A(new_n1023), .B(new_n1024), .C1(new_n565), .C2(new_n510), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(G1981), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(KEYINPUT113), .ZN(new_n1027));
  INV_X1    g602(.A(G1981), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n567), .A2(new_n1028), .A3(new_n568), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT113), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1025), .A2(new_n1030), .A3(G1981), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1027), .A2(new_n1029), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1032), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1022), .B1(new_n1033), .B2(KEYINPUT49), .ZN(new_n1034));
  XOR2_X1   g609(.A(KEYINPUT114), .B(KEYINPUT49), .Z(new_n1035));
  AND3_X1   g610(.A1(new_n1032), .A2(KEYINPUT115), .A3(new_n1035), .ZN(new_n1036));
  AOI21_X1  g611(.A(KEYINPUT115), .B1(new_n1032), .B2(new_n1035), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1034), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n561), .A2(new_n563), .A3(G1976), .ZN(new_n1039));
  INV_X1    g614(.A(G1976), .ZN(new_n1040));
  AOI21_X1  g615(.A(KEYINPUT52), .B1(G288), .B2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1021), .A2(new_n1039), .A3(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT112), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n1021), .A2(KEYINPUT112), .A3(new_n1039), .A4(new_n1041), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1021), .A2(new_n1039), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(KEYINPUT52), .ZN(new_n1048));
  AND3_X1   g623(.A1(new_n1038), .A2(new_n1046), .A3(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT117), .ZN(new_n1050));
  INV_X1    g625(.A(G1384), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n737), .A2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n958), .B1(new_n1052), .B2(new_n955), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1003), .A2(KEYINPUT45), .ZN(new_n1054));
  AOI21_X1  g629(.A(G1971), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n995), .A2(new_n997), .A3(new_n685), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1056), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1050), .B1(new_n1055), .B2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n956), .A2(new_n1054), .A3(new_n959), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(new_n786), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1060), .A2(KEYINPUT117), .A3(new_n1056), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1058), .A2(G8), .A3(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(G303), .A2(G8), .ZN(new_n1063));
  XOR2_X1   g638(.A(new_n1063), .B(KEYINPUT55), .Z(new_n1064));
  INV_X1    g639(.A(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1062), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT111), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n1067), .B(new_n786), .C1(new_n1004), .C2(new_n1005), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(new_n1056), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1067), .B1(new_n1059), .B2(new_n786), .ZN(new_n1070));
  OAI211_X1 g645(.A(G8), .B(new_n1064), .C1(new_n1069), .C2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(G2078), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n956), .A2(new_n1054), .A3(new_n1072), .A4(new_n959), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT53), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1053), .A2(KEYINPUT53), .A3(new_n1072), .A4(new_n1054), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1077), .ZN(new_n1078));
  AND2_X1   g653(.A1(new_n995), .A2(new_n997), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1079), .A2(G1961), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(G301), .B1(new_n1078), .B2(new_n1081), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1049), .A2(new_n1066), .A3(new_n1071), .A4(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1083), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT124), .ZN(new_n1085));
  AOI22_X1  g660(.A1(new_n1012), .A2(new_n1013), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1086));
  OAI211_X1 g661(.A(new_n1085), .B(KEYINPUT62), .C1(new_n1086), .C2(new_n1011), .ZN(new_n1087));
  AND3_X1   g662(.A1(new_n1020), .A2(new_n1084), .A3(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1071), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1038), .A2(new_n1046), .A3(new_n1048), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1007), .A2(G8), .A3(G168), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1092), .ZN(new_n1093));
  OAI21_X1  g668(.A(G8), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(new_n1065), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1091), .A2(KEYINPUT63), .A3(new_n1093), .A4(new_n1095), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1071), .A2(new_n1046), .A3(new_n1048), .A4(new_n1038), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1060), .A2(new_n1056), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n992), .B1(new_n1098), .B2(new_n1050), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1064), .B1(new_n1099), .B2(new_n1061), .ZN(new_n1100));
  NOR3_X1   g675(.A1(new_n1097), .A2(new_n1100), .A3(new_n1092), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1096), .B1(new_n1101), .B2(KEYINPUT63), .ZN(new_n1102));
  NOR2_X1   g677(.A1(G288), .A2(G1976), .ZN(new_n1103));
  AOI22_X1  g678(.A1(new_n1038), .A2(new_n1103), .B1(new_n1028), .B2(new_n774), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1022), .B1(new_n1105), .B2(KEYINPUT116), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT116), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1104), .A2(new_n1107), .ZN(new_n1108));
  AOI22_X1  g683(.A1(new_n1106), .A2(new_n1108), .B1(new_n1089), .B2(new_n1049), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT57), .ZN(new_n1110));
  XNOR2_X1  g685(.A(G299), .B(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n995), .A2(new_n997), .ZN(new_n1112));
  INV_X1    g687(.A(G1956), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  XNOR2_X1  g689(.A(KEYINPUT56), .B(G2072), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n956), .A2(new_n1054), .A3(new_n959), .A4(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1111), .A2(new_n1114), .A3(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(G1348), .B1(new_n995), .B2(new_n997), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1003), .A2(new_n959), .A3(new_n749), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1120), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n590), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1122), .A2(KEYINPUT119), .ZN(new_n1123));
  XNOR2_X1  g698(.A(G299), .B(KEYINPUT57), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1123), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1122), .A2(KEYINPUT119), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1118), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n956), .A2(new_n1054), .A3(new_n969), .A4(new_n959), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT120), .ZN(new_n1130));
  XOR2_X1   g705(.A(KEYINPUT58), .B(G1341), .Z(new_n1131));
  OAI21_X1  g706(.A(new_n1131), .B1(new_n1052), .B2(new_n958), .ZN(new_n1132));
  AND3_X1   g707(.A1(new_n1129), .A2(new_n1130), .A3(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1130), .B1(new_n1129), .B2(new_n1132), .ZN(new_n1134));
  OAI211_X1 g709(.A(KEYINPUT59), .B(new_n541), .C1(new_n1133), .C2(new_n1134), .ZN(new_n1135));
  OAI211_X1 g710(.A(new_n601), .B(new_n1120), .C1(new_n1079), .C2(G1348), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1136), .A2(new_n1122), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n601), .A2(KEYINPUT60), .ZN(new_n1139));
  AOI22_X1  g714(.A1(new_n1137), .A2(KEYINPUT60), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n541), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT59), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1125), .A2(new_n1124), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1144), .A2(KEYINPUT61), .A3(new_n1117), .ZN(new_n1145));
  AND4_X1   g720(.A1(new_n1135), .A2(new_n1140), .A3(new_n1143), .A4(new_n1145), .ZN(new_n1146));
  AOI21_X1  g721(.A(KEYINPUT61), .B1(new_n1144), .B2(new_n1117), .ZN(new_n1147));
  XNOR2_X1  g722(.A(new_n1147), .B(KEYINPUT121), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1128), .B1(new_n1146), .B2(new_n1148), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1097), .A2(new_n1100), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT123), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1075), .A2(new_n1151), .A3(new_n1076), .ZN(new_n1152));
  XOR2_X1   g727(.A(G171), .B(KEYINPUT54), .Z(new_n1153));
  INV_X1    g728(.A(new_n1153), .ZN(new_n1154));
  AOI22_X1  g729(.A1(new_n1078), .A2(new_n1081), .B1(new_n1152), .B2(new_n1154), .ZN(new_n1155));
  NOR4_X1   g730(.A1(new_n1077), .A2(new_n1080), .A3(new_n1151), .A4(new_n1153), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  OAI211_X1 g732(.A(new_n1150), .B(new_n1157), .C1(new_n1011), .C2(new_n1086), .ZN(new_n1158));
  OAI211_X1 g733(.A(new_n1102), .B(new_n1109), .C1(new_n1149), .C2(new_n1158), .ZN(new_n1159));
  OAI211_X1 g734(.A(KEYINPUT125), .B(new_n991), .C1(new_n1088), .C2(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(new_n1108), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1021), .B1(new_n1104), .B2(new_n1107), .ZN(new_n1163));
  OAI22_X1  g738(.A1(new_n1162), .A2(new_n1163), .B1(new_n1071), .B2(new_n1090), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1157), .A2(new_n1091), .A3(new_n1066), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1165), .A2(new_n1018), .ZN(new_n1166));
  INV_X1    g741(.A(new_n1128), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT121), .ZN(new_n1168));
  XNOR2_X1  g743(.A(new_n1147), .B(new_n1168), .ZN(new_n1169));
  NAND4_X1  g744(.A1(new_n1140), .A2(new_n1143), .A3(new_n1135), .A4(new_n1145), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1167), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1164), .B1(new_n1166), .B2(new_n1171), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1020), .A2(new_n1084), .A3(new_n1087), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1172), .A2(new_n1173), .A3(new_n1102), .ZN(new_n1174));
  AOI21_X1  g749(.A(KEYINPUT125), .B1(new_n1174), .B2(new_n991), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n988), .B1(new_n1161), .B2(new_n1175), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g751(.A1(new_n889), .A2(new_n892), .ZN(new_n1178));
  NOR2_X1   g752(.A1(G227), .A2(new_n459), .ZN(new_n1179));
  NAND3_X1  g753(.A1(new_n677), .A2(new_n679), .A3(new_n1179), .ZN(new_n1180));
  NOR2_X1   g754(.A1(new_n1180), .A2(G401), .ZN(new_n1181));
  NAND2_X1  g755(.A1(new_n1178), .A2(new_n1181), .ZN(new_n1182));
  NOR2_X1   g756(.A1(new_n1182), .A2(new_n952), .ZN(G308));
  OAI211_X1 g757(.A(new_n1178), .B(new_n1181), .C1(new_n949), .C2(new_n951), .ZN(G225));
endmodule


