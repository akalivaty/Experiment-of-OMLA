//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 0 0 1 0 0 1 1 0 0 0 0 0 0 1 0 0 1 0 0 0 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 0 1 0 1 1 0 0 0 1 0 0 1 0 0 0 1 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:38 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n713, new_n714, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n742, new_n743,
    new_n744, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n763, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT65), .ZN(new_n188));
  XNOR2_X1  g002(.A(KEYINPUT64), .B(G146), .ZN(new_n189));
  INV_X1    g003(.A(G143), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n188), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT64), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n192), .A2(G146), .ZN(new_n193));
  INV_X1    g007(.A(G146), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n194), .A2(KEYINPUT64), .ZN(new_n195));
  OAI211_X1 g009(.A(KEYINPUT65), .B(G143), .C1(new_n193), .C2(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n191), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT1), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n190), .A2(G146), .ZN(new_n199));
  OR2_X1    g013(.A1(new_n199), .A2(KEYINPUT66), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(KEYINPUT66), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n197), .A2(new_n198), .A3(G128), .A4(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G128), .ZN(new_n204));
  OAI21_X1  g018(.A(G143), .B1(new_n193), .B2(new_n195), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n204), .B1(new_n205), .B2(KEYINPUT1), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n190), .A2(G146), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n207), .B1(new_n189), .B2(new_n190), .ZN(new_n208));
  OAI21_X1  g022(.A(KEYINPUT69), .B1(new_n206), .B2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT69), .ZN(new_n210));
  INV_X1    g024(.A(new_n207), .ZN(new_n211));
  XOR2_X1   g025(.A(KEYINPUT64), .B(G146), .Z(new_n212));
  OAI21_X1  g026(.A(new_n211), .B1(new_n212), .B2(G143), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n198), .B1(new_n212), .B2(G143), .ZN(new_n214));
  OAI211_X1 g028(.A(new_n210), .B(new_n213), .C1(new_n214), .C2(new_n204), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n203), .A2(new_n209), .A3(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G104), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G107), .ZN(new_n218));
  INV_X1    g032(.A(new_n218), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n217), .A2(G107), .ZN(new_n220));
  OAI21_X1  g034(.A(G101), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  OAI21_X1  g035(.A(KEYINPUT3), .B1(new_n217), .B2(G107), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n223));
  INV_X1    g037(.A(G107), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n223), .A2(new_n224), .A3(G104), .ZN(new_n225));
  INV_X1    g039(.A(G101), .ZN(new_n226));
  NAND4_X1  g040(.A1(new_n222), .A2(new_n225), .A3(new_n226), .A4(new_n218), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n221), .A2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT10), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n216), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(KEYINPUT85), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT85), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n216), .A2(new_n233), .A3(new_n230), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n203), .A2(KEYINPUT84), .ZN(new_n236));
  AOI22_X1  g050(.A1(new_n191), .A2(new_n196), .B1(new_n201), .B2(new_n200), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n204), .B1(new_n211), .B2(KEYINPUT1), .ZN(new_n238));
  OR2_X1    g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT84), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n237), .A2(new_n240), .A3(new_n198), .A4(G128), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n236), .A2(new_n239), .A3(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(new_n228), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(new_n229), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n222), .A2(new_n225), .A3(new_n218), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G101), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n247), .A2(KEYINPUT4), .A3(new_n227), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(KEYINPUT83), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT83), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n247), .A2(new_n250), .A3(KEYINPUT4), .A4(new_n227), .ZN(new_n251));
  OAI211_X1 g065(.A(new_n249), .B(new_n251), .C1(KEYINPUT4), .C2(new_n247), .ZN(new_n252));
  AND2_X1   g066(.A1(KEYINPUT0), .A2(G128), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n237), .A2(new_n253), .ZN(new_n254));
  NOR2_X1   g068(.A1(KEYINPUT0), .A2(G128), .ZN(new_n255));
  NOR3_X1   g069(.A1(new_n208), .A2(new_n253), .A3(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n254), .A2(new_n257), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n252), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n235), .A2(new_n245), .A3(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(G137), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G134), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT67), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(KEYINPUT11), .ZN(new_n265));
  OR2_X1    g079(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  OR2_X1    g080(.A1(new_n264), .A2(KEYINPUT11), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n263), .A2(new_n265), .ZN(new_n268));
  INV_X1    g082(.A(G134), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(G137), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n266), .A2(new_n267), .A3(new_n268), .A4(new_n270), .ZN(new_n271));
  XNOR2_X1  g085(.A(new_n271), .B(G131), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n261), .A2(new_n272), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n259), .B1(new_n232), .B2(new_n234), .ZN(new_n274));
  INV_X1    g088(.A(new_n272), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n274), .A2(new_n275), .A3(new_n245), .ZN(new_n276));
  XNOR2_X1  g090(.A(G110), .B(G140), .ZN(new_n277));
  INV_X1    g091(.A(G953), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(G227), .ZN(new_n279));
  XNOR2_X1  g093(.A(new_n277), .B(new_n279), .ZN(new_n280));
  XNOR2_X1  g094(.A(KEYINPUT81), .B(KEYINPUT82), .ZN(new_n281));
  XOR2_X1   g095(.A(new_n280), .B(new_n281), .Z(new_n282));
  NAND3_X1  g096(.A1(new_n273), .A2(new_n276), .A3(new_n282), .ZN(new_n283));
  AND3_X1   g097(.A1(new_n235), .A2(new_n245), .A3(new_n260), .ZN(new_n284));
  AND4_X1   g098(.A1(new_n203), .A2(new_n209), .A3(new_n215), .A4(new_n228), .ZN(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n244), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n287), .A2(KEYINPUT12), .A3(new_n272), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT12), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n285), .B1(new_n242), .B2(new_n243), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n289), .B1(new_n290), .B2(new_n275), .ZN(new_n291));
  AOI22_X1  g105(.A1(new_n284), .A2(new_n275), .B1(new_n288), .B2(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n283), .B1(new_n292), .B2(new_n282), .ZN(new_n293));
  INV_X1    g107(.A(G902), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n187), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  AOI21_X1  g109(.A(KEYINPUT12), .B1(new_n287), .B2(new_n272), .ZN(new_n296));
  NOR3_X1   g110(.A1(new_n290), .A2(new_n289), .A3(new_n275), .ZN(new_n297));
  OAI211_X1 g111(.A(new_n276), .B(new_n282), .C1(new_n296), .C2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n282), .B1(new_n273), .B2(new_n276), .ZN(new_n300));
  OAI211_X1 g114(.A(new_n187), .B(new_n294), .C1(new_n299), .C2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT86), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(new_n282), .ZN(new_n304));
  AND3_X1   g118(.A1(new_n274), .A2(new_n275), .A3(new_n245), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n275), .B1(new_n274), .B2(new_n245), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n304), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  AOI21_X1  g121(.A(G902), .B1(new_n307), .B2(new_n298), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n308), .A2(KEYINPUT86), .A3(new_n187), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n295), .B1(new_n303), .B2(new_n309), .ZN(new_n310));
  XNOR2_X1  g124(.A(KEYINPUT9), .B(G234), .ZN(new_n311));
  OAI21_X1  g125(.A(G221), .B1(new_n311), .B2(G902), .ZN(new_n312));
  XOR2_X1   g126(.A(new_n312), .B(KEYINPUT80), .Z(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  OAI21_X1  g128(.A(KEYINPUT87), .B1(new_n310), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n293), .A2(new_n294), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(G469), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n307), .A2(new_n298), .ZN(new_n318));
  AND4_X1   g132(.A1(KEYINPUT86), .A2(new_n318), .A3(new_n187), .A4(new_n294), .ZN(new_n319));
  AOI21_X1  g133(.A(KEYINPUT86), .B1(new_n308), .B2(new_n187), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n317), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT87), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n321), .A2(new_n322), .A3(new_n313), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n315), .A2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT68), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n263), .A2(new_n270), .A3(new_n325), .ZN(new_n326));
  OAI211_X1 g140(.A(new_n326), .B(G131), .C1(new_n325), .C2(new_n263), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n327), .B1(new_n271), .B2(G131), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n216), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(KEYINPUT72), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n256), .B1(new_n253), .B2(new_n237), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n272), .A2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT72), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n216), .A2(new_n334), .A3(new_n329), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n331), .A2(new_n333), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(KEYINPUT30), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT30), .ZN(new_n338));
  AND3_X1   g152(.A1(new_n330), .A2(new_n338), .A3(new_n333), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n337), .A2(new_n340), .ZN(new_n341));
  XOR2_X1   g155(.A(KEYINPUT2), .B(G113), .Z(new_n342));
  INV_X1    g156(.A(G119), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(G116), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT70), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n345), .B1(new_n343), .B2(G116), .ZN(new_n346));
  INV_X1    g160(.A(G116), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n347), .A2(KEYINPUT70), .A3(G119), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n342), .B1(new_n344), .B2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n342), .A2(new_n349), .A3(new_n344), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n351), .A2(KEYINPUT71), .A3(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT71), .ZN(new_n354));
  INV_X1    g168(.A(new_n352), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n354), .B1(new_n355), .B2(new_n350), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n341), .A2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT31), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n331), .A2(new_n333), .A3(new_n357), .A4(new_n335), .ZN(new_n361));
  NOR2_X1   g175(.A1(G237), .A2(G953), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(G210), .ZN(new_n363));
  XOR2_X1   g177(.A(new_n363), .B(KEYINPUT27), .Z(new_n364));
  XNOR2_X1  g178(.A(new_n364), .B(KEYINPUT26), .ZN(new_n365));
  XNOR2_X1  g179(.A(new_n365), .B(new_n226), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n359), .A2(new_n360), .A3(new_n361), .A4(new_n366), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n339), .B1(new_n336), .B2(KEYINPUT30), .ZN(new_n368));
  OAI211_X1 g182(.A(new_n361), .B(new_n366), .C1(new_n368), .C2(new_n357), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(KEYINPUT31), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n330), .A2(new_n333), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(new_n358), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT28), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n373), .B1(new_n371), .B2(new_n358), .ZN(new_n374));
  OAI211_X1 g188(.A(new_n372), .B(new_n374), .C1(new_n361), .C2(new_n373), .ZN(new_n375));
  INV_X1    g189(.A(new_n366), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n367), .A2(new_n370), .A3(new_n377), .ZN(new_n378));
  NOR2_X1   g192(.A1(G472), .A2(G902), .ZN(new_n379));
  AND3_X1   g193(.A1(new_n378), .A2(KEYINPUT32), .A3(new_n379), .ZN(new_n380));
  AOI21_X1  g194(.A(KEYINPUT32), .B1(new_n378), .B2(new_n379), .ZN(new_n381));
  INV_X1    g195(.A(G472), .ZN(new_n382));
  OR2_X1    g196(.A1(new_n375), .A2(new_n376), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT29), .ZN(new_n384));
  INV_X1    g198(.A(new_n361), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n385), .B1(new_n341), .B2(new_n358), .ZN(new_n386));
  OAI211_X1 g200(.A(new_n383), .B(new_n384), .C1(new_n386), .C2(new_n366), .ZN(new_n387));
  INV_X1    g201(.A(new_n374), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n336), .A2(new_n358), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(new_n361), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n388), .B1(new_n390), .B2(KEYINPUT28), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n376), .A2(new_n384), .ZN(new_n392));
  AOI21_X1  g206(.A(G902), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n382), .B1(new_n387), .B2(new_n393), .ZN(new_n394));
  NOR3_X1   g208(.A1(new_n380), .A2(new_n381), .A3(new_n394), .ZN(new_n395));
  OAI21_X1  g209(.A(KEYINPUT23), .B1(new_n204), .B2(G119), .ZN(new_n396));
  OAI211_X1 g210(.A(new_n396), .B(KEYINPUT74), .C1(new_n343), .C2(G128), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n343), .A2(G128), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT74), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n398), .B1(new_n399), .B2(KEYINPUT23), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n397), .A2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT75), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n397), .A2(KEYINPUT75), .A3(new_n400), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n403), .A2(G110), .A3(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(G140), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(G125), .ZN(new_n407));
  OAI21_X1  g221(.A(KEYINPUT76), .B1(new_n407), .B2(KEYINPUT16), .ZN(new_n408));
  INV_X1    g222(.A(G125), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(G140), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n407), .A2(new_n410), .A3(KEYINPUT16), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT76), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT16), .ZN(new_n413));
  NAND4_X1  g227(.A1(new_n412), .A2(new_n413), .A3(new_n406), .A4(G125), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n408), .A2(new_n411), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(new_n194), .ZN(new_n416));
  NAND4_X1  g230(.A1(new_n408), .A2(new_n411), .A3(G146), .A4(new_n414), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  XOR2_X1   g232(.A(KEYINPUT24), .B(G110), .Z(new_n419));
  XNOR2_X1  g233(.A(G119), .B(G128), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT73), .ZN(new_n422));
  XNOR2_X1  g236(.A(new_n421), .B(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n405), .A2(new_n418), .A3(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT77), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n405), .A2(KEYINPUT77), .A3(new_n423), .A4(new_n418), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT78), .ZN(new_n429));
  XNOR2_X1  g243(.A(new_n417), .B(new_n429), .ZN(new_n430));
  OAI22_X1  g244(.A1(new_n401), .A2(G110), .B1(new_n420), .B2(new_n419), .ZN(new_n431));
  XNOR2_X1  g245(.A(G125), .B(G140), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n212), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n430), .A2(new_n431), .A3(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n278), .A2(G221), .A3(G234), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n435), .B(KEYINPUT22), .ZN(new_n436));
  XNOR2_X1  g250(.A(new_n436), .B(new_n262), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  AND3_X1   g252(.A1(new_n428), .A2(new_n434), .A3(new_n438), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n438), .B1(new_n428), .B2(new_n434), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(G217), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n442), .B1(G234), .B2(new_n294), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n441), .A2(new_n294), .A3(new_n444), .ZN(new_n445));
  XNOR2_X1  g259(.A(new_n445), .B(KEYINPUT79), .ZN(new_n446));
  AOI21_X1  g260(.A(KEYINPUT25), .B1(new_n441), .B2(new_n294), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT25), .ZN(new_n448));
  NOR4_X1   g262(.A1(new_n439), .A2(new_n440), .A3(new_n448), .A4(G902), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n443), .B1(new_n447), .B2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n446), .A2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n395), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n190), .A2(G128), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n204), .A2(G143), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(G134), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n455), .A2(new_n456), .A3(new_n269), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT99), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(G122), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(G116), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n224), .B1(new_n464), .B2(KEYINPUT14), .ZN(new_n465));
  XNOR2_X1  g279(.A(G116), .B(G122), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n465), .B(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n458), .A2(KEYINPUT99), .A3(new_n459), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n462), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT13), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n470), .B1(new_n204), .B2(G143), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n190), .A2(KEYINPUT13), .A3(G128), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n471), .A2(new_n456), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(G134), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(KEYINPUT98), .ZN(new_n475));
  XNOR2_X1  g289(.A(new_n466), .B(new_n224), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT98), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n473), .A2(new_n477), .A3(G134), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n475), .A2(new_n476), .A3(new_n459), .A4(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n469), .A2(new_n479), .ZN(new_n480));
  NOR3_X1   g294(.A1(new_n311), .A2(new_n442), .A3(G953), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n469), .A2(new_n479), .A3(new_n481), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n483), .A2(KEYINPUT100), .A3(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT100), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n480), .A2(new_n486), .A3(new_n482), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n485), .A2(new_n294), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(KEYINPUT101), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT101), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n485), .A2(new_n490), .A3(new_n294), .A4(new_n487), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(G478), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n493), .A2(KEYINPUT15), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n489), .B1(KEYINPUT15), .B2(new_n493), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(G475), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT91), .ZN(new_n499));
  OAI211_X1 g313(.A(new_n433), .B(new_n499), .C1(new_n194), .C2(new_n432), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n407), .A2(new_n410), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n501), .A2(new_n189), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n432), .A2(new_n194), .ZN(new_n503));
  OAI21_X1  g317(.A(KEYINPUT91), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n500), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(KEYINPUT18), .A2(G131), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n506), .B(KEYINPUT92), .ZN(new_n507));
  INV_X1    g321(.A(G237), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n508), .A2(new_n278), .A3(G214), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(new_n190), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n362), .A2(G143), .A3(G214), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n507), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  AND4_X1   g326(.A1(G143), .A2(new_n508), .A3(new_n278), .A4(G214), .ZN(new_n513));
  AOI21_X1  g327(.A(G143), .B1(new_n362), .B2(G214), .ZN(new_n514));
  OAI21_X1  g328(.A(KEYINPUT89), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT89), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n510), .A2(new_n516), .A3(new_n511), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n506), .ZN(new_n519));
  AOI21_X1  g333(.A(KEYINPUT90), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT90), .ZN(new_n521));
  AOI211_X1 g335(.A(new_n521), .B(new_n506), .C1(new_n515), .C2(new_n517), .ZN(new_n522));
  OAI211_X1 g336(.A(new_n505), .B(new_n512), .C1(new_n520), .C2(new_n522), .ZN(new_n523));
  XOR2_X1   g337(.A(G113), .B(G122), .Z(new_n524));
  XNOR2_X1  g338(.A(new_n524), .B(KEYINPUT95), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n525), .B(G104), .ZN(new_n526));
  OAI21_X1  g340(.A(G131), .B1(new_n513), .B2(new_n514), .ZN(new_n527));
  INV_X1    g341(.A(G131), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n510), .A2(new_n528), .A3(new_n511), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  OAI21_X1  g344(.A(KEYINPUT96), .B1(new_n530), .B2(KEYINPUT17), .ZN(new_n531));
  AND2_X1   g345(.A1(new_n416), .A2(new_n417), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT17), .ZN(new_n533));
  OR2_X1    g347(.A1(new_n527), .A2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT96), .ZN(new_n535));
  NAND4_X1  g349(.A1(new_n527), .A2(new_n529), .A3(new_n535), .A4(new_n533), .ZN(new_n536));
  NAND4_X1  g350(.A1(new_n531), .A2(new_n532), .A3(new_n534), .A4(new_n536), .ZN(new_n537));
  AND3_X1   g351(.A1(new_n523), .A2(new_n526), .A3(new_n537), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n526), .B1(new_n523), .B2(new_n537), .ZN(new_n539));
  OR2_X1    g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n498), .B1(new_n540), .B2(new_n294), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n497), .A2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT97), .ZN(new_n543));
  XNOR2_X1  g357(.A(KEYINPUT93), .B(KEYINPUT19), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n432), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(KEYINPUT94), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n501), .A2(KEYINPUT19), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT94), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n432), .A2(new_n544), .A3(new_n548), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n546), .A2(new_n212), .A3(new_n547), .A4(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n430), .A2(new_n530), .A3(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n526), .B1(new_n523), .B2(new_n551), .ZN(new_n552));
  OAI211_X1 g366(.A(new_n498), .B(new_n294), .C1(new_n538), .C2(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n543), .B1(new_n553), .B2(KEYINPUT20), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n553), .A2(new_n543), .A3(KEYINPUT20), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n553), .A2(KEYINPUT20), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n555), .A2(new_n556), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n542), .A2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  OAI21_X1  g375(.A(G214), .B1(G237), .B2(G902), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  AND3_X1   g377(.A1(new_n254), .A2(G125), .A3(new_n257), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n564), .B1(new_n409), .B2(new_n216), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT7), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n344), .A2(KEYINPUT5), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n567), .B(KEYINPUT88), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n349), .A2(KEYINPUT5), .A3(new_n344), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n568), .A2(G113), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(new_n352), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(new_n228), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n570), .A2(new_n352), .A3(new_n243), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  XOR2_X1   g388(.A(G110), .B(G122), .Z(new_n575));
  XOR2_X1   g389(.A(new_n575), .B(KEYINPUT8), .Z(new_n576));
  AOI22_X1  g390(.A1(new_n565), .A2(new_n566), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n216), .A2(new_n409), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n332), .A2(G125), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(G224), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n581), .A2(G953), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n580), .A2(KEYINPUT7), .A3(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n575), .ZN(new_n585));
  OAI211_X1 g399(.A(new_n573), .B(new_n585), .C1(new_n252), .C2(new_n357), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n578), .A2(new_n582), .A3(new_n579), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n577), .A2(new_n584), .A3(new_n586), .A4(new_n587), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n573), .B1(new_n252), .B2(new_n357), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(new_n575), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n590), .A2(KEYINPUT6), .A3(new_n586), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n580), .A2(new_n583), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(new_n587), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT6), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n589), .A2(new_n594), .A3(new_n575), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n591), .A2(new_n593), .A3(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n588), .A2(new_n596), .A3(new_n294), .ZN(new_n597));
  OAI21_X1  g411(.A(G210), .B1(G237), .B2(G902), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n588), .A2(new_n596), .A3(new_n294), .A4(new_n598), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n563), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  AND2_X1   g416(.A1(new_n278), .A2(G952), .ZN(new_n603));
  NAND2_X1  g417(.A1(G234), .A2(G237), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  XOR2_X1   g420(.A(KEYINPUT21), .B(G898), .Z(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n604), .A2(G902), .A3(G953), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n606), .B1(new_n608), .B2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n602), .A2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  NAND4_X1  g428(.A1(new_n324), .A2(new_n454), .A3(new_n561), .A4(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(G101), .ZN(G3));
  INV_X1    g430(.A(new_n541), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n559), .A2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT33), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n485), .A2(new_n619), .A3(new_n487), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n483), .A2(KEYINPUT33), .A3(new_n484), .ZN(new_n621));
  AND2_X1   g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n622), .A2(G478), .A3(new_n294), .ZN(new_n623));
  AND2_X1   g437(.A1(new_n493), .A2(KEYINPUT102), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n493), .A2(KEYINPUT102), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n488), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n623), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n618), .A2(new_n627), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n613), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n378), .A2(new_n294), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(G472), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n378), .A2(new_n379), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n324), .A2(new_n452), .A3(new_n629), .A4(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(G104), .ZN(new_n636));
  XOR2_X1   g450(.A(KEYINPUT103), .B(KEYINPUT34), .Z(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G6));
  XNOR2_X1  g452(.A(new_n557), .B(KEYINPUT104), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n639), .A2(new_n556), .A3(new_n555), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n541), .B1(new_n495), .B2(new_n496), .ZN(new_n641));
  AND4_X1   g455(.A1(new_n612), .A2(new_n640), .A3(new_n602), .A4(new_n641), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n324), .A2(new_n452), .A3(new_n634), .A4(new_n642), .ZN(new_n643));
  XOR2_X1   g457(.A(KEYINPUT35), .B(G107), .Z(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G9));
  AOI21_X1  g459(.A(new_n613), .B1(new_n315), .B2(new_n323), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n428), .A2(new_n434), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n647), .B1(KEYINPUT36), .B2(new_n437), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n437), .A2(KEYINPUT36), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n428), .A2(new_n434), .A3(new_n649), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n648), .A2(new_n294), .A3(new_n444), .A4(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(KEYINPUT105), .ZN(new_n652));
  OR2_X1    g466(.A1(new_n651), .A2(KEYINPUT105), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n450), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n646), .A2(new_n561), .A3(new_n634), .A4(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(KEYINPUT37), .ZN(new_n656));
  XOR2_X1   g470(.A(new_n656), .B(G110), .Z(G12));
  XOR2_X1   g471(.A(KEYINPUT106), .B(G900), .Z(new_n658));
  AOI21_X1  g472(.A(new_n606), .B1(new_n610), .B2(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  AND2_X1   g474(.A1(new_n640), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(new_n641), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n654), .A2(new_n602), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT32), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n632), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n378), .A2(KEYINPUT32), .A3(new_n379), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n387), .A2(new_n393), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(G472), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n666), .A2(new_n667), .A3(new_n669), .ZN(new_n670));
  NOR3_X1   g484(.A1(new_n310), .A2(KEYINPUT87), .A3(new_n314), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n322), .B1(new_n321), .B2(new_n313), .ZN(new_n672));
  OAI211_X1 g486(.A(new_n664), .B(new_n670), .C1(new_n671), .C2(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G128), .ZN(G30));
  XNOR2_X1  g488(.A(new_n659), .B(KEYINPUT107), .ZN(new_n675));
  XOR2_X1   g489(.A(new_n675), .B(KEYINPUT39), .Z(new_n676));
  AOI21_X1  g490(.A(new_n676), .B1(new_n315), .B2(new_n323), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT40), .ZN(new_n678));
  OR2_X1    g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n600), .A2(new_n601), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(KEYINPUT38), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  AND3_X1   g496(.A1(new_n553), .A2(new_n543), .A3(KEYINPUT20), .ZN(new_n683));
  NOR3_X1   g497(.A1(new_n683), .A2(new_n554), .A3(new_n557), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n497), .B1(new_n684), .B2(new_n541), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n677), .A2(new_n678), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n380), .A2(new_n381), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n386), .A2(new_n376), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n294), .B1(new_n390), .B2(new_n366), .ZN(new_n690));
  OAI21_X1  g504(.A(G472), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  NOR3_X1   g507(.A1(new_n693), .A2(new_n563), .A3(new_n654), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n679), .A2(new_n686), .A3(new_n687), .A4(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G143), .ZN(G45));
  NAND3_X1  g510(.A1(new_n618), .A2(new_n627), .A3(new_n660), .ZN(new_n697));
  INV_X1    g511(.A(new_n602), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(KEYINPUT108), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT108), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n701), .B1(new_n697), .B2(new_n698), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n324), .A2(new_n670), .A3(new_n654), .A4(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G146), .ZN(G48));
  OR2_X1    g519(.A1(new_n308), .A2(new_n187), .ZN(new_n706));
  OAI211_X1 g520(.A(new_n312), .B(new_n706), .C1(new_n319), .C2(new_n320), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n454), .A2(new_n629), .A3(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(KEYINPUT41), .B(G113), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n709), .B(new_n710), .ZN(G15));
  NAND4_X1  g525(.A1(new_n708), .A2(new_n670), .A3(new_n452), .A4(new_n642), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT109), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n712), .B(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(new_n347), .ZN(G18));
  AOI21_X1  g529(.A(new_n560), .B1(new_n688), .B2(new_n669), .ZN(new_n716));
  NOR3_X1   g530(.A1(new_n707), .A2(new_n611), .A3(new_n663), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n716), .A2(new_n717), .A3(KEYINPUT110), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT110), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n670), .A2(new_n561), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n308), .A2(new_n187), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n721), .B1(new_n303), .B2(new_n309), .ZN(new_n722));
  AND2_X1   g536(.A1(new_n654), .A2(new_n602), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n722), .A2(new_n723), .A3(new_n312), .A4(new_n612), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n719), .B1(new_n720), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n718), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G119), .ZN(G21));
  INV_X1    g541(.A(KEYINPUT111), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n685), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n618), .A2(KEYINPUT111), .A3(new_n497), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n729), .A2(new_n602), .A3(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(KEYINPUT112), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT112), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n729), .A2(new_n730), .A3(new_n733), .A4(new_n602), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  OAI211_X1 g549(.A(new_n367), .B(new_n370), .C1(new_n366), .C2(new_n391), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(new_n379), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n631), .A2(new_n737), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n738), .A2(new_n453), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n735), .A2(new_n612), .A3(new_n708), .A4(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G122), .ZN(G24));
  INV_X1    g555(.A(new_n654), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n738), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n743), .A2(new_n699), .A3(new_n708), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G125), .ZN(G27));
  OAI21_X1  g559(.A(KEYINPUT113), .B1(new_n380), .B2(new_n381), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT113), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n666), .A2(new_n747), .A3(new_n667), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n746), .A2(new_n748), .A3(new_n669), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n680), .A2(new_n563), .ZN(new_n750));
  INV_X1    g564(.A(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(new_n312), .ZN(new_n752));
  NOR4_X1   g566(.A1(new_n310), .A2(new_n751), .A3(new_n752), .A4(new_n697), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n749), .A2(new_n753), .A3(new_n452), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(KEYINPUT42), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n670), .A2(new_n452), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n321), .A2(new_n312), .A3(new_n750), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n697), .A2(KEYINPUT42), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n755), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(new_n528), .ZN(G33));
  NOR3_X1   g576(.A1(new_n756), .A2(new_n757), .A3(new_n662), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(new_n269), .ZN(G36));
  XNOR2_X1  g578(.A(new_n293), .B(KEYINPUT45), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(G469), .ZN(new_n766));
  NAND2_X1  g580(.A1(G469), .A2(G902), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT46), .ZN(new_n769));
  AOI22_X1  g583(.A1(new_n768), .A2(new_n769), .B1(new_n303), .B2(new_n309), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n770), .B1(new_n769), .B2(new_n768), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(new_n312), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n772), .A2(new_n676), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n559), .A2(new_n617), .A3(new_n627), .ZN(new_n774));
  XOR2_X1   g588(.A(new_n774), .B(KEYINPUT43), .Z(new_n775));
  NAND3_X1  g589(.A1(new_n775), .A2(new_n633), .A3(new_n654), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT44), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n778), .A2(new_n751), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n776), .A2(new_n777), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n773), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G137), .ZN(G39));
  NAND2_X1  g596(.A1(new_n772), .A2(KEYINPUT47), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n670), .A2(new_n452), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT47), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n771), .A2(new_n785), .A3(new_n312), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n751), .A2(new_n697), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n783), .A2(new_n784), .A3(new_n786), .A4(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT114), .ZN(new_n789));
  OR2_X1    g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n788), .A2(new_n789), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G140), .ZN(G42));
  INV_X1    g607(.A(KEYINPUT51), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n722), .A2(new_n314), .ZN(new_n795));
  XOR2_X1   g609(.A(new_n795), .B(KEYINPUT118), .Z(new_n796));
  INV_X1    g610(.A(new_n786), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n785), .B1(new_n771), .B2(new_n312), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n796), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n775), .A2(new_n606), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n800), .A2(new_n739), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n801), .A2(new_n751), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n799), .A2(new_n802), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n801), .A2(new_n707), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n804), .A2(new_n563), .A3(new_n682), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT50), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n804), .A2(KEYINPUT50), .A3(new_n563), .A4(new_n682), .ZN(new_n808));
  AND3_X1   g622(.A1(new_n807), .A2(KEYINPUT119), .A3(new_n808), .ZN(new_n809));
  AOI21_X1  g623(.A(KEYINPUT119), .B1(new_n807), .B2(new_n808), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n803), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n693), .A2(new_n708), .A3(new_n750), .ZN(new_n812));
  NOR3_X1   g626(.A1(new_n812), .A2(new_n453), .A3(new_n605), .ZN(new_n813));
  INV_X1    g627(.A(new_n627), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n813), .A2(new_n559), .A3(new_n617), .A4(new_n814), .ZN(new_n815));
  AND3_X1   g629(.A1(new_n800), .A2(new_n708), .A3(new_n750), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(new_n743), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n794), .B1(new_n811), .B2(new_n818), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n795), .B1(new_n797), .B2(new_n798), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT120), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  OAI211_X1 g636(.A(KEYINPUT120), .B(new_n795), .C1(new_n797), .C2(new_n798), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n822), .A2(new_n802), .A3(new_n823), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n818), .B1(new_n807), .B2(new_n808), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n824), .A2(KEYINPUT51), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n804), .A2(new_n602), .ZN(new_n827));
  AND2_X1   g641(.A1(new_n749), .A2(new_n452), .ZN(new_n828));
  AND2_X1   g642(.A1(new_n816), .A2(new_n828), .ZN(new_n829));
  OAI211_X1 g643(.A(new_n603), .B(new_n827), .C1(new_n829), .C2(KEYINPUT48), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n830), .B1(KEYINPUT48), .B2(new_n829), .ZN(new_n831));
  AND3_X1   g645(.A1(new_n819), .A2(new_n826), .A3(new_n831), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n712), .B(KEYINPUT109), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n833), .A2(new_n615), .A3(new_n709), .A4(new_n740), .ZN(new_n834));
  INV_X1    g648(.A(new_n662), .ZN(new_n835));
  AOI22_X1  g649(.A1(new_n758), .A2(new_n835), .B1(new_n743), .B2(new_n753), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n395), .B1(new_n315), .B2(new_n323), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n661), .A2(new_n542), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n837), .A2(new_n654), .A3(new_n750), .A4(new_n838), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n836), .A2(new_n755), .A3(new_n839), .A4(new_n760), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n602), .A2(new_n559), .A3(new_n612), .A4(new_n641), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT116), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n841), .B(new_n842), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n324), .A2(new_n452), .A3(new_n634), .A4(new_n843), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n655), .A2(new_n726), .A3(new_n635), .A4(new_n844), .ZN(new_n845));
  NOR3_X1   g659(.A1(new_n834), .A2(new_n840), .A3(new_n845), .ZN(new_n846));
  AND3_X1   g660(.A1(new_n704), .A2(new_n673), .A3(new_n744), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n310), .A2(new_n752), .A3(new_n659), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n735), .A2(new_n742), .A3(new_n692), .A4(new_n848), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n847), .A2(KEYINPUT52), .A3(new_n849), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n704), .A2(new_n849), .A3(new_n673), .A4(new_n744), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT52), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT53), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n846), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  AND4_X1   g670(.A1(new_n755), .A2(new_n836), .A3(new_n839), .A4(new_n760), .ZN(new_n857));
  AND4_X1   g671(.A1(new_n635), .A2(new_n655), .A3(new_n726), .A4(new_n844), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n615), .A2(new_n740), .A3(new_n709), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n859), .A2(new_n714), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n857), .A2(new_n858), .A3(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT117), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n853), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n863), .A2(new_n850), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n851), .A2(KEYINPUT117), .A3(new_n852), .ZN(new_n865));
  INV_X1    g679(.A(new_n865), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n861), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n856), .B1(new_n867), .B2(new_n855), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT54), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n846), .A2(new_n854), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n871), .A2(KEYINPUT53), .ZN(new_n872));
  AOI21_X1  g686(.A(KEYINPUT117), .B1(new_n851), .B2(new_n852), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n851), .A2(new_n852), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n846), .B1(new_n875), .B2(new_n865), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n872), .B1(KEYINPUT53), .B2(new_n876), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n832), .B(new_n870), .C1(new_n869), .C2(new_n877), .ZN(new_n878));
  NOR4_X1   g692(.A1(new_n812), .A2(new_n453), .A3(new_n605), .A4(new_n628), .ZN(new_n879));
  OAI22_X1  g693(.A1(new_n878), .A2(new_n879), .B1(G952), .B2(G953), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n452), .A2(new_n313), .A3(new_n562), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT115), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n682), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(new_n722), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n883), .B1(KEYINPUT49), .B2(new_n884), .ZN(new_n885));
  OR2_X1    g699(.A1(new_n884), .A2(KEYINPUT49), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n774), .B1(new_n881), .B2(new_n882), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n885), .A2(new_n693), .A3(new_n886), .A4(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n880), .A2(new_n888), .ZN(G75));
  NAND2_X1  g703(.A1(new_n876), .A2(KEYINPUT53), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n890), .A2(G210), .A3(G902), .A4(new_n856), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT56), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n891), .A2(KEYINPUT122), .A3(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT121), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n891), .A2(new_n894), .A3(new_n892), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n591), .A2(new_n595), .ZN(new_n896));
  XOR2_X1   g710(.A(new_n896), .B(new_n593), .Z(new_n897));
  XNOR2_X1  g711(.A(new_n897), .B(KEYINPUT55), .ZN(new_n898));
  AOI22_X1  g712(.A1(KEYINPUT121), .A2(new_n893), .B1(new_n895), .B2(new_n898), .ZN(new_n899));
  AND3_X1   g713(.A1(new_n893), .A2(KEYINPUT121), .A3(new_n898), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n278), .A2(G952), .ZN(new_n901));
  NOR3_X1   g715(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(G51));
  NOR3_X1   g716(.A1(new_n868), .A2(new_n294), .A3(new_n766), .ZN(new_n903));
  XOR2_X1   g717(.A(new_n767), .B(KEYINPUT57), .Z(new_n904));
  OAI211_X1 g718(.A(KEYINPUT54), .B(new_n856), .C1(new_n867), .C2(new_n855), .ZN(new_n905));
  INV_X1    g719(.A(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(KEYINPUT54), .B1(new_n890), .B2(new_n856), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n904), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n903), .B1(new_n908), .B2(new_n318), .ZN(new_n909));
  OAI21_X1  g723(.A(KEYINPUT123), .B1(new_n909), .B2(new_n901), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT123), .ZN(new_n911));
  INV_X1    g725(.A(new_n901), .ZN(new_n912));
  INV_X1    g726(.A(new_n318), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n870), .A2(new_n905), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n913), .B1(new_n914), .B2(new_n904), .ZN(new_n915));
  OAI211_X1 g729(.A(new_n911), .B(new_n912), .C1(new_n915), .C2(new_n903), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n910), .A2(new_n916), .ZN(G54));
  INV_X1    g731(.A(new_n868), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n918), .A2(KEYINPUT58), .A3(G902), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n538), .A2(new_n552), .ZN(new_n920));
  OR3_X1    g734(.A1(new_n919), .A2(new_n498), .A3(new_n920), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n920), .B1(new_n919), .B2(new_n498), .ZN(new_n922));
  AND3_X1   g736(.A1(new_n921), .A2(new_n912), .A3(new_n922), .ZN(G60));
  OAI21_X1  g737(.A(new_n870), .B1(new_n877), .B2(new_n869), .ZN(new_n924));
  NAND2_X1  g738(.A1(G478), .A2(G902), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n925), .B(KEYINPUT59), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n622), .B1(new_n924), .B2(new_n926), .ZN(new_n927));
  AND3_X1   g741(.A1(new_n914), .A2(new_n622), .A3(new_n926), .ZN(new_n928));
  NOR3_X1   g742(.A1(new_n927), .A2(new_n928), .A3(new_n901), .ZN(G63));
  NAND2_X1  g743(.A1(G217), .A2(G902), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n930), .B(KEYINPUT60), .Z(new_n931));
  NAND2_X1  g745(.A1(new_n918), .A2(new_n931), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n932), .B1(new_n439), .B2(new_n440), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n648), .A2(new_n650), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n934), .B(KEYINPUT124), .Z(new_n935));
  NAND3_X1  g749(.A1(new_n918), .A2(new_n931), .A3(new_n935), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n933), .A2(new_n912), .A3(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT61), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n933), .A2(KEYINPUT61), .A3(new_n912), .A4(new_n936), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n940), .ZN(G66));
  OAI21_X1  g755(.A(G953), .B1(new_n608), .B2(new_n581), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n858), .A2(new_n860), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(KEYINPUT125), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n942), .B1(new_n944), .B2(G953), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n896), .B1(G898), .B2(new_n278), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n946), .B(KEYINPUT126), .Z(new_n947));
  XNOR2_X1  g761(.A(new_n945), .B(new_n947), .ZN(G69));
  NAND3_X1  g762(.A1(new_n546), .A2(new_n547), .A3(new_n549), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n368), .B(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n695), .A2(new_n847), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n951), .B(KEYINPUT62), .ZN(new_n952));
  INV_X1    g766(.A(new_n781), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n677), .A2(new_n454), .A3(new_n560), .ZN(new_n955));
  AOI211_X1 g769(.A(new_n751), .B(new_n955), .C1(new_n618), .C2(new_n814), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n956), .B1(new_n790), .B2(new_n791), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n954), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n950), .B1(new_n958), .B2(new_n278), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n761), .B1(new_n790), .B2(new_n791), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n773), .A2(new_n735), .A3(new_n828), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n781), .A2(new_n961), .A3(new_n847), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n962), .A2(new_n763), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n960), .A2(new_n963), .A3(new_n278), .ZN(new_n964));
  AND2_X1   g778(.A1(new_n964), .A2(new_n950), .ZN(new_n965));
  NAND2_X1  g779(.A1(G900), .A2(G953), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n959), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n278), .B1(G227), .B2(G900), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n964), .A2(new_n950), .A3(new_n966), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n968), .B1(new_n969), .B2(KEYINPUT127), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n967), .B(new_n970), .ZN(G72));
  NAND2_X1  g785(.A1(G472), .A2(G902), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n972), .B(KEYINPUT63), .Z(new_n973));
  INV_X1    g787(.A(new_n973), .ZN(new_n974));
  AND2_X1   g788(.A1(new_n960), .A2(new_n963), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n974), .B1(new_n975), .B2(new_n944), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n386), .A2(new_n376), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n912), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n954), .A2(new_n957), .A3(new_n944), .ZN(new_n979));
  AOI211_X1 g793(.A(new_n386), .B(new_n376), .C1(new_n979), .C2(new_n973), .ZN(new_n980));
  INV_X1    g794(.A(new_n977), .ZN(new_n981));
  NOR4_X1   g795(.A1(new_n877), .A2(new_n689), .A3(new_n974), .A4(new_n981), .ZN(new_n982));
  NOR3_X1   g796(.A1(new_n978), .A2(new_n980), .A3(new_n982), .ZN(G57));
endmodule


