

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769;

  NOR2_X1 U384 ( .A1(n743), .A2(n424), .ZN(n412) );
  XNOR2_X1 U385 ( .A(n598), .B(n597), .ZN(n616) );
  AND2_X1 U386 ( .A1(n453), .A2(n451), .ZN(n450) );
  NAND2_X1 U387 ( .A1(n386), .A2(n385), .ZN(n411) );
  XNOR2_X1 U388 ( .A(n756), .B(G146), .ZN(n524) );
  XNOR2_X1 U389 ( .A(n532), .B(n403), .ZN(n494) );
  AND2_X2 U390 ( .A1(n559), .A2(n365), .ZN(n455) );
  INV_X1 U391 ( .A(n618), .ZN(n700) );
  NOR2_X2 U392 ( .A1(n571), .A2(n572), .ZN(n378) );
  NOR2_X2 U393 ( .A1(n766), .A2(n665), .ZN(n604) );
  XOR2_X2 U394 ( .A(G101), .B(KEYINPUT4), .Z(n522) );
  XNOR2_X2 U395 ( .A(n555), .B(KEYINPUT105), .ZN(n676) );
  XNOR2_X2 U396 ( .A(n607), .B(n606), .ZN(n720) );
  BUF_X1 U397 ( .A(n727), .Z(n736) );
  AND2_X1 U398 ( .A1(n634), .A2(n684), .ZN(n636) );
  XNOR2_X1 U399 ( .A(n430), .B(n581), .ZN(n429) );
  NOR2_X2 U400 ( .A1(n700), .A2(n699), .ZN(n620) );
  XNOR2_X1 U401 ( .A(n387), .B(G146), .ZN(n531) );
  NAND2_X1 U402 ( .A1(n429), .A2(n369), .ZN(n424) );
  OR2_X1 U403 ( .A1(n563), .A2(n564), .ZN(n377) );
  XNOR2_X1 U404 ( .A(n378), .B(KEYINPUT39), .ZN(n582) );
  OR2_X1 U405 ( .A1(n624), .A2(n565), .ZN(n425) );
  AND2_X1 U406 ( .A1(n376), .A2(n602), .ZN(n558) );
  XNOR2_X1 U407 ( .A(n556), .B(n426), .ZN(n694) );
  NAND2_X1 U408 ( .A1(n676), .A2(n673), .ZN(n556) );
  XNOR2_X1 U409 ( .A(n494), .B(n482), .ZN(n756) );
  XNOR2_X1 U410 ( .A(n498), .B(n497), .ZN(n754) );
  XNOR2_X1 U411 ( .A(n531), .B(n420), .ZN(n498) );
  XNOR2_X1 U412 ( .A(G137), .B(G140), .ZN(n497) );
  INV_X2 U413 ( .A(G128), .ZN(n404) );
  XNOR2_X1 U414 ( .A(n486), .B(n485), .ZN(n554) );
  INV_X1 U415 ( .A(KEYINPUT106), .ZN(n426) );
  INV_X1 U416 ( .A(G125), .ZN(n387) );
  XNOR2_X1 U417 ( .A(KEYINPUT45), .B(KEYINPUT85), .ZN(n462) );
  XNOR2_X1 U418 ( .A(G104), .B(G110), .ZN(n748) );
  INV_X1 U419 ( .A(G134), .ZN(n403) );
  XNOR2_X1 U420 ( .A(KEYINPUT8), .B(KEYINPUT67), .ZN(n487) );
  XNOR2_X1 U421 ( .A(n509), .B(n422), .ZN(n421) );
  OR2_X1 U422 ( .A1(n738), .A2(G902), .ZN(n423) );
  XNOR2_X1 U423 ( .A(n508), .B(KEYINPUT97), .ZN(n422) );
  XNOR2_X1 U424 ( .A(n694), .B(KEYINPUT80), .ZN(n624) );
  NAND2_X1 U425 ( .A1(n702), .A2(n365), .ZN(n699) );
  XOR2_X1 U426 ( .A(G902), .B(KEYINPUT15), .Z(n631) );
  XNOR2_X1 U427 ( .A(G128), .B(KEYINPUT95), .ZN(n501) );
  NOR2_X1 U428 ( .A1(n455), .A2(KEYINPUT111), .ZN(n454) );
  OR2_X1 U429 ( .A1(n602), .A2(n448), .ZN(n447) );
  AND2_X1 U430 ( .A1(n690), .A2(n448), .ZN(n445) );
  OR2_X1 U431 ( .A1(n690), .A2(n448), .ZN(n446) );
  AND2_X1 U432 ( .A1(n455), .A2(KEYINPUT111), .ZN(n452) );
  XNOR2_X1 U433 ( .A(n396), .B(n561), .ZN(n594) );
  XNOR2_X1 U434 ( .A(n527), .B(G472), .ZN(n547) );
  NOR2_X1 U435 ( .A1(G902), .A2(n653), .ZN(n527) );
  XNOR2_X1 U436 ( .A(n490), .B(KEYINPUT7), .ZN(n391) );
  XOR2_X1 U437 ( .A(KEYINPUT103), .B(KEYINPUT9), .Z(n490) );
  INV_X1 U438 ( .A(KEYINPUT64), .ZN(n637) );
  XNOR2_X1 U439 ( .A(n398), .B(n530), .ZN(n534) );
  INV_X1 U440 ( .A(KEYINPUT82), .ZN(n402) );
  XNOR2_X1 U441 ( .A(n392), .B(KEYINPUT114), .ZN(n577) );
  XNOR2_X1 U442 ( .A(n547), .B(KEYINPUT109), .ZN(n602) );
  XNOR2_X1 U443 ( .A(n596), .B(KEYINPUT72), .ZN(n597) );
  NAND2_X1 U444 ( .A1(n381), .A2(n371), .ZN(n598) );
  XNOR2_X1 U445 ( .A(n496), .B(n495), .ZN(n575) );
  NAND2_X1 U446 ( .A1(n616), .A2(n617), .ZN(n418) );
  XNOR2_X1 U447 ( .A(G119), .B(G110), .ZN(n504) );
  XNOR2_X1 U448 ( .A(n425), .B(KEYINPUT73), .ZN(n566) );
  NOR2_X1 U449 ( .A1(G953), .A2(G237), .ZN(n525) );
  NAND2_X1 U450 ( .A1(G234), .A2(G237), .ZN(n510) );
  XNOR2_X1 U451 ( .A(n379), .B(KEYINPUT20), .ZN(n515) );
  NAND2_X1 U452 ( .A1(n635), .A2(G234), .ZN(n379) );
  XNOR2_X1 U453 ( .A(n522), .B(n394), .ZN(n393) );
  INV_X1 U454 ( .A(G137), .ZN(n394) );
  XNOR2_X1 U455 ( .A(n580), .B(KEYINPUT86), .ZN(n581) );
  XNOR2_X1 U456 ( .A(n518), .B(n414), .ZN(n537) );
  XNOR2_X1 U457 ( .A(n415), .B(G119), .ZN(n414) );
  INV_X1 U458 ( .A(G113), .ZN(n415) );
  XOR2_X1 U459 ( .A(G104), .B(G122), .Z(n477) );
  XNOR2_X1 U460 ( .A(G143), .B(G113), .ZN(n476) );
  INV_X1 U461 ( .A(KEYINPUT10), .ZN(n420) );
  XNOR2_X1 U462 ( .A(G140), .B(KEYINPUT12), .ZN(n478) );
  XOR2_X1 U463 ( .A(KEYINPUT11), .B(KEYINPUT102), .Z(n479) );
  NAND2_X1 U464 ( .A1(n635), .A2(n461), .ZN(n458) );
  XNOR2_X1 U465 ( .A(n529), .B(KEYINPUT17), .ZN(n398) );
  INV_X1 U466 ( .A(n557), .ZN(n376) );
  NOR2_X1 U467 ( .A1(n397), .A2(n609), .ZN(n409) );
  XNOR2_X1 U468 ( .A(n541), .B(n540), .ZN(n542) );
  INV_X1 U469 ( .A(KEYINPUT93), .ZN(n540) );
  XNOR2_X1 U470 ( .A(n413), .B(n375), .ZN(n622) );
  NOR2_X1 U471 ( .A1(n594), .A2(n593), .ZN(n413) );
  INV_X1 U472 ( .A(KEYINPUT91), .ZN(n465) );
  XNOR2_X1 U473 ( .A(n384), .B(n524), .ZN(n653) );
  XOR2_X1 U474 ( .A(n523), .B(n456), .Z(n384) );
  XNOR2_X1 U475 ( .A(n537), .B(n526), .ZN(n456) );
  XNOR2_X1 U476 ( .A(n521), .B(n393), .ZN(n523) );
  BUF_X1 U477 ( .A(n634), .Z(n743) );
  XOR2_X1 U478 ( .A(KEYINPUT23), .B(KEYINPUT96), .Z(n502) );
  INV_X1 U479 ( .A(KEYINPUT24), .ZN(n500) );
  INV_X1 U480 ( .A(n690), .ZN(n389) );
  XNOR2_X1 U481 ( .A(n419), .B(KEYINPUT35), .ZN(n612) );
  NAND2_X1 U482 ( .A1(n406), .A2(n405), .ZN(n419) );
  NAND2_X1 U483 ( .A1(n410), .A2(n409), .ZN(n405) );
  AND2_X1 U484 ( .A1(n407), .A2(n372), .ZN(n406) );
  NOR2_X1 U485 ( .A1(n442), .A2(n441), .ZN(n440) );
  NOR2_X1 U486 ( .A1(n577), .A2(n594), .ZN(n567) );
  INV_X1 U487 ( .A(n547), .ZN(n706) );
  BUF_X1 U488 ( .A(n622), .Z(n397) );
  XNOR2_X1 U489 ( .A(n536), .B(n391), .ZN(n491) );
  XNOR2_X1 U490 ( .A(n524), .B(n475), .ZN(n729) );
  XNOR2_X1 U491 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U492 ( .A(n645), .B(n468), .ZN(n648) );
  XOR2_X1 U493 ( .A(KEYINPUT92), .B(n641), .Z(n726) );
  INV_X1 U494 ( .A(KEYINPUT84), .ZN(n438) );
  NOR2_X1 U495 ( .A1(n435), .A2(G953), .ZN(n434) );
  NOR2_X1 U496 ( .A1(n363), .A2(n724), .ZN(n435) );
  NOR2_X1 U497 ( .A1(n719), .A2(n577), .ZN(n578) );
  INV_X1 U498 ( .A(n612), .ZN(n765) );
  XNOR2_X1 U499 ( .A(n467), .B(n466), .ZN(n766) );
  XNOR2_X1 U500 ( .A(KEYINPUT32), .B(KEYINPUT77), .ZN(n466) );
  XNOR2_X1 U501 ( .A(n383), .B(KEYINPUT31), .ZN(n675) );
  NOR2_X1 U502 ( .A1(n710), .A2(n397), .ZN(n383) );
  NOR2_X1 U503 ( .A1(n602), .A2(n601), .ZN(n665) );
  NOR2_X1 U504 ( .A1(n575), .A2(n554), .ZN(n555) );
  XNOR2_X1 U505 ( .A(n418), .B(KEYINPUT87), .ZN(n417) );
  XNOR2_X1 U506 ( .A(n737), .B(n738), .ZN(n401) );
  XOR2_X1 U507 ( .A(KEYINPUT123), .B(n723), .Z(n363) );
  AND2_X1 U508 ( .A1(n363), .A2(n724), .ZN(n364) );
  XOR2_X1 U509 ( .A(n516), .B(KEYINPUT21), .Z(n365) );
  XOR2_X1 U510 ( .A(n484), .B(n481), .Z(n366) );
  XNOR2_X1 U511 ( .A(n559), .B(KEYINPUT112), .ZN(n367) );
  AND2_X1 U512 ( .A1(n636), .A2(n461), .ZN(n368) );
  AND2_X1 U513 ( .A1(n588), .A2(n682), .ZN(n369) );
  INV_X1 U514 ( .A(n702), .ZN(n449) );
  NOR2_X1 U515 ( .A1(n557), .A2(n389), .ZN(n370) );
  AND2_X1 U516 ( .A1(n595), .A2(n365), .ZN(n371) );
  AND2_X1 U517 ( .A1(n408), .A2(n610), .ZN(n372) );
  AND2_X1 U518 ( .A1(n702), .A2(n455), .ZN(n373) );
  XOR2_X1 U519 ( .A(KEYINPUT113), .B(KEYINPUT28), .Z(n374) );
  XOR2_X1 U520 ( .A(n465), .B(KEYINPUT0), .Z(n375) );
  INV_X1 U521 ( .A(KEYINPUT111), .ZN(n549) );
  INV_X1 U522 ( .A(G953), .ZN(n761) );
  XNOR2_X1 U523 ( .A(n382), .B(n462), .ZN(n634) );
  NAND2_X1 U524 ( .A1(n615), .A2(n614), .ZN(n464) );
  NOR2_X1 U525 ( .A1(n368), .A2(n400), .ZN(n457) );
  NAND2_X1 U526 ( .A1(n377), .A2(n570), .ZN(n390) );
  NOR2_X1 U527 ( .A1(n454), .A2(n548), .ZN(n453) );
  XNOR2_X1 U528 ( .A(n380), .B(n535), .ZN(n395) );
  XNOR2_X1 U529 ( .A(n533), .B(n534), .ZN(n380) );
  NAND2_X1 U530 ( .A1(n457), .A2(n460), .ZN(n459) );
  NAND2_X1 U531 ( .A1(n463), .A2(n464), .ZN(n382) );
  NAND2_X1 U532 ( .A1(n611), .A2(n765), .ZN(n615) );
  INV_X1 U533 ( .A(n622), .ZN(n381) );
  INV_X1 U534 ( .A(G902), .ZN(n385) );
  INV_X1 U535 ( .A(n729), .ZN(n386) );
  NAND2_X1 U536 ( .A1(n388), .A2(n367), .ZN(n392) );
  XNOR2_X1 U537 ( .A(n558), .B(n374), .ZN(n388) );
  NAND2_X1 U538 ( .A1(n605), .A2(n370), .ZN(n528) );
  XNOR2_X2 U539 ( .A(n411), .B(G469), .ZN(n559) );
  NOR2_X1 U540 ( .A1(n390), .A2(n569), .ZN(n399) );
  XNOR2_X1 U541 ( .A(n395), .B(n746), .ZN(n645) );
  NAND2_X1 U542 ( .A1(n560), .A2(n690), .ZN(n396) );
  NAND2_X1 U543 ( .A1(n399), .A2(n431), .ZN(n430) );
  NAND2_X1 U544 ( .A1(n633), .A2(n458), .ZN(n400) );
  NOR2_X1 U545 ( .A1(n401), .A2(n739), .ZN(G66) );
  XNOR2_X1 U546 ( .A(n636), .B(n402), .ZN(n686) );
  XNOR2_X2 U547 ( .A(n404), .B(G143), .ZN(n532) );
  NAND2_X1 U548 ( .A1(n720), .A2(n609), .ZN(n407) );
  NAND2_X1 U549 ( .A1(n397), .A2(n609), .ZN(n408) );
  INV_X1 U550 ( .A(n720), .ZN(n410) );
  XNOR2_X2 U551 ( .A(n559), .B(KEYINPUT1), .ZN(n618) );
  NAND2_X1 U552 ( .A1(n412), .A2(n630), .ZN(n460) );
  AND2_X1 U553 ( .A1(n412), .A2(KEYINPUT2), .ZN(n687) );
  NAND2_X1 U554 ( .A1(n417), .A2(n416), .ZN(n619) );
  NOR2_X1 U555 ( .A1(n618), .A2(n449), .ZN(n416) );
  XNOR2_X2 U556 ( .A(n423), .B(n421), .ZN(n702) );
  NAND2_X1 U557 ( .A1(n424), .A2(n632), .ZN(n633) );
  NAND2_X1 U558 ( .A1(n424), .A2(n684), .ZN(n685) );
  XNOR2_X1 U559 ( .A(n424), .B(n760), .ZN(n762) );
  XNOR2_X1 U560 ( .A(n427), .B(n366), .ZN(n638) );
  XNOR2_X1 U561 ( .A(n428), .B(n498), .ZN(n427) );
  XNOR2_X1 U562 ( .A(n483), .B(n480), .ZN(n428) );
  NOR2_X1 U563 ( .A1(n769), .A2(n628), .ZN(n463) );
  XNOR2_X1 U564 ( .A(n507), .B(n506), .ZN(n738) );
  XNOR2_X1 U565 ( .A(n579), .B(KEYINPUT46), .ZN(n431) );
  XNOR2_X1 U566 ( .A(n689), .B(n438), .ZN(n437) );
  NAND2_X1 U567 ( .A1(n437), .A2(n364), .ZN(n432) );
  NOR2_X1 U568 ( .A1(n437), .A2(n724), .ZN(n436) );
  NAND2_X1 U569 ( .A1(n432), .A2(n434), .ZN(n433) );
  NOR2_X1 U570 ( .A1(n436), .A2(n433), .ZN(n725) );
  INV_X1 U571 ( .A(G953), .ZN(n439) );
  NAND2_X1 U572 ( .A1(n440), .A2(n450), .ZN(n571) );
  NAND2_X1 U573 ( .A1(n443), .A2(n446), .ZN(n441) );
  NAND2_X1 U574 ( .A1(n447), .A2(n444), .ZN(n442) );
  NAND2_X1 U575 ( .A1(n449), .A2(n549), .ZN(n443) );
  NAND2_X1 U576 ( .A1(n602), .A2(n445), .ZN(n444) );
  INV_X1 U577 ( .A(KEYINPUT30), .ZN(n448) );
  NAND2_X1 U578 ( .A1(n452), .A2(n702), .ZN(n451) );
  XNOR2_X2 U579 ( .A(n459), .B(n637), .ZN(n727) );
  INV_X1 U580 ( .A(KEYINPUT83), .ZN(n461) );
  NAND2_X1 U581 ( .A1(n616), .A2(n599), .ZN(n467) );
  XNOR2_X1 U582 ( .A(n731), .B(n730), .ZN(n732) );
  BUF_X1 U583 ( .A(n560), .Z(n585) );
  XOR2_X1 U584 ( .A(n647), .B(n646), .Z(n468) );
  AND2_X1 U585 ( .A1(G221), .A2(n499), .ZN(n469) );
  INV_X1 U586 ( .A(KEYINPUT33), .ZN(n606) );
  INV_X1 U587 ( .A(KEYINPUT48), .ZN(n580) );
  INV_X1 U588 ( .A(n680), .ZN(n588) );
  XNOR2_X1 U589 ( .A(n501), .B(n500), .ZN(n503) );
  XNOR2_X1 U590 ( .A(n503), .B(n502), .ZN(n505) );
  XNOR2_X1 U591 ( .A(n543), .B(n542), .ZN(n560) );
  XNOR2_X1 U592 ( .A(n754), .B(n469), .ZN(n507) );
  XNOR2_X1 U593 ( .A(n729), .B(n728), .ZN(n730) );
  XNOR2_X1 U594 ( .A(KEYINPUT125), .B(KEYINPUT60), .ZN(n643) );
  XOR2_X1 U595 ( .A(KEYINPUT68), .B(G131), .Z(n482) );
  XNOR2_X1 U596 ( .A(n522), .B(KEYINPUT70), .ZN(n470) );
  XNOR2_X1 U597 ( .A(n470), .B(n748), .ZN(n535) );
  INV_X1 U598 ( .A(n535), .ZN(n474) );
  XNOR2_X1 U599 ( .A(G107), .B(n497), .ZN(n472) );
  NAND2_X1 U600 ( .A1(G227), .A2(n761), .ZN(n471) );
  XNOR2_X1 U601 ( .A(n472), .B(n471), .ZN(n473) );
  XOR2_X1 U602 ( .A(KEYINPUT36), .B(KEYINPUT89), .Z(n545) );
  XNOR2_X1 U603 ( .A(n477), .B(n476), .ZN(n484) );
  XNOR2_X1 U604 ( .A(n479), .B(n478), .ZN(n481) );
  NAND2_X1 U605 ( .A1(G214), .A2(n525), .ZN(n480) );
  XNOR2_X1 U606 ( .A(n482), .B(KEYINPUT101), .ZN(n483) );
  NOR2_X1 U607 ( .A1(G902), .A2(n638), .ZN(n486) );
  XNOR2_X1 U608 ( .A(KEYINPUT13), .B(G475), .ZN(n485) );
  NAND2_X1 U609 ( .A1(n761), .A2(G234), .ZN(n488) );
  XNOR2_X1 U610 ( .A(n488), .B(n487), .ZN(n499) );
  NAND2_X1 U611 ( .A1(n499), .A2(G217), .ZN(n492) );
  XNOR2_X1 U612 ( .A(G116), .B(G122), .ZN(n489) );
  XNOR2_X1 U613 ( .A(n489), .B(G107), .ZN(n536) );
  XNOR2_X1 U614 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U615 ( .A(n494), .B(n493), .ZN(n734) );
  NOR2_X1 U616 ( .A1(G902), .A2(n734), .ZN(n496) );
  XNOR2_X1 U617 ( .A(KEYINPUT104), .B(G478), .ZN(n495) );
  NAND2_X1 U618 ( .A1(n554), .A2(n575), .ZN(n673) );
  INV_X1 U619 ( .A(n631), .ZN(n635) );
  NAND2_X1 U620 ( .A1(n515), .A2(G217), .ZN(n509) );
  XNOR2_X1 U621 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U622 ( .A(KEYINPUT25), .B(KEYINPUT98), .ZN(n508) );
  XNOR2_X1 U623 ( .A(n510), .B(KEYINPUT14), .ZN(n511) );
  NAND2_X1 U624 ( .A1(G952), .A2(n511), .ZN(n718) );
  NOR2_X1 U625 ( .A1(G953), .A2(n718), .ZN(n592) );
  NAND2_X1 U626 ( .A1(G902), .A2(n511), .ZN(n590) );
  NOR2_X1 U627 ( .A1(G900), .A2(n590), .ZN(n512) );
  NAND2_X1 U628 ( .A1(G953), .A2(n512), .ZN(n513) );
  XOR2_X1 U629 ( .A(KEYINPUT110), .B(n513), .Z(n514) );
  NOR2_X1 U630 ( .A1(n592), .A2(n514), .ZN(n548) );
  NOR2_X1 U631 ( .A1(n702), .A2(n548), .ZN(n517) );
  NAND2_X1 U632 ( .A1(n515), .A2(G221), .ZN(n516) );
  NAND2_X1 U633 ( .A1(n517), .A2(n365), .ZN(n557) );
  XNOR2_X1 U634 ( .A(KEYINPUT3), .B(KEYINPUT69), .ZN(n518) );
  XOR2_X1 U635 ( .A(KEYINPUT99), .B(KEYINPUT5), .Z(n520) );
  XNOR2_X1 U636 ( .A(G116), .B(KEYINPUT74), .ZN(n519) );
  XNOR2_X1 U637 ( .A(n520), .B(n519), .ZN(n521) );
  NAND2_X1 U638 ( .A1(n525), .A2(G210), .ZN(n526) );
  XOR2_X1 U639 ( .A(n706), .B(KEYINPUT6), .Z(n605) );
  INV_X1 U640 ( .A(n605), .ZN(n617) );
  OR2_X1 U641 ( .A1(G237), .A2(G902), .ZN(n539) );
  NAND2_X1 U642 ( .A1(G214), .A2(n539), .ZN(n690) );
  NOR2_X1 U643 ( .A1(n673), .A2(n528), .ZN(n583) );
  XOR2_X1 U644 ( .A(KEYINPUT75), .B(KEYINPUT18), .Z(n530) );
  NAND2_X1 U645 ( .A1(G224), .A2(n439), .ZN(n529) );
  XOR2_X1 U646 ( .A(n532), .B(n531), .Z(n533) );
  XNOR2_X1 U647 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U648 ( .A(n538), .B(KEYINPUT16), .ZN(n746) );
  NOR2_X1 U649 ( .A1(n645), .A2(n631), .ZN(n543) );
  NAND2_X1 U650 ( .A1(G210), .A2(n539), .ZN(n541) );
  NAND2_X1 U651 ( .A1(n583), .A2(n585), .ZN(n544) );
  XNOR2_X1 U652 ( .A(n545), .B(n544), .ZN(n546) );
  NOR2_X1 U653 ( .A1(n700), .A2(n546), .ZN(n678) );
  INV_X1 U654 ( .A(n554), .ZN(n574) );
  NOR2_X1 U655 ( .A1(n575), .A2(n574), .ZN(n610) );
  NAND2_X1 U656 ( .A1(n585), .A2(n610), .ZN(n550) );
  NOR2_X1 U657 ( .A1(n571), .A2(n550), .ZN(n669) );
  XNOR2_X1 U658 ( .A(n669), .B(KEYINPUT81), .ZN(n552) );
  INV_X1 U659 ( .A(KEYINPUT47), .ZN(n564) );
  NAND2_X1 U660 ( .A1(KEYINPUT79), .A2(n564), .ZN(n551) );
  NAND2_X1 U661 ( .A1(n552), .A2(n551), .ZN(n553) );
  NOR2_X1 U662 ( .A1(n678), .A2(n553), .ZN(n570) );
  XNOR2_X1 U663 ( .A(KEYINPUT19), .B(KEYINPUT65), .ZN(n561) );
  NOR2_X1 U664 ( .A1(n567), .A2(KEYINPUT79), .ZN(n562) );
  NOR2_X1 U665 ( .A1(n694), .A2(n562), .ZN(n563) );
  XNOR2_X1 U666 ( .A(KEYINPUT66), .B(KEYINPUT47), .ZN(n565) );
  NOR2_X1 U667 ( .A1(KEYINPUT79), .A2(n566), .ZN(n568) );
  INV_X1 U668 ( .A(n567), .ZN(n670) );
  NOR2_X1 U669 ( .A1(n568), .A2(n670), .ZN(n569) );
  XOR2_X1 U670 ( .A(n585), .B(KEYINPUT38), .Z(n691) );
  INV_X1 U671 ( .A(n691), .ZN(n572) );
  NOR2_X1 U672 ( .A1(n582), .A2(n673), .ZN(n573) );
  XNOR2_X1 U673 ( .A(n573), .B(KEYINPUT40), .ZN(n767) );
  NAND2_X1 U674 ( .A1(n691), .A2(n690), .ZN(n695) );
  NAND2_X1 U675 ( .A1(n575), .A2(n574), .ZN(n693) );
  NOR2_X1 U676 ( .A1(n695), .A2(n693), .ZN(n576) );
  XNOR2_X1 U677 ( .A(n576), .B(KEYINPUT41), .ZN(n719) );
  XNOR2_X1 U678 ( .A(n578), .B(KEYINPUT42), .ZN(n768) );
  NOR2_X1 U679 ( .A1(n767), .A2(n768), .ZN(n579) );
  NOR2_X1 U680 ( .A1(n676), .A2(n582), .ZN(n680) );
  NAND2_X1 U681 ( .A1(n700), .A2(n583), .ZN(n584) );
  XNOR2_X1 U682 ( .A(n584), .B(KEYINPUT43), .ZN(n587) );
  INV_X1 U683 ( .A(n585), .ZN(n586) );
  NAND2_X1 U684 ( .A1(n587), .A2(n586), .ZN(n682) );
  NOR2_X1 U685 ( .A1(n702), .A2(n700), .ZN(n589) );
  AND2_X1 U686 ( .A1(n617), .A2(n589), .ZN(n599) );
  INV_X1 U687 ( .A(n693), .ZN(n595) );
  XOR2_X1 U688 ( .A(G898), .B(KEYINPUT94), .Z(n742) );
  NAND2_X1 U689 ( .A1(G953), .A2(n742), .ZN(n750) );
  NOR2_X1 U690 ( .A1(n590), .A2(n750), .ZN(n591) );
  NOR2_X1 U691 ( .A1(n592), .A2(n591), .ZN(n593) );
  INV_X1 U692 ( .A(KEYINPUT22), .ZN(n596) );
  NOR2_X1 U693 ( .A1(n702), .A2(n618), .ZN(n600) );
  NAND2_X1 U694 ( .A1(n616), .A2(n600), .ZN(n601) );
  INV_X1 U695 ( .A(KEYINPUT44), .ZN(n613) );
  NAND2_X1 U696 ( .A1(n613), .A2(KEYINPUT88), .ZN(n603) );
  XNOR2_X1 U697 ( .A(n604), .B(n603), .ZN(n611) );
  NAND2_X1 U698 ( .A1(n605), .A2(n620), .ZN(n607) );
  XOR2_X1 U699 ( .A(KEYINPUT71), .B(KEYINPUT34), .Z(n608) );
  XNOR2_X1 U700 ( .A(KEYINPUT76), .B(n608), .ZN(n609) );
  NAND2_X1 U701 ( .A1(n613), .A2(n612), .ZN(n614) );
  XOR2_X1 U702 ( .A(KEYINPUT108), .B(n619), .Z(n769) );
  NAND2_X1 U703 ( .A1(n620), .A2(n706), .ZN(n621) );
  XNOR2_X1 U704 ( .A(n621), .B(KEYINPUT100), .ZN(n710) );
  NOR2_X1 U705 ( .A1(n706), .A2(n397), .ZN(n623) );
  NAND2_X1 U706 ( .A1(n373), .A2(n623), .ZN(n661) );
  NAND2_X1 U707 ( .A1(n675), .A2(n661), .ZN(n626) );
  INV_X1 U708 ( .A(n624), .ZN(n625) );
  NAND2_X1 U709 ( .A1(n626), .A2(n625), .ZN(n627) );
  XNOR2_X1 U710 ( .A(n627), .B(KEYINPUT107), .ZN(n628) );
  NAND2_X1 U711 ( .A1(KEYINPUT83), .A2(n631), .ZN(n629) );
  INV_X1 U712 ( .A(KEYINPUT2), .ZN(n684) );
  NAND2_X1 U713 ( .A1(n629), .A2(n684), .ZN(n630) );
  NAND2_X1 U714 ( .A1(KEYINPUT2), .A2(n631), .ZN(n632) );
  NAND2_X1 U715 ( .A1(n727), .A2(G475), .ZN(n640) );
  XNOR2_X1 U716 ( .A(n638), .B(KEYINPUT59), .ZN(n639) );
  XNOR2_X1 U717 ( .A(n640), .B(n639), .ZN(n642) );
  NOR2_X1 U718 ( .A1(G952), .A2(n761), .ZN(n641) );
  NAND2_X1 U719 ( .A1(n642), .A2(n726), .ZN(n644) );
  XNOR2_X1 U720 ( .A(n644), .B(n643), .ZN(G60) );
  NAND2_X1 U721 ( .A1(n727), .A2(G210), .ZN(n649) );
  XOR2_X1 U722 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n647) );
  XNOR2_X1 U723 ( .A(KEYINPUT90), .B(KEYINPUT78), .ZN(n646) );
  XNOR2_X1 U724 ( .A(n649), .B(n648), .ZN(n650) );
  NAND2_X1 U725 ( .A1(n650), .A2(n726), .ZN(n652) );
  INV_X1 U726 ( .A(KEYINPUT56), .ZN(n651) );
  XNOR2_X1 U727 ( .A(n652), .B(n651), .ZN(G51) );
  NAND2_X1 U728 ( .A1(n727), .A2(G472), .ZN(n656) );
  XNOR2_X1 U729 ( .A(n653), .B(KEYINPUT115), .ZN(n654) );
  XNOR2_X1 U730 ( .A(n654), .B(KEYINPUT62), .ZN(n655) );
  XNOR2_X1 U731 ( .A(n656), .B(n655), .ZN(n657) );
  NAND2_X1 U732 ( .A1(n657), .A2(n726), .ZN(n658) );
  XNOR2_X1 U733 ( .A(KEYINPUT63), .B(n658), .ZN(G57) );
  NOR2_X1 U734 ( .A1(n673), .A2(n661), .ZN(n659) );
  XOR2_X1 U735 ( .A(KEYINPUT116), .B(n659), .Z(n660) );
  XNOR2_X1 U736 ( .A(G104), .B(n660), .ZN(G6) );
  NOR2_X1 U737 ( .A1(n676), .A2(n661), .ZN(n663) );
  XNOR2_X1 U738 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n662) );
  XNOR2_X1 U739 ( .A(n663), .B(n662), .ZN(n664) );
  XNOR2_X1 U740 ( .A(G107), .B(n664), .ZN(G9) );
  XNOR2_X1 U741 ( .A(G110), .B(n665), .ZN(n666) );
  XNOR2_X1 U742 ( .A(n666), .B(KEYINPUT117), .ZN(G12) );
  NOR2_X1 U743 ( .A1(n676), .A2(n670), .ZN(n668) );
  XNOR2_X1 U744 ( .A(G128), .B(KEYINPUT29), .ZN(n667) );
  XNOR2_X1 U745 ( .A(n668), .B(n667), .ZN(G30) );
  XOR2_X1 U746 ( .A(G143), .B(n669), .Z(G45) );
  NOR2_X1 U747 ( .A1(n673), .A2(n670), .ZN(n671) );
  XOR2_X1 U748 ( .A(KEYINPUT118), .B(n671), .Z(n672) );
  XNOR2_X1 U749 ( .A(G146), .B(n672), .ZN(G48) );
  NOR2_X1 U750 ( .A1(n673), .A2(n675), .ZN(n674) );
  XOR2_X1 U751 ( .A(G113), .B(n674), .Z(G15) );
  NOR2_X1 U752 ( .A1(n676), .A2(n675), .ZN(n677) );
  XOR2_X1 U753 ( .A(G116), .B(n677), .Z(G18) );
  XNOR2_X1 U754 ( .A(G125), .B(n678), .ZN(n679) );
  XNOR2_X1 U755 ( .A(n679), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U756 ( .A(G134), .B(n680), .ZN(n681) );
  XNOR2_X1 U757 ( .A(n681), .B(KEYINPUT119), .ZN(G36) );
  XNOR2_X1 U758 ( .A(G140), .B(KEYINPUT120), .ZN(n683) );
  XNOR2_X1 U759 ( .A(n683), .B(n682), .ZN(G42) );
  NAND2_X1 U760 ( .A1(n686), .A2(n685), .ZN(n688) );
  NOR2_X1 U761 ( .A1(n688), .A2(n687), .ZN(n689) );
  NOR2_X1 U762 ( .A1(n691), .A2(n690), .ZN(n692) );
  NOR2_X1 U763 ( .A1(n693), .A2(n692), .ZN(n697) );
  NOR2_X1 U764 ( .A1(n695), .A2(n694), .ZN(n696) );
  NOR2_X1 U765 ( .A1(n697), .A2(n696), .ZN(n698) );
  NOR2_X1 U766 ( .A1(n698), .A2(n720), .ZN(n715) );
  XNOR2_X1 U767 ( .A(KEYINPUT51), .B(KEYINPUT122), .ZN(n712) );
  NAND2_X1 U768 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U769 ( .A(KEYINPUT50), .B(n701), .ZN(n708) );
  XOR2_X1 U770 ( .A(KEYINPUT49), .B(KEYINPUT121), .Z(n704) );
  OR2_X1 U771 ( .A1(n365), .A2(n702), .ZN(n703) );
  XNOR2_X1 U772 ( .A(n704), .B(n703), .ZN(n705) );
  NOR2_X1 U773 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U774 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U775 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U776 ( .A(n712), .B(n711), .ZN(n713) );
  NOR2_X1 U777 ( .A1(n719), .A2(n713), .ZN(n714) );
  NOR2_X1 U778 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U779 ( .A(n716), .B(KEYINPUT52), .ZN(n717) );
  NOR2_X1 U780 ( .A1(n718), .A2(n717), .ZN(n722) );
  NOR2_X1 U781 ( .A1(n720), .A2(n719), .ZN(n721) );
  NOR2_X1 U782 ( .A1(n722), .A2(n721), .ZN(n723) );
  INV_X1 U783 ( .A(KEYINPUT124), .ZN(n724) );
  XNOR2_X1 U784 ( .A(KEYINPUT53), .B(n725), .ZN(G75) );
  INV_X1 U785 ( .A(n726), .ZN(n739) );
  NAND2_X1 U786 ( .A1(G469), .A2(n727), .ZN(n731) );
  XOR2_X1 U787 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n728) );
  NOR2_X1 U788 ( .A1(n739), .A2(n732), .ZN(G54) );
  NAND2_X1 U789 ( .A1(G478), .A2(n736), .ZN(n733) );
  XNOR2_X1 U790 ( .A(n733), .B(n734), .ZN(n735) );
  NOR2_X1 U791 ( .A1(n739), .A2(n735), .ZN(G63) );
  NAND2_X1 U792 ( .A1(G217), .A2(n736), .ZN(n737) );
  NAND2_X1 U793 ( .A1(G953), .A2(G224), .ZN(n740) );
  XOR2_X1 U794 ( .A(KEYINPUT61), .B(n740), .Z(n741) );
  NOR2_X1 U795 ( .A1(n742), .A2(n741), .ZN(n745) );
  NOR2_X1 U796 ( .A1(G953), .A2(n743), .ZN(n744) );
  NOR2_X1 U797 ( .A1(n745), .A2(n744), .ZN(n753) );
  XOR2_X1 U798 ( .A(n746), .B(KEYINPUT126), .Z(n747) );
  XNOR2_X1 U799 ( .A(n748), .B(n747), .ZN(n749) );
  XNOR2_X1 U800 ( .A(n749), .B(G101), .ZN(n751) );
  NAND2_X1 U801 ( .A1(n751), .A2(n750), .ZN(n752) );
  XNOR2_X1 U802 ( .A(n753), .B(n752), .ZN(G69) );
  XOR2_X1 U803 ( .A(n754), .B(KEYINPUT4), .Z(n755) );
  XOR2_X1 U804 ( .A(n756), .B(n755), .Z(n760) );
  XOR2_X1 U805 ( .A(n760), .B(KEYINPUT127), .Z(n757) );
  XNOR2_X1 U806 ( .A(G227), .B(n757), .ZN(n758) );
  NAND2_X1 U807 ( .A1(G900), .A2(n758), .ZN(n759) );
  NAND2_X1 U808 ( .A1(n759), .A2(G953), .ZN(n764) );
  NAND2_X1 U809 ( .A1(n762), .A2(n761), .ZN(n763) );
  NAND2_X1 U810 ( .A1(n764), .A2(n763), .ZN(G72) );
  XNOR2_X1 U811 ( .A(G122), .B(n765), .ZN(G24) );
  XOR2_X1 U812 ( .A(n766), .B(G119), .Z(G21) );
  XOR2_X1 U813 ( .A(n767), .B(G131), .Z(G33) );
  XOR2_X1 U814 ( .A(n768), .B(G137), .Z(G39) );
  XOR2_X1 U815 ( .A(G101), .B(n769), .Z(G3) );
endmodule

