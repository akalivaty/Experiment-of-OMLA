//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 0 0 0 0 0 0 1 1 0 0 1 0 0 1 0 1 0 1 1 1 1 0 1 0 1 1 1 0 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 1 0 0 0 0 0 0 0 0 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:57 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n748, new_n749,
    new_n750, new_n752, new_n753, new_n754, new_n756, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n787, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n843, new_n844, new_n846, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n886, new_n887, new_n888,
    new_n890, new_n891, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n899, new_n901, new_n902, new_n903, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n939,
    new_n940;
  INV_X1    g000(.A(KEYINPUT87), .ZN(new_n202));
  INV_X1    g001(.A(G169gat), .ZN(new_n203));
  INV_X1    g002(.A(G176gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT67), .ZN(new_n206));
  OAI21_X1  g005(.A(KEYINPUT26), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(G169gat), .A2(G176gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(G169gat), .A2(G176gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT26), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n209), .A2(KEYINPUT67), .A3(new_n210), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n207), .A2(new_n208), .A3(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G190gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(KEYINPUT66), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT66), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(G190gat), .ZN(new_n216));
  INV_X1    g015(.A(G183gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(KEYINPUT27), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT27), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(G183gat), .ZN(new_n220));
  NAND4_X1  g019(.A1(new_n214), .A2(new_n216), .A3(new_n218), .A4(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(KEYINPUT28), .ZN(new_n222));
  NAND2_X1  g021(.A1(G183gat), .A2(G190gat), .ZN(new_n223));
  XNOR2_X1  g022(.A(KEYINPUT66), .B(G190gat), .ZN(new_n224));
  XNOR2_X1  g023(.A(KEYINPUT27), .B(G183gat), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT28), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  NAND4_X1  g026(.A1(new_n212), .A2(new_n222), .A3(new_n223), .A4(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(G226gat), .A2(G233gat), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n203), .A2(new_n204), .A3(KEYINPUT23), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(new_n208), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT64), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n232), .B1(new_n209), .B2(KEYINPUT23), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT23), .ZN(new_n234));
  OAI211_X1 g033(.A(new_n234), .B(KEYINPUT64), .C1(G169gat), .C2(G176gat), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n231), .B1(new_n233), .B2(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n214), .A2(new_n216), .A3(new_n217), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n223), .A2(KEYINPUT65), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(KEYINPUT24), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT24), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n223), .A2(KEYINPUT65), .A3(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n237), .A2(new_n239), .A3(new_n241), .ZN(new_n242));
  AND3_X1   g041(.A1(new_n236), .A2(KEYINPUT25), .A3(new_n242), .ZN(new_n243));
  OAI21_X1  g042(.A(G190gat), .B1(KEYINPUT24), .B2(G183gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n244), .B(new_n245), .ZN(new_n246));
  AOI21_X1  g045(.A(KEYINPUT25), .B1(new_n236), .B2(new_n246), .ZN(new_n247));
  OAI211_X1 g046(.A(new_n228), .B(new_n229), .C1(new_n243), .C2(new_n247), .ZN(new_n248));
  AND3_X1   g047(.A1(new_n222), .A2(new_n223), .A3(new_n227), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT25), .ZN(new_n250));
  AND2_X1   g049(.A1(G169gat), .A2(G176gat), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n251), .B1(KEYINPUT23), .B2(new_n209), .ZN(new_n252));
  AOI21_X1  g051(.A(KEYINPUT64), .B1(new_n205), .B2(new_n234), .ZN(new_n253));
  NOR3_X1   g052(.A1(new_n209), .A2(new_n232), .A3(KEYINPUT23), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n252), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(new_n244), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(new_n245), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n213), .A2(KEYINPUT24), .A3(G183gat), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n250), .B1(new_n255), .B2(new_n259), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n236), .A2(KEYINPUT25), .A3(new_n242), .ZN(new_n261));
  AOI22_X1  g060(.A1(new_n212), .A2(new_n249), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n229), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n263), .A2(KEYINPUT29), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n248), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(G211gat), .B(G218gat), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT72), .ZN(new_n267));
  OR2_X1    g066(.A1(KEYINPUT71), .A2(G197gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(KEYINPUT71), .A2(G197gat), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n268), .A2(G204gat), .A3(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(G204gat), .ZN(new_n271));
  AND2_X1   g070(.A1(KEYINPUT71), .A2(G197gat), .ZN(new_n272));
  NOR2_X1   g071(.A1(KEYINPUT71), .A2(G197gat), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n271), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n270), .A2(new_n274), .ZN(new_n275));
  AOI21_X1  g074(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n267), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  AOI211_X1 g077(.A(KEYINPUT72), .B(new_n276), .C1(new_n270), .C2(new_n274), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n266), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NOR3_X1   g079(.A1(new_n272), .A2(new_n273), .A3(new_n271), .ZN(new_n281));
  AOI21_X1  g080(.A(G204gat), .B1(new_n268), .B2(new_n269), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n277), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(KEYINPUT72), .ZN(new_n284));
  INV_X1    g083(.A(new_n266), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n275), .A2(new_n267), .A3(new_n277), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n284), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n280), .A2(new_n287), .A3(KEYINPUT73), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n280), .A2(new_n287), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT73), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n265), .A2(new_n288), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(KEYINPUT74), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n233), .A2(new_n235), .ZN(new_n294));
  AND3_X1   g093(.A1(new_n294), .A2(KEYINPUT25), .A3(new_n252), .ZN(new_n295));
  NAND4_X1  g094(.A1(new_n294), .A2(new_n252), .A3(new_n258), .A4(new_n257), .ZN(new_n296));
  AOI22_X1  g095(.A1(new_n295), .A2(new_n242), .B1(new_n296), .B2(new_n250), .ZN(new_n297));
  INV_X1    g096(.A(new_n228), .ZN(new_n298));
  OAI22_X1  g097(.A1(new_n297), .A2(new_n298), .B1(KEYINPUT29), .B2(new_n263), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n299), .A2(new_n248), .A3(new_n289), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT74), .ZN(new_n301));
  NAND4_X1  g100(.A1(new_n265), .A2(new_n301), .A3(new_n288), .A4(new_n291), .ZN(new_n302));
  XNOR2_X1  g101(.A(G8gat), .B(G36gat), .ZN(new_n303));
  XNOR2_X1  g102(.A(G64gat), .B(G92gat), .ZN(new_n304));
  XOR2_X1   g103(.A(new_n303), .B(new_n304), .Z(new_n305));
  NAND4_X1  g104(.A1(new_n293), .A2(new_n300), .A3(new_n302), .A4(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT30), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n302), .A2(new_n300), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  NAND4_X1  g109(.A1(new_n310), .A2(KEYINPUT30), .A3(new_n293), .A4(new_n305), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n308), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT75), .ZN(new_n313));
  AND3_X1   g112(.A1(new_n280), .A2(new_n287), .A3(KEYINPUT73), .ZN(new_n314));
  AOI21_X1  g113(.A(KEYINPUT73), .B1(new_n280), .B2(new_n287), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n301), .B1(new_n316), .B2(new_n265), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n313), .B1(new_n309), .B2(new_n317), .ZN(new_n318));
  NAND4_X1  g117(.A1(new_n293), .A2(KEYINPUT75), .A3(new_n300), .A4(new_n302), .ZN(new_n319));
  INV_X1    g118(.A(new_n305), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n318), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(KEYINPUT76), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT76), .ZN(new_n323));
  NAND4_X1  g122(.A1(new_n318), .A2(new_n319), .A3(new_n323), .A4(new_n320), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n312), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(G141gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(G148gat), .ZN(new_n327));
  INV_X1    g126(.A(G148gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(G141gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(G155gat), .A2(G162gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(KEYINPUT2), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(G155gat), .ZN(new_n334));
  INV_X1    g133(.A(G162gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n333), .A2(new_n331), .A3(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT3), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n336), .A2(new_n331), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n330), .A2(new_n339), .A3(new_n332), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n337), .A2(new_n338), .A3(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT29), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n291), .A2(new_n288), .A3(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(G228gat), .ZN(new_n345));
  INV_X1    g144(.A(G233gat), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n337), .A2(new_n340), .ZN(new_n348));
  AOI21_X1  g147(.A(KEYINPUT29), .B1(new_n280), .B2(new_n287), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n348), .B1(new_n349), .B2(KEYINPUT3), .ZN(new_n350));
  AND3_X1   g149(.A1(new_n344), .A2(new_n347), .A3(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n280), .A2(new_n287), .A3(new_n343), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n347), .B1(new_n350), .B2(new_n352), .ZN(new_n353));
  OAI21_X1  g152(.A(G22gat), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n350), .A2(new_n352), .ZN(new_n355));
  INV_X1    g154(.A(new_n347), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n344), .A2(new_n347), .A3(new_n350), .ZN(new_n358));
  INV_X1    g157(.A(G22gat), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n357), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n354), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n289), .A2(new_n342), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(new_n338), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n356), .B1(new_n363), .B2(new_n348), .ZN(new_n364));
  AOI22_X1  g163(.A1(new_n364), .A2(new_n344), .B1(new_n355), .B2(new_n356), .ZN(new_n365));
  AOI21_X1  g164(.A(KEYINPUT82), .B1(new_n365), .B2(new_n359), .ZN(new_n366));
  XNOR2_X1  g165(.A(G78gat), .B(G106gat), .ZN(new_n367));
  XNOR2_X1  g166(.A(KEYINPUT31), .B(G50gat), .ZN(new_n368));
  XNOR2_X1  g167(.A(new_n367), .B(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n361), .B1(new_n366), .B2(new_n370), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n354), .A2(new_n360), .A3(KEYINPUT82), .A4(new_n369), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  OR2_X1    g172(.A1(G113gat), .A2(G120gat), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT1), .ZN(new_n375));
  NAND2_X1  g174(.A1(G113gat), .A2(G120gat), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n374), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  AND2_X1   g176(.A1(G127gat), .A2(G134gat), .ZN(new_n378));
  NOR2_X1   g177(.A1(G127gat), .A2(G134gat), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n377), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n374), .A2(KEYINPUT69), .A3(new_n376), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT69), .ZN(new_n383));
  AND2_X1   g182(.A1(G113gat), .A2(G120gat), .ZN(new_n384));
  NOR2_X1   g183(.A1(G113gat), .A2(G120gat), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n383), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n382), .A2(new_n386), .A3(new_n375), .ZN(new_n387));
  XNOR2_X1  g186(.A(KEYINPUT68), .B(G127gat), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n379), .B1(new_n388), .B2(G134gat), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n381), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n390), .B1(new_n297), .B2(new_n298), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n387), .A2(new_n389), .ZN(new_n392));
  INV_X1    g191(.A(new_n381), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  OAI211_X1 g193(.A(new_n394), .B(new_n228), .C1(new_n243), .C2(new_n247), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n391), .A2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(G227gat), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n397), .A2(new_n346), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n396), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(KEYINPUT34), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT34), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n396), .A2(new_n402), .A3(new_n399), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  XNOR2_X1  g204(.A(G15gat), .B(G43gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(G71gat), .B(G99gat), .ZN(new_n407));
  XNOR2_X1  g206(.A(new_n406), .B(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n391), .A2(new_n398), .A3(new_n395), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n408), .B1(new_n409), .B2(KEYINPUT32), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT33), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT70), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n410), .A2(KEYINPUT70), .A3(new_n412), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  OAI211_X1 g216(.A(new_n409), .B(KEYINPUT32), .C1(new_n411), .C2(new_n408), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n405), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(new_n418), .ZN(new_n420));
  AOI211_X1 g219(.A(new_n404), .B(new_n420), .C1(new_n415), .C2(new_n416), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT35), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n325), .A2(new_n373), .A3(new_n422), .A4(new_n423), .ZN(new_n424));
  AND3_X1   g223(.A1(new_n330), .A2(new_n339), .A3(new_n332), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n339), .B1(new_n332), .B2(new_n330), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n390), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(KEYINPUT4), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT4), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n390), .A2(new_n427), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  OAI21_X1  g231(.A(KEYINPUT3), .B1(new_n425), .B2(new_n426), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n394), .A2(new_n341), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(G225gat), .A2(G233gat), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n436), .A2(KEYINPUT5), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n432), .A2(new_n434), .A3(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT5), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n434), .A2(new_n435), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT77), .ZN(new_n442));
  AOI211_X1 g241(.A(new_n442), .B(new_n430), .C1(new_n390), .C2(new_n427), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n429), .A2(new_n442), .A3(new_n431), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n440), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(new_n428), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n390), .A2(new_n427), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n436), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT78), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n394), .A2(new_n348), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(new_n428), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n453), .A2(KEYINPUT78), .A3(new_n436), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n451), .A2(new_n454), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n439), .B1(new_n446), .B2(new_n455), .ZN(new_n456));
  XOR2_X1   g255(.A(G1gat), .B(G29gat), .Z(new_n457));
  XNOR2_X1  g256(.A(G57gat), .B(G85gat), .ZN(new_n458));
  XNOR2_X1  g257(.A(new_n457), .B(new_n458), .ZN(new_n459));
  XNOR2_X1  g258(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n460));
  XNOR2_X1  g259(.A(new_n459), .B(new_n460), .ZN(new_n461));
  AOI21_X1  g260(.A(KEYINPUT6), .B1(new_n456), .B2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(new_n461), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT83), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n463), .B1(new_n456), .B2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(new_n445), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n435), .B(new_n434), .C1(new_n429), .C2(new_n442), .ZN(new_n467));
  OAI21_X1  g266(.A(KEYINPUT5), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  AOI21_X1  g267(.A(KEYINPUT78), .B1(new_n453), .B2(new_n436), .ZN(new_n469));
  AOI211_X1 g268(.A(new_n450), .B(new_n435), .C1(new_n452), .C2(new_n428), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n438), .B1(new_n468), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n472), .A2(KEYINPUT83), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n462), .B1(new_n465), .B2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT84), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n472), .A2(KEYINPUT6), .A3(new_n463), .ZN(new_n477));
  OAI211_X1 g276(.A(KEYINPUT84), .B(new_n462), .C1(new_n465), .C2(new_n473), .ZN(new_n478));
  AND3_X1   g277(.A1(new_n476), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n202), .B1(new_n424), .B2(new_n479), .ZN(new_n480));
  AND2_X1   g279(.A1(new_n325), .A2(new_n423), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT82), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n360), .A2(new_n482), .ZN(new_n483));
  AOI22_X1  g282(.A1(new_n483), .A2(new_n369), .B1(new_n360), .B2(new_n354), .ZN(new_n484));
  INV_X1    g283(.A(new_n372), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(new_n416), .ZN(new_n487));
  AOI21_X1  g286(.A(KEYINPUT70), .B1(new_n410), .B2(new_n412), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n418), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(new_n404), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n417), .A2(new_n405), .A3(new_n418), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n486), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n476), .A2(new_n477), .A3(new_n478), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n481), .A2(new_n493), .A3(KEYINPUT87), .A4(new_n494), .ZN(new_n495));
  AND2_X1   g294(.A1(new_n480), .A2(new_n495), .ZN(new_n496));
  OAI21_X1  g295(.A(KEYINPUT80), .B1(new_n456), .B2(new_n461), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT80), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n472), .A2(new_n498), .A3(new_n463), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n497), .A2(new_n462), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(new_n477), .ZN(new_n501));
  AOI21_X1  g300(.A(KEYINPUT81), .B1(new_n325), .B2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n325), .A2(KEYINPUT81), .A3(new_n501), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n503), .A2(new_n504), .A3(new_n493), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(KEYINPUT35), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n322), .A2(new_n324), .ZN(new_n507));
  INV_X1    g306(.A(new_n312), .ZN(new_n508));
  AND4_X1   g307(.A1(KEYINPUT81), .A2(new_n507), .A3(new_n501), .A4(new_n508), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n486), .B1(new_n509), .B2(new_n502), .ZN(new_n510));
  AND3_X1   g309(.A1(new_n490), .A2(KEYINPUT36), .A3(new_n491), .ZN(new_n511));
  AOI21_X1  g310(.A(KEYINPUT36), .B1(new_n490), .B2(new_n491), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n507), .A2(new_n508), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n465), .A2(new_n473), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n435), .B1(new_n432), .B2(new_n434), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT39), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n463), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  OAI21_X1  g317(.A(KEYINPUT39), .B1(new_n453), .B2(new_n436), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n518), .B1(new_n516), .B2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT40), .ZN(new_n521));
  AND2_X1   g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n520), .A2(new_n521), .ZN(new_n523));
  NOR3_X1   g322(.A1(new_n515), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n486), .B1(new_n514), .B2(new_n524), .ZN(new_n525));
  AND2_X1   g324(.A1(new_n478), .A2(new_n477), .ZN(new_n526));
  XNOR2_X1  g325(.A(KEYINPUT85), .B(KEYINPUT37), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n293), .A2(new_n300), .A3(new_n302), .A4(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT86), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND4_X1  g329(.A1(new_n310), .A2(KEYINPUT86), .A3(new_n293), .A4(new_n527), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n316), .A2(new_n248), .A3(new_n299), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT37), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n533), .B1(new_n265), .B2(new_n289), .ZN(new_n534));
  AOI21_X1  g333(.A(KEYINPUT38), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n530), .A2(new_n531), .A3(new_n320), .A4(new_n535), .ZN(new_n536));
  AND2_X1   g335(.A1(new_n536), .A2(new_n306), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n530), .A2(new_n531), .A3(new_n320), .ZN(new_n538));
  AND3_X1   g337(.A1(new_n318), .A2(KEYINPUT37), .A3(new_n319), .ZN(new_n539));
  OAI21_X1  g338(.A(KEYINPUT38), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n526), .A2(new_n537), .A3(new_n476), .A4(new_n540), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n513), .B1(new_n525), .B2(new_n541), .ZN(new_n542));
  AOI22_X1  g341(.A1(new_n496), .A2(new_n506), .B1(new_n510), .B2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(G29gat), .ZN(new_n544));
  AND3_X1   g343(.A1(new_n544), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(KEYINPUT14), .B(G29gat), .ZN(new_n546));
  INV_X1    g345(.A(G36gat), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(G43gat), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n549), .A2(G50gat), .ZN(new_n550));
  XNOR2_X1  g349(.A(KEYINPUT89), .B(G50gat), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(new_n549), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n550), .B1(new_n552), .B2(KEYINPUT90), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n553), .B1(KEYINPUT90), .B2(new_n552), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT15), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n548), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(G43gat), .B(G50gat), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT88), .ZN(new_n558));
  AND2_X1   g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n557), .A2(new_n558), .ZN(new_n560));
  NOR3_X1   g359(.A1(new_n559), .A2(new_n560), .A3(new_n555), .ZN(new_n561));
  MUX2_X1   g360(.A(new_n556), .B(new_n548), .S(new_n561), .Z(new_n562));
  XNOR2_X1  g361(.A(G15gat), .B(G22gat), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT16), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n563), .B1(new_n564), .B2(G1gat), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n565), .B1(G1gat), .B2(new_n563), .ZN(new_n566));
  XOR2_X1   g365(.A(new_n566), .B(G8gat), .Z(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n562), .A2(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n569), .B(KEYINPUT91), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT17), .ZN(new_n571));
  OR2_X1    g370(.A1(new_n562), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n562), .A2(new_n571), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n572), .A2(new_n567), .A3(new_n573), .ZN(new_n574));
  AND2_X1   g373(.A1(new_n570), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(G229gat), .A2(G233gat), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT18), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n575), .A2(KEYINPUT18), .A3(new_n576), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n570), .B1(new_n562), .B2(new_n568), .ZN(new_n581));
  XOR2_X1   g380(.A(new_n576), .B(KEYINPUT13), .Z(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n579), .A2(new_n580), .A3(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(G113gat), .B(G141gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(G197gat), .ZN(new_n586));
  XOR2_X1   g385(.A(KEYINPUT11), .B(G169gat), .Z(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  XOR2_X1   g387(.A(new_n588), .B(KEYINPUT12), .Z(new_n589));
  NAND2_X1  g388(.A1(new_n584), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n589), .ZN(new_n591));
  NAND4_X1  g390(.A1(new_n579), .A2(new_n591), .A3(new_n580), .A4(new_n583), .ZN(new_n592));
  AND3_X1   g391(.A1(new_n590), .A2(KEYINPUT92), .A3(new_n592), .ZN(new_n593));
  AOI21_X1  g392(.A(KEYINPUT92), .B1(new_n590), .B2(new_n592), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n543), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(G85gat), .A2(G92gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n597), .B(KEYINPUT7), .ZN(new_n598));
  NAND2_X1  g397(.A1(G99gat), .A2(G106gat), .ZN(new_n599));
  INV_X1    g398(.A(G85gat), .ZN(new_n600));
  INV_X1    g399(.A(G92gat), .ZN(new_n601));
  AOI22_X1  g400(.A1(KEYINPUT8), .A2(new_n599), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n598), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(G99gat), .B(G106gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(G71gat), .A2(G78gat), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT9), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n606), .B1(new_n607), .B2(KEYINPUT93), .ZN(new_n608));
  INV_X1    g407(.A(G71gat), .ZN(new_n609));
  INV_X1    g408(.A(G78gat), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n608), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n607), .B1(new_n609), .B2(new_n610), .ZN(new_n612));
  NAND2_X1  g411(.A1(G57gat), .A2(G64gat), .ZN(new_n613));
  OR2_X1    g412(.A1(G57gat), .A2(G64gat), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n612), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  OR2_X1    g414(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n611), .A2(new_n615), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n605), .B(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT10), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND4_X1  g420(.A1(new_n605), .A2(KEYINPUT10), .A3(new_n616), .A4(new_n617), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(G230gat), .A2(G233gat), .ZN(new_n624));
  AND2_X1   g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n619), .A2(new_n624), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  XOR2_X1   g426(.A(G120gat), .B(G148gat), .Z(new_n628));
  XNOR2_X1  g427(.A(G176gat), .B(G204gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n627), .A2(new_n630), .ZN(new_n631));
  XOR2_X1   g430(.A(new_n631), .B(KEYINPUT99), .Z(new_n632));
  NOR2_X1   g431(.A1(new_n627), .A2(new_n630), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(KEYINPUT100), .ZN(new_n634));
  AND2_X1   g433(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT101), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  AND3_X1   g436(.A1(new_n632), .A2(new_n636), .A3(new_n634), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n605), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n572), .A2(new_n573), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n562), .A2(new_n605), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT41), .ZN(new_n644));
  NAND2_X1  g443(.A1(G232gat), .A2(G233gat), .ZN(new_n645));
  XOR2_X1   g444(.A(new_n645), .B(KEYINPUT96), .Z(new_n646));
  OAI211_X1 g445(.A(new_n642), .B(new_n643), .C1(new_n644), .C2(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(G190gat), .B(G218gat), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n647), .B(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n646), .A2(new_n644), .ZN(new_n650));
  XOR2_X1   g449(.A(G134gat), .B(G162gat), .Z(new_n651));
  XNOR2_X1  g450(.A(new_n650), .B(new_n651), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n652), .A2(KEYINPUT97), .ZN(new_n653));
  OR2_X1    g452(.A1(new_n649), .A2(new_n653), .ZN(new_n654));
  AND2_X1   g453(.A1(new_n652), .A2(KEYINPUT97), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n649), .B1(new_n655), .B2(new_n653), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT21), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n567), .B1(new_n659), .B2(new_n618), .ZN(new_n660));
  XOR2_X1   g459(.A(new_n660), .B(KEYINPUT95), .Z(new_n661));
  NAND2_X1  g460(.A1(G231gat), .A2(G233gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(KEYINPUT94), .ZN(new_n663));
  XOR2_X1   g462(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n664));
  XNOR2_X1  g463(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n661), .B(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n618), .A2(new_n659), .ZN(new_n667));
  XOR2_X1   g466(.A(G127gat), .B(G155gat), .Z(new_n668));
  XNOR2_X1  g467(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XOR2_X1   g468(.A(G183gat), .B(G211gat), .Z(new_n670));
  XNOR2_X1  g469(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n666), .B(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n658), .A2(KEYINPUT98), .A3(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT98), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n675), .B1(new_n657), .B2(new_n672), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n640), .A2(new_n677), .ZN(new_n678));
  AND2_X1   g477(.A1(new_n596), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n501), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n681), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g481(.A1(new_n679), .A2(new_n514), .ZN(new_n683));
  XNOR2_X1  g482(.A(KEYINPUT16), .B(G8gat), .ZN(new_n684));
  OR2_X1    g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT42), .ZN(new_n686));
  OR2_X1    g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT102), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  AND2_X1   g488(.A1(new_n687), .A2(new_n688), .ZN(new_n690));
  AND2_X1   g489(.A1(new_n683), .A2(G8gat), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n685), .B1(new_n691), .B2(new_n686), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n689), .B1(new_n690), .B2(new_n692), .ZN(G1325gat));
  INV_X1    g492(.A(new_n679), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n513), .B(KEYINPUT103), .ZN(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  OAI21_X1  g495(.A(G15gat), .B1(new_n694), .B2(new_n696), .ZN(new_n697));
  OR2_X1    g496(.A1(new_n492), .A2(G15gat), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n697), .B1(new_n694), .B2(new_n698), .ZN(G1326gat));
  NAND2_X1  g498(.A1(new_n679), .A2(new_n486), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(KEYINPUT104), .ZN(new_n701));
  XOR2_X1   g500(.A(KEYINPUT43), .B(G22gat), .Z(new_n702));
  XNOR2_X1  g501(.A(new_n701), .B(new_n702), .ZN(G1327gat));
  NOR2_X1   g502(.A1(KEYINPUT106), .A2(KEYINPUT44), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n704), .B1(new_n543), .B2(new_n658), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n542), .A2(new_n510), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n509), .A2(new_n502), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n423), .B1(new_n707), .B2(new_n493), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n480), .A2(new_n495), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n706), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  XOR2_X1   g509(.A(KEYINPUT106), .B(KEYINPUT44), .Z(new_n711));
  NAND3_X1  g510(.A1(new_n710), .A2(new_n657), .A3(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n705), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n590), .A2(new_n592), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n639), .A2(new_n672), .ZN(new_n716));
  NOR3_X1   g515(.A1(new_n713), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(new_n717), .ZN(new_n718));
  OAI21_X1  g517(.A(G29gat), .B1(new_n718), .B2(new_n501), .ZN(new_n719));
  NOR4_X1   g518(.A1(new_n543), .A2(new_n716), .A3(new_n595), .A4(new_n658), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n720), .A2(new_n544), .A3(new_n680), .ZN(new_n721));
  XOR2_X1   g520(.A(KEYINPUT105), .B(KEYINPUT45), .Z(new_n722));
  XNOR2_X1  g521(.A(new_n721), .B(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n719), .A2(new_n723), .ZN(G1328gat));
  OAI21_X1  g523(.A(G36gat), .B1(new_n718), .B2(new_n325), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n720), .A2(new_n547), .A3(new_n514), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT46), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n727), .A2(KEYINPUT107), .ZN(new_n728));
  AND2_X1   g527(.A1(new_n727), .A2(KEYINPUT107), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n726), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  OAI211_X1 g529(.A(new_n725), .B(new_n730), .C1(new_n728), .C2(new_n726), .ZN(G1329gat));
  INV_X1    g530(.A(new_n513), .ZN(new_n732));
  OAI21_X1  g531(.A(G43gat), .B1(new_n718), .B2(new_n732), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n492), .A2(G43gat), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n720), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n733), .A2(KEYINPUT47), .A3(new_n735), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n549), .B1(new_n717), .B2(new_n695), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n737), .B1(new_n720), .B2(new_n734), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n736), .B1(new_n738), .B2(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g538(.A1(new_n717), .A2(new_n486), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n373), .A2(new_n551), .ZN(new_n741));
  AOI22_X1  g540(.A1(new_n740), .A2(new_n551), .B1(new_n720), .B2(new_n741), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n742), .A2(KEYINPUT108), .ZN(new_n743));
  XOR2_X1   g542(.A(new_n743), .B(KEYINPUT48), .Z(G1331gat));
  NOR4_X1   g543(.A1(new_n543), .A2(new_n677), .A3(new_n714), .A4(new_n639), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(new_n680), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g546(.A1(new_n745), .A2(new_n514), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n748), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n749));
  XOR2_X1   g548(.A(KEYINPUT49), .B(G64gat), .Z(new_n750));
  OAI21_X1  g549(.A(new_n749), .B1(new_n748), .B2(new_n750), .ZN(G1333gat));
  AOI21_X1  g550(.A(new_n609), .B1(new_n745), .B2(new_n695), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n492), .A2(G71gat), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n752), .B1(new_n745), .B2(new_n753), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g554(.A1(new_n745), .A2(new_n486), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g556(.A1(new_n639), .A2(new_n714), .A3(new_n673), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n705), .A2(new_n712), .A3(new_n758), .ZN(new_n759));
  OAI21_X1  g558(.A(G85gat), .B1(new_n759), .B2(new_n501), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT51), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n710), .A2(KEYINPUT109), .A3(new_n657), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n714), .A2(new_n673), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  AOI21_X1  g563(.A(KEYINPUT109), .B1(new_n710), .B2(new_n657), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n761), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT109), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n767), .B1(new_n543), .B2(new_n658), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n768), .A2(KEYINPUT51), .A3(new_n763), .A4(new_n762), .ZN(new_n769));
  AND2_X1   g568(.A1(new_n766), .A2(new_n769), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n640), .A2(new_n600), .A3(new_n680), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n760), .B1(new_n770), .B2(new_n771), .ZN(G1336gat));
  OAI21_X1  g571(.A(G92gat), .B1(new_n759), .B2(new_n325), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT52), .ZN(new_n774));
  NOR3_X1   g573(.A1(new_n639), .A2(G92gat), .A3(new_n325), .ZN(new_n775));
  INV_X1    g574(.A(new_n775), .ZN(new_n776));
  OAI211_X1 g575(.A(new_n773), .B(new_n774), .C1(new_n770), .C2(new_n776), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n766), .A2(KEYINPUT111), .A3(new_n769), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT111), .ZN(new_n779));
  OAI211_X1 g578(.A(new_n779), .B(new_n761), .C1(new_n764), .C2(new_n765), .ZN(new_n780));
  XOR2_X1   g579(.A(new_n775), .B(KEYINPUT110), .Z(new_n781));
  NAND3_X1  g580(.A1(new_n778), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  AND2_X1   g581(.A1(new_n782), .A2(new_n773), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n777), .B1(new_n783), .B2(new_n774), .ZN(G1337gat));
  OAI21_X1  g583(.A(G99gat), .B1(new_n759), .B2(new_n696), .ZN(new_n785));
  OR3_X1    g584(.A1(new_n639), .A2(G99gat), .A3(new_n492), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n785), .B1(new_n770), .B2(new_n786), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n787), .B(KEYINPUT112), .ZN(G1338gat));
  NAND4_X1  g587(.A1(new_n705), .A2(new_n486), .A3(new_n712), .A4(new_n758), .ZN(new_n789));
  AOI21_X1  g588(.A(KEYINPUT53), .B1(new_n789), .B2(G106gat), .ZN(new_n790));
  NOR3_X1   g589(.A1(new_n639), .A2(G106gat), .A3(new_n373), .ZN(new_n791));
  INV_X1    g590(.A(new_n791), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n790), .B1(new_n770), .B2(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT113), .ZN(new_n794));
  AND3_X1   g593(.A1(new_n789), .A2(new_n794), .A3(G106gat), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n794), .B1(new_n789), .B2(G106gat), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  XOR2_X1   g596(.A(new_n791), .B(KEYINPUT114), .Z(new_n798));
  NAND3_X1  g597(.A1(new_n778), .A2(new_n780), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  AOI21_X1  g599(.A(KEYINPUT115), .B1(new_n800), .B2(KEYINPUT53), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT115), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT53), .ZN(new_n803));
  AOI211_X1 g602(.A(new_n802), .B(new_n803), .C1(new_n797), .C2(new_n799), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n793), .B1(new_n801), .B2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT116), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  OAI211_X1 g606(.A(KEYINPUT116), .B(new_n793), .C1(new_n801), .C2(new_n804), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(G1339gat));
  NAND2_X1  g608(.A1(new_n678), .A2(new_n715), .ZN(new_n810));
  OR2_X1    g609(.A1(new_n623), .A2(new_n624), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n623), .A2(new_n624), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n811), .A2(KEYINPUT54), .A3(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT117), .ZN(new_n814));
  XNOR2_X1  g613(.A(new_n813), .B(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT54), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n630), .B1(new_n625), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT55), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT118), .ZN(new_n821));
  XNOR2_X1  g620(.A(new_n820), .B(new_n821), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n575), .A2(new_n576), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n581), .A2(new_n582), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n588), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  AND2_X1   g624(.A1(new_n592), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n815), .A2(KEYINPUT55), .A3(new_n817), .ZN(new_n827));
  AND2_X1   g626(.A1(new_n632), .A2(new_n827), .ZN(new_n828));
  AND4_X1   g627(.A1(new_n657), .A2(new_n822), .A3(new_n826), .A4(new_n828), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n826), .B1(new_n637), .B2(new_n638), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n822), .A2(new_n828), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n830), .B1(new_n831), .B2(new_n715), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n829), .B1(new_n832), .B2(new_n658), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n810), .B1(new_n833), .B2(new_n673), .ZN(new_n834));
  AND2_X1   g633(.A1(new_n834), .A2(new_n493), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n514), .A2(new_n501), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(new_n595), .ZN(new_n839));
  AND3_X1   g638(.A1(new_n838), .A2(G113gat), .A3(new_n839), .ZN(new_n840));
  AOI21_X1  g639(.A(G113gat), .B1(new_n838), .B2(new_n714), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n840), .A2(new_n841), .ZN(G1340gat));
  NOR2_X1   g641(.A1(new_n837), .A2(new_n639), .ZN(new_n843));
  XNOR2_X1  g642(.A(KEYINPUT119), .B(G120gat), .ZN(new_n844));
  XNOR2_X1  g643(.A(new_n843), .B(new_n844), .ZN(G1341gat));
  NAND2_X1  g644(.A1(new_n838), .A2(new_n673), .ZN(new_n846));
  XNOR2_X1  g645(.A(new_n846), .B(new_n388), .ZN(G1342gat));
  NOR2_X1   g646(.A1(new_n658), .A2(new_n514), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n501), .A2(G134gat), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n835), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  XOR2_X1   g649(.A(new_n850), .B(KEYINPUT56), .Z(new_n851));
  OAI21_X1  g650(.A(G134gat), .B1(new_n837), .B2(new_n658), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(G1343gat));
  NAND2_X1  g652(.A1(new_n732), .A2(new_n836), .ZN(new_n854));
  XNOR2_X1  g653(.A(new_n854), .B(KEYINPUT120), .ZN(new_n855));
  INV_X1    g654(.A(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n834), .A2(new_n486), .ZN(new_n857));
  XOR2_X1   g656(.A(KEYINPUT121), .B(KEYINPUT57), .Z(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  OAI211_X1 g658(.A(new_n828), .B(new_n820), .C1(new_n593), .C2(new_n594), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n657), .B1(new_n860), .B2(new_n830), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n672), .B1(new_n861), .B2(new_n829), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(new_n810), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n863), .A2(KEYINPUT57), .A3(new_n486), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n856), .B1(new_n859), .B2(new_n864), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n326), .B1(new_n865), .B2(new_n714), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n857), .A2(new_n695), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(new_n836), .ZN(new_n868));
  NOR3_X1   g667(.A1(new_n868), .A2(G141gat), .A3(new_n595), .ZN(new_n869));
  OAI21_X1  g668(.A(KEYINPUT58), .B1(new_n866), .B2(new_n869), .ZN(new_n870));
  OR2_X1    g669(.A1(new_n869), .A2(KEYINPUT58), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n326), .B1(new_n865), .B2(new_n839), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n870), .B1(new_n871), .B2(new_n872), .ZN(G1344gat));
  INV_X1    g672(.A(new_n858), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n834), .A2(new_n486), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n678), .A2(new_n595), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n373), .B1(new_n862), .B2(new_n876), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n875), .B1(new_n877), .B2(KEYINPUT57), .ZN(new_n878));
  INV_X1    g677(.A(new_n878), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n639), .B1(new_n856), .B2(KEYINPUT122), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n880), .B1(KEYINPUT122), .B2(new_n856), .ZN(new_n881));
  OAI211_X1 g680(.A(KEYINPUT59), .B(G148gat), .C1(new_n879), .C2(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n640), .A2(new_n328), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n328), .B1(new_n865), .B2(new_n640), .ZN(new_n884));
  OAI221_X1 g683(.A(new_n882), .B1(new_n868), .B2(new_n883), .C1(new_n884), .C2(KEYINPUT59), .ZN(G1345gat));
  NAND3_X1  g684(.A1(new_n867), .A2(new_n673), .A3(new_n836), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n673), .A2(G155gat), .ZN(new_n887));
  XNOR2_X1  g686(.A(new_n887), .B(KEYINPUT123), .ZN(new_n888));
  AOI22_X1  g687(.A1(new_n334), .A2(new_n886), .B1(new_n865), .B2(new_n888), .ZN(G1346gat));
  NAND4_X1  g688(.A1(new_n867), .A2(new_n335), .A3(new_n680), .A4(new_n848), .ZN(new_n890));
  AND2_X1   g689(.A1(new_n865), .A2(new_n657), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n890), .B1(new_n891), .B2(new_n335), .ZN(G1347gat));
  NOR4_X1   g691(.A1(new_n325), .A2(new_n486), .A3(new_n680), .A4(new_n492), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n834), .A2(new_n893), .ZN(new_n894));
  NOR3_X1   g693(.A1(new_n894), .A2(new_n203), .A3(new_n595), .ZN(new_n895));
  INV_X1    g694(.A(new_n894), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(new_n714), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n895), .B1(new_n203), .B2(new_n897), .ZN(G1348gat));
  NOR2_X1   g697(.A1(new_n894), .A2(new_n639), .ZN(new_n899));
  XNOR2_X1  g698(.A(new_n899), .B(new_n204), .ZN(G1349gat));
  NAND2_X1  g699(.A1(new_n896), .A2(new_n673), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(new_n217), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n902), .B1(new_n225), .B2(new_n901), .ZN(new_n903));
  XOR2_X1   g702(.A(new_n903), .B(KEYINPUT60), .Z(G1350gat));
  INV_X1    g703(.A(KEYINPUT124), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n894), .A2(new_n658), .ZN(new_n906));
  INV_X1    g705(.A(new_n906), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n905), .B1(new_n907), .B2(G190gat), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT61), .ZN(new_n909));
  AOI22_X1  g708(.A1(new_n908), .A2(new_n909), .B1(new_n224), .B2(new_n906), .ZN(new_n910));
  OR2_X1    g709(.A1(new_n908), .A2(new_n909), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n906), .A2(KEYINPUT124), .A3(new_n213), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n910), .B1(new_n911), .B2(new_n912), .ZN(G1351gat));
  NOR3_X1   g712(.A1(new_n695), .A2(new_n680), .A3(new_n325), .ZN(new_n914));
  AND3_X1   g713(.A1(new_n834), .A2(new_n486), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g714(.A(G197gat), .B1(new_n915), .B2(new_n714), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT125), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n878), .A2(new_n917), .ZN(new_n918));
  OAI211_X1 g717(.A(new_n875), .B(KEYINPUT125), .C1(new_n877), .C2(KEYINPUT57), .ZN(new_n919));
  AND3_X1   g718(.A1(new_n918), .A2(new_n914), .A3(new_n919), .ZN(new_n920));
  AND2_X1   g719(.A1(new_n839), .A2(G197gat), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n916), .B1(new_n920), .B2(new_n921), .ZN(G1352gat));
  XOR2_X1   g721(.A(KEYINPUT126), .B(G204gat), .Z(new_n923));
  NOR2_X1   g722(.A1(new_n639), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n915), .A2(new_n924), .ZN(new_n925));
  XOR2_X1   g724(.A(new_n925), .B(KEYINPUT62), .Z(new_n926));
  NAND4_X1  g725(.A1(new_n918), .A2(new_n640), .A3(new_n914), .A4(new_n919), .ZN(new_n927));
  AND2_X1   g726(.A1(new_n927), .A2(KEYINPUT127), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n923), .B1(new_n927), .B2(KEYINPUT127), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n926), .B1(new_n928), .B2(new_n929), .ZN(G1353gat));
  INV_X1    g729(.A(G211gat), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n915), .A2(new_n931), .A3(new_n673), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n914), .A2(new_n673), .ZN(new_n933));
  INV_X1    g732(.A(new_n933), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n931), .B1(new_n878), .B2(new_n934), .ZN(new_n935));
  AND2_X1   g734(.A1(new_n935), .A2(KEYINPUT63), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n935), .A2(KEYINPUT63), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n932), .B1(new_n936), .B2(new_n937), .ZN(G1354gat));
  AOI21_X1  g737(.A(G218gat), .B1(new_n915), .B2(new_n657), .ZN(new_n939));
  AND2_X1   g738(.A1(new_n657), .A2(G218gat), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n939), .B1(new_n920), .B2(new_n940), .ZN(G1355gat));
endmodule


