//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 0 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 1 1 1 1 1 1 0 0 1 1 1 1 1 0 0 0 1 0 0 1 1 1 0 1 1 1 0 0 1 1 1 0 1 1 0 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:48 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1210, new_n1211, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1258, new_n1259, new_n1260, new_n1261, new_n1262, new_n1263,
    new_n1264, new_n1265, new_n1266, new_n1267, new_n1268, new_n1269,
    new_n1270, new_n1271, new_n1272, new_n1273, new_n1274, new_n1275,
    new_n1276, new_n1277, new_n1278, new_n1279, new_n1280, new_n1281,
    new_n1282, new_n1283, new_n1284;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  NOR2_X1   g0003(.A1(G97), .A2(G107), .ZN(new_n204));
  INV_X1    g0004(.A(new_n204), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n205), .A2(G87), .ZN(G355));
  AOI22_X1  g0006(.A1(G68), .A2(G238), .B1(G97), .B2(G257), .ZN(new_n207));
  NAND2_X1  g0007(.A1(G116), .A2(G270), .ZN(new_n208));
  INV_X1    g0008(.A(G58), .ZN(new_n209));
  INV_X1    g0009(.A(G232), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n207), .B(new_n208), .C1(new_n209), .C2(new_n210), .ZN(new_n211));
  AOI21_X1  g0011(.A(new_n211), .B1(G50), .B2(G226), .ZN(new_n212));
  INV_X1    g0012(.A(G77), .ZN(new_n213));
  INV_X1    g0013(.A(G244), .ZN(new_n214));
  INV_X1    g0014(.A(G87), .ZN(new_n215));
  INV_X1    g0015(.A(G250), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n212), .B1(new_n213), .B2(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  AOI21_X1  g0017(.A(new_n217), .B1(G107), .B2(G264), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G20), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT64), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(KEYINPUT1), .ZN(new_n222));
  INV_X1    g0022(.A(G13), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n220), .A2(new_n223), .ZN(new_n224));
  INV_X1    g0024(.A(new_n224), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n225), .B(G250), .C1(G257), .C2(G264), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT65), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT0), .ZN(new_n228));
  AND2_X1   g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n229), .A2(G20), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n202), .A2(G50), .ZN(new_n231));
  OAI211_X1 g0031(.A(new_n222), .B(new_n228), .C1(new_n230), .C2(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT66), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(new_n210), .ZN(new_n235));
  XOR2_X1   g0035(.A(KEYINPUT2), .B(G226), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G250), .B(G257), .Z(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G68), .B(G77), .Z(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G58), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  INV_X1    g0048(.A(G20), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n249), .A2(G33), .A3(G116), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n249), .A2(G107), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n251), .B(KEYINPUT23), .ZN(new_n252));
  AND2_X1   g0052(.A1(KEYINPUT3), .A2(G33), .ZN(new_n253));
  NOR2_X1   g0053(.A1(KEYINPUT3), .A2(G33), .ZN(new_n254));
  OAI211_X1 g0054(.A(new_n249), .B(G87), .C1(new_n253), .C2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT22), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n256), .A2(KEYINPUT84), .ZN(new_n257));
  AND2_X1   g0057(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n255), .A2(new_n257), .ZN(new_n259));
  OAI211_X1 g0059(.A(new_n250), .B(new_n252), .C1(new_n258), .C2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT24), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g0062(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(G1), .A2(G13), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  XNOR2_X1  g0065(.A(new_n255), .B(new_n257), .ZN(new_n266));
  NAND4_X1  g0066(.A1(new_n266), .A2(KEYINPUT24), .A3(new_n250), .A4(new_n252), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n262), .A2(new_n265), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(KEYINPUT85), .A2(KEYINPUT25), .ZN(new_n269));
  INV_X1    g0069(.A(G1), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n270), .A2(G13), .A3(G20), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G107), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n269), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  OR2_X1    g0074(.A1(KEYINPUT85), .A2(KEYINPUT25), .ZN(new_n275));
  AND4_X1   g0075(.A1(new_n273), .A2(new_n272), .A3(new_n269), .A4(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(new_n265), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n270), .A2(G33), .ZN(new_n278));
  AND3_X1   g0078(.A1(new_n277), .A2(new_n271), .A3(new_n278), .ZN(new_n279));
  AOI211_X1 g0079(.A(new_n274), .B(new_n276), .C1(G107), .C2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n268), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G41), .ZN(new_n282));
  OAI211_X1 g0082(.A(new_n270), .B(G45), .C1(new_n282), .C2(KEYINPUT5), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n282), .A2(KEYINPUT5), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT67), .ZN(new_n286));
  AND2_X1   g0086(.A1(G33), .A2(G41), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n286), .B1(new_n287), .B2(new_n264), .ZN(new_n288));
  NAND2_X1  g0088(.A1(G33), .A2(G41), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n229), .A2(KEYINPUT67), .A3(new_n289), .ZN(new_n290));
  AOI22_X1  g0090(.A1(new_n284), .A2(new_n285), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G1698), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n216), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G257), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(G1698), .ZN(new_n295));
  OAI211_X1 g0095(.A(new_n293), .B(new_n295), .C1(new_n253), .C2(new_n254), .ZN(new_n296));
  INV_X1    g0096(.A(G33), .ZN(new_n297));
  INV_X1    g0097(.A(G294), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n296), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n229), .A2(new_n289), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  AOI22_X1  g0101(.A1(new_n291), .A2(G264), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(new_n285), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n303), .B1(new_n284), .B2(KEYINPUT78), .ZN(new_n304));
  INV_X1    g0104(.A(G274), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n305), .B1(new_n288), .B2(new_n290), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT78), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n283), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n304), .A2(new_n306), .A3(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n302), .A2(G179), .A3(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(G169), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n311), .B1(new_n302), .B2(new_n309), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n310), .B1(new_n312), .B2(KEYINPUT86), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n299), .A2(new_n301), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n288), .A2(new_n290), .ZN(new_n315));
  OAI211_X1 g0115(.A(new_n315), .B(G264), .C1(new_n283), .C2(new_n303), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n309), .A2(new_n314), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(G169), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT86), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n281), .B1(new_n313), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n279), .A2(G97), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n322), .B1(G97), .B2(new_n271), .ZN(new_n323));
  OR2_X1    g0123(.A1(KEYINPUT3), .A2(G33), .ZN(new_n324));
  NAND2_X1  g0124(.A1(KEYINPUT3), .A2(G33), .ZN(new_n325));
  NAND4_X1  g0125(.A1(new_n324), .A2(KEYINPUT7), .A3(new_n249), .A4(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT73), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n253), .A2(new_n254), .ZN(new_n329));
  NAND4_X1  g0129(.A1(new_n329), .A2(KEYINPUT73), .A3(KEYINPUT7), .A4(new_n249), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT7), .ZN(new_n331));
  XNOR2_X1  g0131(.A(KEYINPUT3), .B(G33), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n331), .B1(new_n332), .B2(G20), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n328), .A2(new_n330), .A3(new_n333), .ZN(new_n334));
  NOR2_X1   g0134(.A1(G20), .A2(G33), .ZN(new_n335));
  AOI22_X1  g0135(.A1(new_n334), .A2(G107), .B1(G77), .B2(new_n335), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n273), .A2(KEYINPUT6), .A3(G97), .ZN(new_n337));
  INV_X1    g0137(.A(G97), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n338), .A2(new_n273), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n339), .A2(new_n204), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n337), .B1(new_n340), .B2(KEYINPUT6), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(G20), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n336), .A2(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n323), .B1(new_n343), .B2(new_n265), .ZN(new_n344));
  OAI211_X1 g0144(.A(G244), .B(new_n292), .C1(new_n253), .C2(new_n254), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT4), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND4_X1  g0147(.A1(new_n332), .A2(KEYINPUT4), .A3(G244), .A4(new_n292), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n332), .A2(G250), .A3(G1698), .ZN(new_n349));
  NAND2_X1  g0149(.A1(G33), .A2(G283), .ZN(new_n350));
  NAND4_X1  g0150(.A1(new_n347), .A2(new_n348), .A3(new_n349), .A4(new_n350), .ZN(new_n351));
  AOI22_X1  g0151(.A1(new_n351), .A2(new_n301), .B1(G257), .B2(new_n291), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(new_n309), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n353), .A2(G190), .ZN(new_n354));
  AOI21_X1  g0154(.A(G200), .B1(new_n352), .B2(new_n309), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n344), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(G200), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n317), .A2(new_n357), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n358), .B1(G190), .B2(new_n317), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n359), .A2(new_n280), .A3(new_n268), .ZN(new_n360));
  AND3_X1   g0160(.A1(new_n352), .A2(G179), .A3(new_n309), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n311), .B1(new_n352), .B2(new_n309), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n277), .B1(new_n336), .B2(new_n342), .ZN(new_n363));
  OAI22_X1  g0163(.A1(new_n361), .A2(new_n362), .B1(new_n363), .B2(new_n323), .ZN(new_n364));
  AND4_X1   g0164(.A1(new_n321), .A2(new_n356), .A3(new_n360), .A4(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(G50), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n249), .B1(new_n201), .B2(new_n366), .ZN(new_n367));
  XNOR2_X1  g0167(.A(new_n367), .B(KEYINPUT69), .ZN(new_n368));
  INV_X1    g0168(.A(G150), .ZN(new_n369));
  INV_X1    g0169(.A(new_n335), .ZN(new_n370));
  OR2_X1    g0170(.A1(KEYINPUT8), .A2(G58), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT68), .ZN(new_n372));
  NAND2_X1  g0172(.A1(KEYINPUT8), .A2(G58), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n372), .B1(new_n371), .B2(new_n373), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n297), .A2(G20), .ZN(new_n378));
  INV_X1    g0178(.A(new_n378), .ZN(new_n379));
  OAI221_X1 g0179(.A(new_n368), .B1(new_n369), .B2(new_n370), .C1(new_n377), .C2(new_n379), .ZN(new_n380));
  AOI22_X1  g0180(.A1(new_n380), .A2(new_n265), .B1(new_n366), .B2(new_n272), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n263), .B(new_n264), .C1(G1), .C2(new_n249), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n381), .B1(new_n366), .B2(new_n382), .ZN(new_n383));
  XNOR2_X1  g0183(.A(new_n383), .B(KEYINPUT9), .ZN(new_n384));
  NOR2_X1   g0184(.A1(G222), .A2(G1698), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n292), .A2(G223), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n332), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  OAI211_X1 g0187(.A(new_n387), .B(new_n301), .C1(G77), .C2(new_n332), .ZN(new_n388));
  INV_X1    g0188(.A(G45), .ZN(new_n389));
  AOI21_X1  g0189(.A(G1), .B1(new_n282), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n306), .A2(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n390), .B1(new_n288), .B2(new_n290), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(G226), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n388), .A2(new_n391), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(G200), .ZN(new_n395));
  INV_X1    g0195(.A(G190), .ZN(new_n396));
  OR2_X1    g0196(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n384), .A2(new_n395), .A3(new_n397), .ZN(new_n398));
  XNOR2_X1  g0198(.A(new_n398), .B(KEYINPUT10), .ZN(new_n399));
  INV_X1    g0199(.A(G226), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(new_n292), .ZN(new_n401));
  OAI211_X1 g0201(.A(new_n332), .B(new_n401), .C1(G232), .C2(new_n292), .ZN(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n297), .A2(new_n338), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n301), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n392), .A2(G238), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n405), .A2(new_n391), .A3(new_n406), .ZN(new_n407));
  OR2_X1    g0207(.A1(new_n407), .A2(KEYINPUT13), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n407), .A2(KEYINPUT13), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(G169), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT14), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n412), .A2(KEYINPUT72), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(new_n410), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(G179), .ZN(new_n416));
  OAI211_X1 g0216(.A(new_n410), .B(G169), .C1(KEYINPUT72), .C2(new_n412), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n414), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  OAI22_X1  g0218(.A1(new_n379), .A2(new_n213), .B1(new_n249), .B2(G68), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n370), .A2(new_n366), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n265), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  XNOR2_X1  g0221(.A(new_n421), .B(KEYINPUT11), .ZN(new_n422));
  INV_X1    g0222(.A(G68), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n272), .A2(new_n423), .ZN(new_n424));
  AND2_X1   g0224(.A1(new_n424), .A2(KEYINPUT12), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n424), .A2(KEYINPUT12), .ZN(new_n426));
  OAI221_X1 g0226(.A(new_n422), .B1(new_n423), .B2(new_n382), .C1(new_n425), .C2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT71), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n428), .B1(new_n410), .B2(G200), .ZN(new_n429));
  AOI211_X1 g0229(.A(KEYINPUT71), .B(new_n357), .C1(new_n408), .C2(new_n409), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n427), .B1(new_n415), .B2(G190), .ZN(new_n432));
  AOI22_X1  g0232(.A1(new_n418), .A2(new_n427), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n394), .A2(new_n311), .ZN(new_n434));
  OR2_X1    g0234(.A1(new_n394), .A2(G179), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n383), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n332), .A2(G232), .A3(new_n292), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n332), .A2(G238), .A3(G1698), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n437), .B(new_n438), .C1(new_n273), .C2(new_n332), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(new_n301), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n392), .A2(G244), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n440), .A2(new_n391), .A3(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT70), .ZN(new_n443));
  OR2_X1    g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n442), .A2(new_n443), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(G190), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n444), .A2(G200), .A3(new_n445), .ZN(new_n448));
  NAND2_X1  g0248(.A1(G20), .A2(G77), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n371), .A2(new_n373), .ZN(new_n450));
  XOR2_X1   g0250(.A(KEYINPUT15), .B(G87), .Z(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  OAI221_X1 g0252(.A(new_n449), .B1(new_n370), .B2(new_n450), .C1(new_n452), .C2(new_n379), .ZN(new_n453));
  AOI22_X1  g0253(.A1(new_n453), .A2(new_n265), .B1(new_n213), .B2(new_n272), .ZN(new_n454));
  OR2_X1    g0254(.A1(new_n382), .A2(new_n213), .ZN(new_n455));
  AND2_X1   g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n447), .A2(new_n448), .A3(new_n456), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n399), .A2(new_n433), .A3(new_n436), .A4(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT77), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n382), .B1(new_n375), .B2(new_n376), .ZN(new_n460));
  INV_X1    g0260(.A(new_n376), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n461), .A2(new_n271), .A3(new_n374), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT74), .ZN(new_n463));
  AND3_X1   g0263(.A1(new_n460), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n463), .B1(new_n460), .B2(new_n462), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n209), .A2(new_n423), .ZN(new_n467));
  OAI21_X1  g0267(.A(G20), .B1(new_n467), .B2(new_n201), .ZN(new_n468));
  INV_X1    g0268(.A(G159), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n468), .B1(new_n469), .B2(new_n370), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n470), .B1(new_n334), .B2(G68), .ZN(new_n471));
  OR2_X1    g0271(.A1(new_n471), .A2(KEYINPUT16), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n333), .A2(new_n326), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n470), .B1(new_n473), .B2(G68), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n277), .B1(new_n474), .B2(KEYINPUT16), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n466), .B1(new_n472), .B2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(G223), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(new_n292), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n400), .A2(G1698), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n478), .B(new_n479), .C1(new_n253), .C2(new_n254), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n480), .B1(new_n297), .B2(new_n215), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(new_n301), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n392), .A2(G232), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n482), .A2(new_n391), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(KEYINPUT75), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT75), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n482), .A2(new_n391), .A3(new_n483), .A4(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n485), .A2(new_n357), .A3(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(new_n484), .ZN(new_n489));
  OR2_X1    g0289(.A1(new_n396), .A2(KEYINPUT76), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n396), .A2(KEYINPUT76), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n488), .A2(new_n493), .ZN(new_n494));
  AND3_X1   g0294(.A1(new_n476), .A2(new_n494), .A3(KEYINPUT17), .ZN(new_n495));
  AOI21_X1  g0295(.A(KEYINPUT17), .B1(new_n476), .B2(new_n494), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n459), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n476), .A2(new_n494), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT17), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n476), .A2(new_n494), .A3(KEYINPUT17), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n500), .A2(KEYINPUT77), .A3(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(new_n476), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n485), .A2(new_n311), .A3(new_n487), .ZN(new_n504));
  INV_X1    g0304(.A(G179), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n489), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n503), .A2(new_n508), .A3(KEYINPUT18), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT18), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n510), .B1(new_n476), .B2(new_n507), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n497), .A2(new_n502), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n446), .A2(new_n505), .ZN(new_n514));
  INV_X1    g0314(.A(new_n456), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n444), .A2(new_n311), .A3(new_n445), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(new_n517), .ZN(new_n518));
  OR2_X1    g0318(.A1(new_n513), .A2(new_n518), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n458), .A2(new_n519), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n451), .A2(new_n271), .ZN(new_n521));
  INV_X1    g0321(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n279), .A2(new_n451), .ZN(new_n523));
  AOI21_X1  g0323(.A(G20), .B1(new_n404), .B2(KEYINPUT19), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT80), .ZN(new_n525));
  XNOR2_X1  g0325(.A(KEYINPUT79), .B(G87), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n525), .B1(new_n526), .B2(new_n205), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT79), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n528), .A2(G87), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n215), .A2(KEYINPUT79), .ZN(new_n530));
  OAI211_X1 g0330(.A(KEYINPUT80), .B(new_n204), .C1(new_n529), .C2(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n524), .B1(new_n527), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n332), .A2(new_n249), .A3(G68), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  AOI21_X1  g0334(.A(KEYINPUT19), .B1(new_n378), .B2(G97), .ZN(new_n535));
  NOR3_X1   g0335(.A1(new_n532), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n522), .B(new_n523), .C1(new_n536), .C2(new_n277), .ZN(new_n537));
  OR2_X1    g0337(.A1(G238), .A2(G1698), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n214), .A2(G1698), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n538), .B(new_n539), .C1(new_n253), .C2(new_n254), .ZN(new_n540));
  NAND2_X1  g0340(.A1(G33), .A2(G116), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(new_n301), .ZN(new_n543));
  AOI21_X1  g0343(.A(G250), .B1(new_n270), .B2(G45), .ZN(new_n544));
  INV_X1    g0344(.A(new_n544), .ZN(new_n545));
  NOR3_X1   g0345(.A1(new_n389), .A2(G1), .A3(G274), .ZN(new_n546));
  INV_X1    g0346(.A(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n315), .A2(new_n545), .A3(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n543), .A2(new_n548), .A3(new_n505), .ZN(new_n549));
  AOI211_X1 g0349(.A(new_n544), .B(new_n546), .C1(new_n288), .C2(new_n290), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n300), .B1(new_n540), .B2(new_n541), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n549), .B1(new_n552), .B2(G169), .ZN(new_n553));
  INV_X1    g0353(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n537), .A2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT81), .ZN(new_n556));
  NOR3_X1   g0356(.A1(new_n550), .A2(new_n551), .A3(new_n396), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n357), .B1(new_n543), .B2(new_n548), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(new_n524), .ZN(new_n560));
  NOR3_X1   g0360(.A1(new_n526), .A2(new_n525), .A3(new_n205), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n215), .A2(KEYINPUT79), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n528), .A2(G87), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AOI21_X1  g0364(.A(KEYINPUT80), .B1(new_n564), .B2(new_n204), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n560), .B1(new_n561), .B2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(new_n535), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n566), .A2(new_n533), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n265), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n279), .A2(G87), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n559), .A2(new_n569), .A3(new_n570), .A4(new_n522), .ZN(new_n571));
  AND3_X1   g0371(.A1(new_n555), .A2(new_n556), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n556), .B1(new_n555), .B2(new_n571), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n315), .B(G270), .C1(new_n283), .C2(new_n303), .ZN(new_n575));
  AND2_X1   g0375(.A1(new_n309), .A2(new_n575), .ZN(new_n576));
  OAI211_X1 g0376(.A(G264), .B(G1698), .C1(new_n253), .C2(new_n254), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT82), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n332), .A2(KEYINPUT82), .A3(G264), .A4(G1698), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n332), .A2(G257), .A3(new_n292), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n329), .A2(G303), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n301), .B1(new_n581), .B2(new_n584), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n277), .A2(G116), .A3(new_n271), .A4(new_n278), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n271), .A2(G116), .ZN(new_n587));
  INV_X1    g0387(.A(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(G116), .ZN(new_n589));
  AOI22_X1  g0389(.A1(new_n263), .A2(new_n264), .B1(G20), .B2(new_n589), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n350), .B(new_n249), .C1(G33), .C2(new_n338), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n590), .A2(KEYINPUT20), .A3(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(new_n592), .ZN(new_n593));
  AOI21_X1  g0393(.A(KEYINPUT20), .B1(new_n590), .B2(new_n591), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n586), .B(new_n588), .C1(new_n593), .C2(new_n594), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n576), .A2(G179), .A3(new_n585), .A4(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n585), .A2(new_n309), .A3(new_n575), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n590), .A2(new_n591), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT20), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n587), .B1(new_n600), .B2(new_n592), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n311), .B1(new_n601), .B2(new_n586), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT21), .ZN(new_n603));
  AND3_X1   g0403(.A1(new_n597), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n603), .B1(new_n597), .B2(new_n602), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n596), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(new_n492), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n585), .A2(new_n309), .A3(new_n575), .A4(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(new_n595), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n357), .B1(new_n576), .B2(new_n585), .ZN(new_n611));
  OAI21_X1  g0411(.A(KEYINPUT83), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n597), .A2(G200), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT83), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n613), .A2(new_n614), .A3(new_n609), .A4(new_n608), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n606), .B1(new_n612), .B2(new_n615), .ZN(new_n616));
  AND4_X1   g0416(.A1(new_n365), .A2(new_n520), .A3(new_n574), .A4(new_n616), .ZN(G372));
  OAI211_X1 g0417(.A(new_n570), .B(new_n522), .C1(new_n536), .C2(new_n277), .ZN(new_n618));
  INV_X1    g0418(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n558), .A2(KEYINPUT87), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n543), .A2(new_n548), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(G200), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT87), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n557), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n619), .A2(new_n620), .A3(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n521), .B1(new_n568), .B2(new_n265), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n553), .B1(new_n627), .B2(new_n523), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  AND3_X1   g0429(.A1(new_n356), .A2(new_n364), .A3(new_n360), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n317), .A2(new_n505), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n631), .B1(new_n319), .B2(new_n318), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n312), .A2(KEYINPUT86), .ZN(new_n633));
  AOI22_X1  g0433(.A1(new_n632), .A2(new_n633), .B1(new_n280), .B2(new_n268), .ZN(new_n634));
  OAI211_X1 g0434(.A(new_n629), .B(new_n630), .C1(new_n634), .C2(new_n606), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n361), .A2(new_n362), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT88), .ZN(new_n637));
  XNOR2_X1  g0437(.A(new_n636), .B(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT26), .ZN(new_n639));
  INV_X1    g0439(.A(new_n344), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n629), .A2(new_n638), .A3(new_n639), .A4(new_n640), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n622), .B1(new_n396), .B2(new_n621), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n618), .A2(new_n642), .ZN(new_n643));
  OAI21_X1  g0443(.A(KEYINPUT81), .B1(new_n643), .B2(new_n628), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n555), .A2(new_n571), .A3(new_n556), .ZN(new_n645));
  INV_X1    g0445(.A(new_n364), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n644), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n628), .B1(new_n647), .B2(KEYINPUT26), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n635), .A2(new_n641), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n520), .A2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n436), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n418), .A2(new_n427), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n517), .B1(new_n431), .B2(new_n432), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n497), .A2(new_n502), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n512), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n651), .B1(new_n657), .B2(new_n399), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n650), .A2(new_n658), .ZN(G369));
  INV_X1    g0459(.A(KEYINPUT90), .ZN(new_n660));
  XOR2_X1   g0460(.A(KEYINPUT89), .B(KEYINPUT27), .Z(new_n661));
  NOR3_X1   g0461(.A1(new_n223), .A2(G1), .A3(G20), .ZN(new_n662));
  OR2_X1    g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n661), .A2(new_n662), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n663), .A2(G213), .A3(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(G343), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n616), .B1(new_n609), .B2(new_n668), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n668), .A2(new_n609), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n606), .A2(new_n670), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n660), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  AOI21_X1  g0472(.A(KEYINPUT90), .B1(new_n606), .B2(new_n670), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  AND2_X1   g0475(.A1(new_n321), .A2(new_n360), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n281), .A2(new_n667), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n678), .B1(new_n321), .B2(new_n668), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n675), .A2(G330), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n634), .A2(new_n668), .ZN(new_n681));
  INV_X1    g0481(.A(new_n596), .ZN(new_n682));
  INV_X1    g0482(.A(new_n605), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n597), .A2(new_n602), .A3(new_n603), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n682), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n685), .A2(new_n667), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(new_n676), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n680), .A2(new_n681), .A3(new_n687), .ZN(G399));
  NOR2_X1   g0488(.A1(new_n224), .A2(G41), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(G1), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n527), .A2(new_n589), .A3(new_n531), .ZN(new_n692));
  OAI22_X1  g0492(.A1(new_n691), .A2(new_n692), .B1(new_n231), .B2(new_n690), .ZN(new_n693));
  XNOR2_X1  g0493(.A(new_n693), .B(KEYINPUT28), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n365), .A2(new_n616), .A3(new_n574), .A4(new_n668), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT91), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n612), .A2(new_n615), .ZN(new_n698));
  AND4_X1   g0498(.A1(new_n645), .A2(new_n644), .A3(new_n685), .A4(new_n698), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n699), .A2(KEYINPUT91), .A3(new_n365), .A4(new_n668), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT30), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n631), .A2(new_n352), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n576), .A2(new_n552), .A3(new_n585), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n702), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n597), .A2(new_n621), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n706), .A2(KEYINPUT30), .A3(new_n631), .A4(new_n352), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n552), .A2(G179), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n353), .A2(new_n708), .A3(new_n317), .A4(new_n597), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n705), .A2(new_n707), .A3(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT31), .ZN(new_n711));
  AND3_X1   g0511(.A1(new_n710), .A2(new_n711), .A3(new_n667), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n711), .B1(new_n710), .B2(new_n667), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n701), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(G330), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT29), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n649), .A2(new_n719), .A3(new_n668), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n647), .A2(new_n639), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(KEYINPUT92), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n629), .A2(new_n638), .A3(KEYINPUT26), .A4(new_n640), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT92), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n647), .A2(new_n724), .A3(new_n639), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n722), .A2(new_n723), .A3(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(KEYINPUT93), .B1(new_n634), .B2(new_n606), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT93), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n685), .A2(new_n728), .A3(new_n321), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n626), .B1(new_n727), .B2(new_n729), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n628), .B1(new_n730), .B2(new_n630), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n667), .B1(new_n726), .B2(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n720), .B1(new_n732), .B2(new_n719), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n718), .A2(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n694), .B1(new_n734), .B2(G1), .ZN(G364));
  NOR3_X1   g0535(.A1(new_n223), .A2(new_n389), .A3(G20), .ZN(new_n736));
  OR2_X1    g0536(.A1(new_n736), .A2(KEYINPUT94), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n736), .A2(KEYINPUT94), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n737), .A2(G1), .A3(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n689), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n249), .A2(new_n505), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(G200), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(G190), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  OR2_X1    g0545(.A1(KEYINPUT33), .A2(G317), .ZN(new_n746));
  NAND2_X1  g0546(.A1(KEYINPUT33), .A2(G317), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n745), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n357), .A2(G190), .ZN(new_n749));
  OAI21_X1  g0549(.A(G20), .B1(new_n749), .B2(G179), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT96), .ZN(new_n751));
  OR2_X1    g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n750), .A2(new_n751), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n249), .A2(G179), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n756), .A2(new_n396), .A3(G200), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  AOI22_X1  g0558(.A1(new_n755), .A2(G294), .B1(G283), .B2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n492), .A2(new_n743), .ZN(new_n760));
  XNOR2_X1  g0560(.A(KEYINPUT97), .B(G326), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(G311), .ZN(new_n763));
  NOR2_X1   g0563(.A1(G190), .A2(G200), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n742), .A2(new_n764), .ZN(new_n765));
  OAI211_X1 g0565(.A(new_n759), .B(new_n762), .C1(new_n763), .C2(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n756), .A2(new_n764), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  AOI211_X1 g0568(.A(new_n748), .B(new_n766), .C1(G329), .C2(new_n768), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n756), .A2(G190), .A3(G200), .ZN(new_n770));
  INV_X1    g0570(.A(G303), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n329), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  XNOR2_X1  g0572(.A(new_n772), .B(KEYINPUT98), .ZN(new_n773));
  INV_X1    g0573(.A(G322), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n607), .A2(new_n357), .A3(new_n742), .ZN(new_n775));
  OAI211_X1 g0575(.A(new_n769), .B(new_n773), .C1(new_n774), .C2(new_n775), .ZN(new_n776));
  XOR2_X1   g0576(.A(new_n776), .B(KEYINPUT99), .Z(new_n777));
  NOR2_X1   g0577(.A1(new_n775), .A2(new_n209), .ZN(new_n778));
  AOI22_X1  g0578(.A1(new_n755), .A2(G97), .B1(G50), .B2(new_n760), .ZN(new_n779));
  OAI22_X1  g0579(.A1(new_n745), .A2(new_n423), .B1(new_n765), .B2(new_n213), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n767), .A2(new_n469), .ZN(new_n781));
  INV_X1    g0581(.A(KEYINPUT32), .ZN(new_n782));
  OAI22_X1  g0582(.A1(new_n781), .A2(new_n782), .B1(new_n564), .B2(new_n770), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n780), .A2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n757), .A2(new_n273), .ZN(new_n785));
  AOI211_X1 g0585(.A(new_n329), .B(new_n785), .C1(new_n782), .C2(new_n781), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n779), .A2(new_n784), .A3(new_n786), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n777), .B1(new_n778), .B2(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n264), .B1(G20), .B2(new_n311), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n741), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n224), .A2(new_n329), .ZN(new_n791));
  XNOR2_X1  g0591(.A(new_n791), .B(KEYINPUT95), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(G355), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n231), .A2(G45), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n224), .A2(new_n332), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n795), .B1(new_n247), .B2(new_n389), .ZN(new_n796));
  OAI221_X1 g0596(.A(new_n793), .B1(G116), .B2(new_n225), .C1(new_n794), .C2(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(G13), .A2(G33), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n799), .A2(G20), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n800), .A2(new_n789), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n797), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n800), .ZN(new_n803));
  OAI211_X1 g0603(.A(new_n790), .B(new_n802), .C1(new_n675), .C2(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n675), .A2(G330), .ZN(new_n805));
  INV_X1    g0605(.A(G330), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n674), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n805), .A2(new_n741), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n804), .A2(new_n808), .ZN(G396));
  NAND2_X1  g0609(.A1(new_n649), .A2(new_n668), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n517), .A2(new_n667), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n457), .B1(new_n456), .B2(new_n668), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n811), .B1(new_n812), .B2(new_n517), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n810), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n649), .A2(new_n668), .A3(new_n813), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  XNOR2_X1  g0617(.A(new_n718), .B(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n818), .A2(new_n741), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n814), .A2(new_n798), .ZN(new_n820));
  INV_X1    g0620(.A(new_n775), .ZN(new_n821));
  INV_X1    g0621(.A(new_n765), .ZN(new_n822));
  AOI22_X1  g0622(.A1(new_n821), .A2(G143), .B1(G159), .B2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(G137), .ZN(new_n824));
  INV_X1    g0624(.A(new_n760), .ZN(new_n825));
  OAI221_X1 g0625(.A(new_n823), .B1(new_n824), .B2(new_n825), .C1(new_n369), .C2(new_n745), .ZN(new_n826));
  XNOR2_X1  g0626(.A(new_n826), .B(KEYINPUT34), .ZN(new_n827));
  INV_X1    g0627(.A(G132), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n332), .B1(new_n767), .B2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n770), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n829), .B1(G50), .B2(new_n830), .ZN(new_n831));
  OAI211_X1 g0631(.A(new_n827), .B(new_n831), .C1(new_n423), .C2(new_n757), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n754), .A2(new_n209), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n757), .A2(new_n215), .ZN(new_n834));
  AOI22_X1  g0634(.A1(new_n755), .A2(G97), .B1(G107), .B2(new_n830), .ZN(new_n835));
  INV_X1    g0635(.A(G283), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n835), .B1(new_n836), .B2(new_n745), .C1(new_n298), .C2(new_n775), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n765), .A2(new_n589), .ZN(new_n838));
  OAI22_X1  g0638(.A1(new_n825), .A2(new_n771), .B1(new_n763), .B2(new_n767), .ZN(new_n839));
  OR4_X1    g0639(.A1(new_n834), .A2(new_n837), .A3(new_n838), .A4(new_n839), .ZN(new_n840));
  OAI22_X1  g0640(.A1(new_n832), .A2(new_n833), .B1(new_n840), .B2(new_n332), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(new_n789), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n789), .A2(new_n798), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(new_n213), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n820), .A2(new_n740), .A3(new_n842), .A4(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n819), .A2(new_n845), .ZN(G384));
  OAI211_X1 g0646(.A(G20), .B(new_n229), .C1(new_n341), .C2(KEYINPUT35), .ZN(new_n847));
  AOI211_X1 g0647(.A(new_n589), .B(new_n847), .C1(KEYINPUT35), .C2(new_n341), .ZN(new_n848));
  XOR2_X1   g0648(.A(new_n848), .B(KEYINPUT36), .Z(new_n849));
  OAI21_X1  g0649(.A(G77), .B1(new_n209), .B2(new_n423), .ZN(new_n850));
  OAI22_X1  g0650(.A1(new_n231), .A2(new_n850), .B1(G50), .B2(new_n423), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n851), .A2(G1), .A3(new_n223), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n427), .A2(new_n667), .ZN(new_n853));
  AOI22_X1  g0653(.A1(new_n653), .A2(new_n667), .B1(new_n433), .B2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(KEYINPUT100), .B1(new_n701), .B2(new_n715), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT100), .ZN(new_n857));
  AOI211_X1 g0657(.A(new_n857), .B(new_n714), .C1(new_n697), .C2(new_n700), .ZN(new_n858));
  OAI211_X1 g0658(.A(new_n813), .B(new_n855), .C1(new_n856), .C2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT38), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n503), .A2(new_n508), .ZN(new_n861));
  INV_X1    g0661(.A(new_n665), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n503), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n861), .A2(new_n863), .A3(new_n498), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT37), .ZN(new_n865));
  XNOR2_X1  g0665(.A(new_n864), .B(new_n865), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n495), .A2(new_n496), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n863), .B1(new_n512), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n860), .B1(new_n866), .B2(new_n868), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n475), .B1(KEYINPUT16), .B2(new_n474), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n870), .B1(new_n465), .B2(new_n464), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n513), .A2(new_n862), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n507), .A2(new_n665), .ZN(new_n873));
  AOI22_X1  g0673(.A1(new_n873), .A2(new_n871), .B1(new_n476), .B2(new_n494), .ZN(new_n874));
  OR2_X1    g0674(.A1(new_n874), .A2(new_n865), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n875), .B1(KEYINPUT37), .B2(new_n864), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n872), .A2(KEYINPUT38), .A3(new_n876), .ZN(new_n877));
  AND2_X1   g0677(.A1(new_n869), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g0678(.A(KEYINPUT40), .B1(new_n859), .B2(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n714), .B1(new_n697), .B2(new_n700), .ZN(new_n880));
  XNOR2_X1  g0680(.A(new_n880), .B(KEYINPUT100), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n872), .A2(new_n876), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(new_n860), .ZN(new_n883));
  AOI21_X1  g0683(.A(KEYINPUT40), .B1(new_n883), .B2(new_n877), .ZN(new_n884));
  NAND4_X1  g0684(.A1(new_n881), .A2(new_n884), .A3(new_n813), .A4(new_n855), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n879), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(G330), .ZN(new_n887));
  AND2_X1   g0687(.A1(new_n881), .A2(new_n520), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(G330), .ZN(new_n889));
  AOI22_X1  g0689(.A1(new_n887), .A2(new_n889), .B1(new_n886), .B2(new_n888), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n509), .A2(new_n511), .A3(new_n665), .ZN(new_n891));
  INV_X1    g0691(.A(new_n811), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n854), .B1(new_n816), .B2(new_n892), .ZN(new_n893));
  AND3_X1   g0693(.A1(new_n872), .A2(KEYINPUT38), .A3(new_n876), .ZN(new_n894));
  AOI21_X1  g0694(.A(KEYINPUT38), .B1(new_n872), .B2(new_n876), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n893), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT39), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n897), .B1(new_n883), .B2(new_n877), .ZN(new_n898));
  AND3_X1   g0698(.A1(new_n869), .A2(new_n877), .A3(new_n897), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n652), .A2(new_n667), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n891), .B(new_n896), .C1(new_n900), .C2(new_n902), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n890), .B(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n520), .A2(new_n733), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(new_n658), .ZN(new_n906));
  XOR2_X1   g0706(.A(new_n904), .B(new_n906), .Z(new_n907));
  AOI21_X1  g0707(.A(new_n270), .B1(G13), .B2(new_n249), .ZN(new_n908));
  OAI211_X1 g0708(.A(new_n849), .B(new_n852), .C1(new_n907), .C2(new_n908), .ZN(G367));
  NAND3_X1  g0709(.A1(new_n638), .A2(new_n640), .A3(new_n667), .ZN(new_n910));
  OAI211_X1 g0710(.A(new_n356), .B(new_n364), .C1(new_n344), .C2(new_n668), .ZN(new_n911));
  AND2_X1   g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n687), .A2(new_n681), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  XOR2_X1   g0714(.A(new_n914), .B(KEYINPUT44), .Z(new_n915));
  NOR2_X1   g0715(.A1(new_n912), .A2(new_n913), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n916), .B(KEYINPUT45), .ZN(new_n917));
  AND2_X1   g0717(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(KEYINPUT103), .B1(new_n918), .B2(new_n680), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n915), .A2(new_n917), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n920), .B(new_n680), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n919), .B1(new_n921), .B2(KEYINPUT103), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n687), .B1(new_n679), .B2(new_n686), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n805), .B(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n734), .B1(new_n922), .B2(new_n924), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n689), .B(KEYINPUT41), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT104), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(new_n739), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n925), .A2(KEYINPUT104), .A3(new_n926), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n929), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n364), .B1(new_n912), .B2(new_n321), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(new_n668), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n365), .A2(new_n686), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(KEYINPUT42), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT101), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n937), .B(new_n938), .ZN(new_n939));
  OR2_X1    g0739(.A1(new_n935), .A2(KEYINPUT42), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n629), .B1(new_n619), .B2(new_n668), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n628), .A2(new_n618), .A3(new_n667), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  AOI22_X1  g0743(.A1(new_n939), .A2(new_n940), .B1(KEYINPUT43), .B2(new_n943), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n943), .A2(KEYINPUT43), .ZN(new_n945));
  OR2_X1    g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n944), .A2(new_n945), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(new_n680), .B2(new_n912), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n680), .A2(new_n912), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n946), .A2(new_n950), .A3(new_n947), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(KEYINPUT102), .ZN(new_n952));
  OR2_X1    g0752(.A1(new_n951), .A2(KEYINPUT102), .ZN(new_n953));
  NAND4_X1  g0753(.A1(new_n932), .A2(new_n949), .A3(new_n952), .A4(new_n953), .ZN(new_n954));
  AOI22_X1  g0754(.A1(new_n821), .A2(G303), .B1(G311), .B2(new_n760), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n755), .A2(G107), .ZN(new_n956));
  OAI21_X1  g0756(.A(KEYINPUT105), .B1(new_n770), .B2(new_n589), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n957), .A2(KEYINPUT46), .ZN(new_n958));
  OR2_X1    g0758(.A1(new_n957), .A2(KEYINPUT46), .ZN(new_n959));
  NAND4_X1  g0759(.A1(new_n955), .A2(new_n956), .A3(new_n958), .A4(new_n959), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n757), .A2(new_n338), .ZN(new_n961));
  AOI211_X1 g0761(.A(new_n332), .B(new_n961), .C1(G317), .C2(new_n768), .ZN(new_n962));
  XOR2_X1   g0762(.A(new_n962), .B(KEYINPUT106), .Z(new_n963));
  AOI211_X1 g0763(.A(new_n960), .B(new_n963), .C1(G283), .C2(new_n822), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n744), .A2(G294), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n755), .A2(G68), .ZN(new_n966));
  AOI22_X1  g0766(.A1(new_n760), .A2(G143), .B1(G137), .B2(new_n768), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n967), .B1(new_n369), .B2(new_n775), .ZN(new_n968));
  AOI22_X1  g0768(.A1(new_n744), .A2(G159), .B1(new_n822), .B2(G50), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n969), .B1(new_n209), .B2(new_n770), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n332), .B1(new_n757), .B2(new_n213), .ZN(new_n971));
  NOR3_X1   g0771(.A1(new_n968), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  AOI22_X1  g0772(.A1(new_n964), .A2(new_n965), .B1(new_n966), .B2(new_n972), .ZN(new_n973));
  XOR2_X1   g0773(.A(new_n973), .B(KEYINPUT47), .Z(new_n974));
  NAND2_X1  g0774(.A1(new_n974), .A2(new_n789), .ZN(new_n975));
  INV_X1    g0775(.A(new_n943), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(new_n800), .ZN(new_n977));
  INV_X1    g0777(.A(new_n795), .ZN(new_n978));
  OAI221_X1 g0778(.A(new_n801), .B1(new_n225), .B2(new_n452), .C1(new_n978), .C2(new_n240), .ZN(new_n979));
  NAND4_X1  g0779(.A1(new_n975), .A2(new_n740), .A3(new_n977), .A4(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n954), .A2(new_n980), .ZN(G387));
  NOR2_X1   g0781(.A1(new_n924), .A2(new_n930), .ZN(new_n982));
  INV_X1    g0782(.A(new_n789), .ZN(new_n983));
  AOI22_X1  g0783(.A1(new_n760), .A2(G322), .B1(new_n744), .B2(G311), .ZN(new_n984));
  INV_X1    g0784(.A(G317), .ZN(new_n985));
  OAI221_X1 g0785(.A(new_n984), .B1(new_n771), .B2(new_n765), .C1(new_n985), .C2(new_n775), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n986), .B(KEYINPUT48), .ZN(new_n987));
  OAI221_X1 g0787(.A(new_n987), .B1(new_n836), .B2(new_n754), .C1(new_n298), .C2(new_n770), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n988), .B(KEYINPUT108), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(KEYINPUT49), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n758), .A2(G116), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n768), .A2(new_n761), .ZN(new_n992));
  NAND4_X1  g0792(.A1(new_n990), .A2(new_n329), .A3(new_n991), .A4(new_n992), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n775), .A2(new_n366), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n754), .A2(new_n452), .ZN(new_n995));
  AOI211_X1 g0795(.A(new_n994), .B(new_n995), .C1(G159), .C2(new_n760), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n744), .B1(new_n375), .B2(new_n376), .ZN(new_n997));
  OAI22_X1  g0797(.A1(new_n765), .A2(new_n423), .B1(new_n767), .B2(new_n369), .ZN(new_n998));
  AOI211_X1 g0798(.A(new_n961), .B(new_n998), .C1(G77), .C2(new_n830), .ZN(new_n999));
  NAND4_X1  g0799(.A1(new_n996), .A2(new_n332), .A3(new_n997), .A4(new_n999), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n983), .B1(new_n993), .B2(new_n1000), .ZN(new_n1001));
  NOR3_X1   g0801(.A1(new_n450), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n692), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(G68), .A2(G77), .ZN(new_n1004));
  OAI21_X1  g0804(.A(KEYINPUT50), .B1(new_n450), .B2(G50), .ZN(new_n1005));
  NAND4_X1  g0805(.A1(new_n1003), .A2(new_n389), .A3(new_n1004), .A4(new_n1005), .ZN(new_n1006));
  OAI211_X1 g0806(.A(new_n1006), .B(new_n795), .C1(new_n237), .C2(new_n389), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1007), .B1(G107), .B2(new_n225), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1008), .B1(new_n692), .B2(new_n792), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(KEYINPUT107), .ZN(new_n1010));
  AOI211_X1 g0810(.A(new_n741), .B(new_n1001), .C1(new_n801), .C2(new_n1010), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1011), .B(KEYINPUT109), .ZN(new_n1012));
  OR2_X1    g0812(.A1(new_n679), .A2(new_n803), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n982), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n734), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n1015), .A2(new_n924), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n690), .B1(new_n1015), .B2(new_n924), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1014), .A2(new_n1019), .ZN(G393));
  OR2_X1    g0820(.A1(new_n921), .A2(new_n1016), .ZN(new_n1021));
  OAI211_X1 g0821(.A(new_n1021), .B(new_n689), .C1(new_n922), .C2(new_n1017), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n921), .A2(new_n739), .ZN(new_n1023));
  INV_X1    g0823(.A(KEYINPUT111), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n801), .B1(new_n338), .B2(new_n225), .C1(new_n978), .C2(new_n244), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n469), .A2(new_n775), .B1(new_n825), .B2(new_n369), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT51), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n744), .A2(G50), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n755), .A2(G77), .B1(G143), .B2(new_n768), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n332), .B1(new_n765), .B2(new_n450), .ZN(new_n1030));
  AOI211_X1 g0830(.A(new_n834), .B(new_n1030), .C1(G68), .C2(new_n830), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n1027), .A2(new_n1028), .A3(new_n1029), .A4(new_n1031), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n763), .A2(new_n775), .B1(new_n825), .B2(new_n985), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT52), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n755), .A2(G116), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n329), .B1(new_n765), .B2(new_n298), .ZN(new_n1036));
  AOI211_X1 g0836(.A(new_n785), .B(new_n1036), .C1(G303), .C2(new_n744), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n770), .A2(new_n836), .B1(new_n767), .B2(new_n774), .ZN(new_n1038));
  XOR2_X1   g0838(.A(new_n1038), .B(KEYINPUT110), .Z(new_n1039));
  NAND4_X1  g0839(.A1(new_n1034), .A2(new_n1035), .A3(new_n1037), .A4(new_n1039), .ZN(new_n1040));
  AND2_X1   g0840(.A1(new_n1032), .A2(new_n1040), .ZN(new_n1041));
  OAI211_X1 g0841(.A(new_n740), .B(new_n1025), .C1(new_n1041), .C2(new_n983), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n912), .A2(new_n800), .B1(new_n1024), .B2(new_n1042), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1043), .B1(new_n1024), .B2(new_n1042), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1022), .A2(new_n1023), .A3(new_n1044), .ZN(G390));
  NAND2_X1  g0845(.A1(new_n816), .A2(new_n892), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1046), .A2(new_n855), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1047), .A2(new_n902), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n812), .A2(new_n517), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n1049), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n667), .B(new_n1050), .C1(new_n726), .C2(new_n731), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n855), .B1(new_n1051), .B2(new_n811), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n878), .A2(new_n901), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n900), .A2(new_n1048), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n859), .A2(new_n806), .ZN(new_n1055));
  OR2_X1    g0855(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1053), .A2(new_n1052), .ZN(new_n1057));
  OAI21_X1  g0857(.A(KEYINPUT39), .B1(new_n894), .B2(new_n895), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n869), .A2(new_n877), .A3(new_n897), .ZN(new_n1059));
  OAI211_X1 g0859(.A(new_n1058), .B(new_n1059), .C1(new_n901), .C2(new_n893), .ZN(new_n1060));
  NOR3_X1   g0860(.A1(new_n880), .A2(new_n806), .A3(new_n814), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1061), .A2(new_n855), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n1062), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1057), .A2(new_n1060), .A3(new_n1063), .ZN(new_n1064));
  OAI211_X1 g0864(.A(G330), .B(new_n813), .C1(new_n856), .C2(new_n858), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1063), .B1(new_n854), .B2(new_n1065), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n1051), .A2(new_n811), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT112), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n1068), .B(new_n854), .C1(new_n717), .C2(new_n814), .ZN(new_n1069));
  OAI21_X1  g0869(.A(KEYINPUT112), .B1(new_n1061), .B2(new_n855), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n1069), .B(new_n1070), .C1(new_n806), .C2(new_n859), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n1066), .A2(new_n1067), .B1(new_n1071), .B2(new_n1046), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n906), .B1(G330), .B2(new_n888), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1073), .ZN(new_n1074));
  OAI211_X1 g0874(.A(new_n1056), .B(new_n1064), .C1(new_n1072), .C2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1071), .A2(new_n1046), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1065), .A2(new_n854), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1077), .A2(new_n1067), .A3(new_n1062), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1076), .A2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1064), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1079), .A2(new_n1080), .A3(new_n1073), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1075), .A2(new_n1081), .ZN(new_n1082));
  OAI21_X1  g0882(.A(KEYINPUT113), .B1(new_n1082), .B2(new_n690), .ZN(new_n1083));
  INV_X1    g0883(.A(KEYINPUT113), .ZN(new_n1084));
  NAND4_X1  g0884(.A1(new_n1075), .A2(new_n1084), .A3(new_n689), .A4(new_n1081), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1086));
  AND2_X1   g0886(.A1(new_n1080), .A2(new_n739), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n900), .A2(new_n798), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n758), .A2(G68), .B1(new_n822), .B2(G97), .ZN(new_n1089));
  OAI221_X1 g0889(.A(new_n1089), .B1(new_n825), .B2(new_n836), .C1(new_n754), .C2(new_n213), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(new_n821), .A2(G116), .B1(G294), .B2(new_n768), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1091), .B(new_n329), .C1(new_n215), .C2(new_n770), .ZN(new_n1092));
  AOI211_X1 g0892(.A(new_n1090), .B(new_n1092), .C1(G107), .C2(new_n744), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n760), .A2(G128), .B1(new_n744), .B2(G137), .ZN(new_n1094));
  XOR2_X1   g0894(.A(KEYINPUT54), .B(G143), .Z(new_n1095));
  XNOR2_X1  g0895(.A(new_n1095), .B(KEYINPUT114), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1096), .ZN(new_n1097));
  OAI221_X1 g0897(.A(new_n1094), .B1(new_n828), .B2(new_n775), .C1(new_n1097), .C2(new_n765), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n768), .A2(G125), .ZN(new_n1099));
  OAI221_X1 g0899(.A(new_n1099), .B1(new_n366), .B2(new_n757), .C1(new_n754), .C2(new_n469), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n830), .A2(G150), .ZN(new_n1101));
  AND2_X1   g0901(.A1(new_n1101), .A2(KEYINPUT53), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n332), .B1(new_n1101), .B2(KEYINPUT53), .ZN(new_n1103));
  NOR4_X1   g0903(.A1(new_n1098), .A2(new_n1100), .A3(new_n1102), .A4(new_n1103), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n789), .B1(new_n1093), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n377), .A2(new_n843), .ZN(new_n1106));
  AND4_X1   g0906(.A1(new_n740), .A2(new_n1088), .A3(new_n1105), .A4(new_n1106), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n1087), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1086), .A2(new_n1108), .ZN(G378));
  OR2_X1    g0909(.A1(new_n1073), .A2(KEYINPUT116), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1073), .A2(KEYINPUT116), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1081), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n886), .A2(KEYINPUT115), .A3(G330), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n903), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n383), .A2(new_n862), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1116), .B1(new_n399), .B2(new_n436), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n399), .A2(new_n436), .A3(new_n1116), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1120));
  AND3_X1   g0920(.A1(new_n1118), .A2(new_n1119), .A3(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1120), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n806), .B1(new_n879), .B2(new_n885), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1124), .B1(new_n1125), .B2(KEYINPUT115), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1125), .A2(KEYINPUT115), .A3(new_n903), .ZN(new_n1127));
  AND3_X1   g0927(.A1(new_n1115), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1126), .B1(new_n1115), .B2(new_n1127), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1112), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(KEYINPUT57), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  OAI211_X1 g0932(.A(KEYINPUT57), .B(new_n1112), .C1(new_n1128), .C2(new_n1129), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1132), .A2(new_n689), .A3(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT115), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1123), .B1(new_n887), .B2(new_n1135), .ZN(new_n1136));
  AND3_X1   g0936(.A1(new_n1125), .A2(KEYINPUT115), .A3(new_n903), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n903), .B1(new_n1125), .B2(KEYINPUT115), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1136), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1115), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(new_n739), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1123), .A2(new_n798), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n366), .B1(new_n253), .B2(G41), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n760), .A2(G125), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1145), .B1(new_n754), .B2(new_n369), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n821), .A2(G128), .B1(G132), .B2(new_n744), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1147), .B1(new_n770), .B2(new_n1097), .ZN(new_n1148));
  AOI211_X1 g0948(.A(new_n1146), .B(new_n1148), .C1(G137), .C2(new_n822), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT59), .ZN(new_n1150));
  OR2_X1    g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n758), .A2(G159), .ZN(new_n1152));
  AOI21_X1  g0952(.A(G33), .B1(new_n768), .B2(G124), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n1151), .A2(new_n282), .A3(new_n1152), .A4(new_n1153), .ZN(new_n1154));
  AND2_X1   g0954(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1144), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n757), .A2(new_n209), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(new_n830), .A2(G77), .B1(new_n768), .B2(G283), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n822), .A2(new_n451), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n821), .A2(G107), .ZN(new_n1160));
  NAND4_X1  g0960(.A1(new_n966), .A2(new_n1158), .A3(new_n1159), .A4(new_n1160), .ZN(new_n1161));
  AOI211_X1 g0961(.A(new_n1157), .B(new_n1161), .C1(G116), .C2(new_n760), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n744), .A2(G97), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n1162), .A2(new_n282), .A3(new_n329), .A4(new_n1163), .ZN(new_n1164));
  XOR2_X1   g0964(.A(new_n1164), .B(KEYINPUT58), .Z(new_n1165));
  OAI21_X1  g0965(.A(new_n789), .B1(new_n1156), .B2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n843), .A2(new_n366), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n1143), .A2(new_n740), .A3(new_n1166), .A4(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1142), .A2(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1134), .A2(new_n1170), .ZN(G375));
  NAND2_X1  g0971(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1079), .A2(new_n1073), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1172), .A2(new_n1173), .A3(new_n926), .ZN(new_n1174));
  OAI221_X1 g0974(.A(new_n329), .B1(new_n273), .B2(new_n765), .C1(new_n745), .C2(new_n589), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n995), .B1(G294), .B2(new_n760), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n830), .A2(G97), .B1(new_n758), .B2(G77), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n1176), .B(new_n1177), .C1(new_n836), .C2(new_n775), .ZN(new_n1178));
  AOI211_X1 g0978(.A(new_n1175), .B(new_n1178), .C1(G303), .C2(new_n768), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1157), .B1(new_n755), .B2(G50), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1180), .B1(new_n469), .B2(new_n770), .ZN(new_n1181));
  OAI221_X1 g0981(.A(new_n332), .B1(new_n828), .B2(new_n825), .C1(new_n1097), .C2(new_n745), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n765), .A2(new_n369), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n768), .A2(G128), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1184), .B1(new_n775), .B2(new_n824), .ZN(new_n1185));
  NOR4_X1   g0985(.A1(new_n1181), .A2(new_n1182), .A3(new_n1183), .A4(new_n1185), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n789), .B1(new_n1179), .B2(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(KEYINPUT118), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n741), .B1(new_n423), .B2(new_n843), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1187), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n855), .A2(new_n799), .ZN(new_n1191));
  AOI211_X1 g0991(.A(new_n1190), .B(new_n1191), .C1(new_n1188), .C2(new_n1189), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(new_n739), .B(KEYINPUT117), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1192), .B1(new_n1079), .B2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1174), .A2(new_n1194), .ZN(G381));
  INV_X1    g0995(.A(new_n1133), .ZN(new_n1196));
  AOI21_X1  g0996(.A(KEYINPUT57), .B1(new_n1141), .B2(new_n1112), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1169), .B1(new_n1198), .B2(new_n689), .ZN(new_n1199));
  XNOR2_X1  g0999(.A(new_n1199), .B(KEYINPUT119), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1108), .B1(new_n1082), .B2(new_n690), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(G387), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(G393), .A2(G396), .ZN(new_n1204));
  INV_X1    g1004(.A(G384), .ZN(new_n1205));
  INV_X1    g1005(.A(G390), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1204), .A2(new_n1205), .A3(new_n1206), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n1207), .A2(G381), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1202), .A2(new_n1203), .A3(new_n1208), .ZN(G407));
  NAND2_X1  g1009(.A1(new_n1202), .A2(new_n666), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(G407), .A2(G213), .A3(new_n1210), .ZN(new_n1211));
  XOR2_X1   g1011(.A(new_n1211), .B(KEYINPUT120), .Z(G409));
  AOI22_X1  g1012(.A1(new_n1014), .A2(new_n1019), .B1(new_n804), .B2(new_n808), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n1204), .A2(new_n1213), .ZN(new_n1214));
  AND2_X1   g1014(.A1(new_n1214), .A2(KEYINPUT123), .ZN(new_n1215));
  AND3_X1   g1015(.A1(new_n1215), .A2(new_n1203), .A3(G390), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(G387), .A2(new_n1206), .A3(new_n1214), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n1203), .A2(G390), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1217), .B1(new_n1218), .B2(new_n1215), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1203), .A2(G390), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1216), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(G378), .A2(new_n1134), .A3(new_n1170), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1141), .A2(new_n926), .A3(new_n1112), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1141), .A2(new_n1193), .ZN(new_n1224));
  AND3_X1   g1024(.A1(new_n1223), .A2(new_n1168), .A3(new_n1224), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1222), .B1(new_n1201), .B2(new_n1225), .ZN(new_n1226));
  OR2_X1    g1026(.A1(new_n1226), .A2(KEYINPUT121), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n666), .A2(G213), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1226), .A2(KEYINPUT121), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1227), .A2(new_n1228), .A3(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT60), .ZN(new_n1231));
  OAI211_X1 g1031(.A(new_n689), .B(new_n1173), .C1(new_n1172), .C2(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(KEYINPUT60), .B1(new_n1072), .B2(new_n1074), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1194), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1234));
  XNOR2_X1  g1034(.A(new_n1234), .B(new_n1205), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n666), .A2(G213), .A3(G2897), .ZN(new_n1236));
  XOR2_X1   g1036(.A(new_n1235), .B(new_n1236), .Z(new_n1237));
  INV_X1    g1037(.A(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1221), .B1(new_n1230), .B2(new_n1238), .ZN(new_n1239));
  AND2_X1   g1039(.A1(new_n1226), .A2(new_n1228), .ZN(new_n1240));
  AND2_X1   g1040(.A1(new_n1240), .A2(KEYINPUT63), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1235), .ZN(new_n1242));
  AOI21_X1  g1042(.A(KEYINPUT61), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1227), .A2(new_n1242), .A3(new_n1228), .A4(new_n1229), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT63), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT122), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1244), .A2(KEYINPUT122), .A3(new_n1245), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1239), .A2(new_n1243), .A3(new_n1248), .A4(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT62), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(new_n1235), .A2(new_n1251), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(new_n1244), .A2(new_n1251), .B1(new_n1240), .B2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT61), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1254), .B1(new_n1240), .B2(new_n1237), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1221), .B1(new_n1253), .B2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1250), .A2(new_n1256), .ZN(G405));
  INV_X1    g1057(.A(new_n1221), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT126), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT125), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT124), .ZN(new_n1261));
  AND3_X1   g1061(.A1(G378), .A2(new_n1134), .A3(new_n1170), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1201), .B1(new_n1134), .B2(new_n1170), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1261), .B1(new_n1262), .B2(new_n1263), .ZN(new_n1264));
  OAI211_X1 g1064(.A(KEYINPUT124), .B(new_n1222), .C1(new_n1199), .C2(new_n1201), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1260), .B1(new_n1266), .B2(new_n1242), .ZN(new_n1267));
  AOI211_X1 g1067(.A(KEYINPUT125), .B(new_n1235), .C1(new_n1264), .C2(new_n1265), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1201), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(G375), .A2(new_n1270), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1271), .A2(new_n1235), .A3(new_n1222), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1259), .B1(new_n1269), .B2(new_n1272), .ZN(new_n1273));
  NOR3_X1   g1073(.A1(new_n1262), .A2(new_n1263), .A3(new_n1261), .ZN(new_n1274));
  AOI21_X1  g1074(.A(KEYINPUT124), .B1(new_n1271), .B2(new_n1222), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1242), .B1(new_n1274), .B2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(KEYINPUT125), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1266), .A2(new_n1260), .A3(new_n1242), .ZN(new_n1278));
  AND4_X1   g1078(.A1(new_n1259), .A2(new_n1277), .A3(new_n1272), .A4(new_n1278), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1258), .B1(new_n1273), .B2(new_n1279), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1269), .A2(new_n1259), .A3(new_n1272), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1277), .A2(new_n1272), .A3(new_n1278), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(KEYINPUT126), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1281), .A2(new_n1283), .A3(new_n1221), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1280), .A2(new_n1284), .ZN(G402));
endmodule


