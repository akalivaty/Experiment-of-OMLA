

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582;

  XNOR2_X1 U323 ( .A(n333), .B(n332), .ZN(n337) );
  XNOR2_X1 U324 ( .A(n331), .B(n330), .ZN(n332) );
  XNOR2_X1 U325 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n392) );
  XNOR2_X1 U326 ( .A(n393), .B(n392), .ZN(n532) );
  XNOR2_X1 U327 ( .A(KEYINPUT58), .B(G190GAT), .ZN(n457) );
  XNOR2_X1 U328 ( .A(n458), .B(n457), .ZN(G1351GAT) );
  XOR2_X1 U329 ( .A(KEYINPUT120), .B(KEYINPUT54), .Z(n395) );
  XOR2_X1 U330 ( .A(G183GAT), .B(KEYINPUT82), .Z(n305) );
  XOR2_X1 U331 ( .A(KEYINPUT96), .B(n305), .Z(n292) );
  NAND2_X1 U332 ( .A1(G226GAT), .A2(G233GAT), .ZN(n291) );
  XNOR2_X1 U333 ( .A(n292), .B(n291), .ZN(n298) );
  XOR2_X1 U334 ( .A(G36GAT), .B(G190GAT), .Z(n325) );
  XNOR2_X1 U335 ( .A(G176GAT), .B(G92GAT), .ZN(n293) );
  XNOR2_X1 U336 ( .A(n293), .B(G64GAT), .ZN(n353) );
  XOR2_X1 U337 ( .A(n325), .B(n353), .Z(n296) );
  XOR2_X1 U338 ( .A(G169GAT), .B(G8GAT), .Z(n367) );
  XNOR2_X1 U339 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n294) );
  XNOR2_X1 U340 ( .A(n294), .B(KEYINPUT17), .ZN(n442) );
  XNOR2_X1 U341 ( .A(n367), .B(n442), .ZN(n295) );
  XNOR2_X1 U342 ( .A(n296), .B(n295), .ZN(n297) );
  XNOR2_X1 U343 ( .A(n298), .B(n297), .ZN(n302) );
  XOR2_X1 U344 ( .A(G211GAT), .B(G218GAT), .Z(n300) );
  XNOR2_X1 U345 ( .A(KEYINPUT21), .B(G204GAT), .ZN(n299) );
  XNOR2_X1 U346 ( .A(n300), .B(n299), .ZN(n301) );
  XNOR2_X1 U347 ( .A(G197GAT), .B(n301), .ZN(n432) );
  XOR2_X1 U348 ( .A(n302), .B(n432), .Z(n522) );
  INV_X1 U349 ( .A(n522), .ZN(n466) );
  XOR2_X1 U350 ( .A(KEYINPUT85), .B(KEYINPUT86), .Z(n304) );
  XNOR2_X1 U351 ( .A(KEYINPUT12), .B(KEYINPUT87), .ZN(n303) );
  XNOR2_X1 U352 ( .A(n304), .B(n303), .ZN(n324) );
  XOR2_X1 U353 ( .A(G22GAT), .B(G155GAT), .Z(n420) );
  XOR2_X1 U354 ( .A(n305), .B(n420), .Z(n307) );
  XNOR2_X1 U355 ( .A(G127GAT), .B(G71GAT), .ZN(n306) );
  XNOR2_X1 U356 ( .A(n307), .B(n306), .ZN(n320) );
  XOR2_X1 U357 ( .A(G64GAT), .B(G78GAT), .Z(n309) );
  XNOR2_X1 U358 ( .A(G8GAT), .B(G211GAT), .ZN(n308) );
  XNOR2_X1 U359 ( .A(n309), .B(n308), .ZN(n313) );
  XOR2_X1 U360 ( .A(KEYINPUT15), .B(KEYINPUT84), .Z(n311) );
  XNOR2_X1 U361 ( .A(KEYINPUT83), .B(KEYINPUT14), .ZN(n310) );
  XNOR2_X1 U362 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U363 ( .A(n313), .B(n312), .Z(n318) );
  XNOR2_X1 U364 ( .A(G15GAT), .B(G1GAT), .ZN(n314) );
  XNOR2_X1 U365 ( .A(n314), .B(KEYINPUT69), .ZN(n368) );
  XOR2_X1 U366 ( .A(KEYINPUT13), .B(KEYINPUT70), .Z(n316) );
  XNOR2_X1 U367 ( .A(G57GAT), .B(KEYINPUT71), .ZN(n315) );
  XNOR2_X1 U368 ( .A(n316), .B(n315), .ZN(n360) );
  XNOR2_X1 U369 ( .A(n368), .B(n360), .ZN(n317) );
  XNOR2_X1 U370 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U371 ( .A(n320), .B(n319), .Z(n322) );
  NAND2_X1 U372 ( .A1(G231GAT), .A2(G233GAT), .ZN(n321) );
  XNOR2_X1 U373 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U374 ( .A(n324), .B(n323), .Z(n554) );
  XOR2_X1 U375 ( .A(KEYINPUT9), .B(n325), .Z(n327) );
  XOR2_X1 U376 ( .A(G99GAT), .B(G85GAT), .Z(n354) );
  XNOR2_X1 U377 ( .A(G218GAT), .B(n354), .ZN(n326) );
  XNOR2_X1 U378 ( .A(n327), .B(n326), .ZN(n333) );
  XOR2_X1 U379 ( .A(KEYINPUT11), .B(KEYINPUT81), .Z(n329) );
  XNOR2_X1 U380 ( .A(G106GAT), .B(G92GAT), .ZN(n328) );
  XOR2_X1 U381 ( .A(n329), .B(n328), .Z(n331) );
  NAND2_X1 U382 ( .A1(G232GAT), .A2(G233GAT), .ZN(n330) );
  XOR2_X1 U383 ( .A(KEYINPUT80), .B(KEYINPUT10), .Z(n335) );
  XNOR2_X1 U384 ( .A(G134GAT), .B(KEYINPUT79), .ZN(n334) );
  XOR2_X1 U385 ( .A(n335), .B(n334), .Z(n336) );
  XNOR2_X1 U386 ( .A(n337), .B(n336), .ZN(n342) );
  XOR2_X1 U387 ( .A(G29GAT), .B(G43GAT), .Z(n339) );
  XNOR2_X1 U388 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n338) );
  XNOR2_X1 U389 ( .A(n339), .B(n338), .ZN(n372) );
  XNOR2_X1 U390 ( .A(G50GAT), .B(KEYINPUT78), .ZN(n340) );
  XNOR2_X1 U391 ( .A(n340), .B(G162GAT), .ZN(n427) );
  XNOR2_X1 U392 ( .A(n372), .B(n427), .ZN(n341) );
  XNOR2_X1 U393 ( .A(n342), .B(n341), .ZN(n557) );
  XOR2_X1 U394 ( .A(KEYINPUT36), .B(KEYINPUT103), .Z(n343) );
  XNOR2_X1 U395 ( .A(n557), .B(n343), .ZN(n580) );
  AND2_X1 U396 ( .A1(n554), .A2(n580), .ZN(n345) );
  XNOR2_X1 U397 ( .A(KEYINPUT45), .B(KEYINPUT113), .ZN(n344) );
  XNOR2_X1 U398 ( .A(n345), .B(n344), .ZN(n365) );
  XOR2_X1 U399 ( .A(KEYINPUT72), .B(KEYINPUT75), .Z(n347) );
  XNOR2_X1 U400 ( .A(KEYINPUT74), .B(KEYINPUT77), .ZN(n346) );
  XNOR2_X1 U401 ( .A(n347), .B(n346), .ZN(n364) );
  XOR2_X1 U402 ( .A(KEYINPUT31), .B(KEYINPUT73), .Z(n349) );
  XNOR2_X1 U403 ( .A(KEYINPUT33), .B(KEYINPUT32), .ZN(n348) );
  XNOR2_X1 U404 ( .A(n349), .B(n348), .ZN(n350) );
  XNOR2_X1 U405 ( .A(n350), .B(KEYINPUT76), .ZN(n352) );
  XOR2_X1 U406 ( .A(G120GAT), .B(G71GAT), .Z(n438) );
  XOR2_X1 U407 ( .A(n438), .B(G204GAT), .Z(n351) );
  XOR2_X1 U408 ( .A(n352), .B(n351), .Z(n358) );
  XOR2_X1 U409 ( .A(n354), .B(n353), .Z(n356) );
  NAND2_X1 U410 ( .A1(G230GAT), .A2(G233GAT), .ZN(n355) );
  XNOR2_X1 U411 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U412 ( .A(n358), .B(n357), .ZN(n362) );
  XNOR2_X1 U413 ( .A(G106GAT), .B(G78GAT), .ZN(n359) );
  XNOR2_X1 U414 ( .A(n359), .B(G148GAT), .ZN(n419) );
  XNOR2_X1 U415 ( .A(n419), .B(n360), .ZN(n361) );
  XNOR2_X1 U416 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U417 ( .A(n364), .B(n363), .ZN(n571) );
  NOR2_X1 U418 ( .A1(n365), .A2(n571), .ZN(n366) );
  XNOR2_X1 U419 ( .A(n366), .B(KEYINPUT114), .ZN(n383) );
  XOR2_X1 U420 ( .A(n368), .B(n367), .Z(n370) );
  NAND2_X1 U421 ( .A1(G229GAT), .A2(G233GAT), .ZN(n369) );
  XNOR2_X1 U422 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U423 ( .A(n371), .B(KEYINPUT29), .Z(n374) );
  XNOR2_X1 U424 ( .A(n372), .B(KEYINPUT67), .ZN(n373) );
  XNOR2_X1 U425 ( .A(n374), .B(n373), .ZN(n382) );
  XOR2_X1 U426 ( .A(G141GAT), .B(G113GAT), .Z(n376) );
  XNOR2_X1 U427 ( .A(G36GAT), .B(G50GAT), .ZN(n375) );
  XNOR2_X1 U428 ( .A(n376), .B(n375), .ZN(n380) );
  XOR2_X1 U429 ( .A(KEYINPUT68), .B(KEYINPUT30), .Z(n378) );
  XNOR2_X1 U430 ( .A(G197GAT), .B(G22GAT), .ZN(n377) );
  XNOR2_X1 U431 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U432 ( .A(n380), .B(n379), .Z(n381) );
  XNOR2_X1 U433 ( .A(n382), .B(n381), .ZN(n561) );
  INV_X1 U434 ( .A(n561), .ZN(n567) );
  NAND2_X1 U435 ( .A1(n383), .A2(n567), .ZN(n391) );
  INV_X1 U436 ( .A(KEYINPUT41), .ZN(n384) );
  XNOR2_X1 U437 ( .A(n571), .B(n384), .ZN(n459) );
  NAND2_X1 U438 ( .A1(n459), .A2(n561), .ZN(n386) );
  XNOR2_X1 U439 ( .A(KEYINPUT46), .B(KEYINPUT112), .ZN(n385) );
  XNOR2_X1 U440 ( .A(n386), .B(n385), .ZN(n387) );
  INV_X1 U441 ( .A(n554), .ZN(n576) );
  NAND2_X1 U442 ( .A1(n387), .A2(n576), .ZN(n388) );
  NOR2_X1 U443 ( .A1(n388), .A2(n557), .ZN(n389) );
  XNOR2_X1 U444 ( .A(KEYINPUT47), .B(n389), .ZN(n390) );
  NAND2_X1 U445 ( .A1(n391), .A2(n390), .ZN(n393) );
  NAND2_X1 U446 ( .A1(n466), .A2(n532), .ZN(n394) );
  XNOR2_X1 U447 ( .A(n395), .B(n394), .ZN(n417) );
  XOR2_X1 U448 ( .A(KEYINPUT95), .B(KEYINPUT4), .Z(n397) );
  XNOR2_X1 U449 ( .A(KEYINPUT5), .B(KEYINPUT1), .ZN(n396) );
  XNOR2_X1 U450 ( .A(n397), .B(n396), .ZN(n416) );
  XOR2_X1 U451 ( .A(G85GAT), .B(G162GAT), .Z(n399) );
  XNOR2_X1 U452 ( .A(G29GAT), .B(G120GAT), .ZN(n398) );
  XNOR2_X1 U453 ( .A(n399), .B(n398), .ZN(n403) );
  XOR2_X1 U454 ( .A(KEYINPUT6), .B(G148GAT), .Z(n401) );
  XNOR2_X1 U455 ( .A(G1GAT), .B(G155GAT), .ZN(n400) );
  XNOR2_X1 U456 ( .A(n401), .B(n400), .ZN(n402) );
  XOR2_X1 U457 ( .A(n403), .B(n402), .Z(n414) );
  XNOR2_X1 U458 ( .A(G127GAT), .B(KEYINPUT88), .ZN(n404) );
  XNOR2_X1 U459 ( .A(n404), .B(KEYINPUT0), .ZN(n405) );
  XOR2_X1 U460 ( .A(n405), .B(KEYINPUT89), .Z(n407) );
  XNOR2_X1 U461 ( .A(G113GAT), .B(G134GAT), .ZN(n406) );
  XNOR2_X1 U462 ( .A(n407), .B(n406), .ZN(n450) );
  XOR2_X1 U463 ( .A(KEYINPUT2), .B(KEYINPUT3), .Z(n409) );
  XNOR2_X1 U464 ( .A(G141GAT), .B(KEYINPUT93), .ZN(n408) );
  XNOR2_X1 U465 ( .A(n409), .B(n408), .ZN(n426) );
  XOR2_X1 U466 ( .A(n426), .B(G57GAT), .Z(n411) );
  NAND2_X1 U467 ( .A1(G225GAT), .A2(G233GAT), .ZN(n410) );
  XNOR2_X1 U468 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U469 ( .A(n450), .B(n412), .ZN(n413) );
  XNOR2_X1 U470 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U471 ( .A(n416), .B(n415), .ZN(n477) );
  INV_X1 U472 ( .A(n477), .ZN(n519) );
  NAND2_X1 U473 ( .A1(n417), .A2(n519), .ZN(n418) );
  XNOR2_X1 U474 ( .A(n418), .B(KEYINPUT65), .ZN(n565) );
  XOR2_X1 U475 ( .A(n419), .B(KEYINPUT24), .Z(n422) );
  XNOR2_X1 U476 ( .A(n420), .B(KEYINPUT22), .ZN(n421) );
  XNOR2_X1 U477 ( .A(n422), .B(n421), .ZN(n431) );
  XOR2_X1 U478 ( .A(KEYINPUT94), .B(KEYINPUT92), .Z(n424) );
  NAND2_X1 U479 ( .A1(G228GAT), .A2(G233GAT), .ZN(n423) );
  XNOR2_X1 U480 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U481 ( .A(n425), .B(KEYINPUT23), .Z(n429) );
  XNOR2_X1 U482 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U483 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U484 ( .A(n431), .B(n430), .ZN(n433) );
  XNOR2_X1 U485 ( .A(n433), .B(n432), .ZN(n470) );
  NAND2_X1 U486 ( .A1(n565), .A2(n470), .ZN(n435) );
  XOR2_X1 U487 ( .A(KEYINPUT121), .B(KEYINPUT55), .Z(n434) );
  XNOR2_X1 U488 ( .A(n435), .B(n434), .ZN(n453) );
  XOR2_X1 U489 ( .A(KEYINPUT91), .B(KEYINPUT20), .Z(n437) );
  XNOR2_X1 U490 ( .A(G190GAT), .B(G99GAT), .ZN(n436) );
  XNOR2_X1 U491 ( .A(n437), .B(n436), .ZN(n439) );
  XOR2_X1 U492 ( .A(n439), .B(n438), .Z(n441) );
  XNOR2_X1 U493 ( .A(G43GAT), .B(G15GAT), .ZN(n440) );
  XNOR2_X1 U494 ( .A(n441), .B(n440), .ZN(n446) );
  XOR2_X1 U495 ( .A(n442), .B(G169GAT), .Z(n444) );
  NAND2_X1 U496 ( .A1(G227GAT), .A2(G233GAT), .ZN(n443) );
  XNOR2_X1 U497 ( .A(n444), .B(n443), .ZN(n445) );
  XOR2_X1 U498 ( .A(n446), .B(n445), .Z(n452) );
  XOR2_X1 U499 ( .A(G176GAT), .B(KEYINPUT66), .Z(n448) );
  XNOR2_X1 U500 ( .A(G183GAT), .B(KEYINPUT90), .ZN(n447) );
  XNOR2_X1 U501 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U502 ( .A(n450), .B(n449), .ZN(n451) );
  XOR2_X1 U503 ( .A(n452), .B(n451), .Z(n534) );
  INV_X1 U504 ( .A(n534), .ZN(n471) );
  NAND2_X1 U505 ( .A1(n453), .A2(n471), .ZN(n454) );
  XOR2_X1 U506 ( .A(KEYINPUT122), .B(n454), .Z(n560) );
  NAND2_X1 U507 ( .A1(n560), .A2(n554), .ZN(n456) );
  XNOR2_X1 U508 ( .A(KEYINPUT124), .B(G183GAT), .ZN(n455) );
  XNOR2_X1 U509 ( .A(n456), .B(n455), .ZN(G1350GAT) );
  NAND2_X1 U510 ( .A1(n560), .A2(n557), .ZN(n458) );
  NAND2_X1 U511 ( .A1(n560), .A2(n459), .ZN(n463) );
  XOR2_X1 U512 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n461) );
  XOR2_X1 U513 ( .A(G176GAT), .B(KEYINPUT56), .Z(n460) );
  XNOR2_X1 U514 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U515 ( .A(n463), .B(n462), .ZN(G1349GAT) );
  NOR2_X1 U516 ( .A1(n567), .A2(n571), .ZN(n498) );
  XNOR2_X1 U517 ( .A(KEYINPUT28), .B(n470), .ZN(n531) );
  XNOR2_X1 U518 ( .A(KEYINPUT27), .B(n522), .ZN(n474) );
  NOR2_X1 U519 ( .A1(n519), .A2(n474), .ZN(n533) );
  NAND2_X1 U520 ( .A1(n531), .A2(n533), .ZN(n464) );
  XOR2_X1 U521 ( .A(KEYINPUT97), .B(n464), .Z(n465) );
  NOR2_X1 U522 ( .A1(n471), .A2(n465), .ZN(n480) );
  NAND2_X1 U523 ( .A1(n471), .A2(n466), .ZN(n467) );
  XOR2_X1 U524 ( .A(KEYINPUT99), .B(n467), .Z(n468) );
  NAND2_X1 U525 ( .A1(n468), .A2(n470), .ZN(n469) );
  XNOR2_X1 U526 ( .A(n469), .B(KEYINPUT25), .ZN(n476) );
  NOR2_X1 U527 ( .A1(n471), .A2(n470), .ZN(n473) );
  XNOR2_X1 U528 ( .A(KEYINPUT98), .B(KEYINPUT26), .ZN(n472) );
  XOR2_X1 U529 ( .A(n473), .B(n472), .Z(n563) );
  NOR2_X1 U530 ( .A1(n563), .A2(n474), .ZN(n475) );
  NOR2_X1 U531 ( .A1(n476), .A2(n475), .ZN(n478) );
  NOR2_X1 U532 ( .A1(n478), .A2(n477), .ZN(n479) );
  NOR2_X1 U533 ( .A1(n480), .A2(n479), .ZN(n494) );
  NOR2_X1 U534 ( .A1(n557), .A2(n576), .ZN(n481) );
  XOR2_X1 U535 ( .A(KEYINPUT16), .B(n481), .Z(n482) );
  NOR2_X1 U536 ( .A1(n494), .A2(n482), .ZN(n483) );
  XNOR2_X1 U537 ( .A(KEYINPUT100), .B(n483), .ZN(n508) );
  NAND2_X1 U538 ( .A1(n498), .A2(n508), .ZN(n490) );
  NOR2_X1 U539 ( .A1(n519), .A2(n490), .ZN(n484) );
  XOR2_X1 U540 ( .A(G1GAT), .B(n484), .Z(n485) );
  XNOR2_X1 U541 ( .A(KEYINPUT34), .B(n485), .ZN(G1324GAT) );
  NOR2_X1 U542 ( .A1(n522), .A2(n490), .ZN(n486) );
  XOR2_X1 U543 ( .A(G8GAT), .B(n486), .Z(G1325GAT) );
  NOR2_X1 U544 ( .A1(n534), .A2(n490), .ZN(n488) );
  XNOR2_X1 U545 ( .A(KEYINPUT101), .B(KEYINPUT35), .ZN(n487) );
  XNOR2_X1 U546 ( .A(n488), .B(n487), .ZN(n489) );
  XOR2_X1 U547 ( .A(G15GAT), .B(n489), .Z(G1326GAT) );
  NOR2_X1 U548 ( .A1(n531), .A2(n490), .ZN(n491) );
  XOR2_X1 U549 ( .A(KEYINPUT102), .B(n491), .Z(n492) );
  XNOR2_X1 U550 ( .A(G22GAT), .B(n492), .ZN(G1327GAT) );
  XNOR2_X1 U551 ( .A(G29GAT), .B(KEYINPUT105), .ZN(n493) );
  XNOR2_X1 U552 ( .A(n493), .B(KEYINPUT39), .ZN(n501) );
  XNOR2_X1 U553 ( .A(KEYINPUT104), .B(KEYINPUT37), .ZN(n497) );
  NOR2_X1 U554 ( .A1(n554), .A2(n494), .ZN(n495) );
  NAND2_X1 U555 ( .A1(n495), .A2(n580), .ZN(n496) );
  XNOR2_X1 U556 ( .A(n497), .B(n496), .ZN(n517) );
  NAND2_X1 U557 ( .A1(n517), .A2(n498), .ZN(n499) );
  XNOR2_X1 U558 ( .A(n499), .B(KEYINPUT38), .ZN(n505) );
  NOR2_X1 U559 ( .A1(n519), .A2(n505), .ZN(n500) );
  XOR2_X1 U560 ( .A(n501), .B(n500), .Z(G1328GAT) );
  NOR2_X1 U561 ( .A1(n522), .A2(n505), .ZN(n502) );
  XOR2_X1 U562 ( .A(G36GAT), .B(n502), .Z(G1329GAT) );
  NOR2_X1 U563 ( .A1(n505), .A2(n534), .ZN(n503) );
  XOR2_X1 U564 ( .A(KEYINPUT40), .B(n503), .Z(n504) );
  XNOR2_X1 U565 ( .A(G43GAT), .B(n504), .ZN(G1330GAT) );
  NOR2_X1 U566 ( .A1(n531), .A2(n505), .ZN(n506) );
  XOR2_X1 U567 ( .A(KEYINPUT106), .B(n506), .Z(n507) );
  XNOR2_X1 U568 ( .A(G50GAT), .B(n507), .ZN(G1331GAT) );
  AND2_X1 U569 ( .A1(n459), .A2(n567), .ZN(n518) );
  NAND2_X1 U570 ( .A1(n518), .A2(n508), .ZN(n513) );
  NOR2_X1 U571 ( .A1(n519), .A2(n513), .ZN(n509) );
  XOR2_X1 U572 ( .A(G57GAT), .B(n509), .Z(n510) );
  XNOR2_X1 U573 ( .A(KEYINPUT42), .B(n510), .ZN(G1332GAT) );
  NOR2_X1 U574 ( .A1(n522), .A2(n513), .ZN(n511) );
  XOR2_X1 U575 ( .A(G64GAT), .B(n511), .Z(G1333GAT) );
  NOR2_X1 U576 ( .A1(n534), .A2(n513), .ZN(n512) );
  XOR2_X1 U577 ( .A(G71GAT), .B(n512), .Z(G1334GAT) );
  NOR2_X1 U578 ( .A1(n531), .A2(n513), .ZN(n515) );
  XNOR2_X1 U579 ( .A(KEYINPUT107), .B(KEYINPUT43), .ZN(n514) );
  XNOR2_X1 U580 ( .A(n515), .B(n514), .ZN(n516) );
  XOR2_X1 U581 ( .A(G78GAT), .B(n516), .Z(G1335GAT) );
  NAND2_X1 U582 ( .A1(n518), .A2(n517), .ZN(n528) );
  NOR2_X1 U583 ( .A1(n519), .A2(n528), .ZN(n520) );
  XOR2_X1 U584 ( .A(G85GAT), .B(n520), .Z(n521) );
  XNOR2_X1 U585 ( .A(KEYINPUT108), .B(n521), .ZN(G1336GAT) );
  NOR2_X1 U586 ( .A1(n522), .A2(n528), .ZN(n523) );
  XOR2_X1 U587 ( .A(G92GAT), .B(n523), .Z(G1337GAT) );
  NOR2_X1 U588 ( .A1(n534), .A2(n528), .ZN(n525) );
  XNOR2_X1 U589 ( .A(G99GAT), .B(KEYINPUT109), .ZN(n524) );
  XNOR2_X1 U590 ( .A(n525), .B(n524), .ZN(G1338GAT) );
  XOR2_X1 U591 ( .A(KEYINPUT110), .B(KEYINPUT111), .Z(n527) );
  XNOR2_X1 U592 ( .A(G106GAT), .B(KEYINPUT44), .ZN(n526) );
  XNOR2_X1 U593 ( .A(n527), .B(n526), .ZN(n530) );
  NOR2_X1 U594 ( .A1(n531), .A2(n528), .ZN(n529) );
  XOR2_X1 U595 ( .A(n530), .B(n529), .Z(G1339GAT) );
  INV_X1 U596 ( .A(n531), .ZN(n537) );
  NAND2_X1 U597 ( .A1(n533), .A2(n532), .ZN(n548) );
  NOR2_X1 U598 ( .A1(n534), .A2(n548), .ZN(n535) );
  XNOR2_X1 U599 ( .A(n535), .B(KEYINPUT115), .ZN(n536) );
  NOR2_X1 U600 ( .A1(n537), .A2(n536), .ZN(n545) );
  NAND2_X1 U601 ( .A1(n545), .A2(n561), .ZN(n538) );
  XNOR2_X1 U602 ( .A(G113GAT), .B(n538), .ZN(G1340GAT) );
  XOR2_X1 U603 ( .A(G120GAT), .B(KEYINPUT49), .Z(n540) );
  NAND2_X1 U604 ( .A1(n545), .A2(n459), .ZN(n539) );
  XNOR2_X1 U605 ( .A(n540), .B(n539), .ZN(G1341GAT) );
  XNOR2_X1 U606 ( .A(G127GAT), .B(KEYINPUT117), .ZN(n544) );
  XOR2_X1 U607 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n542) );
  NAND2_X1 U608 ( .A1(n545), .A2(n554), .ZN(n541) );
  XNOR2_X1 U609 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U610 ( .A(n544), .B(n543), .ZN(G1342GAT) );
  XOR2_X1 U611 ( .A(G134GAT), .B(KEYINPUT51), .Z(n547) );
  NAND2_X1 U612 ( .A1(n545), .A2(n557), .ZN(n546) );
  XNOR2_X1 U613 ( .A(n547), .B(n546), .ZN(G1343GAT) );
  NOR2_X1 U614 ( .A1(n563), .A2(n548), .ZN(n558) );
  NAND2_X1 U615 ( .A1(n558), .A2(n561), .ZN(n549) );
  XNOR2_X1 U616 ( .A(G141GAT), .B(n549), .ZN(G1344GAT) );
  XNOR2_X1 U617 ( .A(G148GAT), .B(KEYINPUT118), .ZN(n553) );
  XOR2_X1 U618 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n551) );
  NAND2_X1 U619 ( .A1(n558), .A2(n459), .ZN(n550) );
  XNOR2_X1 U620 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U621 ( .A(n553), .B(n552), .ZN(G1345GAT) );
  XOR2_X1 U622 ( .A(G155GAT), .B(KEYINPUT119), .Z(n556) );
  NAND2_X1 U623 ( .A1(n558), .A2(n554), .ZN(n555) );
  XNOR2_X1 U624 ( .A(n556), .B(n555), .ZN(G1346GAT) );
  NAND2_X1 U625 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n559), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U628 ( .A(G169GAT), .B(n562), .ZN(G1348GAT) );
  INV_X1 U629 ( .A(n563), .ZN(n564) );
  NAND2_X1 U630 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U631 ( .A(KEYINPUT125), .B(n566), .ZN(n579) );
  INV_X1 U632 ( .A(n579), .ZN(n575) );
  NOR2_X1 U633 ( .A1(n567), .A2(n575), .ZN(n569) );
  XNOR2_X1 U634 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U636 ( .A(G197GAT), .B(n570), .ZN(G1352GAT) );
  AND2_X1 U637 ( .A1(n571), .A2(n579), .ZN(n573) );
  XNOR2_X1 U638 ( .A(KEYINPUT126), .B(KEYINPUT61), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n573), .B(n572), .ZN(n574) );
  XNOR2_X1 U640 ( .A(G204GAT), .B(n574), .ZN(G1353GAT) );
  NOR2_X1 U641 ( .A1(n576), .A2(n575), .ZN(n578) );
  XNOR2_X1 U642 ( .A(G211GAT), .B(KEYINPUT127), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(G1354GAT) );
  NAND2_X1 U644 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U645 ( .A(n581), .B(KEYINPUT62), .ZN(n582) );
  XNOR2_X1 U646 ( .A(G218GAT), .B(n582), .ZN(G1355GAT) );
endmodule

