//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 1 1 0 0 1 0 1 1 0 1 1 0 1 1 0 1 0 1 0 0 1 1 0 1 0 1 0 0 1 0 1 1 1 1 1 1 1 0 1 0 1 1 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:29 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n559, new_n561, new_n562, new_n563, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n628, new_n629, new_n630,
    new_n631, new_n634, new_n635, new_n637, new_n638, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1221;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT65), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT66), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  NAND2_X1  g035(.A1(KEYINPUT67), .A2(G2104), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g038(.A1(KEYINPUT67), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AOI22_X1  g040(.A1(new_n465), .A2(G137), .B1(G101), .B2(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n466), .A2(G2105), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(KEYINPUT3), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n462), .A2(G2104), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n470), .A2(new_n471), .A3(G125), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n468), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n467), .A2(new_n474), .ZN(G160));
  XNOR2_X1  g050(.A(new_n465), .B(KEYINPUT68), .ZN(new_n476));
  AND2_X1   g051(.A1(new_n476), .A2(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  XNOR2_X1  g053(.A(new_n478), .B(KEYINPUT69), .ZN(new_n479));
  OAI21_X1  g054(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n480));
  INV_X1    g055(.A(G112), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n480), .B1(new_n481), .B2(G2105), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n476), .A2(new_n468), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n482), .B1(new_n484), .B2(G136), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n479), .A2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G162));
  NAND4_X1  g062(.A1(new_n470), .A2(new_n471), .A3(G138), .A4(new_n468), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(G126), .A2(G2105), .ZN(new_n491));
  NAND2_X1  g066(.A1(KEYINPUT4), .A2(G138), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n491), .B1(new_n492), .B2(G2105), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n465), .A2(new_n493), .ZN(new_n494));
  OR2_X1    g069(.A1(new_n468), .A2(G114), .ZN(new_n495));
  OAI21_X1  g070(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n490), .A2(new_n494), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(KEYINPUT70), .ZN(new_n500));
  AOI22_X1  g075(.A1(new_n465), .A2(new_n493), .B1(new_n495), .B2(new_n497), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT70), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n501), .A2(new_n502), .A3(new_n490), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n500), .A2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(G164));
  INV_X1    g080(.A(G62), .ZN(new_n506));
  NAND2_X1  g081(.A1(KEYINPUT71), .A2(G543), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT5), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g084(.A1(KEYINPUT71), .A2(KEYINPUT5), .A3(G543), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n506), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(G75), .A2(G543), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(new_n513));
  OAI21_X1  g088(.A(G651), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  OR2_X1    g089(.A1(KEYINPUT6), .A2(G651), .ZN(new_n515));
  NAND2_X1  g090(.A1(KEYINPUT6), .A2(G651), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n509), .A2(new_n510), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G88), .ZN(new_n518));
  INV_X1    g093(.A(G543), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n519), .B1(new_n515), .B2(new_n516), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G50), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n514), .A2(new_n518), .A3(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT72), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND4_X1  g099(.A1(new_n514), .A2(new_n518), .A3(KEYINPUT72), .A4(new_n521), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(new_n525), .ZN(G166));
  NAND2_X1  g101(.A1(new_n520), .A2(G51), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n509), .A2(new_n510), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n528), .A2(G63), .A3(G651), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n530), .B(KEYINPUT7), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n527), .A2(new_n529), .A3(new_n531), .ZN(new_n532));
  AND2_X1   g107(.A1(new_n517), .A2(G89), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n532), .A2(new_n533), .ZN(G168));
  AOI22_X1  g109(.A1(new_n528), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  INV_X1    g110(.A(G651), .ZN(new_n536));
  OR2_X1    g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n515), .A2(new_n516), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n538), .A2(G52), .A3(G543), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n528), .A2(new_n538), .ZN(new_n540));
  INV_X1    g115(.A(G90), .ZN(new_n541));
  OAI211_X1 g116(.A(new_n539), .B(KEYINPUT73), .C1(new_n540), .C2(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n517), .A2(G90), .ZN(new_n544));
  AOI21_X1  g119(.A(KEYINPUT73), .B1(new_n544), .B2(new_n539), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n537), .B1(new_n543), .B2(new_n545), .ZN(G301));
  INV_X1    g121(.A(G301), .ZN(G171));
  INV_X1    g122(.A(G56), .ZN(new_n548));
  AOI21_X1  g123(.A(new_n548), .B1(new_n509), .B2(new_n510), .ZN(new_n549));
  INV_X1    g124(.A(KEYINPUT74), .ZN(new_n550));
  AND2_X1   g125(.A1(G68), .A2(G543), .ZN(new_n551));
  OR3_X1    g126(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n550), .B1(new_n549), .B2(new_n551), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n552), .A2(G651), .A3(new_n553), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n517), .A2(G81), .B1(new_n520), .B2(G43), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(G153));
  NAND4_X1  g133(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n559));
  XOR2_X1   g134(.A(new_n559), .B(KEYINPUT75), .Z(G176));
  NAND2_X1  g135(.A1(G1), .A2(G3), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT76), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT8), .ZN(new_n563));
  NAND4_X1  g138(.A1(G319), .A2(G483), .A3(G661), .A4(new_n563), .ZN(G188));
  NAND3_X1  g139(.A1(new_n538), .A2(G53), .A3(G543), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(KEYINPUT9), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT9), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n520), .A2(new_n567), .A3(G53), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(G65), .ZN(new_n570));
  AOI21_X1  g145(.A(new_n570), .B1(new_n509), .B2(new_n510), .ZN(new_n571));
  AND2_X1   g146(.A1(G78), .A2(G543), .ZN(new_n572));
  OAI21_X1  g147(.A(G651), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n517), .A2(G91), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n569), .A2(new_n573), .A3(new_n574), .ZN(G299));
  INV_X1    g150(.A(G168), .ZN(G286));
  INV_X1    g151(.A(G166), .ZN(G303));
  NAND3_X1  g152(.A1(new_n538), .A2(G49), .A3(G543), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT77), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n520), .A2(KEYINPUT77), .A3(G49), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(G74), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n509), .A2(new_n583), .A3(new_n510), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n517), .A2(G87), .B1(new_n584), .B2(G651), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n582), .A2(new_n585), .ZN(G288));
  INV_X1    g161(.A(new_n510), .ZN(new_n587));
  AOI21_X1  g162(.A(KEYINPUT5), .B1(KEYINPUT71), .B2(G543), .ZN(new_n588));
  OAI21_X1  g163(.A(G61), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(G73), .A2(G543), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n591), .A2(G651), .B1(new_n520), .B2(G48), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n517), .A2(G86), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT78), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n517), .A2(KEYINPUT78), .A3(G86), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n592), .A2(new_n595), .A3(new_n596), .ZN(G305));
  NAND2_X1  g172(.A1(G72), .A2(G543), .ZN(new_n598));
  INV_X1    g173(.A(new_n528), .ZN(new_n599));
  INV_X1    g174(.A(G60), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n598), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT79), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n536), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n603), .B1(new_n602), .B2(new_n601), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n517), .A2(G85), .B1(new_n520), .B2(G47), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n604), .A2(new_n605), .ZN(G290));
  NAND2_X1  g181(.A1(G301), .A2(G868), .ZN(new_n607));
  XNOR2_X1  g182(.A(KEYINPUT80), .B(KEYINPUT10), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(G92), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n540), .B2(new_n610), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n517), .A2(G92), .A3(new_n608), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n611), .A2(new_n612), .B1(G54), .B2(new_n520), .ZN(new_n613));
  NAND2_X1  g188(.A1(G79), .A2(G543), .ZN(new_n614));
  INV_X1    g189(.A(KEYINPUT81), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n614), .B(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(KEYINPUT82), .ZN(new_n617));
  INV_X1    g192(.A(G66), .ZN(new_n618));
  OAI211_X1 g193(.A(new_n616), .B(new_n617), .C1(new_n599), .C2(new_n618), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n614), .B(KEYINPUT81), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n618), .B1(new_n509), .B2(new_n510), .ZN(new_n621));
  OAI21_X1  g196(.A(KEYINPUT82), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n619), .A2(new_n622), .A3(G651), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n613), .A2(new_n623), .ZN(new_n624));
  INV_X1    g199(.A(new_n624), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n607), .B1(new_n625), .B2(G868), .ZN(G284));
  OAI21_X1  g201(.A(new_n607), .B1(new_n625), .B2(G868), .ZN(G321));
  INV_X1    g202(.A(G868), .ZN(new_n628));
  NOR2_X1   g203(.A1(G286), .A2(new_n628), .ZN(new_n629));
  AND3_X1   g204(.A1(new_n569), .A2(new_n573), .A3(new_n574), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT83), .ZN(new_n631));
  AOI21_X1  g206(.A(new_n629), .B1(new_n631), .B2(new_n628), .ZN(G297));
  AOI21_X1  g207(.A(new_n629), .B1(new_n631), .B2(new_n628), .ZN(G280));
  INV_X1    g208(.A(G860), .ZN(new_n634));
  AOI21_X1  g209(.A(new_n624), .B1(G559), .B2(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT84), .ZN(G148));
  NAND2_X1  g211(.A1(new_n556), .A2(new_n628), .ZN(new_n637));
  NOR2_X1   g212(.A1(new_n624), .A2(G559), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n637), .B1(new_n638), .B2(new_n628), .ZN(G323));
  XNOR2_X1  g214(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g215(.A1(new_n484), .A2(G135), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n477), .A2(G123), .ZN(new_n642));
  OR2_X1    g217(.A1(G99), .A2(G2105), .ZN(new_n643));
  OAI211_X1 g218(.A(new_n643), .B(G2104), .C1(G111), .C2(new_n468), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n641), .A2(new_n642), .A3(new_n644), .ZN(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(new_n646));
  INV_X1    g221(.A(G2096), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n645), .A2(G2096), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n468), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n650), .B(KEYINPUT12), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT13), .ZN(new_n652));
  INV_X1    g227(.A(G2100), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n648), .A2(new_n649), .A3(new_n654), .ZN(G156));
  XOR2_X1   g230(.A(G2451), .B(G2454), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT16), .ZN(new_n657));
  XNOR2_X1  g232(.A(G1341), .B(G1348), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  INV_X1    g234(.A(KEYINPUT14), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2427), .B(G2438), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(G2430), .ZN(new_n662));
  XNOR2_X1  g237(.A(KEYINPUT15), .B(G2435), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n660), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n664), .B1(new_n663), .B2(new_n662), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n659), .B(new_n665), .Z(new_n666));
  XNOR2_X1  g241(.A(G2443), .B(G2446), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n666), .A2(new_n667), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n668), .A2(new_n669), .A3(G14), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n670), .B(KEYINPUT85), .Z(G401));
  INV_X1    g246(.A(KEYINPUT18), .ZN(new_n672));
  XOR2_X1   g247(.A(G2084), .B(G2090), .Z(new_n673));
  XNOR2_X1  g248(.A(G2067), .B(G2678), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n675), .A2(KEYINPUT17), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n673), .A2(new_n674), .ZN(new_n677));
  OAI21_X1  g252(.A(new_n672), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(new_n653), .ZN(new_n679));
  XOR2_X1   g254(.A(G2072), .B(G2078), .Z(new_n680));
  AOI21_X1  g255(.A(new_n680), .B1(new_n675), .B2(KEYINPUT18), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(new_n647), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n679), .B(new_n682), .ZN(G227));
  XOR2_X1   g258(.A(G1971), .B(G1976), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT19), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1956), .B(G2474), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1961), .B(G1966), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  AND2_X1   g263(.A1(new_n686), .A2(new_n687), .ZN(new_n689));
  NOR3_X1   g264(.A1(new_n685), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n685), .A2(new_n688), .ZN(new_n691));
  XOR2_X1   g266(.A(new_n691), .B(KEYINPUT20), .Z(new_n692));
  AOI211_X1 g267(.A(new_n690), .B(new_n692), .C1(new_n685), .C2(new_n689), .ZN(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1991), .B(G1996), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1981), .B(G1986), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(G229));
  INV_X1    g275(.A(G29), .ZN(new_n701));
  AND2_X1   g276(.A1(new_n701), .A2(G35), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n702), .B1(new_n486), .B2(G29), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT29), .ZN(new_n704));
  INV_X1    g279(.A(G2090), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  XOR2_X1   g281(.A(new_n706), .B(KEYINPUT95), .Z(new_n707));
  NAND2_X1  g282(.A1(new_n646), .A2(G29), .ZN(new_n708));
  INV_X1    g283(.A(G16), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G5), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(G171), .B2(new_n709), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(G1961), .ZN(new_n712));
  INV_X1    g287(.A(G28), .ZN(new_n713));
  OR2_X1    g288(.A1(new_n713), .A2(KEYINPUT30), .ZN(new_n714));
  AOI21_X1  g289(.A(G29), .B1(new_n713), .B2(KEYINPUT30), .ZN(new_n715));
  OR2_X1    g290(.A1(KEYINPUT31), .A2(G11), .ZN(new_n716));
  NAND2_X1  g291(.A1(KEYINPUT31), .A2(G11), .ZN(new_n717));
  AOI22_X1  g292(.A1(new_n714), .A2(new_n715), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n709), .A2(G21), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(G168), .B2(new_n709), .ZN(new_n720));
  INV_X1    g295(.A(G1966), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  NAND4_X1  g297(.A1(new_n708), .A2(new_n712), .A3(new_n718), .A4(new_n722), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n723), .A2(KEYINPUT94), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n701), .A2(G26), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT28), .ZN(new_n726));
  OAI21_X1  g301(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n727));
  INV_X1    g302(.A(G116), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n727), .B1(new_n728), .B2(G2105), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(new_n477), .B2(G128), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n484), .A2(G140), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n732), .A2(G29), .ZN(new_n733));
  AND2_X1   g308(.A1(new_n733), .A2(KEYINPUT89), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n733), .A2(KEYINPUT89), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n726), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(G2067), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(new_n705), .B2(new_n704), .ZN(new_n738));
  NOR2_X1   g313(.A1(G29), .A2(G33), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT90), .ZN(new_n740));
  NAND3_X1  g315(.A1(new_n470), .A2(new_n471), .A3(G127), .ZN(new_n741));
  INV_X1    g316(.A(G115), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n741), .B1(new_n742), .B2(new_n469), .ZN(new_n743));
  INV_X1    g318(.A(KEYINPUT25), .ZN(new_n744));
  NAND2_X1  g319(.A1(G103), .A2(G2104), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n744), .B1(new_n745), .B2(G2105), .ZN(new_n746));
  NAND4_X1  g321(.A1(new_n468), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n747));
  AOI22_X1  g322(.A1(new_n743), .A2(G2105), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(G139), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n748), .B1(new_n483), .B2(new_n749), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT91), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n740), .B1(new_n751), .B2(new_n701), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(G2072), .Z(new_n753));
  NAND2_X1  g328(.A1(G164), .A2(G29), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(G27), .B2(G29), .ZN(new_n755));
  INV_X1    g330(.A(G2078), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n755), .A2(new_n756), .ZN(new_n758));
  INV_X1    g333(.A(G34), .ZN(new_n759));
  AND2_X1   g334(.A1(new_n759), .A2(KEYINPUT24), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n759), .A2(KEYINPUT24), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n701), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G160), .B2(new_n701), .ZN(new_n763));
  INV_X1    g338(.A(G2084), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n758), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n709), .A2(G20), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT23), .Z(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(G299), .B2(G16), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(G1956), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n557), .A2(G16), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(G16), .B2(G19), .ZN(new_n772));
  INV_X1    g347(.A(G1341), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n770), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NOR4_X1   g349(.A1(new_n753), .A2(new_n757), .A3(new_n766), .A4(new_n774), .ZN(new_n775));
  NOR2_X1   g350(.A1(G4), .A2(G16), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(new_n625), .B2(G16), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(G1348), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n772), .A2(new_n773), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G1961), .B2(new_n711), .ZN(new_n780));
  AOI211_X1 g355(.A(new_n778), .B(new_n780), .C1(KEYINPUT94), .C2(new_n723), .ZN(new_n781));
  NAND3_X1  g356(.A1(new_n738), .A2(new_n775), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n701), .A2(G32), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n484), .A2(G141), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(KEYINPUT92), .Z(new_n785));
  NAND3_X1  g360(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n786));
  INV_X1    g361(.A(KEYINPUT26), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  NAND3_X1  g363(.A1(new_n468), .A2(G105), .A3(G2104), .ZN(new_n789));
  AOI21_X1  g364(.A(KEYINPUT93), .B1(new_n477), .B2(G129), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n476), .A2(G2105), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT93), .ZN(new_n792));
  INV_X1    g367(.A(G129), .ZN(new_n793));
  NOR3_X1   g368(.A1(new_n791), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  OAI211_X1 g369(.A(new_n788), .B(new_n789), .C1(new_n790), .C2(new_n794), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n785), .A2(new_n795), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n783), .B1(new_n796), .B2(new_n701), .ZN(new_n797));
  XOR2_X1   g372(.A(KEYINPUT27), .B(G1996), .Z(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  NOR4_X1   g374(.A1(new_n707), .A2(new_n724), .A3(new_n782), .A4(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n709), .A2(G6), .ZN(new_n801));
  INV_X1    g376(.A(G305), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n801), .B1(new_n802), .B2(new_n709), .ZN(new_n803));
  XNOR2_X1  g378(.A(KEYINPUT32), .B(G1981), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n709), .A2(G22), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT88), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(G166), .B2(new_n709), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n805), .B1(G1971), .B2(new_n808), .ZN(new_n809));
  NOR2_X1   g384(.A1(G16), .A2(G23), .ZN(new_n810));
  XOR2_X1   g385(.A(new_n810), .B(KEYINPUT86), .Z(new_n811));
  INV_X1    g386(.A(KEYINPUT87), .ZN(new_n812));
  NAND2_X1  g387(.A1(G288), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n582), .A2(KEYINPUT87), .A3(new_n585), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n811), .B1(new_n815), .B2(new_n709), .ZN(new_n816));
  XOR2_X1   g391(.A(KEYINPUT33), .B(G1976), .Z(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  OAI211_X1 g393(.A(new_n809), .B(new_n818), .C1(G1971), .C2(new_n808), .ZN(new_n819));
  OR2_X1    g394(.A1(new_n819), .A2(KEYINPUT34), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n819), .A2(KEYINPUT34), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n484), .A2(G131), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n477), .A2(G119), .ZN(new_n823));
  OR2_X1    g398(.A1(G95), .A2(G2105), .ZN(new_n824));
  OAI211_X1 g399(.A(new_n824), .B(G2104), .C1(G107), .C2(new_n468), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n822), .A2(new_n823), .A3(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n827), .A2(G29), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n828), .B1(G25), .B2(G29), .ZN(new_n829));
  XOR2_X1   g404(.A(KEYINPUT35), .B(G1991), .Z(new_n830));
  NOR2_X1   g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(G1986), .ZN(new_n832));
  AND2_X1   g407(.A1(new_n604), .A2(new_n605), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n833), .A2(new_n709), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n834), .B1(new_n709), .B2(G24), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n831), .B1(new_n832), .B2(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(new_n835), .ZN(new_n837));
  AOI22_X1  g412(.A1(new_n829), .A2(new_n830), .B1(new_n837), .B2(G1986), .ZN(new_n838));
  NAND4_X1  g413(.A1(new_n820), .A2(new_n821), .A3(new_n836), .A4(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT36), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n800), .A2(new_n840), .ZN(G150));
  INV_X1    g416(.A(G150), .ZN(G311));
  NAND2_X1  g417(.A1(new_n517), .A2(G93), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n520), .A2(G55), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n528), .A2(G67), .ZN(new_n846));
  NAND2_X1  g421(.A1(G80), .A2(G543), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n536), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g423(.A(KEYINPUT96), .B1(new_n845), .B2(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(G67), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n850), .B1(new_n509), .B2(new_n510), .ZN(new_n851));
  INV_X1    g426(.A(new_n847), .ZN(new_n852));
  OAI21_X1  g427(.A(G651), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT96), .ZN(new_n854));
  NAND4_X1  g429(.A1(new_n853), .A2(new_n843), .A3(new_n854), .A4(new_n844), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n849), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n856), .A2(new_n556), .ZN(new_n857));
  NAND4_X1  g432(.A1(new_n849), .A2(new_n554), .A3(new_n555), .A4(new_n855), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  XOR2_X1   g434(.A(new_n859), .B(KEYINPUT38), .Z(new_n860));
  NAND2_X1  g435(.A1(new_n625), .A2(G559), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n860), .B(new_n861), .ZN(new_n862));
  OR2_X1    g437(.A1(new_n862), .A2(KEYINPUT39), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(KEYINPUT39), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n863), .A2(new_n634), .A3(new_n864), .ZN(new_n865));
  OAI21_X1  g440(.A(G860), .B1(new_n845), .B2(new_n848), .ZN(new_n866));
  XOR2_X1   g441(.A(new_n866), .B(KEYINPUT37), .Z(new_n867));
  NAND2_X1  g442(.A1(new_n865), .A2(new_n867), .ZN(G145));
  INV_X1    g443(.A(G37), .ZN(new_n869));
  OAI21_X1  g444(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n870));
  OR2_X1    g445(.A1(new_n870), .A2(KEYINPUT99), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(KEYINPUT99), .ZN(new_n872));
  OR3_X1    g447(.A1(new_n468), .A2(KEYINPUT98), .A3(G118), .ZN(new_n873));
  OAI21_X1  g448(.A(KEYINPUT98), .B1(new_n468), .B2(G118), .ZN(new_n874));
  NAND4_X1  g449(.A1(new_n871), .A2(new_n872), .A3(new_n873), .A4(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(G130), .ZN(new_n876));
  INV_X1    g451(.A(G142), .ZN(new_n877));
  OAI221_X1 g452(.A(new_n875), .B1(new_n791), .B2(new_n876), .C1(new_n877), .C2(new_n483), .ZN(new_n878));
  AND2_X1   g453(.A1(new_n878), .A2(new_n651), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n878), .A2(new_n651), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n881), .A2(new_n827), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n826), .B1(new_n879), .B2(new_n880), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n732), .A2(new_n499), .ZN(new_n885));
  INV_X1    g460(.A(new_n499), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n730), .A2(new_n886), .A3(new_n731), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n796), .A2(new_n888), .ZN(new_n889));
  OAI211_X1 g464(.A(new_n887), .B(new_n885), .C1(new_n785), .C2(new_n795), .ZN(new_n890));
  OR2_X1    g465(.A1(new_n751), .A2(KEYINPUT97), .ZN(new_n891));
  AND3_X1   g466(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n751), .A2(KEYINPUT97), .ZN(new_n893));
  AOI22_X1  g468(.A1(new_n889), .A2(new_n890), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  OAI211_X1 g469(.A(KEYINPUT100), .B(new_n884), .C1(new_n892), .C2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n889), .A2(new_n890), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n891), .A2(new_n893), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n884), .A2(KEYINPUT100), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT100), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n882), .A2(new_n901), .A3(new_n883), .ZN(new_n902));
  NAND4_X1  g477(.A1(new_n898), .A2(new_n899), .A3(new_n900), .A4(new_n902), .ZN(new_n903));
  OR2_X1    g478(.A1(new_n486), .A2(G160), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n486), .A2(G160), .ZN(new_n905));
  AND3_X1   g480(.A1(new_n904), .A2(new_n646), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n646), .B1(new_n904), .B2(new_n905), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n895), .A2(new_n903), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n908), .B1(new_n895), .B2(new_n903), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n910), .A2(KEYINPUT101), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT101), .ZN(new_n912));
  AOI211_X1 g487(.A(new_n912), .B(new_n908), .C1(new_n895), .C2(new_n903), .ZN(new_n913));
  OAI211_X1 g488(.A(new_n869), .B(new_n909), .C1(new_n911), .C2(new_n913), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n914), .B(KEYINPUT40), .ZN(G395));
  OAI21_X1  g490(.A(new_n628), .B1(new_n845), .B2(new_n848), .ZN(new_n916));
  XOR2_X1   g491(.A(new_n859), .B(new_n638), .Z(new_n917));
  NAND2_X1  g492(.A1(new_n624), .A2(new_n630), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT102), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g495(.A1(G299), .A2(new_n613), .A3(new_n623), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n624), .A2(KEYINPUT102), .A3(new_n630), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n920), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n917), .A2(new_n923), .ZN(new_n924));
  XOR2_X1   g499(.A(new_n924), .B(KEYINPUT103), .Z(new_n925));
  INV_X1    g500(.A(KEYINPUT41), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n922), .A2(new_n921), .ZN(new_n927));
  AOI21_X1  g502(.A(KEYINPUT102), .B1(new_n624), .B2(new_n630), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n926), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT104), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n923), .A2(KEYINPUT104), .A3(new_n926), .ZN(new_n932));
  XNOR2_X1  g507(.A(KEYINPUT105), .B(KEYINPUT41), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  NAND4_X1  g509(.A1(new_n920), .A2(new_n921), .A3(new_n922), .A4(new_n934), .ZN(new_n935));
  AND3_X1   g510(.A1(new_n931), .A2(new_n932), .A3(new_n935), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n925), .B1(new_n917), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n833), .A2(G166), .ZN(new_n938));
  NAND2_X1  g513(.A1(G290), .A2(G303), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  XNOR2_X1  g515(.A(new_n815), .B(new_n802), .ZN(new_n941));
  AND2_X1   g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n940), .A2(new_n941), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n944), .A2(KEYINPUT106), .ZN(new_n945));
  XOR2_X1   g520(.A(new_n945), .B(KEYINPUT42), .Z(new_n946));
  XNOR2_X1  g521(.A(new_n937), .B(new_n946), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n916), .B1(new_n947), .B2(new_n628), .ZN(G295));
  OAI21_X1  g523(.A(new_n916), .B1(new_n947), .B2(new_n628), .ZN(G331));
  INV_X1    g524(.A(KEYINPUT43), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT110), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT109), .ZN(new_n952));
  NAND2_X1  g527(.A1(G301), .A2(G286), .ZN(new_n953));
  OAI211_X1 g528(.A(G168), .B(new_n537), .C1(new_n545), .C2(new_n543), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n859), .A2(new_n955), .ZN(new_n956));
  NAND4_X1  g531(.A1(new_n857), .A2(new_n953), .A3(new_n858), .A4(new_n954), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n956), .A2(KEYINPUT107), .A3(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT107), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n859), .A2(new_n955), .A3(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  AOI22_X1  g536(.A1(new_n923), .A2(new_n934), .B1(new_n956), .B2(new_n957), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n923), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(KEYINPUT41), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(new_n944), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n952), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  AOI211_X1 g542(.A(KEYINPUT109), .B(new_n944), .C1(new_n963), .C2(new_n964), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n923), .A2(new_n956), .A3(new_n957), .ZN(new_n970));
  OAI211_X1 g545(.A(new_n944), .B(new_n970), .C1(new_n936), .C2(new_n961), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(KEYINPUT108), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n931), .A2(new_n932), .A3(new_n935), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n973), .A2(new_n960), .A3(new_n958), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT108), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n974), .A2(new_n975), .A3(new_n944), .A4(new_n970), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n972), .A2(new_n869), .A3(new_n976), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n951), .B1(new_n969), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n923), .A2(new_n934), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n956), .A2(new_n957), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n981), .A2(new_n960), .A3(new_n958), .ZN(new_n982));
  AOI22_X1  g557(.A1(new_n982), .A2(new_n923), .B1(KEYINPUT41), .B2(new_n962), .ZN(new_n983));
  OAI21_X1  g558(.A(KEYINPUT109), .B1(new_n983), .B2(new_n944), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n965), .A2(new_n952), .A3(new_n966), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(G37), .B1(new_n971), .B2(KEYINPUT108), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n986), .A2(KEYINPUT110), .A3(new_n976), .A4(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n950), .B1(new_n978), .B2(new_n988), .ZN(new_n989));
  AND2_X1   g564(.A1(new_n974), .A2(new_n970), .ZN(new_n990));
  OAI211_X1 g565(.A(new_n987), .B(new_n976), .C1(new_n944), .C2(new_n990), .ZN(new_n991));
  AND2_X1   g566(.A1(new_n991), .A2(new_n950), .ZN(new_n992));
  OAI21_X1  g567(.A(KEYINPUT44), .B1(new_n989), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n991), .A2(KEYINPUT43), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n986), .A2(new_n976), .A3(new_n987), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n994), .B1(new_n995), .B2(KEYINPUT43), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT44), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n993), .A2(new_n998), .ZN(G397));
  INV_X1    g574(.A(G1384), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n499), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(new_n474), .ZN(new_n1003));
  OAI211_X1 g578(.A(new_n1003), .B(G40), .C1(new_n466), .C2(G2105), .ZN(new_n1004));
  NOR3_X1   g579(.A1(new_n1002), .A2(new_n1004), .A3(KEYINPUT45), .ZN(new_n1005));
  XNOR2_X1  g580(.A(new_n796), .B(G1996), .ZN(new_n1006));
  INV_X1    g581(.A(G2067), .ZN(new_n1007));
  XNOR2_X1  g582(.A(new_n732), .B(new_n1007), .ZN(new_n1008));
  XNOR2_X1  g583(.A(new_n826), .B(new_n830), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1006), .A2(new_n1008), .A3(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n833), .A2(new_n832), .ZN(new_n1011));
  NAND2_X1  g586(.A1(G290), .A2(G1986), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1005), .B1(new_n1010), .B2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n524), .A2(new_n525), .A3(G8), .ZN(new_n1015));
  XNOR2_X1  g590(.A(new_n1015), .B(KEYINPUT55), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1016), .ZN(new_n1017));
  AND3_X1   g592(.A1(new_n501), .A2(new_n502), .A3(new_n490), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n502), .B1(new_n501), .B2(new_n490), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1000), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT45), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g597(.A(KEYINPUT111), .B1(new_n1001), .B2(new_n1021), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1004), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1020), .A2(KEYINPUT111), .A3(new_n1021), .ZN(new_n1025));
  AOI21_X1  g600(.A(G1971), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(G40), .ZN(new_n1027));
  NOR3_X1   g602(.A1(new_n467), .A2(new_n1027), .A3(new_n474), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1028), .B1(KEYINPUT50), .B2(new_n1001), .ZN(new_n1029));
  AOI21_X1  g604(.A(G1384), .B1(new_n500), .B2(new_n503), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT50), .ZN(new_n1031));
  OAI21_X1  g606(.A(KEYINPUT112), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT112), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1020), .A2(new_n1033), .A3(KEYINPUT50), .ZN(new_n1034));
  AOI211_X1 g609(.A(G2090), .B(new_n1029), .C1(new_n1032), .C2(new_n1034), .ZN(new_n1035));
  OAI211_X1 g610(.A(G8), .B(new_n1017), .C1(new_n1026), .C2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n813), .A2(G1976), .A3(new_n814), .ZN(new_n1037));
  OAI21_X1  g612(.A(G8), .B1(new_n1004), .B2(new_n1001), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(G1976), .ZN(new_n1040));
  AOI21_X1  g615(.A(KEYINPUT52), .B1(G288), .B2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1037), .A2(new_n1039), .A3(new_n1041), .ZN(new_n1042));
  AND3_X1   g617(.A1(new_n582), .A2(KEYINPUT87), .A3(new_n585), .ZN(new_n1043));
  AOI21_X1  g618(.A(KEYINPUT87), .B1(new_n582), .B2(new_n585), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1038), .B1(new_n1045), .B2(G1976), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT52), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1042), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT113), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n520), .A2(G48), .ZN(new_n1050));
  AOI22_X1  g625(.A1(new_n528), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n1051));
  OAI211_X1 g626(.A(new_n593), .B(new_n1050), .C1(new_n1051), .C2(new_n536), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1049), .B1(new_n1052), .B2(G1981), .ZN(new_n1053));
  INV_X1    g628(.A(G1981), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n592), .A2(new_n1054), .A3(new_n595), .A4(new_n596), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1053), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT49), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1052), .A2(new_n1049), .A3(G1981), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1056), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(KEYINPUT114), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT114), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1056), .A2(new_n1061), .A3(new_n1057), .A4(new_n1058), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1060), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1038), .B1(new_n1064), .B2(KEYINPUT49), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1048), .B1(new_n1063), .B2(new_n1065), .ZN(new_n1066));
  AND2_X1   g641(.A1(new_n1036), .A2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1029), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1030), .A2(KEYINPUT45), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1004), .B1(new_n1021), .B2(new_n1001), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  AOI22_X1  g646(.A1(new_n1068), .A2(new_n764), .B1(new_n721), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(G8), .ZN(new_n1073));
  NOR3_X1   g648(.A1(new_n1072), .A2(new_n1073), .A3(G286), .ZN(new_n1074));
  OAI21_X1  g649(.A(G8), .B1(new_n1026), .B2(new_n1035), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(new_n1016), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1067), .A2(KEYINPUT63), .A3(new_n1074), .A4(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT116), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1036), .A2(new_n1066), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT115), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1004), .B1(KEYINPUT50), .B2(new_n1001), .ZN(new_n1081));
  OAI211_X1 g656(.A(new_n1031), .B(new_n1000), .C1(new_n1018), .C2(new_n1019), .ZN(new_n1082));
  AND3_X1   g657(.A1(new_n1081), .A2(new_n705), .A3(new_n1082), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1080), .B1(new_n1026), .B2(new_n1083), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1023), .B1(new_n1030), .B2(KEYINPUT45), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1085), .A2(new_n1028), .A3(new_n1025), .ZN(new_n1086));
  INV_X1    g661(.A(G1971), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1083), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(KEYINPUT115), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1084), .A2(new_n1089), .A3(G8), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1079), .B1(new_n1016), .B2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1078), .B1(new_n1091), .B2(new_n1074), .ZN(new_n1092));
  OAI21_X1  g667(.A(G8), .B1(new_n1088), .B2(KEYINPUT115), .ZN(new_n1093));
  AOI211_X1 g668(.A(new_n1080), .B(new_n1083), .C1(new_n1086), .C2(new_n1087), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1016), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1067), .A2(new_n1095), .A3(new_n1078), .A4(new_n1074), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT63), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1077), .B1(new_n1092), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT117), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n582), .A2(new_n1040), .A3(new_n585), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1055), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1036), .ZN(new_n1105));
  AOI22_X1  g680(.A1(new_n1104), .A2(new_n1039), .B1(new_n1105), .B2(new_n1066), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1099), .A2(new_n1100), .A3(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1071), .A2(new_n721), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1029), .ZN(new_n1109));
  NOR3_X1   g684(.A1(new_n1030), .A2(KEYINPUT112), .A3(new_n1031), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1033), .B1(new_n1020), .B2(KEYINPUT50), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1109), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  OAI211_X1 g687(.A(new_n1108), .B(G168), .C1(new_n1112), .C2(G2084), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(G8), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1068), .A2(new_n764), .ZN(new_n1115));
  AOI21_X1  g690(.A(G168), .B1(new_n1115), .B2(new_n1108), .ZN(new_n1116));
  OAI21_X1  g691(.A(KEYINPUT51), .B1(new_n1114), .B2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT62), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT51), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1113), .A2(new_n1119), .A3(G8), .ZN(new_n1120));
  AND3_X1   g695(.A1(new_n1117), .A2(new_n1118), .A3(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1118), .B1(new_n1117), .B2(new_n1120), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1024), .A2(new_n756), .A3(new_n1025), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT53), .ZN(new_n1124));
  XNOR2_X1  g699(.A(KEYINPUT127), .B(G1961), .ZN(new_n1125));
  AOI22_X1  g700(.A1(new_n1123), .A2(new_n1124), .B1(new_n1112), .B2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1069), .A2(new_n756), .A3(new_n1070), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT126), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1124), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1129), .B1(new_n1128), .B2(new_n1127), .ZN(new_n1130));
  AOI21_X1  g705(.A(G301), .B1(new_n1126), .B2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1067), .A2(new_n1095), .A3(new_n1131), .ZN(new_n1132));
  NOR3_X1   g707(.A1(new_n1121), .A2(new_n1122), .A3(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1028), .A2(new_n1007), .A3(new_n1002), .ZN(new_n1134));
  OAI211_X1 g709(.A(KEYINPUT60), .B(new_n1134), .C1(new_n1068), .C2(G1348), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT124), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n625), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(G1348), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1112), .A2(new_n1139), .ZN(new_n1140));
  XNOR2_X1  g715(.A(new_n624), .B(new_n1136), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1140), .A2(KEYINPUT60), .A3(new_n1134), .A4(new_n1141), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1134), .B1(new_n1068), .B2(G1348), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT60), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1138), .A2(new_n1142), .A3(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT125), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1138), .A2(new_n1142), .A3(KEYINPUT125), .A4(new_n1145), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT61), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT119), .ZN(new_n1152));
  XOR2_X1   g727(.A(KEYINPUT56), .B(G2072), .Z(new_n1153));
  OAI21_X1  g728(.A(new_n1152), .B1(new_n1086), .B2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1153), .ZN(new_n1155));
  NAND4_X1  g730(.A1(new_n1024), .A2(KEYINPUT119), .A3(new_n1025), .A4(new_n1155), .ZN(new_n1156));
  AND2_X1   g731(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1157));
  OR2_X1    g732(.A1(new_n1157), .A2(G1956), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1154), .A2(new_n1156), .A3(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT57), .ZN(new_n1160));
  AOI21_X1  g735(.A(G299), .B1(KEYINPUT118), .B2(new_n1160), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1161), .B1(KEYINPUT118), .B2(new_n1160), .ZN(new_n1162));
  OR3_X1    g737(.A1(new_n630), .A2(KEYINPUT118), .A3(new_n1160), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1159), .A2(KEYINPUT123), .A3(new_n1164), .ZN(new_n1165));
  AND2_X1   g740(.A1(new_n1159), .A2(new_n1164), .ZN(new_n1166));
  INV_X1    g741(.A(new_n1164), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1154), .A2(new_n1167), .A3(new_n1158), .A4(new_n1156), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT123), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  OAI211_X1 g745(.A(new_n1151), .B(new_n1165), .C1(new_n1166), .C2(new_n1170), .ZN(new_n1171));
  XOR2_X1   g746(.A(KEYINPUT121), .B(G1996), .Z(new_n1172));
  NAND4_X1  g747(.A1(new_n1085), .A2(new_n1028), .A3(new_n1025), .A4(new_n1172), .ZN(new_n1173));
  XOR2_X1   g748(.A(KEYINPUT58), .B(G1341), .Z(new_n1174));
  OAI21_X1  g749(.A(new_n1174), .B1(new_n1004), .B2(new_n1001), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1173), .A2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n556), .B1(KEYINPUT122), .B2(KEYINPUT59), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  NOR2_X1   g753(.A1(KEYINPUT122), .A2(KEYINPUT59), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  OAI211_X1 g755(.A(new_n1176), .B(new_n1177), .C1(KEYINPUT122), .C2(KEYINPUT59), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1164), .A2(KEYINPUT120), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT120), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1162), .A2(new_n1184), .A3(new_n1163), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1183), .A2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1151), .B1(new_n1159), .B2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1182), .B1(new_n1168), .B2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1150), .A2(new_n1171), .A3(new_n1188), .ZN(new_n1189));
  AND2_X1   g764(.A1(new_n1159), .A2(new_n1186), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n624), .B1(new_n1140), .B2(new_n1134), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1168), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1189), .A2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1117), .A2(new_n1120), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1126), .A2(new_n1130), .ZN(new_n1195));
  XNOR2_X1  g770(.A(G301), .B(KEYINPUT54), .ZN(new_n1196));
  AOI211_X1 g771(.A(new_n1124), .B(G2078), .C1(new_n1002), .C2(KEYINPUT45), .ZN(new_n1197));
  AOI21_X1  g772(.A(new_n1196), .B1(new_n1070), .B2(new_n1197), .ZN(new_n1198));
  AOI22_X1  g773(.A1(new_n1195), .A2(new_n1196), .B1(new_n1126), .B2(new_n1198), .ZN(new_n1199));
  AND3_X1   g774(.A1(new_n1091), .A2(new_n1194), .A3(new_n1199), .ZN(new_n1200));
  AOI21_X1  g775(.A(new_n1133), .B1(new_n1193), .B2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1107), .A2(new_n1201), .ZN(new_n1202));
  AOI21_X1  g777(.A(new_n1100), .B1(new_n1099), .B2(new_n1106), .ZN(new_n1203));
  OAI21_X1  g778(.A(new_n1014), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  AND4_X1   g779(.A1(new_n827), .A2(new_n1006), .A3(new_n830), .A4(new_n1008), .ZN(new_n1205));
  NOR2_X1   g780(.A1(new_n732), .A2(G2067), .ZN(new_n1206));
  OAI21_X1  g781(.A(new_n1005), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  INV_X1    g782(.A(G1996), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1005), .A2(new_n1208), .ZN(new_n1209));
  XOR2_X1   g784(.A(new_n1209), .B(KEYINPUT46), .Z(new_n1210));
  NAND2_X1  g785(.A1(new_n796), .A2(new_n1008), .ZN(new_n1211));
  AOI21_X1  g786(.A(new_n1210), .B1(new_n1211), .B2(new_n1005), .ZN(new_n1212));
  XOR2_X1   g787(.A(new_n1212), .B(KEYINPUT47), .Z(new_n1213));
  NAND2_X1  g788(.A1(new_n1207), .A2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1010), .A2(new_n1005), .ZN(new_n1215));
  NAND3_X1  g790(.A1(new_n833), .A2(new_n1005), .A3(new_n832), .ZN(new_n1216));
  XNOR2_X1  g791(.A(new_n1216), .B(KEYINPUT48), .ZN(new_n1217));
  AOI21_X1  g792(.A(new_n1214), .B1(new_n1215), .B2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g793(.A1(new_n1204), .A2(new_n1218), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g794(.A1(G401), .A2(new_n459), .A3(G227), .ZN(new_n1221));
  NAND4_X1  g795(.A1(new_n996), .A2(new_n914), .A3(new_n699), .A4(new_n1221), .ZN(G225));
  INV_X1    g796(.A(G225), .ZN(G308));
endmodule


