

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591;

  NOR2_X1 U326 ( .A1(n554), .A2(n441), .ZN(n576) );
  XNOR2_X1 U327 ( .A(KEYINPUT100), .B(n473), .ZN(n554) );
  XNOR2_X1 U328 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U329 ( .A(n439), .B(n438), .ZN(n553) );
  XNOR2_X1 U330 ( .A(n422), .B(n421), .ZN(n426) );
  XNOR2_X1 U331 ( .A(KEYINPUT123), .B(n460), .ZN(n572) );
  NOR2_X1 U332 ( .A1(n521), .A2(n509), .ZN(n517) );
  XNOR2_X1 U333 ( .A(n458), .B(n457), .ZN(n537) );
  XNOR2_X1 U334 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U335 ( .A(n464), .B(n463), .ZN(G1349GAT) );
  XOR2_X1 U336 ( .A(G148GAT), .B(KEYINPUT22), .Z(n297) );
  XOR2_X1 U337 ( .A(G50GAT), .B(KEYINPUT76), .Z(n357) );
  XOR2_X1 U338 ( .A(G78GAT), .B(G204GAT), .Z(n295) );
  XNOR2_X1 U339 ( .A(G106GAT), .B(KEYINPUT73), .ZN(n294) );
  XNOR2_X1 U340 ( .A(n295), .B(n294), .ZN(n424) );
  XNOR2_X1 U341 ( .A(n357), .B(n424), .ZN(n296) );
  XNOR2_X1 U342 ( .A(n297), .B(n296), .ZN(n301) );
  XOR2_X1 U343 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n299) );
  NAND2_X1 U344 ( .A1(G228GAT), .A2(G233GAT), .ZN(n298) );
  XNOR2_X1 U345 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U346 ( .A(n301), .B(n300), .Z(n307) );
  XNOR2_X1 U347 ( .A(G155GAT), .B(KEYINPUT93), .ZN(n302) );
  XNOR2_X1 U348 ( .A(n302), .B(KEYINPUT3), .ZN(n303) );
  XOR2_X1 U349 ( .A(n303), .B(KEYINPUT2), .Z(n305) );
  XNOR2_X1 U350 ( .A(G141GAT), .B(G162GAT), .ZN(n304) );
  XNOR2_X1 U351 ( .A(n305), .B(n304), .ZN(n320) );
  XNOR2_X1 U352 ( .A(G22GAT), .B(n320), .ZN(n306) );
  XNOR2_X1 U353 ( .A(n307), .B(n306), .ZN(n311) );
  XOR2_X1 U354 ( .A(KEYINPUT92), .B(G218GAT), .Z(n309) );
  XNOR2_X1 U355 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n308) );
  XNOR2_X1 U356 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U357 ( .A(G197GAT), .B(n310), .ZN(n335) );
  XNOR2_X1 U358 ( .A(n311), .B(n335), .ZN(n475) );
  XNOR2_X1 U359 ( .A(G29GAT), .B(G134GAT), .ZN(n312) );
  XNOR2_X1 U360 ( .A(n312), .B(KEYINPUT82), .ZN(n346) );
  XNOR2_X1 U361 ( .A(G120GAT), .B(G148GAT), .ZN(n313) );
  XNOR2_X1 U362 ( .A(n313), .B(G57GAT), .ZN(n408) );
  XNOR2_X1 U363 ( .A(n346), .B(n408), .ZN(n330) );
  XOR2_X1 U364 ( .A(KEYINPUT97), .B(KEYINPUT1), .Z(n315) );
  XNOR2_X1 U365 ( .A(KEYINPUT6), .B(KEYINPUT95), .ZN(n314) );
  XNOR2_X1 U366 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U367 ( .A(KEYINPUT4), .B(n316), .Z(n318) );
  NAND2_X1 U368 ( .A1(G225GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U369 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U370 ( .A(n319), .B(KEYINPUT98), .Z(n322) );
  XNOR2_X1 U371 ( .A(n320), .B(KEYINPUT96), .ZN(n321) );
  XNOR2_X1 U372 ( .A(n322), .B(n321), .ZN(n326) );
  XOR2_X1 U373 ( .A(KEYINPUT5), .B(KEYINPUT94), .Z(n324) );
  XNOR2_X1 U374 ( .A(G85GAT), .B(KEYINPUT99), .ZN(n323) );
  XNOR2_X1 U375 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U376 ( .A(n326), .B(n325), .Z(n328) );
  XOR2_X1 U377 ( .A(G113GAT), .B(KEYINPUT0), .Z(n446) );
  XOR2_X1 U378 ( .A(G1GAT), .B(G127GAT), .Z(n373) );
  XNOR2_X1 U379 ( .A(n446), .B(n373), .ZN(n327) );
  XNOR2_X1 U380 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U381 ( .A(n330), .B(n329), .ZN(n473) );
  XNOR2_X1 U382 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n331) );
  XNOR2_X1 U383 ( .A(n331), .B(KEYINPUT90), .ZN(n332) );
  XOR2_X1 U384 ( .A(n332), .B(KEYINPUT19), .Z(n334) );
  XNOR2_X1 U385 ( .A(G169GAT), .B(KEYINPUT89), .ZN(n333) );
  XNOR2_X1 U386 ( .A(n334), .B(n333), .ZN(n456) );
  INV_X1 U387 ( .A(n335), .ZN(n336) );
  XNOR2_X1 U388 ( .A(n456), .B(n336), .ZN(n344) );
  XNOR2_X1 U389 ( .A(G36GAT), .B(G190GAT), .ZN(n337) );
  XNOR2_X1 U390 ( .A(n337), .B(G92GAT), .ZN(n345) );
  XOR2_X1 U391 ( .A(G176GAT), .B(G64GAT), .Z(n407) );
  XOR2_X1 U392 ( .A(n345), .B(n407), .Z(n339) );
  NAND2_X1 U393 ( .A1(G226GAT), .A2(G233GAT), .ZN(n338) );
  XNOR2_X1 U394 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U395 ( .A(G8GAT), .B(G183GAT), .Z(n370) );
  XOR2_X1 U396 ( .A(n340), .B(n370), .Z(n342) );
  XNOR2_X1 U397 ( .A(G204GAT), .B(KEYINPUT101), .ZN(n341) );
  XNOR2_X1 U398 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U399 ( .A(n344), .B(n343), .ZN(n469) );
  XNOR2_X1 U400 ( .A(n346), .B(n345), .ZN(n365) );
  XOR2_X1 U401 ( .A(KEYINPUT11), .B(KEYINPUT10), .Z(n348) );
  XNOR2_X1 U402 ( .A(G162GAT), .B(KEYINPUT80), .ZN(n347) );
  XNOR2_X1 U403 ( .A(n348), .B(n347), .ZN(n352) );
  XOR2_X1 U404 ( .A(KEYINPUT77), .B(KEYINPUT9), .Z(n350) );
  XNOR2_X1 U405 ( .A(KEYINPUT79), .B(KEYINPUT81), .ZN(n349) );
  XNOR2_X1 U406 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U407 ( .A(n352), .B(n351), .Z(n363) );
  XNOR2_X1 U408 ( .A(G43GAT), .B(KEYINPUT8), .ZN(n353) );
  XNOR2_X1 U409 ( .A(n353), .B(KEYINPUT7), .ZN(n404) );
  XOR2_X1 U410 ( .A(G106GAT), .B(n404), .Z(n355) );
  NAND2_X1 U411 ( .A1(G232GAT), .A2(G233GAT), .ZN(n354) );
  XNOR2_X1 U412 ( .A(n355), .B(n354), .ZN(n361) );
  XNOR2_X1 U413 ( .A(G99GAT), .B(G85GAT), .ZN(n356) );
  XNOR2_X1 U414 ( .A(n356), .B(KEYINPUT74), .ZN(n416) );
  XOR2_X1 U415 ( .A(KEYINPUT78), .B(n416), .Z(n359) );
  XNOR2_X1 U416 ( .A(G218GAT), .B(n357), .ZN(n358) );
  XNOR2_X1 U417 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U418 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U419 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U420 ( .A(n365), .B(n364), .ZN(n570) );
  XOR2_X1 U421 ( .A(KEYINPUT13), .B(KEYINPUT70), .Z(n367) );
  XNOR2_X1 U422 ( .A(G71GAT), .B(KEYINPUT71), .ZN(n366) );
  XNOR2_X1 U423 ( .A(n367), .B(n366), .ZN(n423) );
  XOR2_X1 U424 ( .A(KEYINPUT12), .B(n423), .Z(n369) );
  NAND2_X1 U425 ( .A1(G231GAT), .A2(G233GAT), .ZN(n368) );
  XNOR2_X1 U426 ( .A(n369), .B(n368), .ZN(n371) );
  XOR2_X1 U427 ( .A(n371), .B(n370), .Z(n375) );
  XNOR2_X1 U428 ( .A(G22GAT), .B(G15GAT), .ZN(n372) );
  XNOR2_X1 U429 ( .A(n372), .B(KEYINPUT69), .ZN(n403) );
  XNOR2_X1 U430 ( .A(n403), .B(n373), .ZN(n374) );
  XNOR2_X1 U431 ( .A(n375), .B(n374), .ZN(n379) );
  XOR2_X1 U432 ( .A(G64GAT), .B(G78GAT), .Z(n377) );
  XNOR2_X1 U433 ( .A(G211GAT), .B(G155GAT), .ZN(n376) );
  XNOR2_X1 U434 ( .A(n377), .B(n376), .ZN(n378) );
  XOR2_X1 U435 ( .A(n379), .B(n378), .Z(n387) );
  XOR2_X1 U436 ( .A(KEYINPUT86), .B(KEYINPUT85), .Z(n381) );
  XNOR2_X1 U437 ( .A(KEYINPUT84), .B(KEYINPUT14), .ZN(n380) );
  XNOR2_X1 U438 ( .A(n381), .B(n380), .ZN(n385) );
  XOR2_X1 U439 ( .A(KEYINPUT83), .B(KEYINPUT87), .Z(n383) );
  XNOR2_X1 U440 ( .A(G57GAT), .B(KEYINPUT15), .ZN(n382) );
  XNOR2_X1 U441 ( .A(n383), .B(n382), .ZN(n384) );
  XNOR2_X1 U442 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U443 ( .A(n387), .B(n386), .ZN(n561) );
  NAND2_X1 U444 ( .A1(n570), .A2(n561), .ZN(n431) );
  XNOR2_X1 U445 ( .A(KEYINPUT46), .B(KEYINPUT116), .ZN(n429) );
  XOR2_X1 U446 ( .A(G197GAT), .B(G36GAT), .Z(n389) );
  XNOR2_X1 U447 ( .A(G50GAT), .B(G29GAT), .ZN(n388) );
  XNOR2_X1 U448 ( .A(n389), .B(n388), .ZN(n393) );
  XOR2_X1 U449 ( .A(G8GAT), .B(G113GAT), .Z(n391) );
  XNOR2_X1 U450 ( .A(G169GAT), .B(G141GAT), .ZN(n390) );
  XNOR2_X1 U451 ( .A(n391), .B(n390), .ZN(n392) );
  XOR2_X1 U452 ( .A(n393), .B(n392), .Z(n398) );
  XOR2_X1 U453 ( .A(KEYINPUT30), .B(KEYINPUT68), .Z(n395) );
  NAND2_X1 U454 ( .A1(G229GAT), .A2(G233GAT), .ZN(n394) );
  XNOR2_X1 U455 ( .A(n395), .B(n394), .ZN(n396) );
  XNOR2_X1 U456 ( .A(KEYINPUT67), .B(n396), .ZN(n397) );
  XNOR2_X1 U457 ( .A(n398), .B(n397), .ZN(n402) );
  XOR2_X1 U458 ( .A(KEYINPUT66), .B(KEYINPUT29), .Z(n400) );
  XNOR2_X1 U459 ( .A(G1GAT), .B(KEYINPUT65), .ZN(n399) );
  XNOR2_X1 U460 ( .A(n400), .B(n399), .ZN(n401) );
  XOR2_X1 U461 ( .A(n402), .B(n401), .Z(n406) );
  XNOR2_X1 U462 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U463 ( .A(n406), .B(n405), .ZN(n565) );
  XNOR2_X1 U464 ( .A(n408), .B(n407), .ZN(n412) );
  INV_X1 U465 ( .A(n412), .ZN(n410) );
  AND2_X1 U466 ( .A1(G230GAT), .A2(G233GAT), .ZN(n411) );
  INV_X1 U467 ( .A(n411), .ZN(n409) );
  NAND2_X1 U468 ( .A1(n410), .A2(n409), .ZN(n414) );
  NAND2_X1 U469 ( .A1(n412), .A2(n411), .ZN(n413) );
  NAND2_X1 U470 ( .A1(n414), .A2(n413), .ZN(n415) );
  XNOR2_X1 U471 ( .A(n415), .B(KEYINPUT72), .ZN(n422) );
  XOR2_X1 U472 ( .A(n416), .B(KEYINPUT31), .Z(n420) );
  XOR2_X1 U473 ( .A(KEYINPUT75), .B(KEYINPUT32), .Z(n418) );
  XNOR2_X1 U474 ( .A(G92GAT), .B(KEYINPUT33), .ZN(n417) );
  XNOR2_X1 U475 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U476 ( .A(n424), .B(n423), .Z(n425) );
  XNOR2_X1 U477 ( .A(n426), .B(n425), .ZN(n581) );
  INV_X1 U478 ( .A(KEYINPUT41), .ZN(n427) );
  XNOR2_X1 U479 ( .A(n581), .B(n427), .ZN(n539) );
  NAND2_X1 U480 ( .A1(n565), .A2(n539), .ZN(n428) );
  XOR2_X1 U481 ( .A(n429), .B(n428), .Z(n430) );
  NOR2_X1 U482 ( .A1(n431), .A2(n430), .ZN(n432) );
  XNOR2_X1 U483 ( .A(n432), .B(KEYINPUT47), .ZN(n437) );
  XNOR2_X1 U484 ( .A(KEYINPUT36), .B(n570), .ZN(n589) );
  NOR2_X1 U485 ( .A1(n561), .A2(n589), .ZN(n433) );
  XOR2_X1 U486 ( .A(KEYINPUT45), .B(n433), .Z(n434) );
  NOR2_X1 U487 ( .A1(n581), .A2(n434), .ZN(n435) );
  INV_X1 U488 ( .A(n565), .ZN(n577) );
  NAND2_X1 U489 ( .A1(n435), .A2(n577), .ZN(n436) );
  NAND2_X1 U490 ( .A1(n437), .A2(n436), .ZN(n439) );
  XNOR2_X1 U491 ( .A(KEYINPUT117), .B(KEYINPUT48), .ZN(n438) );
  NOR2_X1 U492 ( .A1(n469), .A2(n553), .ZN(n440) );
  XOR2_X1 U493 ( .A(KEYINPUT54), .B(n440), .Z(n441) );
  NAND2_X1 U494 ( .A1(n475), .A2(n576), .ZN(n442) );
  XNOR2_X1 U495 ( .A(KEYINPUT55), .B(n442), .ZN(n459) );
  XOR2_X1 U496 ( .A(G99GAT), .B(G190GAT), .Z(n444) );
  XNOR2_X1 U497 ( .A(G43GAT), .B(G134GAT), .ZN(n443) );
  XNOR2_X1 U498 ( .A(n444), .B(n443), .ZN(n445) );
  XOR2_X1 U499 ( .A(n446), .B(n445), .Z(n448) );
  NAND2_X1 U500 ( .A1(G227GAT), .A2(G233GAT), .ZN(n447) );
  XNOR2_X1 U501 ( .A(n448), .B(n447), .ZN(n452) );
  XOR2_X1 U502 ( .A(G183GAT), .B(KEYINPUT20), .Z(n450) );
  XNOR2_X1 U503 ( .A(G127GAT), .B(G176GAT), .ZN(n449) );
  XNOR2_X1 U504 ( .A(n450), .B(n449), .ZN(n451) );
  XOR2_X1 U505 ( .A(n452), .B(n451), .Z(n458) );
  XOR2_X1 U506 ( .A(KEYINPUT91), .B(G71GAT), .Z(n454) );
  XNOR2_X1 U507 ( .A(G15GAT), .B(G120GAT), .ZN(n453) );
  XNOR2_X1 U508 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U509 ( .A(n456), .B(n455), .ZN(n457) );
  NAND2_X1 U510 ( .A1(n459), .A2(n537), .ZN(n460) );
  NAND2_X1 U511 ( .A1(n572), .A2(n539), .ZN(n464) );
  XOR2_X1 U512 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n462) );
  XNOR2_X1 U513 ( .A(G176GAT), .B(KEYINPUT126), .ZN(n461) );
  NOR2_X1 U514 ( .A1(n581), .A2(n577), .ZN(n497) );
  INV_X1 U515 ( .A(n469), .ZN(n525) );
  NAND2_X1 U516 ( .A1(n537), .A2(n525), .ZN(n465) );
  NAND2_X1 U517 ( .A1(n475), .A2(n465), .ZN(n466) );
  XNOR2_X1 U518 ( .A(KEYINPUT25), .B(n466), .ZN(n471) );
  XNOR2_X1 U519 ( .A(KEYINPUT26), .B(KEYINPUT102), .ZN(n468) );
  NOR2_X1 U520 ( .A1(n537), .A2(n475), .ZN(n467) );
  XNOR2_X1 U521 ( .A(n468), .B(n467), .ZN(n575) );
  XOR2_X1 U522 ( .A(n469), .B(KEYINPUT27), .Z(n474) );
  NAND2_X1 U523 ( .A1(n575), .A2(n474), .ZN(n552) );
  XNOR2_X1 U524 ( .A(KEYINPUT103), .B(n552), .ZN(n470) );
  NOR2_X1 U525 ( .A1(n471), .A2(n470), .ZN(n472) );
  NOR2_X1 U526 ( .A1(n473), .A2(n472), .ZN(n480) );
  INV_X1 U527 ( .A(n474), .ZN(n477) );
  XOR2_X1 U528 ( .A(n475), .B(KEYINPUT64), .Z(n476) );
  XNOR2_X1 U529 ( .A(KEYINPUT28), .B(n476), .ZN(n532) );
  NOR2_X1 U530 ( .A1(n477), .A2(n532), .ZN(n478) );
  NAND2_X1 U531 ( .A1(n478), .A2(n554), .ZN(n535) );
  NOR2_X1 U532 ( .A1(n537), .A2(n535), .ZN(n479) );
  NOR2_X1 U533 ( .A1(n480), .A2(n479), .ZN(n493) );
  INV_X1 U534 ( .A(n561), .ZN(n584) );
  NAND2_X1 U535 ( .A1(n584), .A2(n570), .ZN(n481) );
  XNOR2_X1 U536 ( .A(n481), .B(KEYINPUT88), .ZN(n482) );
  XNOR2_X1 U537 ( .A(n482), .B(KEYINPUT16), .ZN(n483) );
  NOR2_X1 U538 ( .A1(n493), .A2(n483), .ZN(n508) );
  AND2_X1 U539 ( .A1(n497), .A2(n508), .ZN(n491) );
  NAND2_X1 U540 ( .A1(n554), .A2(n491), .ZN(n487) );
  XOR2_X1 U541 ( .A(KEYINPUT104), .B(KEYINPUT34), .Z(n485) );
  XNOR2_X1 U542 ( .A(G1GAT), .B(KEYINPUT105), .ZN(n484) );
  XNOR2_X1 U543 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U544 ( .A(n487), .B(n486), .ZN(G1324GAT) );
  NAND2_X1 U545 ( .A1(n525), .A2(n491), .ZN(n488) );
  XNOR2_X1 U546 ( .A(n488), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U547 ( .A(G15GAT), .B(KEYINPUT35), .Z(n490) );
  NAND2_X1 U548 ( .A1(n491), .A2(n537), .ZN(n489) );
  XNOR2_X1 U549 ( .A(n490), .B(n489), .ZN(G1326GAT) );
  NAND2_X1 U550 ( .A1(n532), .A2(n491), .ZN(n492) );
  XNOR2_X1 U551 ( .A(n492), .B(G22GAT), .ZN(G1327GAT) );
  NOR2_X1 U552 ( .A1(n493), .A2(n589), .ZN(n494) );
  NAND2_X1 U553 ( .A1(n561), .A2(n494), .ZN(n496) );
  XNOR2_X1 U554 ( .A(KEYINPUT106), .B(KEYINPUT37), .ZN(n495) );
  XNOR2_X1 U555 ( .A(n496), .B(n495), .ZN(n520) );
  NAND2_X1 U556 ( .A1(n520), .A2(n497), .ZN(n498) );
  XOR2_X1 U557 ( .A(KEYINPUT38), .B(n498), .Z(n506) );
  NAND2_X1 U558 ( .A1(n554), .A2(n506), .ZN(n500) );
  XOR2_X1 U559 ( .A(G29GAT), .B(KEYINPUT39), .Z(n499) );
  XNOR2_X1 U560 ( .A(n500), .B(n499), .ZN(G1328GAT) );
  NAND2_X1 U561 ( .A1(n506), .A2(n525), .ZN(n501) );
  XNOR2_X1 U562 ( .A(n501), .B(G36GAT), .ZN(G1329GAT) );
  XNOR2_X1 U563 ( .A(G43GAT), .B(KEYINPUT108), .ZN(n505) );
  XOR2_X1 U564 ( .A(KEYINPUT40), .B(KEYINPUT107), .Z(n503) );
  NAND2_X1 U565 ( .A1(n537), .A2(n506), .ZN(n502) );
  XNOR2_X1 U566 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U567 ( .A(n505), .B(n504), .ZN(G1330GAT) );
  NAND2_X1 U568 ( .A1(n506), .A2(n532), .ZN(n507) );
  XNOR2_X1 U569 ( .A(n507), .B(G50GAT), .ZN(G1331GAT) );
  NAND2_X1 U570 ( .A1(n539), .A2(n577), .ZN(n521) );
  INV_X1 U571 ( .A(n508), .ZN(n509) );
  NAND2_X1 U572 ( .A1(n554), .A2(n517), .ZN(n513) );
  XOR2_X1 U573 ( .A(KEYINPUT109), .B(KEYINPUT42), .Z(n511) );
  XNOR2_X1 U574 ( .A(G57GAT), .B(KEYINPUT110), .ZN(n510) );
  XNOR2_X1 U575 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U576 ( .A(n513), .B(n512), .ZN(G1332GAT) );
  XOR2_X1 U577 ( .A(G64GAT), .B(KEYINPUT111), .Z(n515) );
  NAND2_X1 U578 ( .A1(n517), .A2(n525), .ZN(n514) );
  XNOR2_X1 U579 ( .A(n515), .B(n514), .ZN(G1333GAT) );
  NAND2_X1 U580 ( .A1(n517), .A2(n537), .ZN(n516) );
  XNOR2_X1 U581 ( .A(n516), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U582 ( .A(G78GAT), .B(KEYINPUT43), .Z(n519) );
  NAND2_X1 U583 ( .A1(n517), .A2(n532), .ZN(n518) );
  XNOR2_X1 U584 ( .A(n519), .B(n518), .ZN(G1335GAT) );
  XNOR2_X1 U585 ( .A(G85GAT), .B(KEYINPUT112), .ZN(n524) );
  INV_X1 U586 ( .A(n520), .ZN(n522) );
  NOR2_X1 U587 ( .A1(n522), .A2(n521), .ZN(n531) );
  NAND2_X1 U588 ( .A1(n531), .A2(n554), .ZN(n523) );
  XNOR2_X1 U589 ( .A(n524), .B(n523), .ZN(G1336GAT) );
  XOR2_X1 U590 ( .A(G92GAT), .B(KEYINPUT113), .Z(n527) );
  NAND2_X1 U591 ( .A1(n531), .A2(n525), .ZN(n526) );
  XNOR2_X1 U592 ( .A(n527), .B(n526), .ZN(G1337GAT) );
  XOR2_X1 U593 ( .A(KEYINPUT114), .B(KEYINPUT115), .Z(n529) );
  NAND2_X1 U594 ( .A1(n531), .A2(n537), .ZN(n528) );
  XNOR2_X1 U595 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U596 ( .A(G99GAT), .B(n530), .ZN(G1338GAT) );
  NAND2_X1 U597 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U598 ( .A(n533), .B(KEYINPUT44), .ZN(n534) );
  XNOR2_X1 U599 ( .A(G106GAT), .B(n534), .ZN(G1339GAT) );
  NOR2_X1 U600 ( .A1(n553), .A2(n535), .ZN(n536) );
  NAND2_X1 U601 ( .A1(n537), .A2(n536), .ZN(n547) );
  NOR2_X1 U602 ( .A1(n577), .A2(n547), .ZN(n538) );
  XOR2_X1 U603 ( .A(G113GAT), .B(n538), .Z(G1340GAT) );
  INV_X1 U604 ( .A(n539), .ZN(n557) );
  NOR2_X1 U605 ( .A1(n547), .A2(n557), .ZN(n543) );
  XOR2_X1 U606 ( .A(KEYINPUT118), .B(KEYINPUT49), .Z(n541) );
  XNOR2_X1 U607 ( .A(G120GAT), .B(KEYINPUT119), .ZN(n540) );
  XNOR2_X1 U608 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U609 ( .A(n543), .B(n542), .ZN(G1341GAT) );
  NOR2_X1 U610 ( .A1(n561), .A2(n547), .ZN(n545) );
  XNOR2_X1 U611 ( .A(KEYINPUT120), .B(KEYINPUT50), .ZN(n544) );
  XNOR2_X1 U612 ( .A(n545), .B(n544), .ZN(n546) );
  XOR2_X1 U613 ( .A(G127GAT), .B(n546), .Z(G1342GAT) );
  NOR2_X1 U614 ( .A1(n547), .A2(n570), .ZN(n551) );
  XOR2_X1 U615 ( .A(KEYINPUT121), .B(KEYINPUT51), .Z(n549) );
  XNOR2_X1 U616 ( .A(G134GAT), .B(KEYINPUT122), .ZN(n548) );
  XNOR2_X1 U617 ( .A(n549), .B(n548), .ZN(n550) );
  XNOR2_X1 U618 ( .A(n551), .B(n550), .ZN(G1343GAT) );
  NOR2_X1 U619 ( .A1(n553), .A2(n552), .ZN(n555) );
  NAND2_X1 U620 ( .A1(n555), .A2(n554), .ZN(n563) );
  NOR2_X1 U621 ( .A1(n577), .A2(n563), .ZN(n556) );
  XOR2_X1 U622 ( .A(G141GAT), .B(n556), .Z(G1344GAT) );
  NOR2_X1 U623 ( .A1(n557), .A2(n563), .ZN(n559) );
  XNOR2_X1 U624 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U626 ( .A(G148GAT), .B(n560), .ZN(G1345GAT) );
  NOR2_X1 U627 ( .A1(n561), .A2(n563), .ZN(n562) );
  XOR2_X1 U628 ( .A(G155GAT), .B(n562), .Z(G1346GAT) );
  NOR2_X1 U629 ( .A1(n570), .A2(n563), .ZN(n564) );
  XOR2_X1 U630 ( .A(G162GAT), .B(n564), .Z(G1347GAT) );
  NAND2_X1 U631 ( .A1(n572), .A2(n565), .ZN(n568) );
  XOR2_X1 U632 ( .A(G169GAT), .B(KEYINPUT124), .Z(n566) );
  XNOR2_X1 U633 ( .A(KEYINPUT125), .B(n566), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(G1348GAT) );
  NAND2_X1 U635 ( .A1(n584), .A2(n572), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n569), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U637 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n574) );
  INV_X1 U638 ( .A(n570), .ZN(n571) );
  NAND2_X1 U639 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(G1351GAT) );
  NAND2_X1 U641 ( .A1(n576), .A2(n575), .ZN(n588) );
  NOR2_X1 U642 ( .A1(n577), .A2(n588), .ZN(n579) );
  XNOR2_X1 U643 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U645 ( .A(G197GAT), .B(n580), .ZN(G1352GAT) );
  XOR2_X1 U646 ( .A(G204GAT), .B(KEYINPUT61), .Z(n583) );
  INV_X1 U647 ( .A(n588), .ZN(n585) );
  NAND2_X1 U648 ( .A1(n585), .A2(n581), .ZN(n582) );
  XNOR2_X1 U649 ( .A(n583), .B(n582), .ZN(G1353GAT) );
  XOR2_X1 U650 ( .A(G211GAT), .B(KEYINPUT127), .Z(n587) );
  NAND2_X1 U651 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U652 ( .A(n587), .B(n586), .ZN(G1354GAT) );
  NOR2_X1 U653 ( .A1(n589), .A2(n588), .ZN(n590) );
  XOR2_X1 U654 ( .A(KEYINPUT62), .B(n590), .Z(n591) );
  XNOR2_X1 U655 ( .A(G218GAT), .B(n591), .ZN(G1355GAT) );
endmodule

