//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 0 0 1 1 1 0 0 0 0 0 1 0 0 0 1 0 1 1 0 0 1 1 0 1 0 0 0 0 0 0 0 0 1 0 1 1 1 0 1 1 0 0 0 0 1 1 1 1 1 1 0 1 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:14 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n446, new_n448, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n587,
    new_n588, new_n589, new_n591, new_n592, new_n593, new_n594, new_n595,
    new_n596, new_n597, new_n598, new_n599, new_n600, new_n601, new_n602,
    new_n605, new_n606, new_n607, new_n608, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n649, new_n652, new_n653,
    new_n655, new_n656, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XOR2_X1   g017(.A(new_n442), .B(KEYINPUT64), .Z(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  NAND2_X1  g020(.A1(G94), .A2(G452), .ZN(new_n446));
  XNOR2_X1  g021(.A(new_n446), .B(KEYINPUT65), .ZN(G173));
  XNOR2_X1  g022(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n448));
  AND2_X1   g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n448), .B(new_n449), .ZN(G223));
  NAND2_X1  g025(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n449), .A2(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n455), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n457), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n464), .A2(G101), .A3(G2104), .ZN(new_n465));
  XNOR2_X1  g040(.A(KEYINPUT3), .B(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(new_n464), .ZN(new_n467));
  INV_X1    g042(.A(G137), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n465), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n466), .A2(G125), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n464), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n469), .A2(new_n472), .ZN(G160));
  INV_X1    g048(.A(KEYINPUT67), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n467), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n466), .A2(KEYINPUT67), .A3(new_n464), .ZN(new_n476));
  AND2_X1   g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G136), .ZN(new_n478));
  OR2_X1    g053(.A1(G100), .A2(G2105), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n479), .B(G2104), .C1(G112), .C2(new_n464), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n466), .A2(G2105), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT68), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n482), .B(new_n483), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n481), .B1(G124), .B2(new_n484), .ZN(G162));
  INV_X1    g060(.A(KEYINPUT70), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n466), .A2(G126), .A3(G2105), .ZN(new_n487));
  OAI21_X1  g062(.A(KEYINPUT69), .B1(new_n464), .B2(G114), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT69), .ZN(new_n489));
  INV_X1    g064(.A(G114), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n489), .A2(new_n490), .A3(G2105), .ZN(new_n491));
  OR2_X1    g066(.A1(G102), .A2(G2105), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n488), .A2(new_n491), .A3(G2104), .A4(new_n492), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n487), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n466), .A2(G138), .A3(new_n464), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT4), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n466), .A2(new_n497), .A3(G138), .A4(new_n464), .ZN(new_n498));
  AOI22_X1  g073(.A1(new_n486), .A2(new_n494), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n494), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(KEYINPUT70), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(G164));
  INV_X1    g078(.A(G543), .ZN(new_n504));
  OAI21_X1  g079(.A(KEYINPUT72), .B1(new_n504), .B2(KEYINPUT5), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT72), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT5), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n506), .A2(new_n507), .A3(G543), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n505), .A2(new_n508), .B1(KEYINPUT5), .B2(new_n504), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n509), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n510));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(KEYINPUT71), .A2(G651), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT6), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g090(.A1(KEYINPUT71), .A2(KEYINPUT6), .A3(G651), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n504), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G50), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n515), .A2(new_n516), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n509), .A2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(G88), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n518), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  OR2_X1    g097(.A1(new_n512), .A2(new_n522), .ZN(G303));
  INV_X1    g098(.A(G303), .ZN(G166));
  NAND2_X1  g099(.A1(new_n505), .A2(new_n508), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n504), .A2(KEYINPUT5), .ZN(new_n526));
  AND2_X1   g101(.A1(KEYINPUT75), .A2(G89), .ZN(new_n527));
  NOR2_X1   g102(.A1(KEYINPUT75), .A2(G89), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND4_X1  g104(.A1(new_n525), .A2(new_n519), .A3(new_n526), .A4(new_n529), .ZN(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n531), .B(KEYINPUT7), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT76), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n530), .A2(KEYINPUT76), .A3(new_n532), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n506), .B1(new_n507), .B2(G543), .ZN(new_n537));
  NOR3_X1   g112(.A1(new_n504), .A2(KEYINPUT72), .A3(KEYINPUT5), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n526), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(KEYINPUT73), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT73), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n525), .A2(new_n541), .A3(new_n526), .ZN(new_n542));
  AND2_X1   g117(.A1(G63), .A2(G651), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n540), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n504), .B1(new_n519), .B2(KEYINPUT74), .ZN(new_n545));
  INV_X1    g120(.A(KEYINPUT74), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n515), .A2(new_n546), .A3(new_n516), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n545), .A2(G51), .A3(new_n547), .ZN(new_n548));
  NAND4_X1  g123(.A1(new_n535), .A2(new_n536), .A3(new_n544), .A4(new_n548), .ZN(G286));
  INV_X1    g124(.A(G286), .ZN(G168));
  NAND3_X1  g125(.A1(new_n509), .A2(G90), .A3(new_n519), .ZN(new_n551));
  INV_X1    g126(.A(new_n516), .ZN(new_n552));
  AOI21_X1  g127(.A(KEYINPUT6), .B1(KEYINPUT71), .B2(G651), .ZN(new_n553));
  OAI21_X1  g128(.A(KEYINPUT74), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND4_X1  g129(.A1(new_n554), .A2(G52), .A3(new_n547), .A4(G543), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT77), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n551), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(new_n557), .ZN(new_n558));
  AOI21_X1  g133(.A(new_n556), .B1(new_n551), .B2(new_n555), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n540), .A2(G64), .A3(new_n542), .ZN(new_n561));
  NAND2_X1  g136(.A1(G77), .A2(G543), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n511), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n560), .A2(new_n563), .ZN(G171));
  AND3_X1   g139(.A1(new_n525), .A2(new_n541), .A3(new_n526), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n541), .B1(new_n525), .B2(new_n526), .ZN(new_n566));
  INV_X1    g141(.A(G56), .ZN(new_n567));
  NOR3_X1   g142(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(G68), .ZN(new_n569));
  NOR2_X1   g144(.A1(new_n569), .A2(new_n504), .ZN(new_n570));
  OAI21_X1  g145(.A(G651), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n554), .A2(G543), .A3(new_n547), .ZN(new_n572));
  INV_X1    g147(.A(G43), .ZN(new_n573));
  INV_X1    g148(.A(G81), .ZN(new_n574));
  OAI22_X1  g149(.A1(new_n572), .A2(new_n573), .B1(new_n520), .B2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n571), .A2(KEYINPUT78), .A3(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT78), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n540), .A2(G56), .A3(new_n542), .ZN(new_n579));
  INV_X1    g154(.A(new_n570), .ZN(new_n580));
  AOI21_X1  g155(.A(new_n511), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n578), .B1(new_n581), .B2(new_n575), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n577), .A2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n584), .A2(G860), .ZN(G153));
  NAND4_X1  g160(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g161(.A1(G1), .A2(G3), .ZN(new_n587));
  XNOR2_X1  g162(.A(new_n587), .B(KEYINPUT8), .ZN(new_n588));
  NAND4_X1  g163(.A1(G319), .A2(G483), .A3(G661), .A4(new_n588), .ZN(new_n589));
  XNOR2_X1  g164(.A(new_n589), .B(KEYINPUT79), .ZN(G188));
  NAND2_X1  g165(.A1(G78), .A2(G543), .ZN(new_n591));
  INV_X1    g166(.A(G65), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n539), .B2(new_n592), .ZN(new_n593));
  AND2_X1   g168(.A1(new_n509), .A2(new_n519), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n593), .A2(G651), .B1(new_n594), .B2(G91), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT9), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n596), .A2(KEYINPUT80), .ZN(new_n597));
  INV_X1    g172(.A(G53), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n572), .B2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(new_n597), .ZN(new_n600));
  NAND4_X1  g175(.A1(new_n545), .A2(G53), .A3(new_n547), .A4(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n595), .A2(new_n602), .ZN(G299));
  INV_X1    g178(.A(G171), .ZN(G301));
  NAND3_X1  g179(.A1(new_n509), .A2(G87), .A3(new_n519), .ZN(new_n605));
  NAND4_X1  g180(.A1(new_n554), .A2(G49), .A3(new_n547), .A4(G543), .ZN(new_n606));
  AND2_X1   g181(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  AOI21_X1  g182(.A(G74), .B1(new_n540), .B2(new_n542), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n608), .B2(new_n511), .ZN(G288));
  NAND2_X1  g184(.A1(G73), .A2(G543), .ZN(new_n610));
  INV_X1    g185(.A(G61), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n539), .B2(new_n611), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n612), .A2(G651), .B1(G48), .B2(new_n517), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n594), .A2(G86), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(new_n614), .ZN(G305));
  INV_X1    g190(.A(G60), .ZN(new_n616));
  NOR3_X1   g191(.A1(new_n565), .A2(new_n566), .A3(new_n616), .ZN(new_n617));
  INV_X1    g192(.A(G72), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n618), .A2(new_n504), .ZN(new_n619));
  OAI21_X1  g194(.A(KEYINPUT81), .B1(new_n617), .B2(new_n619), .ZN(new_n620));
  NAND3_X1  g195(.A1(new_n540), .A2(G60), .A3(new_n542), .ZN(new_n621));
  INV_X1    g196(.A(KEYINPUT81), .ZN(new_n622));
  INV_X1    g197(.A(new_n619), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n620), .A2(G651), .A3(new_n624), .ZN(new_n625));
  NAND4_X1  g200(.A1(new_n554), .A2(G47), .A3(new_n547), .A4(G543), .ZN(new_n626));
  INV_X1    g201(.A(KEYINPUT82), .ZN(new_n627));
  NAND4_X1  g202(.A1(new_n525), .A2(new_n519), .A3(G85), .A4(new_n526), .ZN(new_n628));
  AND3_X1   g203(.A1(new_n626), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n627), .B1(new_n626), .B2(new_n628), .ZN(new_n630));
  NOR2_X1   g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g206(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n625), .A2(new_n632), .ZN(G290));
  NAND2_X1  g208(.A1(G79), .A2(G543), .ZN(new_n634));
  INV_X1    g209(.A(G66), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n634), .B1(new_n539), .B2(new_n635), .ZN(new_n636));
  AND3_X1   g211(.A1(new_n554), .A2(G543), .A3(new_n547), .ZN(new_n637));
  AOI22_X1  g212(.A1(G651), .A2(new_n636), .B1(new_n637), .B2(G54), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n509), .A2(G92), .A3(new_n519), .ZN(new_n639));
  INV_X1    g214(.A(KEYINPUT10), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND4_X1  g216(.A1(new_n509), .A2(KEYINPUT10), .A3(G92), .A4(new_n519), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n638), .A2(new_n643), .ZN(new_n644));
  INV_X1    g219(.A(G868), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n646), .B1(G171), .B2(new_n645), .ZN(G284));
  OAI21_X1  g222(.A(new_n646), .B1(G171), .B2(new_n645), .ZN(G321));
  NAND2_X1  g223(.A1(G299), .A2(new_n645), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n649), .B1(new_n645), .B2(G168), .ZN(G297));
  OAI21_X1  g225(.A(new_n649), .B1(new_n645), .B2(G168), .ZN(G280));
  INV_X1    g226(.A(new_n644), .ZN(new_n652));
  INV_X1    g227(.A(G559), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n652), .B1(new_n653), .B2(G860), .ZN(G148));
  NAND2_X1  g229(.A1(new_n652), .A2(new_n653), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n655), .A2(G868), .ZN(new_n656));
  OAI21_X1  g231(.A(new_n656), .B1(new_n584), .B2(G868), .ZN(G323));
  XNOR2_X1  g232(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g233(.A1(new_n484), .A2(G123), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n477), .A2(G135), .ZN(new_n660));
  OR2_X1    g235(.A1(G99), .A2(G2105), .ZN(new_n661));
  OAI211_X1 g236(.A(new_n661), .B(G2104), .C1(G111), .C2(new_n464), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n659), .A2(new_n660), .A3(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(G2096), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n464), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n667), .B(KEYINPUT12), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT13), .ZN(new_n669));
  INV_X1    g244(.A(G2100), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n663), .A2(G2096), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n666), .A2(new_n671), .A3(new_n672), .ZN(G156));
  XOR2_X1   g248(.A(KEYINPUT15), .B(G2435), .Z(new_n674));
  XNOR2_X1  g249(.A(KEYINPUT83), .B(G2438), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G2427), .B(G2430), .ZN(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  OR2_X1    g254(.A1(new_n674), .A2(new_n675), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n674), .A2(new_n675), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n680), .A2(new_n677), .A3(new_n681), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n679), .A2(KEYINPUT14), .A3(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(G2443), .B(G2446), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(G1341), .B(G1348), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(G2451), .B(G2454), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT16), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT84), .ZN(new_n690));
  OR2_X1    g265(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n687), .A2(new_n690), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n691), .A2(G14), .A3(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(G401));
  INV_X1    g269(.A(KEYINPUT18), .ZN(new_n695));
  XOR2_X1   g270(.A(G2084), .B(G2090), .Z(new_n696));
  XNOR2_X1  g271(.A(G2067), .B(G2678), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(KEYINPUT17), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n696), .A2(new_n697), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n695), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(new_n670), .ZN(new_n702));
  XOR2_X1   g277(.A(G2072), .B(G2078), .Z(new_n703));
  AOI21_X1  g278(.A(new_n703), .B1(new_n698), .B2(KEYINPUT18), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(new_n665), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n702), .B(new_n705), .ZN(G227));
  XOR2_X1   g281(.A(G1991), .B(G1996), .Z(new_n707));
  XNOR2_X1  g282(.A(G1961), .B(G1966), .ZN(new_n708));
  OR2_X1    g283(.A1(new_n708), .A2(KEYINPUT86), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n708), .A2(KEYINPUT86), .ZN(new_n710));
  XOR2_X1   g285(.A(G1956), .B(G2474), .Z(new_n711));
  NAND3_X1  g286(.A1(new_n709), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(G1971), .B(G1976), .ZN(new_n713));
  XNOR2_X1  g288(.A(KEYINPUT85), .B(KEYINPUT19), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n712), .A2(new_n715), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(KEYINPUT20), .Z(new_n717));
  NAND2_X1  g292(.A1(new_n712), .A2(new_n715), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n709), .A2(new_n710), .ZN(new_n719));
  INV_X1    g294(.A(new_n711), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  MUX2_X1   g296(.A(new_n715), .B(new_n718), .S(new_n721), .Z(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n717), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(new_n724), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n723), .B1(new_n717), .B2(new_n722), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n707), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(new_n726), .ZN(new_n728));
  INV_X1    g303(.A(new_n707), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n728), .A2(new_n729), .A3(new_n724), .ZN(new_n730));
  XNOR2_X1  g305(.A(G1981), .B(G1986), .ZN(new_n731));
  AND3_X1   g306(.A1(new_n727), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n731), .B1(new_n727), .B2(new_n730), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n732), .A2(new_n733), .ZN(G229));
  INV_X1    g309(.A(G16), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n735), .A2(G23), .ZN(new_n736));
  INV_X1    g311(.A(G288), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n736), .B1(new_n737), .B2(new_n735), .ZN(new_n738));
  XOR2_X1   g313(.A(KEYINPUT33), .B(G1976), .Z(new_n739));
  AND2_X1   g314(.A1(new_n735), .A2(G6), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(G305), .B2(G16), .ZN(new_n741));
  XOR2_X1   g316(.A(KEYINPUT32), .B(G1981), .Z(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT89), .ZN(new_n743));
  AOI22_X1  g318(.A1(new_n738), .A2(new_n739), .B1(new_n741), .B2(new_n743), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(new_n741), .B2(new_n743), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n735), .A2(G22), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(G166), .B2(new_n735), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(G1971), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n738), .A2(new_n739), .ZN(new_n749));
  OR3_X1    g324(.A1(new_n745), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  AND2_X1   g325(.A1(new_n750), .A2(KEYINPUT34), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n484), .A2(G119), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n475), .A2(G131), .A3(new_n476), .ZN(new_n753));
  OR2_X1    g328(.A1(G95), .A2(G2105), .ZN(new_n754));
  OAI211_X1 g329(.A(new_n754), .B(G2104), .C1(G107), .C2(new_n464), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT87), .Z(new_n756));
  NAND3_X1  g331(.A1(new_n752), .A2(new_n753), .A3(new_n756), .ZN(new_n757));
  MUX2_X1   g332(.A(G25), .B(new_n757), .S(G29), .Z(new_n758));
  XOR2_X1   g333(.A(KEYINPUT35), .B(G1991), .Z(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(new_n750), .B2(KEYINPUT34), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n735), .A2(G24), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT88), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(G290), .B2(G16), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(G1986), .Z(new_n765));
  NOR3_X1   g340(.A1(new_n751), .A2(new_n761), .A3(new_n765), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT36), .ZN(new_n767));
  INV_X1    g342(.A(KEYINPUT30), .ZN(new_n768));
  AND2_X1   g343(.A1(new_n768), .A2(G28), .ZN(new_n769));
  INV_X1    g344(.A(G29), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(new_n768), .B2(G28), .ZN(new_n771));
  AND2_X1   g346(.A1(KEYINPUT31), .A2(G11), .ZN(new_n772));
  NOR2_X1   g347(.A1(KEYINPUT31), .A2(G11), .ZN(new_n773));
  OAI22_X1  g348(.A1(new_n769), .A2(new_n771), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  AND2_X1   g349(.A1(KEYINPUT24), .A2(G34), .ZN(new_n775));
  NOR2_X1   g350(.A1(KEYINPUT24), .A2(G34), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n770), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT94), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(G160), .B2(G29), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n774), .B1(new_n779), .B2(G2084), .ZN(new_n780));
  INV_X1    g355(.A(KEYINPUT99), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n779), .A2(G2084), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n484), .A2(G129), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n477), .A2(G141), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n464), .A2(G105), .A3(G2104), .ZN(new_n785));
  NAND3_X1  g360(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT95), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT26), .ZN(new_n788));
  NAND4_X1  g363(.A1(new_n783), .A2(new_n784), .A3(new_n785), .A4(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n790), .A2(new_n770), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(new_n770), .B2(G32), .ZN(new_n792));
  XNOR2_X1  g367(.A(KEYINPUT27), .B(G1996), .ZN(new_n793));
  OAI221_X1 g368(.A(new_n780), .B1(new_n781), .B2(new_n782), .C1(new_n792), .C2(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n664), .A2(G29), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n795), .A2(KEYINPUT97), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n795), .A2(KEYINPUT97), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n782), .A2(new_n781), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n770), .A2(G27), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(G164), .B2(new_n770), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(G2078), .ZN(new_n802));
  NOR4_X1   g377(.A1(new_n794), .A2(new_n796), .A3(new_n799), .A4(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n770), .A2(G26), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT92), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT28), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n484), .A2(G128), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n477), .A2(G140), .ZN(new_n808));
  OAI21_X1  g383(.A(KEYINPUT90), .B1(G104), .B2(G2105), .ZN(new_n809));
  INV_X1    g384(.A(new_n809), .ZN(new_n810));
  NOR3_X1   g385(.A1(KEYINPUT90), .A2(G104), .A3(G2105), .ZN(new_n811));
  OAI221_X1 g386(.A(G2104), .B1(G116), .B2(new_n464), .C1(new_n810), .C2(new_n811), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n807), .A2(new_n808), .A3(new_n812), .ZN(new_n813));
  AND3_X1   g388(.A1(new_n813), .A2(KEYINPUT91), .A3(G29), .ZN(new_n814));
  AOI21_X1  g389(.A(KEYINPUT91), .B1(new_n813), .B2(G29), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n806), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(G2067), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n803), .A2(new_n818), .ZN(new_n819));
  NOR2_X1   g394(.A1(G29), .A2(G35), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n820), .B1(G162), .B2(G29), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT29), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(G2090), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n735), .A2(G4), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n824), .B1(new_n652), .B2(new_n735), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(G1348), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n466), .A2(G127), .ZN(new_n827));
  NAND2_X1  g402(.A1(G115), .A2(G2104), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n464), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT93), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT25), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n832), .B1(new_n477), .B2(G139), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n830), .A2(new_n833), .ZN(new_n834));
  MUX2_X1   g409(.A(G33), .B(new_n834), .S(G29), .Z(new_n835));
  AOI22_X1  g410(.A1(new_n792), .A2(new_n793), .B1(G2072), .B2(new_n835), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n836), .B1(G2072), .B2(new_n835), .ZN(new_n837));
  NOR4_X1   g412(.A1(new_n819), .A2(new_n823), .A3(new_n826), .A4(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n735), .A2(G21), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n839), .B1(G168), .B2(new_n735), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT96), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(G1966), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n735), .A2(G19), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n843), .B1(new_n584), .B2(new_n735), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n844), .B(G1341), .Z(new_n845));
  NOR2_X1   g420(.A1(G5), .A2(G16), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT98), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n847), .B1(G301), .B2(new_n735), .ZN(new_n848));
  INV_X1    g423(.A(G1961), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n848), .B(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(KEYINPUT100), .B(KEYINPUT23), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n735), .A2(G20), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n851), .B(new_n852), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n853), .B1(G299), .B2(G16), .ZN(new_n854));
  INV_X1    g429(.A(G1956), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n854), .B(new_n855), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n850), .A2(new_n856), .ZN(new_n857));
  NAND4_X1  g432(.A1(new_n838), .A2(new_n842), .A3(new_n845), .A4(new_n857), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n767), .A2(new_n858), .ZN(G311));
  OR2_X1    g434(.A1(new_n767), .A2(new_n858), .ZN(G150));
  XOR2_X1   g435(.A(KEYINPUT102), .B(G55), .Z(new_n861));
  NAND2_X1  g436(.A1(new_n637), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n594), .A2(G93), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n540), .A2(G67), .A3(new_n542), .ZN(new_n865));
  NAND2_X1  g440(.A1(G80), .A2(G543), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n864), .B1(new_n867), .B2(G651), .ZN(new_n868));
  XOR2_X1   g443(.A(KEYINPUT103), .B(G860), .Z(new_n869));
  NOR2_X1   g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(KEYINPUT37), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n868), .B1(new_n577), .B2(new_n582), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n867), .A2(G651), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n873), .A2(new_n863), .A3(new_n862), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n571), .A2(new_n576), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n872), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n644), .A2(new_n653), .ZN(new_n878));
  XOR2_X1   g453(.A(KEYINPUT101), .B(KEYINPUT38), .Z(new_n879));
  XNOR2_X1  g454(.A(new_n878), .B(new_n879), .ZN(new_n880));
  XOR2_X1   g455(.A(new_n877), .B(new_n880), .Z(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n882), .A2(KEYINPUT39), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT39), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n869), .B1(new_n881), .B2(new_n884), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n871), .B1(new_n883), .B2(new_n885), .ZN(G145));
  INV_X1    g461(.A(KEYINPUT107), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n757), .A2(new_n887), .ZN(new_n888));
  NAND4_X1  g463(.A1(new_n752), .A2(KEYINPUT107), .A3(new_n753), .A4(new_n756), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n890), .A2(new_n668), .ZN(new_n891));
  INV_X1    g466(.A(new_n668), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n888), .A2(new_n892), .A3(new_n889), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT106), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n789), .A2(new_n834), .A3(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n789), .B1(new_n834), .B2(new_n894), .ZN(new_n897));
  OAI211_X1 g472(.A(new_n891), .B(new_n893), .C1(new_n896), .C2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n897), .ZN(new_n899));
  AND3_X1   g474(.A1(new_n888), .A2(new_n892), .A3(new_n889), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n892), .B1(new_n888), .B2(new_n889), .ZN(new_n901));
  OAI211_X1 g476(.A(new_n899), .B(new_n895), .C1(new_n900), .C2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n898), .A2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT104), .ZN(new_n904));
  AND3_X1   g479(.A1(new_n496), .A2(new_n904), .A3(new_n498), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n904), .B1(new_n496), .B2(new_n498), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n500), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT105), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  OAI211_X1 g484(.A(KEYINPUT105), .B(new_n500), .C1(new_n905), .C2(new_n906), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n813), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n484), .A2(G130), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n477), .A2(G142), .ZN(new_n915));
  OR2_X1    g490(.A1(G106), .A2(G2105), .ZN(new_n916));
  OAI211_X1 g491(.A(new_n916), .B(G2104), .C1(G118), .C2(new_n464), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n914), .A2(new_n915), .A3(new_n917), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n909), .A2(new_n813), .A3(new_n910), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n913), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n918), .B1(new_n913), .B2(new_n919), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n903), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(new_n922), .ZN(new_n924));
  NAND4_X1  g499(.A1(new_n924), .A2(new_n920), .A3(new_n898), .A4(new_n902), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n663), .B(G160), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n927), .B(G162), .ZN(new_n928));
  AOI21_X1  g503(.A(G37), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(new_n928), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n923), .A2(new_n930), .A3(new_n925), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  XNOR2_X1  g507(.A(KEYINPUT108), .B(KEYINPUT40), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n932), .B(new_n933), .ZN(G395));
  XNOR2_X1  g509(.A(new_n877), .B(new_n655), .ZN(new_n935));
  NAND2_X1  g510(.A1(G299), .A2(new_n644), .ZN(new_n936));
  NAND4_X1  g511(.A1(new_n595), .A2(new_n638), .A3(new_n602), .A4(new_n643), .ZN(new_n937));
  AOI21_X1  g512(.A(KEYINPUT41), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  AND3_X1   g513(.A1(new_n936), .A2(KEYINPUT41), .A3(new_n937), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n935), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n936), .A2(new_n937), .ZN(new_n941));
  INV_X1    g516(.A(new_n941), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n940), .B1(new_n942), .B2(new_n935), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT109), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n621), .A2(new_n623), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n511), .B1(new_n945), .B2(KEYINPUT81), .ZN(new_n946));
  AOI211_X1 g521(.A(G288), .B(new_n631), .C1(new_n946), .C2(new_n624), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n737), .B1(new_n625), .B2(new_n632), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n944), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  AND3_X1   g524(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n622), .B1(new_n621), .B2(new_n623), .ZN(new_n951));
  NOR3_X1   g526(.A1(new_n950), .A2(new_n951), .A3(new_n511), .ZN(new_n952));
  OAI21_X1  g527(.A(G288), .B1(new_n952), .B2(new_n631), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n625), .A2(new_n632), .A3(new_n737), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n953), .A2(KEYINPUT109), .A3(new_n954), .ZN(new_n955));
  XNOR2_X1  g530(.A(G303), .B(G305), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n949), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(new_n956), .ZN(new_n958));
  OAI211_X1 g533(.A(new_n958), .B(new_n944), .C1(new_n948), .C2(new_n947), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT110), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n960), .A2(new_n961), .A3(KEYINPUT42), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(KEYINPUT42), .ZN(new_n963));
  OR2_X1    g538(.A1(new_n961), .A2(KEYINPUT42), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n957), .A2(new_n959), .A3(new_n963), .A4(new_n964), .ZN(new_n965));
  AND3_X1   g540(.A1(new_n943), .A2(new_n962), .A3(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n943), .B1(new_n965), .B2(new_n962), .ZN(new_n967));
  OAI21_X1  g542(.A(G868), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n968), .B1(G868), .B2(new_n868), .ZN(G295));
  OAI21_X1  g544(.A(new_n968), .B1(G868), .B2(new_n868), .ZN(G331));
  AOI21_X1  g545(.A(KEYINPUT78), .B1(new_n571), .B2(new_n576), .ZN(new_n971));
  NOR3_X1   g546(.A1(new_n581), .A2(new_n578), .A3(new_n575), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n874), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n868), .A2(new_n571), .A3(new_n576), .ZN(new_n974));
  INV_X1    g549(.A(new_n563), .ZN(new_n975));
  INV_X1    g550(.A(new_n559), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(new_n557), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n975), .A2(new_n977), .A3(G286), .ZN(new_n978));
  OAI21_X1  g553(.A(G168), .B1(new_n563), .B2(new_n560), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n973), .A2(new_n974), .A3(new_n978), .A4(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n978), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n981), .B1(new_n872), .B2(new_n876), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n941), .B1(new_n980), .B2(new_n982), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n939), .A2(new_n938), .ZN(new_n984));
  AND3_X1   g559(.A1(new_n980), .A2(new_n984), .A3(new_n982), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n960), .B1(new_n983), .B2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(G37), .ZN(new_n987));
  NOR3_X1   g562(.A1(new_n981), .A2(new_n872), .A3(new_n876), .ZN(new_n988));
  AOI22_X1  g563(.A1(new_n973), .A2(new_n974), .B1(new_n978), .B2(new_n979), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n942), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n980), .A2(new_n984), .A3(new_n982), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n990), .A2(new_n957), .A3(new_n959), .A4(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n986), .A2(new_n987), .A3(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(KEYINPUT43), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT43), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n986), .A2(new_n992), .A3(new_n995), .A4(new_n987), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n994), .A2(KEYINPUT44), .A3(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT111), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n994), .A2(new_n998), .A3(new_n996), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n993), .A2(KEYINPUT111), .A3(KEYINPUT43), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n997), .B1(new_n1001), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g577(.A(G1996), .ZN(new_n1003));
  XNOR2_X1  g578(.A(new_n789), .B(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g579(.A(new_n813), .B(new_n817), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(new_n759), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n757), .A2(new_n1007), .ZN(new_n1008));
  AND2_X1   g583(.A1(new_n757), .A2(new_n1007), .ZN(new_n1009));
  OR3_X1    g584(.A1(new_n1006), .A2(new_n1008), .A3(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1010), .B1(G1986), .B2(G290), .ZN(new_n1011));
  OR2_X1    g586(.A1(G290), .A2(G1986), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(KEYINPUT112), .B1(new_n911), .B2(G1384), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT45), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT112), .ZN(new_n1016));
  INV_X1    g591(.A(G1384), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n909), .A2(new_n1016), .A3(new_n1017), .A4(new_n910), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1014), .A2(new_n1015), .A3(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(G160), .A2(G40), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1013), .A2(new_n1021), .ZN(new_n1022));
  XOR2_X1   g597(.A(KEYINPUT122), .B(KEYINPUT54), .Z(new_n1023));
  NAND2_X1  g598(.A1(new_n502), .A2(new_n1017), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT113), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1024), .A2(new_n1025), .A3(new_n1015), .ZN(new_n1026));
  AOI21_X1  g601(.A(G1384), .B1(new_n499), .B2(new_n501), .ZN(new_n1027));
  OAI21_X1  g602(.A(KEYINPUT113), .B1(new_n1027), .B2(KEYINPUT45), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(G2078), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n909), .A2(KEYINPUT45), .A3(new_n1017), .A4(new_n910), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1020), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n1029), .A2(new_n1030), .A3(new_n1031), .A4(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT53), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1020), .B1(new_n1024), .B2(KEYINPUT50), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT50), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n907), .A2(new_n1036), .A3(new_n1017), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1035), .A2(new_n1037), .ZN(new_n1038));
  AOI22_X1  g613(.A1(new_n1033), .A2(new_n1034), .B1(new_n849), .B2(new_n1038), .ZN(new_n1039));
  NOR3_X1   g614(.A1(new_n1020), .A2(new_n1034), .A3(G2078), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1019), .A2(new_n1031), .A3(new_n1040), .ZN(new_n1041));
  AND3_X1   g616(.A1(new_n1039), .A2(new_n1041), .A3(G301), .ZN(new_n1042));
  AOI21_X1  g617(.A(KEYINPUT45), .B1(new_n907), .B2(new_n1017), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1020), .B1(new_n1027), .B2(KEYINPUT45), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1044), .A2(new_n1030), .A3(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT123), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1044), .A2(KEYINPUT123), .A3(new_n1045), .A4(new_n1030), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1048), .A2(KEYINPUT53), .A3(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(G301), .B1(new_n1039), .B2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1023), .B1(new_n1042), .B2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1039), .A2(new_n1050), .A3(G301), .ZN(new_n1053));
  AND2_X1   g628(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1054));
  OAI211_X1 g629(.A(KEYINPUT54), .B(new_n1053), .C1(new_n1054), .C2(G301), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT49), .ZN(new_n1056));
  INV_X1    g631(.A(G1981), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n613), .A2(new_n1057), .A3(new_n614), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1058), .ZN(new_n1059));
  XNOR2_X1  g634(.A(KEYINPUT117), .B(G86), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n594), .A2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1057), .B1(new_n613), .B2(new_n1061), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1056), .B1(new_n1059), .B2(new_n1062), .ZN(new_n1063));
  AND2_X1   g638(.A1(new_n613), .A2(new_n1061), .ZN(new_n1064));
  OAI211_X1 g639(.A(KEYINPUT49), .B(new_n1058), .C1(new_n1064), .C2(new_n1057), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1032), .A2(new_n907), .A3(new_n1017), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1063), .A2(new_n1065), .A3(G8), .A4(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n737), .A2(G1976), .ZN(new_n1068));
  INV_X1    g643(.A(G1976), .ZN(new_n1069));
  AOI21_X1  g644(.A(KEYINPUT52), .B1(G288), .B2(new_n1069), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1068), .A2(new_n1066), .A3(new_n1070), .A4(G8), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1067), .A2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1068), .A2(new_n1066), .A3(G8), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(KEYINPUT52), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(KEYINPUT116), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT116), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1073), .A2(new_n1076), .A3(KEYINPUT52), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1072), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1078));
  OAI211_X1 g653(.A(KEYINPUT55), .B(G8), .C1(new_n512), .C2(new_n522), .ZN(new_n1079));
  XNOR2_X1  g654(.A(new_n1079), .B(KEYINPUT114), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT115), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  OR2_X1    g657(.A1(new_n1079), .A2(KEYINPUT114), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1079), .A2(KEYINPUT114), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1083), .A2(KEYINPUT115), .A3(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT55), .ZN(new_n1086));
  INV_X1    g661(.A(G8), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1086), .B1(G166), .B2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1082), .A2(new_n1085), .A3(new_n1088), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1020), .B1(new_n1026), .B2(new_n1028), .ZN(new_n1090));
  AOI21_X1  g665(.A(G1971), .B1(new_n1090), .B2(new_n1031), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1038), .A2(G2090), .ZN(new_n1092));
  OAI211_X1 g667(.A(new_n1089), .B(G8), .C1(new_n1091), .C2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1029), .A2(new_n1032), .A3(new_n1031), .ZN(new_n1094));
  INV_X1    g669(.A(G1971), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1027), .A2(new_n1036), .ZN(new_n1097));
  XNOR2_X1  g672(.A(new_n1097), .B(KEYINPUT118), .ZN(new_n1098));
  INV_X1    g673(.A(G2090), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n907), .A2(new_n1017), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1020), .B1(new_n1100), .B2(KEYINPUT50), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1098), .A2(new_n1099), .A3(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1087), .B1(new_n1096), .B2(new_n1102), .ZN(new_n1103));
  OAI211_X1 g678(.A(new_n1078), .B(new_n1093), .C1(new_n1103), .C2(new_n1089), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(G1966), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1032), .B1(new_n1024), .B2(new_n1015), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1106), .B1(new_n1107), .B2(new_n1043), .ZN(new_n1108));
  INV_X1    g683(.A(G2084), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1035), .A2(new_n1109), .A3(new_n1037), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1108), .A2(G168), .A3(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1111), .A2(G8), .ZN(new_n1112));
  AOI21_X1  g687(.A(G168), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1113));
  OAI21_X1  g688(.A(KEYINPUT51), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT51), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1111), .A2(new_n1115), .A3(G8), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1052), .A2(new_n1055), .A3(new_n1105), .A4(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT118), .ZN(new_n1119));
  XNOR2_X1  g694(.A(new_n1097), .B(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1101), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n855), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  XOR2_X1   g697(.A(G299), .B(KEYINPUT57), .Z(new_n1123));
  XNOR2_X1  g698(.A(KEYINPUT56), .B(G2072), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1090), .A2(new_n1031), .A3(new_n1124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1122), .A2(new_n1123), .A3(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1123), .B1(new_n1122), .B2(new_n1125), .ZN(new_n1128));
  OAI21_X1  g703(.A(KEYINPUT120), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(KEYINPUT61), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1066), .ZN(new_n1131));
  XNOR2_X1  g706(.A(KEYINPUT58), .B(G1341), .ZN(new_n1132));
  OAI22_X1  g707(.A1(new_n1094), .A2(G1996), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1133), .A2(new_n584), .ZN(new_n1134));
  XNOR2_X1  g709(.A(new_n1134), .B(KEYINPUT59), .ZN(new_n1135));
  INV_X1    g710(.A(G1348), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1038), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1131), .A2(new_n817), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT60), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n644), .A2(KEYINPUT121), .ZN(new_n1142));
  OR2_X1    g717(.A1(new_n644), .A2(KEYINPUT121), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1141), .A2(new_n1142), .A3(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1145));
  OAI211_X1 g720(.A(new_n1144), .B(new_n1145), .C1(new_n1141), .C2(new_n1142), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT61), .ZN(new_n1147));
  OAI211_X1 g722(.A(KEYINPUT120), .B(new_n1147), .C1(new_n1127), .C2(new_n1128), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1130), .A2(new_n1135), .A3(new_n1146), .A4(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n644), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1126), .B1(new_n1128), .B2(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT119), .ZN(new_n1152));
  XNOR2_X1  g727(.A(new_n1151), .B(new_n1152), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1118), .B1(new_n1149), .B2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT124), .ZN(new_n1155));
  AND3_X1   g730(.A1(new_n1111), .A2(new_n1115), .A3(G8), .ZN(new_n1156));
  AND3_X1   g731(.A1(new_n1035), .A2(new_n1109), .A3(new_n1037), .ZN(new_n1157));
  AOI21_X1  g732(.A(G1966), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1158));
  OAI21_X1  g733(.A(G286), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1159), .A2(G8), .A3(new_n1111), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1156), .B1(KEYINPUT51), .B2(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT62), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1155), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1051), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1104), .A2(new_n1164), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1117), .A2(KEYINPUT124), .A3(KEYINPUT62), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1163), .A2(new_n1165), .A3(new_n1166), .A4(new_n1167), .ZN(new_n1168));
  AND3_X1   g743(.A1(new_n1067), .A2(new_n1069), .A3(new_n737), .ZN(new_n1169));
  OAI211_X1 g744(.A(G8), .B(new_n1066), .C1(new_n1169), .C2(new_n1059), .ZN(new_n1170));
  INV_X1    g745(.A(new_n1078), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1170), .B1(new_n1171), .B2(new_n1093), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT63), .ZN(new_n1173));
  OAI211_X1 g748(.A(G8), .B(G168), .C1(new_n1157), .C2(new_n1158), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1173), .B1(new_n1104), .B2(new_n1174), .ZN(new_n1175));
  OAI21_X1  g750(.A(G8), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1176));
  NAND4_X1  g751(.A1(new_n1176), .A2(new_n1085), .A3(new_n1088), .A4(new_n1082), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n1174), .A2(new_n1173), .ZN(new_n1178));
  NAND4_X1  g753(.A1(new_n1177), .A2(new_n1093), .A3(new_n1078), .A4(new_n1178), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1172), .B1(new_n1175), .B2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1168), .A2(new_n1180), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1022), .B1(new_n1154), .B2(new_n1181), .ZN(new_n1182));
  INV_X1    g757(.A(new_n1021), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT48), .ZN(new_n1184));
  OR3_X1    g759(.A1(new_n1183), .A2(new_n1184), .A3(new_n1012), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1184), .B1(new_n1183), .B2(new_n1012), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1010), .A2(new_n1021), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1185), .A2(new_n1186), .A3(new_n1187), .ZN(new_n1188));
  INV_X1    g763(.A(new_n1006), .ZN(new_n1189));
  OAI21_X1  g764(.A(new_n1008), .B1(new_n1183), .B2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n912), .A2(new_n817), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1190), .A2(KEYINPUT125), .A3(new_n1191), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1192), .A2(new_n1021), .ZN(new_n1193));
  AOI21_X1  g768(.A(KEYINPUT125), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1188), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  INV_X1    g770(.A(KEYINPUT46), .ZN(new_n1196));
  OAI211_X1 g771(.A(new_n1005), .B(new_n790), .C1(new_n1196), .C2(G1996), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1021), .A2(new_n1197), .ZN(new_n1198));
  INV_X1    g773(.A(KEYINPUT126), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1021), .A2(new_n1003), .ZN(new_n1200));
  AOI21_X1  g775(.A(new_n1199), .B1(new_n1200), .B2(new_n1196), .ZN(new_n1201));
  AOI211_X1 g776(.A(KEYINPUT126), .B(KEYINPUT46), .C1(new_n1021), .C2(new_n1003), .ZN(new_n1202));
  OAI21_X1  g777(.A(new_n1198), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1203), .A2(KEYINPUT47), .ZN(new_n1204));
  OR2_X1    g779(.A1(new_n1203), .A2(KEYINPUT47), .ZN(new_n1205));
  AOI21_X1  g780(.A(new_n1195), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1182), .A2(new_n1206), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g782(.A1(G227), .A2(new_n462), .ZN(new_n1209));
  OAI211_X1 g783(.A(new_n693), .B(new_n1209), .C1(new_n732), .C2(new_n733), .ZN(new_n1210));
  AOI21_X1  g784(.A(new_n1210), .B1(new_n929), .B2(new_n931), .ZN(new_n1211));
  NAND3_X1  g785(.A1(new_n999), .A2(new_n1000), .A3(new_n1211), .ZN(new_n1212));
  NAND2_X1  g786(.A1(new_n1212), .A2(KEYINPUT127), .ZN(new_n1213));
  INV_X1    g787(.A(KEYINPUT127), .ZN(new_n1214));
  NAND4_X1  g788(.A1(new_n999), .A2(new_n1211), .A3(new_n1214), .A4(new_n1000), .ZN(new_n1215));
  AND2_X1   g789(.A1(new_n1213), .A2(new_n1215), .ZN(G308));
  NAND2_X1  g790(.A1(new_n1213), .A2(new_n1215), .ZN(G225));
endmodule


