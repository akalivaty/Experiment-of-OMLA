//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 0 0 1 1 0 1 0 0 1 0 1 0 1 1 0 0 0 1 1 1 0 1 0 0 0 0 1 0 1 0 1 0 1 1 1 0 1 0 0 0 0 1 1 0 0 1 1 0 1 1 0 1 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:33 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n708, new_n709, new_n710,
    new_n711, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n729, new_n730, new_n731, new_n732, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n748, new_n749, new_n750,
    new_n751, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n765, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n964, new_n965, new_n966, new_n967, new_n968, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  XNOR2_X1  g001(.A(new_n187), .B(KEYINPUT83), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G104), .ZN(new_n190));
  OAI21_X1  g004(.A(KEYINPUT3), .B1(new_n190), .B2(G107), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT3), .ZN(new_n192));
  INV_X1    g006(.A(G107), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n192), .A2(new_n193), .A3(G104), .ZN(new_n194));
  INV_X1    g008(.A(G101), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n190), .A2(G107), .ZN(new_n196));
  NAND4_X1  g010(.A1(new_n191), .A2(new_n194), .A3(new_n195), .A4(new_n196), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n190), .A2(G107), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n193), .A2(G104), .ZN(new_n199));
  OAI21_X1  g013(.A(G101), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n197), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G119), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G116), .ZN(new_n203));
  INV_X1    g017(.A(G116), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G119), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n203), .A2(new_n205), .A3(KEYINPUT5), .ZN(new_n206));
  OAI211_X1 g020(.A(new_n206), .B(G113), .C1(KEYINPUT5), .C2(new_n203), .ZN(new_n207));
  NAND2_X1  g021(.A1(KEYINPUT2), .A2(G113), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(KEYINPUT66), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT66), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n210), .A2(KEYINPUT2), .A3(G113), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT2), .ZN(new_n212));
  INV_X1    g026(.A(G113), .ZN(new_n213));
  AOI22_X1  g027(.A1(new_n209), .A2(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  XNOR2_X1  g028(.A(G116), .B(G119), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n201), .A2(new_n207), .A3(new_n216), .ZN(new_n217));
  XNOR2_X1  g031(.A(G110), .B(G122), .ZN(new_n218));
  XNOR2_X1  g032(.A(KEYINPUT86), .B(KEYINPUT8), .ZN(new_n219));
  XNOR2_X1  g033(.A(new_n218), .B(new_n219), .ZN(new_n220));
  OAI21_X1  g034(.A(G113), .B1(new_n203), .B2(KEYINPUT5), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT87), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n221), .B1(new_n222), .B2(new_n206), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n215), .A2(KEYINPUT87), .A3(KEYINPUT5), .ZN(new_n224));
  AOI22_X1  g038(.A1(new_n223), .A2(new_n224), .B1(new_n214), .B2(new_n215), .ZN(new_n225));
  OAI211_X1 g039(.A(new_n217), .B(new_n220), .C1(new_n225), .C2(new_n201), .ZN(new_n226));
  INV_X1    g040(.A(G146), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(G143), .ZN(new_n228));
  INV_X1    g042(.A(G143), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(G146), .ZN(new_n230));
  AND2_X1   g044(.A1(KEYINPUT0), .A2(G128), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n228), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  XNOR2_X1  g046(.A(G143), .B(G146), .ZN(new_n233));
  XNOR2_X1  g047(.A(KEYINPUT0), .B(G128), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n232), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G125), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT88), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  XOR2_X1   g052(.A(KEYINPUT85), .B(G224), .Z(new_n239));
  INV_X1    g053(.A(G953), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(KEYINPUT7), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n228), .A2(new_n230), .ZN(new_n243));
  XNOR2_X1  g057(.A(KEYINPUT65), .B(G128), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT1), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n245), .B1(G143), .B2(new_n227), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n243), .B1(new_n244), .B2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(G125), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n233), .A2(new_n245), .A3(G128), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n247), .A2(new_n248), .A3(new_n249), .ZN(new_n250));
  AOI22_X1  g064(.A1(new_n238), .A2(new_n242), .B1(new_n236), .B2(new_n250), .ZN(new_n251));
  AND4_X1   g065(.A1(KEYINPUT88), .A2(new_n250), .A3(new_n236), .A4(new_n242), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n226), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT89), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  AND2_X1   g069(.A1(new_n197), .A2(new_n200), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n256), .A2(new_n216), .A3(new_n207), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n191), .A2(new_n194), .A3(new_n196), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n258), .A2(new_n259), .A3(G101), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n209), .A2(new_n211), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n212), .A2(new_n213), .ZN(new_n262));
  AND3_X1   g076(.A1(new_n261), .A2(new_n262), .A3(new_n215), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n215), .B1(new_n261), .B2(new_n262), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n260), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n258), .A2(G101), .ZN(new_n266));
  AND3_X1   g080(.A1(new_n266), .A2(KEYINPUT4), .A3(new_n197), .ZN(new_n267));
  OAI211_X1 g081(.A(new_n218), .B(new_n257), .C1(new_n265), .C2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT84), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(new_n264), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(new_n216), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n266), .A2(KEYINPUT4), .A3(new_n197), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n272), .A2(new_n273), .A3(new_n260), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n274), .A2(KEYINPUT84), .A3(new_n218), .A4(new_n257), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n270), .A2(new_n275), .ZN(new_n276));
  OAI211_X1 g090(.A(new_n226), .B(KEYINPUT89), .C1(new_n251), .C2(new_n252), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n255), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(G902), .ZN(new_n279));
  AND2_X1   g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n218), .B1(new_n274), .B2(new_n257), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT6), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n281), .B1(new_n270), .B2(new_n275), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n284), .B1(new_n285), .B2(new_n283), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n250), .A2(new_n236), .ZN(new_n287));
  XNOR2_X1  g101(.A(new_n287), .B(new_n241), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n286), .A2(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(G210), .B1(G237), .B2(G902), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n280), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n291), .B1(new_n280), .B2(new_n290), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n189), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  XNOR2_X1  g110(.A(G113), .B(G122), .ZN(new_n297));
  XNOR2_X1  g111(.A(new_n297), .B(new_n190), .ZN(new_n298));
  INV_X1    g112(.A(G140), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(G125), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n248), .A2(G140), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  XNOR2_X1  g116(.A(new_n302), .B(G146), .ZN(new_n303));
  XNOR2_X1  g117(.A(new_n303), .B(KEYINPUT90), .ZN(new_n304));
  INV_X1    g118(.A(G237), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n305), .A2(new_n240), .A3(G214), .ZN(new_n306));
  XNOR2_X1  g120(.A(new_n306), .B(G143), .ZN(new_n307));
  NAND2_X1  g121(.A1(KEYINPUT18), .A2(G131), .ZN(new_n308));
  XOR2_X1   g122(.A(new_n307), .B(new_n308), .Z(new_n309));
  NAND2_X1  g123(.A1(new_n304), .A2(new_n309), .ZN(new_n310));
  NAND4_X1  g124(.A1(new_n300), .A2(new_n301), .A3(KEYINPUT73), .A4(KEYINPUT16), .ZN(new_n311));
  AND3_X1   g125(.A1(new_n300), .A2(new_n301), .A3(KEYINPUT16), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT16), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n313), .A2(new_n299), .A3(G125), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT73), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n311), .B1(new_n312), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(G146), .ZN(new_n318));
  OAI211_X1 g132(.A(new_n227), .B(new_n311), .C1(new_n312), .C2(new_n316), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n318), .A2(KEYINPUT74), .A3(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT91), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT74), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n317), .A2(new_n322), .A3(G146), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n320), .A2(new_n321), .A3(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(new_n307), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n325), .A2(KEYINPUT17), .A3(G131), .ZN(new_n326));
  AND2_X1   g140(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n319), .A2(KEYINPUT74), .ZN(new_n328));
  OAI211_X1 g142(.A(new_n315), .B(new_n314), .C1(new_n302), .C2(new_n313), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n227), .B1(new_n329), .B2(new_n311), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(new_n323), .ZN(new_n332));
  OAI21_X1  g146(.A(KEYINPUT91), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  AOI21_X1  g147(.A(KEYINPUT92), .B1(new_n327), .B2(new_n333), .ZN(new_n334));
  NAND4_X1  g148(.A1(new_n333), .A2(KEYINPUT92), .A3(new_n326), .A4(new_n324), .ZN(new_n335));
  INV_X1    g149(.A(G131), .ZN(new_n336));
  XNOR2_X1  g150(.A(new_n307), .B(new_n336), .ZN(new_n337));
  OR2_X1    g151(.A1(new_n337), .A2(KEYINPUT17), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n335), .A2(new_n338), .ZN(new_n339));
  OAI211_X1 g153(.A(new_n298), .B(new_n310), .C1(new_n334), .C2(new_n339), .ZN(new_n340));
  XNOR2_X1  g154(.A(new_n302), .B(KEYINPUT19), .ZN(new_n341));
  OAI211_X1 g155(.A(new_n337), .B(new_n318), .C1(G146), .C2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n310), .A2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(new_n298), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n340), .A2(new_n345), .ZN(new_n346));
  NOR2_X1   g160(.A1(G475), .A2(G902), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(KEYINPUT20), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT20), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n346), .A2(new_n350), .A3(new_n347), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  OAI21_X1  g166(.A(G478), .B1(KEYINPUT97), .B2(KEYINPUT15), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n353), .B1(KEYINPUT97), .B2(KEYINPUT15), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT98), .ZN(new_n356));
  XNOR2_X1  g170(.A(KEYINPUT9), .B(G234), .ZN(new_n357));
  INV_X1    g171(.A(G217), .ZN(new_n358));
  NOR3_X1   g172(.A1(new_n357), .A2(new_n358), .A3(G953), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n204), .A2(G122), .ZN(new_n361));
  XNOR2_X1  g175(.A(new_n361), .B(KEYINPUT95), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT96), .ZN(new_n363));
  AND2_X1   g177(.A1(KEYINPUT94), .A2(G122), .ZN(new_n364));
  NOR2_X1   g178(.A1(KEYINPUT94), .A2(G122), .ZN(new_n365));
  OAI21_X1  g179(.A(G116), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  AND3_X1   g180(.A1(new_n362), .A2(new_n363), .A3(new_n366), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n363), .B1(new_n362), .B2(new_n366), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n193), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT95), .ZN(new_n370));
  XNOR2_X1  g184(.A(new_n361), .B(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT14), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n366), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n362), .A2(KEYINPUT14), .ZN(new_n374));
  OAI21_X1  g188(.A(G107), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n244), .A2(G143), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n229), .A2(G128), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  XNOR2_X1  g192(.A(new_n378), .B(G134), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n369), .A2(new_n375), .A3(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n362), .A2(new_n366), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(KEYINPUT96), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n362), .A2(new_n363), .A3(new_n366), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n383), .A2(G107), .A3(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(new_n376), .ZN(new_n386));
  OAI21_X1  g200(.A(G134), .B1(new_n386), .B2(KEYINPUT13), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(new_n378), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n376), .A2(KEYINPUT13), .A3(G134), .A4(new_n377), .ZN(new_n389));
  AOI22_X1  g203(.A1(new_n369), .A2(new_n385), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n360), .B1(new_n381), .B2(new_n390), .ZN(new_n391));
  AND2_X1   g205(.A1(new_n369), .A2(new_n385), .ZN(new_n392));
  AND2_X1   g206(.A1(new_n388), .A2(new_n389), .ZN(new_n393));
  OAI211_X1 g207(.A(new_n380), .B(new_n359), .C1(new_n392), .C2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n391), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n356), .B1(new_n395), .B2(new_n279), .ZN(new_n396));
  AOI211_X1 g210(.A(KEYINPUT98), .B(G902), .C1(new_n391), .C2(new_n394), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n355), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n395), .A2(new_n356), .A3(new_n279), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(new_n354), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n240), .A2(G952), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n402), .B1(G234), .B2(G237), .ZN(new_n403));
  AOI211_X1 g217(.A(new_n279), .B(new_n240), .C1(G234), .C2(G237), .ZN(new_n404));
  XNOR2_X1  g218(.A(KEYINPUT21), .B(G898), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n403), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n401), .A2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT92), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n324), .A2(new_n326), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n321), .B1(new_n320), .B2(new_n323), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n408), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n411), .A2(new_n338), .A3(new_n335), .ZN(new_n412));
  AND3_X1   g226(.A1(new_n412), .A2(new_n298), .A3(new_n310), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n298), .B1(new_n412), .B2(new_n310), .ZN(new_n414));
  NOR3_X1   g228(.A1(new_n413), .A2(new_n414), .A3(KEYINPUT93), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n412), .A2(new_n310), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n416), .A2(KEYINPUT93), .A3(new_n344), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(new_n279), .ZN(new_n418));
  OAI21_X1  g232(.A(G475), .B1(new_n415), .B2(new_n418), .ZN(new_n419));
  AND4_X1   g233(.A1(new_n296), .A2(new_n352), .A3(new_n407), .A4(new_n419), .ZN(new_n420));
  OAI21_X1  g234(.A(G221), .B1(new_n357), .B2(G902), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  XNOR2_X1  g236(.A(G110), .B(G140), .ZN(new_n423));
  INV_X1    g237(.A(G227), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n424), .A2(G953), .ZN(new_n425));
  XNOR2_X1  g239(.A(new_n423), .B(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(new_n249), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n228), .A2(KEYINPUT1), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n233), .B1(G128), .B2(new_n428), .ZN(new_n429));
  OAI211_X1 g243(.A(new_n197), .B(new_n200), .C1(new_n427), .C2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT10), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n431), .B1(new_n247), .B2(new_n249), .ZN(new_n432));
  AOI22_X1  g246(.A1(new_n430), .A2(new_n431), .B1(new_n256), .B2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT67), .ZN(new_n434));
  OAI211_X1 g248(.A(new_n232), .B(new_n434), .C1(new_n233), .C2(new_n234), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(KEYINPUT0), .A2(G128), .ZN(new_n437));
  OR2_X1    g251(.A1(KEYINPUT0), .A2(G128), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n229), .A2(G146), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n227), .A2(G143), .ZN(new_n440));
  OAI211_X1 g254(.A(new_n437), .B(new_n438), .C1(new_n439), .C2(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n434), .B1(new_n441), .B2(new_n232), .ZN(new_n442));
  OAI211_X1 g256(.A(new_n273), .B(new_n260), .C1(new_n436), .C2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n433), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(KEYINPUT80), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT11), .ZN(new_n446));
  INV_X1    g260(.A(G134), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n446), .B1(new_n447), .B2(G137), .ZN(new_n448));
  INV_X1    g262(.A(G137), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n449), .A2(KEYINPUT11), .A3(G134), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n447), .A2(G137), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n448), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(G131), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n448), .A2(new_n450), .A3(new_n336), .A4(new_n451), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT80), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n433), .A2(new_n456), .A3(new_n443), .ZN(new_n457));
  AND3_X1   g271(.A1(new_n445), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n430), .A2(new_n431), .ZN(new_n459));
  INV_X1    g273(.A(new_n455), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n432), .A2(new_n256), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n459), .A2(new_n443), .A3(new_n460), .A4(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(KEYINPUT79), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT79), .ZN(new_n464));
  NAND4_X1  g278(.A1(new_n433), .A2(new_n464), .A3(new_n460), .A4(new_n443), .ZN(new_n465));
  AND2_X1   g279(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n426), .B1(new_n458), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n463), .A2(new_n465), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT81), .ZN(new_n469));
  INV_X1    g283(.A(new_n426), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n247), .A2(new_n249), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n430), .B1(new_n472), .B2(new_n256), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(new_n455), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT12), .ZN(new_n475));
  XNOR2_X1  g289(.A(new_n474), .B(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n471), .A2(new_n476), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n426), .B1(new_n463), .B2(new_n465), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n478), .A2(new_n469), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n467), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(G469), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n480), .A2(new_n481), .A3(new_n279), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(KEYINPUT82), .ZN(new_n483));
  XNOR2_X1  g297(.A(new_n474), .B(KEYINPUT12), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n484), .B1(new_n478), .B2(new_n469), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n468), .A2(new_n470), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(KEYINPUT81), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(G902), .B1(new_n488), .B2(new_n467), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT82), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n489), .A2(new_n490), .A3(new_n481), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n483), .A2(new_n491), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n466), .A2(new_n484), .ZN(new_n493));
  OAI22_X1  g307(.A1(new_n493), .A2(new_n470), .B1(new_n486), .B2(new_n458), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n481), .B1(new_n494), .B2(new_n279), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n422), .B1(new_n492), .B2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT77), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n302), .A2(G146), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n330), .A2(new_n499), .ZN(new_n500));
  XOR2_X1   g314(.A(KEYINPUT24), .B(G110), .Z(new_n501));
  NAND2_X1  g315(.A1(new_n244), .A2(G119), .ZN(new_n502));
  INV_X1    g316(.A(G128), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n502), .B1(G119), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(KEYINPUT72), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT72), .ZN(new_n506));
  OAI211_X1 g320(.A(new_n502), .B(new_n506), .C1(G119), .C2(new_n503), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n501), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(KEYINPUT23), .B1(new_n503), .B2(G119), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n509), .B1(new_n202), .B2(G128), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT23), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n510), .B1(new_n502), .B2(new_n511), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n512), .A2(G110), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n500), .B1(new_n508), .B2(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n505), .A2(new_n507), .A3(new_n501), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n512), .A2(G110), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n320), .A2(new_n515), .A3(new_n323), .A4(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n514), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n240), .A2(G221), .A3(G234), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n519), .B(KEYINPUT75), .ZN(new_n520));
  XNOR2_X1  g334(.A(KEYINPUT22), .B(G137), .ZN(new_n521));
  XNOR2_X1  g335(.A(new_n520), .B(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n518), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n514), .A2(new_n517), .A3(new_n522), .ZN(new_n525));
  AOI21_X1  g339(.A(G902), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  XNOR2_X1  g340(.A(KEYINPUT76), .B(KEYINPUT25), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n498), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  AND3_X1   g343(.A1(new_n514), .A2(new_n517), .A3(new_n522), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n522), .B1(new_n514), .B2(new_n517), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  OAI211_X1 g346(.A(KEYINPUT77), .B(new_n527), .C1(new_n532), .C2(G902), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n526), .A2(KEYINPUT25), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n529), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n358), .B1(G234), .B2(new_n279), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(new_n532), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n536), .A2(G902), .ZN(new_n539));
  XOR2_X1   g353(.A(new_n539), .B(KEYINPUT78), .Z(new_n540));
  NAND2_X1  g354(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n537), .A2(new_n541), .ZN(new_n542));
  NOR2_X1   g356(.A1(G472), .A2(G902), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n455), .B1(new_n436), .B2(new_n442), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n447), .A2(G137), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n449), .A2(G134), .ZN(new_n546));
  OAI21_X1  g360(.A(G131), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  AND2_X1   g361(.A1(new_n454), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(new_n472), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n544), .A2(KEYINPUT30), .A3(new_n549), .ZN(new_n550));
  XOR2_X1   g364(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n551));
  NAND2_X1  g365(.A1(new_n454), .A2(new_n547), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n552), .B1(new_n247), .B2(new_n249), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n235), .B1(new_n453), .B2(new_n454), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n551), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n550), .A2(new_n272), .A3(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n305), .A2(new_n240), .A3(G210), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n557), .B(KEYINPUT27), .ZN(new_n558));
  XNOR2_X1  g372(.A(KEYINPUT26), .B(G101), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n558), .B(new_n559), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n263), .A2(new_n264), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n544), .A2(new_n561), .A3(new_n549), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n556), .A2(new_n560), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(KEYINPUT31), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT31), .ZN(new_n565));
  NAND4_X1  g379(.A1(new_n556), .A2(new_n565), .A3(new_n560), .A4(new_n562), .ZN(new_n566));
  OAI211_X1 g380(.A(KEYINPUT68), .B(new_n272), .C1(new_n553), .C2(new_n554), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n562), .A2(new_n567), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n549), .B1(new_n460), .B2(new_n235), .ZN(new_n569));
  AOI21_X1  g383(.A(KEYINPUT68), .B1(new_n569), .B2(new_n272), .ZN(new_n570));
  OAI21_X1  g384(.A(KEYINPUT28), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT28), .ZN(new_n572));
  AND2_X1   g386(.A1(new_n562), .A2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n560), .B1(new_n571), .B2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT69), .ZN(new_n576));
  OAI211_X1 g390(.A(new_n564), .B(new_n566), .C1(new_n575), .C2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n571), .A2(new_n574), .ZN(new_n578));
  INV_X1    g392(.A(new_n560), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n578), .A2(new_n576), .A3(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n543), .B1(new_n577), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(KEYINPUT32), .ZN(new_n583));
  AND2_X1   g397(.A1(new_n564), .A2(new_n566), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT68), .ZN(new_n585));
  INV_X1    g399(.A(new_n235), .ZN(new_n586));
  AOI22_X1  g400(.A1(new_n455), .A2(new_n586), .B1(new_n548), .B2(new_n472), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n585), .B1(new_n587), .B2(new_n561), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n588), .A2(new_n562), .A3(new_n567), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n573), .B1(new_n589), .B2(KEYINPUT28), .ZN(new_n590));
  OAI21_X1  g404(.A(KEYINPUT69), .B1(new_n590), .B2(new_n560), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n584), .A2(new_n580), .A3(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT32), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n592), .A2(new_n593), .A3(new_n543), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n583), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n544), .A2(new_n549), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(new_n272), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT70), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n597), .A2(new_n598), .A3(new_n562), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n596), .A2(KEYINPUT70), .A3(new_n272), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n599), .A2(KEYINPUT28), .A3(new_n600), .ZN(new_n601));
  AND2_X1   g415(.A1(new_n560), .A2(KEYINPUT29), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n601), .A2(new_n574), .A3(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n603), .B(KEYINPUT71), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n590), .A2(new_n560), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n560), .B1(new_n556), .B2(new_n562), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n606), .A2(KEYINPUT29), .ZN(new_n607));
  AOI21_X1  g421(.A(G902), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(G472), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n542), .B1(new_n595), .B2(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n420), .A2(new_n497), .A3(new_n611), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n612), .B(G101), .ZN(G3));
  AOI21_X1  g427(.A(new_n495), .B1(new_n483), .B2(new_n491), .ZN(new_n614));
  INV_X1    g428(.A(G472), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n615), .B1(new_n592), .B2(new_n279), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  AOI22_X1  g431(.A1(new_n535), .A2(new_n536), .B1(new_n538), .B2(new_n540), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n617), .A2(new_n618), .A3(new_n582), .ZN(new_n619));
  NOR3_X1   g433(.A1(new_n614), .A2(new_n619), .A3(new_n422), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n350), .B1(new_n346), .B2(new_n347), .ZN(new_n621));
  INV_X1    g435(.A(new_n347), .ZN(new_n622));
  AOI211_X1 g436(.A(KEYINPUT20), .B(new_n622), .C1(new_n340), .C2(new_n345), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(G475), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n416), .A2(new_n344), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT93), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n626), .A2(new_n627), .A3(new_n340), .ZN(new_n628));
  AOI21_X1  g442(.A(G902), .B1(new_n414), .B2(KEYINPUT93), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n625), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n624), .A2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(G478), .ZN(new_n632));
  OAI21_X1  g446(.A(KEYINPUT100), .B1(new_n381), .B2(new_n390), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(KEYINPUT33), .ZN(new_n634));
  OR2_X1    g448(.A1(new_n395), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(new_n395), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n632), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n395), .A2(new_n632), .A3(new_n279), .ZN(new_n638));
  NAND2_X1  g452(.A1(G478), .A2(G902), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n637), .A2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n631), .A2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n291), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n276), .A2(new_n282), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(KEYINPUT6), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n288), .B1(new_n646), .B2(new_n284), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n278), .A2(new_n279), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n644), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n649), .A2(KEYINPUT99), .A3(new_n292), .ZN(new_n650));
  INV_X1    g464(.A(new_n187), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT99), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n651), .B1(new_n294), .B2(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n406), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n650), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  AOI21_X1  g470(.A(KEYINPUT101), .B1(new_n643), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n352), .A2(new_n419), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(new_n641), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT101), .ZN(new_n660));
  NOR3_X1   g474(.A1(new_n659), .A2(new_n660), .A3(new_n655), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n620), .B1(new_n657), .B2(new_n661), .ZN(new_n662));
  XOR2_X1   g476(.A(KEYINPUT34), .B(G104), .Z(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G6));
  NAND3_X1  g478(.A1(new_n352), .A2(new_n419), .A3(new_n401), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  AOI21_X1  g480(.A(KEYINPUT102), .B1(new_n666), .B2(new_n656), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT102), .ZN(new_n668));
  NOR3_X1   g482(.A1(new_n665), .A2(new_n668), .A3(new_n655), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n620), .B1(new_n667), .B2(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(new_n193), .ZN(new_n671));
  XNOR2_X1  g485(.A(KEYINPUT103), .B(KEYINPUT35), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(G9));
  AOI21_X1  g487(.A(new_n616), .B1(new_n543), .B2(new_n592), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n522), .A2(KEYINPUT36), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n518), .B(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(new_n540), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n537), .A2(new_n677), .ZN(new_n678));
  AND2_X1   g492(.A1(new_n674), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n420), .A2(new_n497), .A3(new_n679), .ZN(new_n680));
  XOR2_X1   g494(.A(KEYINPUT37), .B(G110), .Z(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(G12));
  INV_X1    g496(.A(G900), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n403), .B1(new_n404), .B2(new_n683), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n665), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n650), .A2(new_n653), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  AND2_X1   g501(.A1(new_n537), .A2(new_n677), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n688), .B1(new_n595), .B2(new_n610), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n685), .A2(new_n497), .A3(new_n687), .A4(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G128), .ZN(G30));
  XOR2_X1   g505(.A(new_n684), .B(KEYINPUT39), .Z(new_n692));
  NAND2_X1  g506(.A1(new_n497), .A2(new_n692), .ZN(new_n693));
  OR2_X1    g507(.A1(new_n693), .A2(KEYINPUT40), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n649), .A2(new_n292), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(KEYINPUT38), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n696), .A2(new_n187), .A3(new_n401), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n599), .A2(new_n600), .ZN(new_n698));
  AOI21_X1  g512(.A(G902), .B1(new_n698), .B2(new_n579), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n556), .A2(new_n562), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(new_n560), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n615), .B1(new_n699), .B2(new_n701), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n702), .B1(new_n583), .B2(new_n594), .ZN(new_n703));
  NOR4_X1   g517(.A1(new_n697), .A2(new_n631), .A3(new_n678), .A4(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n693), .A2(KEYINPUT40), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n694), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G143), .ZN(G45));
  INV_X1    g521(.A(new_n684), .ZN(new_n708));
  OAI211_X1 g522(.A(new_n641), .B(new_n708), .C1(new_n624), .C2(new_n630), .ZN(new_n709));
  INV_X1    g523(.A(new_n709), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n710), .A2(new_n689), .A3(new_n497), .A4(new_n687), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G146), .ZN(G48));
  NAND3_X1  g526(.A1(new_n445), .A2(new_n455), .A3(new_n457), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n470), .B1(new_n713), .B2(new_n468), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n714), .B1(new_n485), .B2(new_n487), .ZN(new_n715));
  OAI21_X1  g529(.A(KEYINPUT104), .B1(new_n715), .B2(G902), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT104), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n481), .B1(new_n489), .B2(new_n717), .ZN(new_n718));
  AOI22_X1  g532(.A1(new_n716), .A2(new_n718), .B1(new_n483), .B2(new_n491), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n719), .A2(new_n611), .A3(new_n421), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n643), .A2(KEYINPUT101), .A3(new_n656), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n660), .B1(new_n659), .B2(new_n655), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n720), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  XOR2_X1   g537(.A(KEYINPUT41), .B(G113), .Z(new_n724));
  XNOR2_X1  g538(.A(new_n723), .B(new_n724), .ZN(G15));
  INV_X1    g539(.A(new_n720), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n726), .B1(new_n667), .B2(new_n669), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G116), .ZN(G18));
  NAND3_X1  g542(.A1(new_n719), .A2(new_n421), .A3(new_n687), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n595), .A2(new_n610), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n730), .A2(new_n631), .A3(new_n407), .A4(new_n678), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(new_n202), .ZN(G21));
  NAND3_X1  g547(.A1(new_n480), .A2(new_n717), .A3(new_n279), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n716), .A2(new_n734), .A3(G469), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n492), .A2(new_n421), .A3(new_n735), .ZN(new_n736));
  AND2_X1   g550(.A1(new_n601), .A2(new_n574), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n584), .B1(new_n737), .B2(new_n560), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n543), .B(KEYINPUT105), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n616), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(new_n618), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n736), .A2(new_n741), .ZN(new_n742));
  AND3_X1   g556(.A1(new_n650), .A2(new_n653), .A3(new_n401), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n658), .A2(new_n743), .A3(new_n654), .ZN(new_n744));
  INV_X1    g558(.A(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n742), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G122), .ZN(G24));
  NOR2_X1   g561(.A1(new_n736), .A2(new_n686), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n740), .A2(new_n678), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n709), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G125), .ZN(G27));
  INV_X1    g566(.A(KEYINPUT42), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n490), .B1(new_n489), .B2(new_n481), .ZN(new_n754));
  NOR4_X1   g568(.A1(new_n715), .A2(KEYINPUT82), .A3(G469), .A4(G902), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n496), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n649), .A2(new_n292), .A3(new_n187), .ZN(new_n757));
  INV_X1    g571(.A(new_n757), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n611), .A2(new_n756), .A3(new_n758), .A4(new_n421), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n753), .B1(new_n759), .B2(new_n709), .ZN(new_n760));
  NOR3_X1   g574(.A1(new_n614), .A2(new_n422), .A3(new_n757), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n761), .A2(KEYINPUT42), .A3(new_n611), .A4(new_n710), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G131), .ZN(G33));
  NAND3_X1  g578(.A1(new_n761), .A2(new_n611), .A3(new_n685), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G134), .ZN(G36));
  NOR2_X1   g580(.A1(new_n481), .A2(new_n279), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT45), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n494), .A2(new_n768), .ZN(new_n769));
  OAI221_X1 g583(.A(KEYINPUT45), .B1(new_n486), .B2(new_n458), .C1(new_n493), .C2(new_n470), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n769), .A2(G469), .A3(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT106), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n769), .A2(KEYINPUT106), .A3(new_n770), .A4(G469), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n767), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  AND2_X1   g589(.A1(new_n775), .A2(KEYINPUT46), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n492), .B1(new_n775), .B2(KEYINPUT46), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n421), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(new_n692), .ZN(new_n779));
  OR2_X1    g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(new_n780), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n658), .A2(new_n642), .ZN(new_n782));
  OR2_X1    g596(.A1(new_n782), .A2(KEYINPUT43), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(KEYINPUT43), .ZN(new_n784));
  AOI211_X1 g598(.A(new_n674), .B(new_n688), .C1(new_n783), .C2(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(KEYINPUT44), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n781), .A2(new_n786), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n758), .B1(new_n785), .B2(KEYINPUT44), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(new_n449), .ZN(G39));
  INV_X1    g604(.A(KEYINPUT47), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n778), .A2(new_n791), .ZN(new_n792));
  OAI211_X1 g606(.A(KEYINPUT47), .B(new_n421), .C1(new_n776), .C2(new_n777), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n730), .A2(new_n618), .A3(new_n757), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n794), .A2(new_n710), .A3(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT107), .ZN(new_n797));
  OR2_X1    g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n796), .A2(new_n797), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(G140), .ZN(G42));
  OR2_X1    g615(.A1(G952), .A2(G953), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT119), .ZN(new_n803));
  INV_X1    g617(.A(new_n403), .ZN(new_n804));
  NOR3_X1   g618(.A1(new_n736), .A2(new_n804), .A3(new_n757), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n703), .A2(new_n618), .ZN(new_n806));
  INV_X1    g620(.A(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n808), .A2(KEYINPUT115), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT115), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n805), .A2(new_n810), .A3(new_n807), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n809), .A2(new_n631), .A3(new_n642), .A4(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n782), .B(KEYINPUT43), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n813), .A2(new_n678), .A3(new_n740), .A4(new_n805), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n804), .B1(new_n783), .B2(new_n784), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n738), .A2(new_n739), .ZN(new_n816));
  AND3_X1   g630(.A1(new_n618), .A2(new_n617), .A3(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n719), .A2(new_n817), .A3(new_n421), .ZN(new_n818));
  NOR3_X1   g632(.A1(new_n818), .A2(new_n187), .A3(new_n696), .ZN(new_n819));
  AND3_X1   g633(.A1(new_n815), .A2(KEYINPUT50), .A3(new_n819), .ZN(new_n820));
  AOI21_X1  g634(.A(KEYINPUT50), .B1(new_n815), .B2(new_n819), .ZN(new_n821));
  OAI211_X1 g635(.A(new_n812), .B(new_n814), .C1(new_n820), .C2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n813), .A2(new_n403), .A3(new_n817), .A4(new_n758), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT113), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(new_n719), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n827), .A2(new_n421), .ZN(new_n828));
  INV_X1    g642(.A(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n792), .A2(new_n793), .A3(new_n829), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n815), .A2(KEYINPUT113), .A3(new_n817), .A4(new_n758), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n826), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n823), .A2(KEYINPUT116), .A3(KEYINPUT51), .A4(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT116), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n832), .A2(KEYINPUT51), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n834), .B1(new_n835), .B2(new_n822), .ZN(new_n836));
  AND2_X1   g650(.A1(new_n833), .A2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT51), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n826), .A2(new_n831), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n828), .B1(new_n794), .B2(KEYINPUT114), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT114), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n792), .A2(new_n841), .A3(new_n793), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n839), .B1(new_n840), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n838), .B1(new_n843), .B2(new_n822), .ZN(new_n844));
  AND3_X1   g658(.A1(new_n813), .A2(new_n611), .A3(new_n805), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT48), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(KEYINPUT118), .ZN(new_n847));
  OR2_X1    g661(.A1(new_n846), .A2(KEYINPUT118), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n845), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n849), .B1(new_n847), .B2(new_n845), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n809), .A2(new_n643), .A3(new_n811), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n815), .A2(new_n748), .A3(new_n817), .ZN(new_n852));
  XNOR2_X1  g666(.A(new_n402), .B(KEYINPUT117), .ZN(new_n853));
  NOR4_X1   g667(.A1(new_n850), .A2(new_n851), .A3(new_n852), .A4(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n844), .A2(new_n854), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n803), .B1(new_n837), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n833), .A2(new_n836), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n857), .A2(new_n844), .A3(KEYINPUT119), .A4(new_n854), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT111), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT52), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n658), .A2(new_n743), .ZN(new_n862));
  INV_X1    g676(.A(new_n702), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n592), .A2(new_n593), .A3(new_n543), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n593), .B1(new_n592), .B2(new_n543), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n863), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n866), .A2(new_n688), .A3(new_n708), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n862), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g682(.A(KEYINPUT109), .B1(new_n868), .B2(new_n497), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n703), .A2(new_n678), .A3(new_n684), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n650), .A2(new_n653), .A3(new_n401), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n871), .B1(new_n419), .B2(new_n352), .ZN(new_n872));
  AND4_X1   g686(.A1(KEYINPUT109), .A2(new_n870), .A3(new_n497), .A4(new_n872), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n869), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n751), .A2(new_n690), .A3(new_n711), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n861), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  AND3_X1   g690(.A1(new_n751), .A2(new_n690), .A3(new_n711), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n870), .A2(new_n872), .A3(new_n497), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT109), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n868), .A2(KEYINPUT109), .A3(new_n497), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n877), .A2(KEYINPUT52), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n876), .A2(new_n883), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n726), .B1(new_n657), .B2(new_n661), .ZN(new_n885));
  INV_X1    g699(.A(new_n731), .ZN(new_n886));
  AOI22_X1  g700(.A1(new_n886), .A2(new_n748), .B1(new_n742), .B2(new_n745), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n763), .A2(new_n885), .A3(new_n887), .A4(new_n727), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n398), .A2(new_n400), .A3(new_n708), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n757), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n890), .A2(new_n419), .A3(new_n352), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT108), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n890), .A2(new_n352), .A3(KEYINPUT108), .A4(new_n419), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n893), .A2(new_n497), .A3(new_n689), .A4(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n750), .A2(new_n761), .ZN(new_n896));
  AND3_X1   g710(.A1(new_n895), .A2(new_n765), .A3(new_n896), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n665), .B1(new_n631), .B2(new_n642), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n295), .A2(new_n406), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n620), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  OAI211_X1 g714(.A(new_n420), .B(new_n497), .C1(new_n679), .C2(new_n611), .ZN(new_n901));
  AND2_X1   g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n897), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n888), .A2(new_n903), .ZN(new_n904));
  AND2_X1   g718(.A1(new_n884), .A2(new_n904), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n860), .B1(new_n905), .B2(KEYINPUT53), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n876), .A2(KEYINPUT110), .A3(new_n883), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT110), .ZN(new_n908));
  OAI211_X1 g722(.A(new_n908), .B(new_n861), .C1(new_n874), .C2(new_n875), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT112), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n888), .A2(new_n911), .ZN(new_n912));
  OAI22_X1  g726(.A1(new_n729), .A2(new_n731), .B1(new_n818), .B2(new_n744), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n723), .A2(new_n913), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n914), .A2(KEYINPUT112), .A3(new_n727), .A4(new_n763), .ZN(new_n915));
  AND3_X1   g729(.A1(new_n897), .A2(KEYINPUT53), .A3(new_n902), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n912), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  OR2_X1    g731(.A1(new_n910), .A2(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT54), .ZN(new_n919));
  AOI21_X1  g733(.A(KEYINPUT53), .B1(new_n884), .B2(new_n904), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(KEYINPUT111), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n906), .A2(new_n918), .A3(new_n919), .A4(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT53), .ZN(new_n923));
  OR2_X1    g737(.A1(new_n905), .A2(new_n923), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n907), .A2(new_n923), .A3(new_n904), .A4(new_n909), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n924), .A2(KEYINPUT54), .A3(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n922), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n802), .B1(new_n859), .B2(new_n927), .ZN(new_n928));
  OR2_X1    g742(.A1(new_n827), .A2(KEYINPUT49), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n618), .A2(new_n421), .A3(new_n189), .ZN(new_n930));
  NOR3_X1   g744(.A1(new_n696), .A2(new_n866), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n827), .A2(KEYINPUT49), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n929), .A2(new_n931), .A3(new_n782), .A4(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n928), .A2(new_n933), .ZN(G75));
  NOR2_X1   g748(.A1(new_n240), .A2(G952), .ZN(new_n935));
  INV_X1    g749(.A(new_n935), .ZN(new_n936));
  OAI22_X1  g750(.A1(new_n920), .A2(KEYINPUT111), .B1(new_n910), .B2(new_n917), .ZN(new_n937));
  AOI211_X1 g751(.A(new_n860), .B(KEYINPUT53), .C1(new_n884), .C2(new_n904), .ZN(new_n938));
  OAI211_X1 g752(.A(G210), .B(G902), .C1(new_n937), .C2(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT56), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n286), .B(KEYINPUT120), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(KEYINPUT55), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(new_n289), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n936), .B1(new_n941), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n941), .A2(new_n944), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(KEYINPUT121), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT121), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n941), .A2(new_n948), .A3(new_n944), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n945), .B1(new_n947), .B2(new_n949), .ZN(G51));
  OAI21_X1  g764(.A(KEYINPUT54), .B1(new_n937), .B2(new_n938), .ZN(new_n951));
  AND2_X1   g765(.A1(new_n922), .A2(new_n951), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n767), .B(KEYINPUT57), .Z(new_n953));
  OAI21_X1  g767(.A(new_n480), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n906), .A2(new_n918), .A3(new_n921), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n955), .A2(G902), .A3(new_n773), .A4(new_n774), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n935), .B1(new_n954), .B2(new_n956), .ZN(G54));
  NAND2_X1  g771(.A1(KEYINPUT58), .A2(G475), .ZN(new_n958));
  INV_X1    g772(.A(new_n958), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n955), .A2(G902), .A3(new_n959), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n960), .A2(new_n340), .A3(new_n345), .ZN(new_n961));
  NAND4_X1  g775(.A1(new_n955), .A2(G902), .A3(new_n346), .A4(new_n959), .ZN(new_n962));
  AND3_X1   g776(.A1(new_n961), .A2(new_n936), .A3(new_n962), .ZN(G60));
  AND2_X1   g777(.A1(new_n635), .A2(new_n636), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n639), .B(KEYINPUT59), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n936), .B1(new_n952), .B2(new_n966), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n964), .B1(new_n927), .B2(new_n965), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n967), .A2(new_n968), .ZN(G63));
  NOR2_X1   g783(.A1(new_n937), .A2(new_n938), .ZN(new_n970));
  NAND2_X1  g784(.A1(G217), .A2(G902), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n971), .B(KEYINPUT60), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n532), .B1(new_n970), .B2(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(new_n972), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n955), .A2(new_n676), .A3(new_n974), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n973), .A2(new_n936), .A3(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT61), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n973), .A2(new_n975), .A3(KEYINPUT61), .A4(new_n936), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n978), .A2(new_n979), .ZN(G66));
  INV_X1    g794(.A(new_n239), .ZN(new_n981));
  OAI21_X1  g795(.A(G953), .B1(new_n981), .B2(new_n405), .ZN(new_n982));
  AND3_X1   g796(.A1(new_n914), .A2(new_n727), .A3(new_n902), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n982), .B1(new_n983), .B2(G953), .ZN(new_n984));
  INV_X1    g798(.A(G898), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n942), .B1(new_n985), .B2(G953), .ZN(new_n986));
  XOR2_X1   g800(.A(new_n984), .B(new_n986), .Z(G69));
  NAND2_X1  g801(.A1(new_n550), .A2(new_n555), .ZN(new_n988));
  XOR2_X1   g802(.A(new_n988), .B(KEYINPUT122), .Z(new_n989));
  XOR2_X1   g803(.A(new_n989), .B(new_n341), .Z(new_n990));
  NAND2_X1  g804(.A1(new_n990), .A2(KEYINPUT125), .ZN(new_n991));
  OAI211_X1 g805(.A(new_n991), .B(G953), .C1(new_n424), .C2(new_n683), .ZN(new_n992));
  XOR2_X1   g806(.A(new_n992), .B(KEYINPUT126), .Z(new_n993));
  INV_X1    g807(.A(new_n993), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n877), .B1(new_n787), .B2(new_n788), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n995), .B(KEYINPUT124), .ZN(new_n996));
  INV_X1    g810(.A(new_n611), .ZN(new_n997));
  NOR2_X1   g811(.A1(new_n997), .A2(new_n862), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n781), .A2(new_n998), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n999), .A2(new_n763), .A3(new_n765), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n1000), .B1(new_n798), .B2(new_n799), .ZN(new_n1001));
  INV_X1    g815(.A(new_n1001), .ZN(new_n1002));
  OAI211_X1 g816(.A(new_n240), .B(new_n990), .C1(new_n996), .C2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n683), .A2(G953), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n898), .B(KEYINPUT123), .ZN(new_n1006));
  NOR3_X1   g820(.A1(new_n1006), .A2(new_n779), .A3(new_n759), .ZN(new_n1007));
  NOR2_X1   g821(.A1(new_n789), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n706), .A2(new_n877), .ZN(new_n1009));
  XOR2_X1   g823(.A(new_n1009), .B(KEYINPUT62), .Z(new_n1010));
  NAND3_X1  g824(.A1(new_n800), .A2(new_n1008), .A3(new_n1010), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n990), .B1(new_n1011), .B2(new_n240), .ZN(new_n1012));
  OAI21_X1  g826(.A(new_n994), .B1(new_n1005), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g827(.A(new_n1012), .ZN(new_n1014));
  NAND4_X1  g828(.A1(new_n1014), .A2(new_n1003), .A3(new_n993), .A4(new_n1004), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1013), .A2(new_n1015), .ZN(G72));
  INV_X1    g830(.A(KEYINPUT124), .ZN(new_n1017));
  AND2_X1   g831(.A1(new_n995), .A2(new_n1017), .ZN(new_n1018));
  OAI211_X1 g832(.A(KEYINPUT124), .B(new_n877), .C1(new_n787), .C2(new_n788), .ZN(new_n1019));
  INV_X1    g833(.A(new_n1019), .ZN(new_n1020));
  OAI211_X1 g834(.A(new_n1001), .B(new_n983), .C1(new_n1018), .C2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g835(.A1(G472), .A2(G902), .ZN(new_n1022));
  XOR2_X1   g836(.A(new_n1022), .B(KEYINPUT63), .Z(new_n1023));
  XOR2_X1   g837(.A(new_n1023), .B(KEYINPUT127), .Z(new_n1024));
  AOI211_X1 g838(.A(new_n560), .B(new_n700), .C1(new_n1021), .C2(new_n1024), .ZN(new_n1025));
  NAND4_X1  g839(.A1(new_n800), .A2(new_n1008), .A3(new_n983), .A4(new_n1010), .ZN(new_n1026));
  AOI21_X1  g840(.A(new_n701), .B1(new_n1026), .B2(new_n1024), .ZN(new_n1027));
  INV_X1    g841(.A(new_n563), .ZN(new_n1028));
  OR2_X1    g842(.A1(new_n1028), .A2(new_n606), .ZN(new_n1029));
  AND4_X1   g843(.A1(new_n924), .A2(new_n925), .A3(new_n1023), .A4(new_n1029), .ZN(new_n1030));
  NOR4_X1   g844(.A1(new_n1025), .A2(new_n1027), .A3(new_n935), .A4(new_n1030), .ZN(G57));
endmodule


