//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 1 1 0 1 1 1 0 1 1 1 0 1 1 1 0 0 1 0 1 1 1 1 0 1 0 1 0 0 1 0 1 1 1 1 0 1 0 0 1 1 1 1 0 0 0 1 1 0 1 1 0 0 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:29 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1210, new_n1211, new_n1213,
    new_n1214, new_n1215, new_n1216, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G68), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G250), .ZN(new_n206));
  INV_X1    g0006(.A(KEYINPUT64), .ZN(new_n207));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  OAI21_X1  g0011(.A(new_n207), .B1(new_n211), .B2(G13), .ZN(new_n212));
  INV_X1    g0012(.A(G13), .ZN(new_n213));
  NAND3_X1  g0013(.A1(new_n210), .A2(KEYINPUT64), .A3(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(G257), .ZN(new_n217));
  INV_X1    g0017(.A(G264), .ZN(new_n218));
  AOI211_X1 g0018(.A(new_n206), .B(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  XNOR2_X1  g0019(.A(KEYINPUT65), .B(G20), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G1), .A2(G13), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(G50), .B1(G58), .B2(G68), .ZN(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(new_n219), .A2(KEYINPUT0), .B1(new_n222), .B2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n225), .B1(KEYINPUT0), .B2(new_n219), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n227));
  INV_X1    g0027(.A(G77), .ZN(new_n228));
  INV_X1    g0028(.A(G244), .ZN(new_n229));
  INV_X1    g0029(.A(G107), .ZN(new_n230));
  OAI221_X1 g0030(.A(new_n227), .B1(new_n228), .B2(new_n229), .C1(new_n230), .C2(new_n218), .ZN(new_n231));
  AOI22_X1  g0031(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n232));
  INV_X1    g0032(.A(G232), .ZN(new_n233));
  INV_X1    g0033(.A(G97), .ZN(new_n234));
  OAI221_X1 g0034(.A(new_n232), .B1(new_n202), .B2(new_n233), .C1(new_n234), .C2(new_n217), .ZN(new_n235));
  OAI21_X1  g0035(.A(new_n211), .B1(new_n231), .B2(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT1), .ZN(new_n237));
  NOR2_X1   g0037(.A1(new_n226), .A2(new_n237), .ZN(G361));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(KEYINPUT2), .B(G226), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G264), .B(G270), .Z(new_n243));
  XNOR2_X1  g0043(.A(G250), .B(G257), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G358));
  XOR2_X1   g0046(.A(G68), .B(G77), .Z(new_n247));
  XNOR2_X1  g0047(.A(G50), .B(G58), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(G87), .B(G97), .Z(new_n250));
  XNOR2_X1  g0050(.A(G107), .B(G116), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n249), .B(new_n252), .ZN(G351));
  AOI21_X1  g0053(.A(new_n221), .B1(G33), .B2(G41), .ZN(new_n254));
  INV_X1    g0054(.A(G274), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n256));
  NOR3_X1   g0056(.A1(new_n254), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(new_n256), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n254), .A2(new_n258), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n257), .B1(G226), .B2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  AND2_X1   g0061(.A1(KEYINPUT3), .A2(G33), .ZN(new_n262));
  NOR2_X1   g0062(.A1(KEYINPUT3), .A2(G33), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n264), .A2(G1698), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G222), .ZN(new_n266));
  OR2_X1    g0066(.A1(KEYINPUT3), .A2(G33), .ZN(new_n267));
  NAND2_X1  g0067(.A1(KEYINPUT3), .A2(G33), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G223), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(G1698), .ZN(new_n271));
  OAI221_X1 g0071(.A(new_n266), .B1(new_n228), .B2(new_n269), .C1(new_n270), .C2(new_n271), .ZN(new_n272));
  OR2_X1    g0072(.A1(new_n272), .A2(KEYINPUT66), .ZN(new_n273));
  INV_X1    g0073(.A(new_n254), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n274), .B1(new_n272), .B2(KEYINPUT66), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n261), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G190), .ZN(new_n277));
  NOR2_X1   g0077(.A1(G20), .A2(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G150), .ZN(new_n279));
  OAI21_X1  g0079(.A(G20), .B1(new_n203), .B2(G68), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n220), .A2(G33), .ZN(new_n281));
  XNOR2_X1  g0081(.A(KEYINPUT8), .B(G58), .ZN(new_n282));
  OAI211_X1 g0082(.A(new_n279), .B(new_n280), .C1(new_n281), .C2(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(new_n221), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  NOR3_X1   g0086(.A1(new_n213), .A2(new_n209), .A3(G1), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n287), .A2(new_n285), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n208), .A2(G20), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G50), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  AOI22_X1  g0091(.A1(new_n288), .A2(new_n291), .B1(new_n201), .B2(new_n287), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT71), .ZN(new_n293));
  OR2_X1    g0093(.A1(new_n293), .A2(KEYINPUT9), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n286), .A2(new_n292), .A3(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n293), .A2(KEYINPUT9), .ZN(new_n296));
  XOR2_X1   g0096(.A(new_n295), .B(new_n296), .Z(new_n297));
  INV_X1    g0097(.A(G200), .ZN(new_n298));
  OAI211_X1 g0098(.A(new_n277), .B(new_n297), .C1(new_n298), .C2(new_n276), .ZN(new_n299));
  XNOR2_X1  g0099(.A(new_n299), .B(KEYINPUT10), .ZN(new_n300));
  INV_X1    g0100(.A(G179), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n276), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n286), .A2(new_n292), .ZN(new_n303));
  OAI211_X1 g0103(.A(new_n302), .B(new_n303), .C1(G169), .C2(new_n276), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n300), .A2(new_n304), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n213), .A2(G1), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(G20), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n307), .A2(G68), .ZN(new_n308));
  XNOR2_X1  g0108(.A(new_n308), .B(KEYINPUT12), .ZN(new_n309));
  INV_X1    g0109(.A(new_n285), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n220), .A2(G33), .A3(G77), .ZN(new_n311));
  INV_X1    g0111(.A(G68), .ZN(new_n312));
  AOI22_X1  g0112(.A1(new_n278), .A2(G50), .B1(G20), .B2(new_n312), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n310), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n309), .B1(new_n314), .B2(KEYINPUT11), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n310), .A2(new_n307), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT68), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n288), .A2(KEYINPUT68), .ZN(new_n319));
  AND2_X1   g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n320), .A2(G68), .A3(new_n289), .ZN(new_n321));
  OR2_X1    g0121(.A1(new_n314), .A2(KEYINPUT11), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n315), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT14), .ZN(new_n324));
  NAND2_X1  g0124(.A1(G33), .A2(G97), .ZN(new_n325));
  INV_X1    g0125(.A(G1698), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n269), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(G226), .ZN(new_n328));
  OAI221_X1 g0128(.A(new_n325), .B1(new_n327), .B2(new_n328), .C1(new_n233), .C2(new_n271), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(new_n254), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT13), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n257), .B1(G238), .B2(new_n259), .ZN(new_n332));
  AND3_X1   g0132(.A1(new_n330), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n331), .B1(new_n330), .B2(new_n332), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n324), .B(G169), .C1(new_n333), .C2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n330), .A2(new_n332), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(KEYINPUT13), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n330), .A2(new_n331), .A3(new_n332), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n337), .A2(G179), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n335), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n337), .A2(new_n338), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n324), .B1(new_n341), .B2(G169), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n323), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  OAI21_X1  g0143(.A(G200), .B1(new_n333), .B2(new_n334), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n337), .A2(G190), .A3(new_n338), .ZN(new_n345));
  INV_X1    g0145(.A(new_n323), .ZN(new_n346));
  AND3_X1   g0146(.A1(new_n344), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n343), .A2(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n257), .B1(G244), .B2(new_n259), .ZN(new_n350));
  INV_X1    g0150(.A(G238), .ZN(new_n351));
  OAI22_X1  g0151(.A1(new_n271), .A2(new_n351), .B1(new_n230), .B2(new_n269), .ZN(new_n352));
  OR3_X1    g0152(.A1(new_n327), .A2(KEYINPUT67), .A3(new_n233), .ZN(new_n353));
  OAI21_X1  g0153(.A(KEYINPUT67), .B1(new_n327), .B2(new_n233), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n352), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n350), .B1(new_n355), .B2(new_n274), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT70), .ZN(new_n357));
  OR3_X1    g0157(.A1(new_n356), .A2(new_n357), .A3(G179), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n357), .B1(new_n356), .B2(G179), .ZN(new_n359));
  INV_X1    g0159(.A(G169), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n320), .A2(G77), .A3(new_n289), .ZN(new_n361));
  INV_X1    g0161(.A(new_n282), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n209), .A2(KEYINPUT65), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT65), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(G20), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  AOI22_X1  g0166(.A1(new_n362), .A2(new_n278), .B1(new_n366), .B2(G77), .ZN(new_n367));
  XNOR2_X1  g0167(.A(KEYINPUT15), .B(G87), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n367), .B1(new_n281), .B2(new_n368), .ZN(new_n369));
  AOI22_X1  g0169(.A1(new_n369), .A2(new_n285), .B1(new_n228), .B2(new_n287), .ZN(new_n370));
  AOI22_X1  g0170(.A1(new_n356), .A2(new_n360), .B1(new_n361), .B2(new_n370), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n358), .A2(new_n359), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n370), .A2(new_n361), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n373), .B1(G200), .B2(new_n356), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT69), .ZN(new_n375));
  INV_X1    g0175(.A(G190), .ZN(new_n376));
  OAI22_X1  g0176(.A1(new_n374), .A2(new_n375), .B1(new_n376), .B2(new_n356), .ZN(new_n377));
  AND2_X1   g0177(.A1(new_n374), .A2(new_n375), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n372), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NOR3_X1   g0179(.A1(new_n305), .A2(new_n349), .A3(new_n379), .ZN(new_n380));
  XNOR2_X1  g0180(.A(G58), .B(G68), .ZN(new_n381));
  AOI22_X1  g0181(.A1(new_n381), .A2(G20), .B1(G159), .B2(new_n278), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n264), .A2(new_n220), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT7), .ZN(new_n384));
  NOR3_X1   g0184(.A1(new_n262), .A2(new_n263), .A3(G20), .ZN(new_n385));
  XNOR2_X1  g0185(.A(KEYINPUT72), .B(KEYINPUT7), .ZN(new_n386));
  AOI22_X1  g0186(.A1(new_n383), .A2(new_n384), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n382), .B1(new_n387), .B2(new_n312), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT16), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n285), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT73), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n391), .B1(new_n385), .B2(new_n386), .ZN(new_n392));
  XOR2_X1   g0192(.A(KEYINPUT72), .B(KEYINPUT7), .Z(new_n393));
  NAND3_X1  g0193(.A1(new_n267), .A2(new_n209), .A3(new_n268), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n393), .A2(new_n394), .A3(KEYINPUT73), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n264), .A2(new_n220), .A3(KEYINPUT7), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n392), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(G68), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT74), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n397), .A2(KEYINPUT74), .A3(G68), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n400), .A2(new_n382), .A3(new_n401), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n390), .B1(new_n402), .B2(new_n389), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n362), .A2(new_n289), .ZN(new_n405));
  OAI22_X1  g0205(.A1(new_n405), .A2(new_n316), .B1(new_n307), .B2(new_n362), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n257), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n274), .A2(G232), .A3(new_n256), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n328), .A2(G1698), .ZN(new_n411));
  OAI211_X1 g0211(.A(new_n269), .B(new_n411), .C1(G223), .C2(G1698), .ZN(new_n412));
  NAND2_X1  g0212(.A1(G33), .A2(G87), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n274), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n410), .A2(new_n414), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n415), .A2(new_n298), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n416), .B1(new_n415), .B2(G190), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n404), .A2(KEYINPUT17), .A3(new_n407), .A4(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(new_n382), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n419), .B1(new_n398), .B2(new_n399), .ZN(new_n420));
  AOI21_X1  g0220(.A(KEYINPUT16), .B1(new_n420), .B2(new_n401), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n417), .B(new_n407), .C1(new_n421), .C2(new_n390), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT17), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n418), .A2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT76), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT18), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n412), .A2(new_n413), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(new_n254), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n257), .B1(G232), .B2(new_n259), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n429), .A2(G179), .A3(new_n430), .ZN(new_n431));
  OAI21_X1  g0231(.A(G169), .B1(new_n410), .B2(new_n414), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT75), .ZN(new_n433));
  AND3_X1   g0233(.A1(new_n431), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n433), .B1(new_n431), .B2(new_n432), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  OAI211_X1 g0236(.A(new_n427), .B(new_n436), .C1(new_n403), .C2(new_n406), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n407), .B1(new_n421), .B2(new_n390), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n427), .B1(new_n439), .B2(new_n436), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n426), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n436), .B1(new_n403), .B2(new_n406), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(KEYINPUT18), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n443), .A2(KEYINPUT76), .A3(new_n437), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n425), .B1(new_n441), .B2(new_n444), .ZN(new_n445));
  AND2_X1   g0245(.A1(new_n380), .A2(new_n445), .ZN(new_n446));
  XOR2_X1   g0246(.A(KEYINPUT80), .B(KEYINPUT19), .Z(new_n447));
  OAI21_X1  g0247(.A(new_n220), .B1(new_n447), .B2(new_n325), .ZN(new_n448));
  INV_X1    g0248(.A(G87), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n449), .A2(new_n234), .A3(new_n230), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n447), .B1(new_n281), .B2(new_n234), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n269), .A2(new_n220), .A3(G68), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n451), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT81), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n310), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n451), .A2(KEYINPUT81), .A3(new_n452), .A4(new_n453), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n208), .A2(G33), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n288), .A2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n368), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n462), .A2(new_n307), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n458), .A2(new_n463), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(KEYINPUT82), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n464), .B1(new_n456), .B2(new_n457), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT82), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n468), .A2(new_n469), .A3(new_n463), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n269), .A2(G238), .A3(new_n326), .ZN(new_n472));
  INV_X1    g0272(.A(G33), .ZN(new_n473));
  INV_X1    g0273(.A(G116), .ZN(new_n474));
  OAI221_X1 g0274(.A(new_n472), .B1(new_n473), .B2(new_n474), .C1(new_n271), .C2(new_n229), .ZN(new_n475));
  INV_X1    g0275(.A(G45), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n476), .A2(G1), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(new_n255), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n477), .A2(G250), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n479), .A2(new_n254), .ZN(new_n480));
  AOI22_X1  g0280(.A1(new_n475), .A2(new_n254), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n481), .A2(G169), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n482), .B1(new_n301), .B2(new_n481), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n468), .B1(new_n449), .B2(new_n460), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(new_n481), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(G200), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n481), .A2(G190), .ZN(new_n488));
  AND2_X1   g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  AOI22_X1  g0289(.A1(new_n471), .A2(new_n483), .B1(new_n485), .B2(new_n489), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n474), .B1(new_n208), .B2(G33), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n320), .A2(KEYINPUT83), .A3(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n318), .A2(new_n319), .A3(new_n491), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT83), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(G33), .A2(G283), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n220), .B(new_n497), .C1(G33), .C2(new_n234), .ZN(new_n498));
  AOI22_X1  g0298(.A1(new_n284), .A2(new_n221), .B1(G20), .B2(new_n474), .ZN(new_n499));
  AND3_X1   g0299(.A1(new_n498), .A2(KEYINPUT20), .A3(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(KEYINPUT20), .B1(new_n498), .B2(new_n499), .ZN(new_n501));
  OAI22_X1  g0301(.A1(new_n500), .A2(new_n501), .B1(G116), .B2(new_n307), .ZN(new_n502));
  INV_X1    g0302(.A(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n496), .A2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT21), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n269), .A2(G257), .A3(new_n326), .ZN(new_n506));
  INV_X1    g0306(.A(G303), .ZN(new_n507));
  OAI221_X1 g0307(.A(new_n506), .B1(new_n507), .B2(new_n269), .C1(new_n271), .C2(new_n218), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(new_n254), .ZN(new_n509));
  XNOR2_X1  g0309(.A(KEYINPUT5), .B(G41), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(new_n477), .ZN(new_n511));
  NOR3_X1   g0311(.A1(new_n511), .A2(new_n255), .A3(new_n254), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n274), .ZN(new_n513));
  INV_X1    g0313(.A(new_n513), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n512), .B1(new_n514), .B2(G270), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n360), .B1(new_n509), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n504), .A2(new_n505), .A3(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n502), .B1(new_n492), .B2(new_n495), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n509), .A2(new_n515), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(G169), .ZN(new_n520));
  OAI21_X1  g0320(.A(KEYINPUT21), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n517), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n509), .A2(new_n515), .A3(G179), .ZN(new_n523));
  INV_X1    g0323(.A(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n504), .A2(KEYINPUT84), .A3(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT84), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n526), .B1(new_n518), .B2(new_n523), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n519), .A2(G200), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n518), .B(new_n529), .C1(new_n376), .C2(new_n519), .ZN(new_n530));
  AND3_X1   g0330(.A1(new_n522), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n278), .A2(G77), .ZN(new_n532));
  XNOR2_X1  g0332(.A(new_n532), .B(KEYINPUT77), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT6), .ZN(new_n534));
  NOR3_X1   g0334(.A1(new_n534), .A2(new_n234), .A3(G107), .ZN(new_n535));
  XNOR2_X1  g0335(.A(G97), .B(G107), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n535), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n533), .B1(new_n220), .B2(new_n537), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n538), .B1(G107), .B2(new_n397), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n539), .A2(new_n310), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n287), .A2(new_n234), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n541), .B1(new_n460), .B2(new_n234), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n269), .A2(G244), .A3(new_n326), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT78), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n545), .A2(KEYINPUT4), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(new_n546), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n269), .A2(new_n548), .A3(G244), .A4(new_n326), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n269), .A2(G250), .A3(G1698), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n547), .A2(new_n497), .A3(new_n549), .A4(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(new_n254), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n274), .A2(G274), .A3(new_n477), .A4(new_n510), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n553), .B1(new_n513), .B2(new_n217), .ZN(new_n554));
  INV_X1    g0354(.A(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n552), .A2(new_n555), .A3(new_n301), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n554), .B1(new_n551), .B2(new_n254), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n556), .B1(G169), .B2(new_n557), .ZN(new_n558));
  OAI21_X1  g0358(.A(KEYINPUT79), .B1(new_n543), .B2(new_n558), .ZN(new_n559));
  OAI221_X1 g0359(.A(new_n541), .B1(new_n234), .B2(new_n460), .C1(new_n539), .C2(new_n310), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT79), .ZN(new_n561));
  INV_X1    g0361(.A(new_n557), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(new_n360), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n560), .A2(new_n561), .A3(new_n563), .A4(new_n556), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n562), .A2(G200), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n557), .A2(G190), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n543), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n559), .A2(new_n564), .A3(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n269), .A2(G257), .A3(G1698), .ZN(new_n569));
  NAND2_X1  g0369(.A1(G33), .A2(G294), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n569), .B(new_n570), .C1(new_n327), .C2(new_n206), .ZN(new_n571));
  AOI22_X1  g0371(.A1(new_n571), .A2(new_n254), .B1(new_n514), .B2(G264), .ZN(new_n572));
  AOI21_X1  g0372(.A(G169), .B1(new_n572), .B2(new_n553), .ZN(new_n573));
  AND2_X1   g0373(.A1(new_n572), .A2(new_n553), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n573), .B1(new_n301), .B2(new_n574), .ZN(new_n575));
  NOR2_X1   g0375(.A1(KEYINPUT23), .A2(G107), .ZN(new_n576));
  AND3_X1   g0376(.A1(new_n366), .A2(KEYINPUT85), .A3(new_n576), .ZN(new_n577));
  AOI21_X1  g0377(.A(KEYINPUT85), .B1(new_n366), .B2(new_n576), .ZN(new_n578));
  NOR3_X1   g0378(.A1(new_n473), .A2(new_n474), .A3(G20), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT23), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n580), .B1(G20), .B2(new_n230), .ZN(new_n581));
  NOR4_X1   g0381(.A1(new_n577), .A2(new_n578), .A3(new_n579), .A4(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n269), .A2(new_n220), .A3(G87), .ZN(new_n583));
  XNOR2_X1  g0383(.A(new_n583), .B(KEYINPUT22), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(KEYINPUT24), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT24), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n582), .A2(new_n584), .A3(new_n587), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n310), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n306), .A2(G20), .A3(new_n230), .ZN(new_n590));
  XNOR2_X1  g0390(.A(new_n590), .B(KEYINPUT25), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n591), .B1(new_n461), .B2(G107), .ZN(new_n592));
  INV_X1    g0392(.A(new_n592), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n575), .B1(new_n589), .B2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(new_n588), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n587), .B1(new_n582), .B2(new_n584), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n285), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n298), .B1(new_n572), .B2(new_n553), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n571), .A2(new_n254), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n514), .A2(G264), .ZN(new_n600));
  AND4_X1   g0400(.A1(G190), .A2(new_n599), .A3(new_n553), .A4(new_n600), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n597), .A2(new_n602), .A3(new_n592), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n594), .A2(new_n603), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n568), .A2(new_n604), .ZN(new_n605));
  AND4_X1   g0405(.A1(new_n446), .A2(new_n490), .A3(new_n531), .A4(new_n605), .ZN(G372));
  INV_X1    g0406(.A(new_n470), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n469), .B1(new_n468), .B2(new_n463), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n483), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n485), .A2(new_n489), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n559), .A2(new_n564), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  XOR2_X1   g0412(.A(KEYINPUT87), .B(KEYINPUT26), .Z(new_n613));
  NOR2_X1   g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT26), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT86), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n486), .A2(new_n616), .A3(G200), .ZN(new_n617));
  OAI21_X1  g0417(.A(KEYINPUT86), .B1(new_n481), .B2(new_n298), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n617), .A2(new_n618), .A3(new_n488), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n484), .A2(new_n619), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n620), .B1(new_n471), .B2(new_n483), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n543), .A2(new_n558), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n614), .B1(new_n615), .B2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n603), .ZN(new_n625));
  NOR3_X1   g0425(.A1(new_n568), .A2(new_n625), .A3(new_n620), .ZN(new_n626));
  AND2_X1   g0426(.A1(new_n522), .A2(new_n528), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(new_n594), .ZN(new_n628));
  AOI22_X1  g0428(.A1(new_n626), .A2(new_n628), .B1(new_n471), .B2(new_n483), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n446), .B1(new_n624), .B2(new_n630), .ZN(new_n631));
  OR2_X1    g0431(.A1(new_n347), .A2(new_n372), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n425), .B1(new_n632), .B2(new_n343), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n431), .A2(new_n432), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n634), .B1(new_n403), .B2(new_n406), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(KEYINPUT18), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n439), .A2(new_n427), .A3(new_n634), .ZN(new_n637));
  AND2_X1   g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n300), .B1(new_n633), .B2(new_n639), .ZN(new_n640));
  AND2_X1   g0440(.A1(new_n640), .A2(new_n304), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n631), .A2(new_n641), .ZN(G369));
  NAND2_X1  g0442(.A1(new_n220), .A2(new_n306), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(KEYINPUT27), .ZN(new_n644));
  XNOR2_X1  g0444(.A(new_n644), .B(KEYINPUT88), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n643), .A2(KEYINPUT27), .ZN(new_n646));
  INV_X1    g0446(.A(G213), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n650), .A2(KEYINPUT89), .A3(G343), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT89), .ZN(new_n652));
  INV_X1    g0452(.A(G343), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n652), .B1(new_n649), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(new_n504), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n531), .A2(new_n656), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n657), .B1(new_n627), .B2(new_n656), .ZN(new_n658));
  XOR2_X1   g0458(.A(KEYINPUT90), .B(G330), .Z(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  AND2_X1   g0460(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n604), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n655), .B1(new_n589), .B2(new_n593), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  AND2_X1   g0464(.A1(new_n651), .A2(new_n654), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n664), .B1(new_n594), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n661), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n627), .A2(new_n655), .ZN(new_n668));
  INV_X1    g0468(.A(new_n594), .ZN(new_n669));
  XNOR2_X1  g0469(.A(new_n655), .B(KEYINPUT91), .ZN(new_n670));
  AOI22_X1  g0470(.A1(new_n668), .A2(new_n662), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n667), .A2(new_n671), .ZN(G399));
  NOR2_X1   g0472(.A1(new_n216), .A2(G41), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n450), .A2(G116), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NOR3_X1   g0475(.A1(new_n673), .A2(new_n208), .A3(new_n675), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n676), .B1(new_n224), .B2(new_n673), .ZN(new_n677));
  XNOR2_X1  g0477(.A(new_n677), .B(KEYINPUT92), .ZN(new_n678));
  XOR2_X1   g0478(.A(new_n678), .B(KEYINPUT28), .Z(new_n679));
  OR2_X1    g0479(.A1(new_n484), .A2(new_n619), .ZN(new_n680));
  NAND4_X1  g0480(.A1(new_n609), .A2(KEYINPUT26), .A3(new_n680), .A4(new_n622), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT94), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n621), .A2(KEYINPUT94), .A3(KEYINPUT26), .A4(new_n622), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n612), .A2(new_n613), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n683), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(new_n629), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n687), .A2(KEYINPUT29), .A3(new_n665), .ZN(new_n688));
  XNOR2_X1  g0488(.A(new_n665), .B(KEYINPUT91), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n623), .A2(new_n615), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n690), .B1(new_n612), .B2(new_n613), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n689), .B1(new_n691), .B2(new_n629), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n688), .B1(new_n692), .B2(KEYINPUT29), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT31), .ZN(new_n694));
  AND2_X1   g0494(.A1(new_n481), .A2(new_n572), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT30), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n695), .A2(new_n524), .A3(new_n696), .A4(new_n557), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n557), .A2(new_n481), .A3(new_n572), .ZN(new_n698));
  OAI21_X1  g0498(.A(KEYINPUT30), .B1(new_n698), .B2(new_n523), .ZN(new_n699));
  AND3_X1   g0499(.A1(new_n519), .A2(new_n486), .A3(new_n301), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n574), .A2(new_n557), .ZN(new_n701));
  AOI22_X1  g0501(.A1(new_n697), .A2(new_n699), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  NOR3_X1   g0502(.A1(new_n670), .A2(new_n694), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n697), .A2(new_n699), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n700), .A2(new_n701), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  AOI21_X1  g0506(.A(KEYINPUT31), .B1(new_n706), .B2(new_n655), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(KEYINPUT93), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n694), .B1(new_n702), .B2(new_n665), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT93), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n703), .B1(new_n708), .B2(new_n711), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n605), .A2(new_n490), .A3(new_n531), .A4(new_n670), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n659), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n693), .A2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n679), .B1(new_n717), .B2(G1), .ZN(G364));
  NOR2_X1   g0518(.A1(new_n366), .A2(new_n213), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n208), .B1(new_n719), .B2(G45), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n673), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n661), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n723), .B1(new_n660), .B2(new_n658), .ZN(new_n724));
  INV_X1    g0524(.A(new_n722), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n216), .A2(new_n269), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n224), .A2(new_n476), .ZN(new_n727));
  OAI211_X1 g0527(.A(new_n726), .B(new_n727), .C1(new_n476), .C2(new_n249), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n216), .A2(new_n264), .ZN(new_n729));
  AOI22_X1  g0529(.A1(new_n729), .A2(G355), .B1(new_n474), .B2(new_n216), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n360), .A2(KEYINPUT95), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n209), .B1(KEYINPUT95), .B2(new_n360), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n221), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(G13), .A2(G33), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(G20), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n735), .A2(new_n738), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n725), .B1(new_n731), .B2(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(KEYINPUT96), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n740), .A2(KEYINPUT96), .ZN(new_n742));
  INV_X1    g0542(.A(new_n735), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n298), .A2(G179), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n366), .A2(new_n376), .A3(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(new_n230), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n744), .A2(G20), .A3(G190), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(G87), .ZN(new_n749));
  NOR3_X1   g0549(.A1(new_n376), .A2(G179), .A3(G200), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n220), .A2(new_n750), .ZN(new_n751));
  OAI211_X1 g0551(.A(new_n749), .B(new_n269), .C1(new_n234), .C2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n220), .A2(new_n301), .ZN(new_n753));
  NOR2_X1   g0553(.A1(G190), .A2(G200), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  AOI211_X1 g0556(.A(new_n746), .B(new_n752), .C1(G77), .C2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n376), .A2(G200), .ZN(new_n758));
  AND3_X1   g0558(.A1(new_n753), .A2(KEYINPUT97), .A3(new_n758), .ZN(new_n759));
  AOI21_X1  g0559(.A(KEYINPUT97), .B1(new_n753), .B2(new_n758), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(G58), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n753), .A2(G200), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(new_n376), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n764), .A2(G190), .ZN(new_n766));
  AOI22_X1  g0566(.A1(G50), .A2(new_n765), .B1(new_n766), .B2(G68), .ZN(new_n767));
  NOR4_X1   g0567(.A1(new_n220), .A2(G179), .A3(G190), .A4(G200), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(G159), .ZN(new_n769));
  XOR2_X1   g0569(.A(new_n769), .B(KEYINPUT32), .Z(new_n770));
  NAND4_X1  g0570(.A1(new_n757), .A2(new_n763), .A3(new_n767), .A4(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n762), .A2(G322), .ZN(new_n772));
  INV_X1    g0572(.A(G294), .ZN(new_n773));
  OAI221_X1 g0573(.A(new_n264), .B1(new_n507), .B2(new_n747), .C1(new_n751), .C2(new_n773), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n774), .B1(G329), .B2(new_n768), .ZN(new_n775));
  INV_X1    g0575(.A(new_n745), .ZN(new_n776));
  AOI22_X1  g0576(.A1(new_n756), .A2(G311), .B1(G283), .B2(new_n776), .ZN(new_n777));
  XNOR2_X1  g0577(.A(KEYINPUT33), .B(G317), .ZN(new_n778));
  AOI22_X1  g0578(.A1(G326), .A2(new_n765), .B1(new_n766), .B2(new_n778), .ZN(new_n779));
  NAND4_X1  g0579(.A1(new_n772), .A2(new_n775), .A3(new_n777), .A4(new_n779), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n743), .B1(new_n771), .B2(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n742), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n738), .ZN(new_n783));
  OAI211_X1 g0583(.A(new_n741), .B(new_n782), .C1(new_n658), .C2(new_n783), .ZN(new_n784));
  AND2_X1   g0584(.A1(new_n724), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(G396));
  NAND2_X1  g0586(.A1(new_n655), .A2(new_n373), .ZN(new_n787));
  OAI211_X1 g0587(.A(new_n372), .B(new_n787), .C1(new_n377), .C2(new_n378), .ZN(new_n788));
  OR2_X1    g0588(.A1(new_n372), .A2(new_n787), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n692), .B(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n722), .B1(new_n791), .B2(new_n715), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n792), .B1(new_n715), .B2(new_n791), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n735), .A2(new_n736), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n722), .B1(G77), .B2(new_n795), .ZN(new_n796));
  AOI22_X1  g0596(.A1(new_n765), .A2(G137), .B1(new_n756), .B2(G159), .ZN(new_n797));
  INV_X1    g0597(.A(G150), .ZN(new_n798));
  INV_X1    g0598(.A(new_n766), .ZN(new_n799));
  XNOR2_X1  g0599(.A(KEYINPUT98), .B(G143), .ZN(new_n800));
  OAI221_X1 g0600(.A(new_n797), .B1(new_n798), .B2(new_n799), .C1(new_n761), .C2(new_n800), .ZN(new_n801));
  XNOR2_X1  g0601(.A(new_n801), .B(KEYINPUT34), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n745), .A2(new_n312), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  OAI221_X1 g0604(.A(new_n269), .B1(new_n201), .B2(new_n747), .C1(new_n751), .C2(new_n202), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n805), .B1(G132), .B2(new_n768), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n802), .A2(new_n804), .A3(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n761), .A2(new_n773), .ZN(new_n808));
  AOI22_X1  g0608(.A1(G283), .A2(new_n766), .B1(new_n765), .B2(G303), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n264), .B1(new_n747), .B2(new_n230), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n751), .A2(new_n234), .ZN(new_n811));
  AOI211_X1 g0611(.A(new_n810), .B(new_n811), .C1(G311), .C2(new_n768), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n756), .A2(G116), .B1(G87), .B2(new_n776), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n809), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n807), .B1(new_n808), .B2(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n796), .B1(new_n815), .B2(new_n735), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n816), .B1(new_n737), .B2(new_n790), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n793), .A2(new_n817), .ZN(G384));
  NOR2_X1   g0618(.A1(new_n719), .A2(new_n208), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n655), .A2(new_n323), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n343), .A2(new_n348), .A3(new_n820), .ZN(new_n821));
  OAI21_X1  g0621(.A(G169), .B1(new_n333), .B2(new_n334), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n822), .A2(KEYINPUT14), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n823), .A2(new_n339), .A3(new_n335), .ZN(new_n824));
  OAI211_X1 g0624(.A(new_n323), .B(new_n655), .C1(new_n824), .C2(new_n347), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n821), .A2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  OAI211_X1 g0627(.A(new_n670), .B(new_n790), .C1(new_n624), .C2(new_n630), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n372), .A2(new_n655), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n827), .B1(new_n828), .B2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n439), .A2(new_n650), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT37), .ZN(new_n834));
  NAND4_X1  g0634(.A1(new_n833), .A2(new_n442), .A3(new_n834), .A4(new_n422), .ZN(new_n835));
  AND2_X1   g0635(.A1(new_n388), .A2(new_n389), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n407), .B1(new_n836), .B2(new_n390), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n837), .B1(new_n634), .B2(new_n650), .ZN(new_n838));
  AND2_X1   g0638(.A1(new_n422), .A2(new_n838), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n835), .B1(new_n834), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n837), .A2(new_n650), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n840), .B1(new_n445), .B2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT38), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  OAI211_X1 g0644(.A(KEYINPUT38), .B(new_n840), .C1(new_n445), .C2(new_n841), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n844), .A2(KEYINPUT99), .A3(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT99), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n842), .A2(new_n847), .A3(new_n843), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  OAI22_X1  g0649(.A1(new_n832), .A2(new_n849), .B1(new_n638), .B2(new_n650), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT39), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n851), .B1(new_n846), .B2(new_n848), .ZN(new_n852));
  NAND4_X1  g0652(.A1(new_n636), .A2(new_n418), .A3(new_n424), .A4(new_n637), .ZN(new_n853));
  INV_X1    g0653(.A(new_n833), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT100), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n833), .A2(new_n422), .A3(new_n635), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(KEYINPUT37), .ZN(new_n858));
  AOI22_X1  g0658(.A1(new_n855), .A2(new_n856), .B1(new_n835), .B2(new_n858), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n853), .A2(KEYINPUT100), .A3(new_n854), .ZN(new_n860));
  AOI21_X1  g0660(.A(KEYINPUT38), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(KEYINPUT39), .B1(new_n862), .B2(new_n845), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n824), .A2(new_n323), .A3(new_n665), .ZN(new_n864));
  NOR3_X1   g0664(.A1(new_n852), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n850), .A2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  OAI211_X1 g0667(.A(new_n446), .B(new_n688), .C1(new_n692), .C2(KEYINPUT29), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(new_n641), .ZN(new_n869));
  XNOR2_X1  g0669(.A(new_n869), .B(KEYINPUT101), .ZN(new_n870));
  XNOR2_X1  g0670(.A(new_n867), .B(new_n870), .ZN(new_n871));
  NOR3_X1   g0671(.A1(new_n702), .A2(new_n694), .A3(new_n665), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n707), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n713), .A2(new_n873), .ZN(new_n874));
  AOI22_X1  g0674(.A1(new_n821), .A2(new_n825), .B1(new_n788), .B2(new_n789), .ZN(new_n875));
  AND3_X1   g0675(.A1(new_n874), .A2(KEYINPUT40), .A3(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n845), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n876), .B1(new_n861), .B2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT103), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  OAI211_X1 g0680(.A(new_n876), .B(KEYINPUT103), .C1(new_n861), .C2(new_n877), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT102), .ZN(new_n882));
  AND3_X1   g0682(.A1(new_n874), .A2(new_n882), .A3(new_n875), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n882), .B1(new_n874), .B2(new_n875), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n846), .A2(new_n885), .A3(new_n848), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT40), .ZN(new_n887));
  AOI22_X1  g0687(.A1(new_n880), .A2(new_n881), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n446), .A2(new_n874), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n659), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n891), .B1(new_n890), .B2(new_n889), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n819), .B1(new_n871), .B2(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n893), .B1(new_n871), .B2(new_n892), .ZN(new_n894));
  INV_X1    g0694(.A(new_n537), .ZN(new_n895));
  OR2_X1    g0695(.A1(new_n895), .A2(KEYINPUT35), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(KEYINPUT35), .ZN(new_n897));
  NAND4_X1  g0697(.A1(new_n896), .A2(G116), .A3(new_n222), .A4(new_n897), .ZN(new_n898));
  XNOR2_X1  g0698(.A(new_n898), .B(KEYINPUT36), .ZN(new_n899));
  OAI21_X1  g0699(.A(G77), .B1(new_n202), .B2(new_n312), .ZN(new_n900));
  OAI22_X1  g0700(.A1(new_n900), .A2(new_n223), .B1(G50), .B2(new_n312), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n901), .A2(G1), .A3(new_n213), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n894), .A2(new_n899), .A3(new_n902), .ZN(G367));
  NAND2_X1  g0703(.A1(new_n689), .A2(new_n622), .ZN(new_n904));
  INV_X1    g0704(.A(new_n568), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n905), .B1(new_n670), .B2(new_n543), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n908), .A2(new_n594), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n670), .B1(new_n909), .B2(new_n611), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n907), .A2(new_n662), .A3(new_n668), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(KEYINPUT42), .ZN(new_n912));
  OR2_X1    g0712(.A1(new_n911), .A2(KEYINPUT42), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n910), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n485), .A2(new_n665), .ZN(new_n915));
  INV_X1    g0715(.A(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n621), .A2(new_n916), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n917), .B1(new_n609), .B2(new_n916), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(KEYINPUT43), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n919), .B(KEYINPUT104), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n914), .A2(new_n920), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n918), .A2(KEYINPUT43), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n921), .A2(new_n922), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n667), .A2(new_n908), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n926), .B(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n671), .A2(new_n907), .ZN(new_n929));
  XOR2_X1   g0729(.A(new_n929), .B(KEYINPUT45), .Z(new_n930));
  NOR2_X1   g0730(.A1(new_n671), .A2(new_n907), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n931), .B(KEYINPUT44), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(new_n667), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n930), .A2(new_n667), .A3(new_n932), .ZN(new_n936));
  AND2_X1   g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n668), .A2(new_n662), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT105), .ZN(new_n939));
  OAI221_X1 g0739(.A(new_n938), .B1(new_n666), .B2(new_n668), .C1(new_n661), .C2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n661), .A2(new_n939), .ZN(new_n941));
  XOR2_X1   g0741(.A(new_n940), .B(new_n941), .Z(new_n942));
  AOI21_X1  g0742(.A(new_n716), .B1(new_n937), .B2(new_n942), .ZN(new_n943));
  XOR2_X1   g0743(.A(new_n673), .B(KEYINPUT41), .Z(new_n944));
  OAI21_X1  g0744(.A(new_n720), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n928), .A2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(new_n726), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n947), .A2(new_n245), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n739), .B1(new_n215), .B2(new_n368), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n722), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n776), .A2(G97), .ZN(new_n951));
  INV_X1    g0751(.A(G283), .ZN(new_n952));
  INV_X1    g0752(.A(new_n768), .ZN(new_n953));
  INV_X1    g0753(.A(G317), .ZN(new_n954));
  OAI221_X1 g0754(.A(new_n951), .B1(new_n952), .B2(new_n755), .C1(new_n953), .C2(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n748), .A2(G116), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n956), .B(KEYINPUT46), .ZN(new_n957));
  OAI211_X1 g0757(.A(new_n957), .B(new_n264), .C1(new_n230), .C2(new_n751), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n958), .B1(G311), .B2(new_n765), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n959), .B1(new_n773), .B2(new_n799), .ZN(new_n960));
  AOI211_X1 g0760(.A(new_n955), .B(new_n960), .C1(G303), .C2(new_n762), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n762), .A2(G150), .ZN(new_n962));
  INV_X1    g0762(.A(G159), .ZN(new_n963));
  INV_X1    g0763(.A(new_n765), .ZN(new_n964));
  OAI22_X1  g0764(.A1(new_n963), .A2(new_n799), .B1(new_n964), .B2(new_n800), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n776), .A2(G77), .ZN(new_n966));
  INV_X1    g0766(.A(new_n751), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(G68), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n264), .B1(new_n748), .B2(G58), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n966), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(G137), .ZN(new_n971));
  OAI22_X1  g0771(.A1(new_n953), .A2(new_n971), .B1(new_n201), .B2(new_n755), .ZN(new_n972));
  NOR3_X1   g0772(.A1(new_n965), .A2(new_n970), .A3(new_n972), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n961), .B1(new_n962), .B2(new_n973), .ZN(new_n974));
  XOR2_X1   g0774(.A(new_n974), .B(KEYINPUT47), .Z(new_n975));
  AOI21_X1  g0775(.A(new_n950), .B1(new_n975), .B2(new_n735), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n976), .B1(new_n783), .B2(new_n918), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n946), .A2(new_n977), .ZN(G387));
  AOI22_X1  g0778(.A1(new_n729), .A2(new_n675), .B1(new_n230), .B2(new_n216), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n242), .A2(new_n476), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n362), .A2(new_n201), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n981), .B(KEYINPUT50), .ZN(new_n982));
  OAI211_X1 g0782(.A(new_n674), .B(new_n476), .C1(new_n312), .C2(new_n228), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n726), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n979), .B1(new_n980), .B2(new_n984), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n985), .A2(KEYINPUT106), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(KEYINPUT106), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n987), .A2(new_n739), .ZN(new_n988));
  OAI221_X1 g0788(.A(new_n722), .B1(new_n986), .B2(new_n988), .C1(new_n666), .C2(new_n783), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n967), .A2(new_n462), .ZN(new_n990));
  OAI221_X1 g0790(.A(new_n990), .B1(new_n312), .B2(new_n755), .C1(new_n964), .C2(new_n963), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n991), .B1(new_n362), .B2(new_n766), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n264), .B1(new_n748), .B2(G77), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n951), .B(new_n993), .C1(new_n953), .C2(new_n798), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n994), .B(KEYINPUT107), .Z(new_n995));
  OAI211_X1 g0795(.A(new_n992), .B(new_n995), .C1(new_n201), .C2(new_n761), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n269), .B1(new_n768), .B2(G326), .ZN(new_n997));
  OAI22_X1  g0797(.A1(new_n751), .A2(new_n952), .B1(new_n773), .B2(new_n747), .ZN(new_n998));
  AOI22_X1  g0798(.A1(new_n766), .A2(G311), .B1(new_n756), .B2(G303), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n765), .A2(G322), .ZN(new_n1000));
  OAI211_X1 g0800(.A(new_n999), .B(new_n1000), .C1(new_n954), .C2(new_n761), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT48), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n998), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n1003), .B1(new_n1002), .B2(new_n1001), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT49), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n997), .B1(new_n474), .B2(new_n745), .C1(new_n1004), .C2(new_n1005), .ZN(new_n1006));
  AND2_X1   g0806(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n996), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n989), .B1(new_n735), .B2(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(KEYINPUT108), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1010), .B1(new_n942), .B2(new_n721), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n942), .A2(new_n717), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1012), .A2(new_n673), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n942), .A2(new_n717), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1011), .B1(new_n1013), .B2(new_n1014), .ZN(G393));
  NAND3_X1  g0815(.A1(new_n937), .A2(new_n717), .A3(new_n942), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n935), .A2(new_n936), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1012), .A2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1016), .A2(new_n673), .A3(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n937), .A2(new_n721), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT111), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n947), .A2(new_n252), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n739), .B1(new_n215), .B2(new_n234), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n722), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n953), .A2(new_n800), .B1(new_n282), .B2(new_n755), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n967), .A2(G77), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n264), .B1(new_n748), .B2(G68), .ZN(new_n1027));
  OAI211_X1 g0827(.A(new_n1026), .B(new_n1027), .C1(new_n449), .C2(new_n745), .ZN(new_n1028));
  AOI211_X1 g0828(.A(new_n1025), .B(new_n1028), .C1(G50), .C2(new_n766), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(new_n762), .A2(G159), .B1(G150), .B2(new_n765), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT51), .ZN(new_n1031));
  AND2_X1   g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1029), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT109), .ZN(new_n1035));
  OR2_X1    g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n762), .A2(G311), .B1(G317), .B2(new_n765), .ZN(new_n1037));
  XOR2_X1   g0837(.A(new_n1037), .B(KEYINPUT52), .Z(new_n1038));
  OAI21_X1  g0838(.A(new_n264), .B1(new_n747), .B2(new_n952), .ZN(new_n1039));
  AOI211_X1 g0839(.A(new_n1039), .B(new_n746), .C1(G322), .C2(new_n768), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT110), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n766), .A2(G303), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n756), .A2(G294), .B1(G116), .B2(new_n967), .ZN(new_n1043));
  NAND4_X1  g0843(.A1(new_n1038), .A2(new_n1041), .A3(new_n1042), .A4(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1036), .A2(new_n1044), .A3(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1024), .B1(new_n1046), .B2(new_n735), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(new_n907), .B2(new_n783), .ZN(new_n1048));
  AND3_X1   g0848(.A1(new_n1020), .A2(new_n1021), .A3(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1021), .B1(new_n1020), .B2(new_n1048), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1019), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(KEYINPUT112), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  OAI211_X1 g0853(.A(KEYINPUT112), .B(new_n1019), .C1(new_n1049), .C2(new_n1050), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1053), .A2(new_n1054), .ZN(G390));
  AND3_X1   g0855(.A1(new_n714), .A2(new_n790), .A3(new_n826), .ZN(new_n1056));
  AND2_X1   g0856(.A1(new_n874), .A2(G330), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n826), .B1(new_n1057), .B2(new_n790), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n790), .ZN(new_n1060));
  AOI211_X1 g0860(.A(new_n655), .B(new_n1060), .C1(new_n686), .C2(new_n629), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n1061), .A2(new_n829), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n828), .A2(new_n830), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1057), .A2(new_n875), .ZN(new_n1064));
  AOI211_X1 g0864(.A(new_n659), .B(new_n1060), .C1(new_n712), .C2(new_n713), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1064), .B1(new_n1065), .B2(new_n826), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n1059), .A2(new_n1062), .B1(new_n1063), .B2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n446), .A2(new_n1057), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n868), .A2(new_n641), .A3(new_n1068), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n1070), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n826), .B1(new_n1061), .B2(new_n829), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n862), .A2(new_n845), .ZN(new_n1073));
  XOR2_X1   g0873(.A(new_n864), .B(KEYINPUT113), .Z(new_n1074));
  AND3_X1   g0874(.A1(new_n1072), .A2(new_n1073), .A3(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n849), .A2(KEYINPUT39), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n863), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n864), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n831), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1075), .B1(new_n1078), .B2(new_n1081), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n1082), .A2(new_n1064), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1072), .A2(new_n1073), .A3(new_n1074), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1056), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n852), .A2(new_n863), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n1084), .B(new_n1085), .C1(new_n1086), .C2(new_n1080), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1087), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1071), .B1(new_n1083), .B2(new_n1088), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n1087), .B(new_n1070), .C1(new_n1082), .C2(new_n1064), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1089), .A2(new_n673), .A3(new_n1090), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n722), .B1(new_n362), .B2(new_n795), .ZN(new_n1092));
  XOR2_X1   g0892(.A(new_n1092), .B(KEYINPUT114), .Z(new_n1093));
  NOR2_X1   g0893(.A1(new_n799), .A2(new_n971), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n747), .A2(new_n798), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(new_n1095), .B(KEYINPUT53), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n1096), .B(new_n269), .C1(new_n963), .C2(new_n751), .ZN(new_n1097));
  AOI211_X1 g0897(.A(new_n1094), .B(new_n1097), .C1(G128), .C2(new_n765), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(G125), .A2(new_n768), .B1(new_n776), .B2(G50), .ZN(new_n1099));
  XOR2_X1   g0899(.A(KEYINPUT54), .B(G143), .Z(new_n1100));
  NAND2_X1  g0900(.A1(new_n756), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1102), .B1(G132), .B2(new_n762), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n762), .A2(G116), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n230), .A2(new_n799), .B1(new_n964), .B2(new_n952), .ZN(new_n1105));
  NAND4_X1  g0905(.A1(new_n804), .A2(new_n264), .A3(new_n1026), .A4(new_n749), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n953), .A2(new_n773), .B1(new_n234), .B2(new_n755), .ZN(new_n1107));
  NOR3_X1   g0907(.A1(new_n1105), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n1098), .A2(new_n1103), .B1(new_n1104), .B2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1093), .B1(new_n1109), .B2(new_n743), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1110), .B1(new_n1078), .B2(new_n736), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n1083), .A2(new_n1088), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1111), .B1(new_n1112), .B2(new_n721), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1091), .A2(new_n1113), .ZN(G378));
  INV_X1    g0914(.A(new_n1069), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1090), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n880), .A2(new_n881), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n886), .A2(new_n887), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1117), .A2(new_n1118), .A3(G330), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n650), .A2(new_n303), .ZN(new_n1120));
  XNOR2_X1  g0920(.A(new_n305), .B(new_n1120), .ZN(new_n1121));
  XNOR2_X1  g0921(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(new_n1121), .B(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1119), .A2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n888), .A2(G330), .A3(new_n1123), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(KEYINPUT118), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1128), .B1(new_n850), .B2(new_n865), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n849), .ZN(new_n1130));
  AOI22_X1  g0930(.A1(new_n1130), .A2(new_n831), .B1(new_n639), .B2(new_n649), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1076), .A2(new_n1077), .A3(new_n1079), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1131), .A2(new_n1132), .A3(KEYINPUT118), .ZN(new_n1133));
  NAND4_X1  g0933(.A1(new_n1127), .A2(KEYINPUT119), .A3(new_n1129), .A4(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1123), .B1(new_n888), .B2(G330), .ZN(new_n1135));
  AND4_X1   g0935(.A1(G330), .A2(new_n1117), .A3(new_n1118), .A4(new_n1123), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1129), .A2(new_n1133), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1125), .A2(new_n1126), .A3(new_n866), .ZN(new_n1140));
  INV_X1    g0940(.A(KEYINPUT119), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n1116), .B(new_n1134), .C1(new_n1139), .C2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(KEYINPUT57), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n673), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1144), .B1(new_n1090), .B2(new_n1115), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1127), .A2(new_n867), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1148), .A2(new_n1140), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1146), .B1(new_n1147), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1145), .A2(new_n1150), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n721), .B(new_n1134), .C1(new_n1139), .C2(new_n1142), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n722), .B1(G50), .B2(new_n795), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(G33), .A2(G41), .ZN(new_n1154));
  INV_X1    g0954(.A(G41), .ZN(new_n1155));
  AOI211_X1 g0955(.A(G50), .B(new_n1154), .C1(new_n264), .C2(new_n1155), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n745), .A2(new_n202), .ZN(new_n1157));
  AOI211_X1 g0957(.A(G41), .B(new_n269), .C1(new_n748), .C2(G77), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n1158), .B(new_n968), .C1(new_n368), .C2(new_n755), .ZN(new_n1159));
  AOI211_X1 g0959(.A(new_n1157), .B(new_n1159), .C1(G283), .C2(new_n768), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(G97), .A2(new_n766), .B1(new_n765), .B2(G116), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n1160), .B(new_n1161), .C1(new_n230), .C2(new_n761), .ZN(new_n1162));
  INV_X1    g0962(.A(KEYINPUT58), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1156), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(new_n765), .A2(G125), .B1(G150), .B2(new_n967), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(new_n1165), .B(KEYINPUT115), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n762), .A2(G128), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n766), .A2(G132), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n756), .A2(G137), .B1(new_n748), .B2(new_n1100), .ZN(new_n1169));
  NAND4_X1  g0969(.A1(new_n1166), .A2(new_n1167), .A3(new_n1168), .A4(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1170), .A2(KEYINPUT59), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1154), .ZN(new_n1172));
  XOR2_X1   g0972(.A(KEYINPUT116), .B(G124), .Z(new_n1173));
  AOI21_X1  g0973(.A(new_n1172), .B1(new_n768), .B2(new_n1173), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n1171), .B(new_n1174), .C1(new_n963), .C2(new_n745), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n1170), .A2(KEYINPUT59), .ZN(new_n1176));
  OAI221_X1 g0976(.A(new_n1164), .B1(new_n1163), .B2(new_n1162), .C1(new_n1175), .C2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1153), .B1(new_n1177), .B2(new_n735), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1178), .B1(new_n1123), .B2(new_n737), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(new_n1179), .B(KEYINPUT117), .ZN(new_n1180));
  AND2_X1   g0980(.A1(new_n1152), .A2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1151), .A2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1182), .A2(KEYINPUT120), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT120), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1151), .A2(new_n1184), .A3(new_n1181), .ZN(new_n1185));
  AND2_X1   g0985(.A1(new_n1183), .A2(new_n1185), .ZN(G375));
  NAND2_X1  g0986(.A1(new_n1059), .A2(new_n1062), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1066), .A2(new_n1063), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n827), .A2(new_n736), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n722), .B1(G68), .B2(new_n795), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n269), .B1(new_n747), .B2(new_n963), .ZN(new_n1192));
  AOI211_X1 g0992(.A(new_n1192), .B(new_n1157), .C1(G128), .C2(new_n768), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(G132), .A2(new_n765), .B1(new_n766), .B2(new_n1100), .ZN(new_n1194));
  OAI211_X1 g0994(.A(new_n1193), .B(new_n1194), .C1(new_n971), .C2(new_n761), .ZN(new_n1195));
  OAI22_X1  g0995(.A1(new_n755), .A2(new_n798), .B1(new_n201), .B2(new_n751), .ZN(new_n1196));
  XOR2_X1   g0996(.A(new_n1196), .B(KEYINPUT121), .Z(new_n1197));
  AOI22_X1  g0997(.A1(G116), .A2(new_n766), .B1(new_n765), .B2(G294), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n269), .B1(new_n748), .B2(G97), .ZN(new_n1199));
  AND3_X1   g0999(.A1(new_n966), .A2(new_n990), .A3(new_n1199), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n756), .A2(G107), .B1(G303), .B2(new_n768), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1198), .A2(new_n1200), .A3(new_n1201), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n761), .A2(new_n952), .ZN(new_n1203));
  OAI22_X1  g1003(.A1(new_n1195), .A2(new_n1197), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1191), .B1(new_n1204), .B2(new_n735), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(new_n1189), .A2(new_n721), .B1(new_n1190), .B2(new_n1205), .ZN(new_n1206));
  OR2_X1    g1006(.A1(new_n1070), .A2(new_n944), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n1189), .A2(new_n1115), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1206), .B1(new_n1207), .B2(new_n1208), .ZN(G381));
  OR2_X1    g1009(.A1(G393), .A2(G396), .ZN(new_n1210));
  OR4_X1    g1010(.A1(G384), .A2(G387), .A3(new_n1210), .A4(G381), .ZN(new_n1211));
  OR4_X1    g1011(.A1(G390), .A2(G375), .A3(G378), .A4(new_n1211), .ZN(G407));
  AOI21_X1  g1012(.A(G378), .B1(new_n1183), .B2(new_n1185), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n647), .A2(G343), .ZN(new_n1214));
  XOR2_X1   g1014(.A(new_n1214), .B(KEYINPUT122), .Z(new_n1215));
  NAND2_X1  g1015(.A1(new_n1213), .A2(new_n1215), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(G407), .A2(G213), .A3(new_n1216), .ZN(G409));
  INV_X1    g1017(.A(KEYINPUT127), .ZN(new_n1218));
  XNOR2_X1  g1018(.A(G393), .B(new_n785), .ZN(new_n1219));
  AOI21_X1  g1019(.A(G387), .B1(new_n1054), .B2(new_n1053), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1219), .B1(new_n1220), .B2(KEYINPUT125), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(G390), .A2(new_n946), .A3(new_n977), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(G387), .A2(new_n1053), .A3(new_n1054), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1221), .A2(new_n1224), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n1222), .A2(KEYINPUT125), .A3(new_n1223), .A4(new_n1219), .ZN(new_n1226));
  AND2_X1   g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1151), .A2(G378), .A3(new_n1181), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1149), .A2(new_n721), .ZN(new_n1229));
  OAI211_X1 g1029(.A(new_n1179), .B(new_n1229), .C1(new_n1143), .C2(new_n944), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1230), .A2(new_n1091), .A3(new_n1113), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1228), .A2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1214), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT123), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n673), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT60), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1236), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1237), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1067), .A2(new_n1236), .A3(new_n1069), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1235), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(G384), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1206), .ZN(new_n1242));
  NOR3_X1   g1042(.A1(new_n1240), .A2(new_n1241), .A3(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1239), .ZN(new_n1244));
  OAI211_X1 g1044(.A(new_n1071), .B(new_n673), .C1(new_n1244), .C2(new_n1237), .ZN(new_n1245));
  AOI21_X1  g1045(.A(G384), .B1(new_n1245), .B2(new_n1206), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1234), .B1(new_n1243), .B2(new_n1246), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1241), .B1(new_n1240), .B2(new_n1242), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1245), .A2(G384), .A3(new_n1206), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1248), .A2(new_n1249), .A3(KEYINPUT123), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1247), .A2(new_n1250), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1232), .A2(new_n1233), .A3(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT62), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1215), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1253), .B1(new_n1247), .B2(new_n1250), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1232), .A2(new_n1255), .A3(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT126), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1215), .B1(new_n1228), .B2(new_n1231), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1260), .A2(KEYINPUT126), .A3(new_n1256), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1254), .A2(new_n1259), .A3(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT61), .ZN(new_n1263));
  INV_X1    g1063(.A(G2897), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1233), .A2(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1265), .B1(new_n1247), .B2(new_n1250), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1267), .A2(G2897), .A3(new_n1215), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  OAI21_X1  g1069(.A(KEYINPUT124), .B1(new_n1266), .B2(new_n1269), .ZN(new_n1270));
  AND3_X1   g1070(.A1(new_n1248), .A2(KEYINPUT123), .A3(new_n1249), .ZN(new_n1271));
  AOI21_X1  g1071(.A(KEYINPUT123), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1272));
  OAI22_X1  g1072(.A1(new_n1271), .A2(new_n1272), .B1(new_n1264), .B2(new_n1233), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT124), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1273), .A2(new_n1274), .A3(new_n1268), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1270), .A2(new_n1275), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1263), .B1(new_n1276), .B2(new_n1260), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1227), .B1(new_n1262), .B2(new_n1278), .ZN(new_n1279));
  AND3_X1   g1079(.A1(new_n1225), .A2(new_n1263), .A3(new_n1226), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1281), .A2(new_n1275), .A3(new_n1270), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT63), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1252), .A2(new_n1283), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1260), .A2(KEYINPUT63), .A3(new_n1251), .ZN(new_n1285));
  NAND4_X1  g1085(.A1(new_n1280), .A2(new_n1282), .A3(new_n1284), .A4(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1286), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1218), .B1(new_n1279), .B2(new_n1287), .ZN(new_n1288));
  AOI22_X1  g1088(.A1(new_n1258), .A2(new_n1257), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1277), .B1(new_n1289), .B2(new_n1261), .ZN(new_n1290));
  OAI211_X1 g1090(.A(KEYINPUT127), .B(new_n1286), .C1(new_n1290), .C2(new_n1227), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1288), .A2(new_n1291), .ZN(G405));
  AND2_X1   g1092(.A1(new_n1182), .A2(G378), .ZN(new_n1293));
  NOR2_X1   g1093(.A1(new_n1213), .A2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1294), .A2(new_n1251), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1267), .B1(new_n1213), .B2(new_n1293), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  XOR2_X1   g1097(.A(new_n1297), .B(new_n1227), .Z(G402));
endmodule


