

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U549 ( .A1(n785), .A2(n691), .ZN(n694) );
  NOR2_X2 U550 ( .A1(G164), .A2(G1384), .ZN(n785) );
  INV_X1 U551 ( .A(KEYINPUT17), .ZN(n518) );
  NOR2_X1 U552 ( .A1(G651), .A2(G543), .ZN(n656) );
  INV_X1 U553 ( .A(n694), .ZN(n713) );
  NOR2_X1 U554 ( .A1(n694), .A2(n919), .ZN(n696) );
  NOR2_X1 U555 ( .A1(G2104), .A2(G2105), .ZN(n519) );
  INV_X1 U556 ( .A(KEYINPUT66), .ZN(n521) );
  NAND2_X1 U557 ( .A1(n873), .A2(G138), .ZN(n534) );
  XNOR2_X1 U558 ( .A(n523), .B(n522), .ZN(n525) );
  NOR2_X2 U559 ( .A1(G2104), .A2(n526), .ZN(n531) );
  AND2_X1 U560 ( .A1(n829), .A2(n956), .ZN(n515) );
  XNOR2_X1 U561 ( .A(KEYINPUT65), .B(n527), .ZN(n516) );
  OR2_X1 U562 ( .A1(n777), .A2(n776), .ZN(n517) );
  INV_X1 U563 ( .A(KEYINPUT26), .ZN(n695) );
  XNOR2_X1 U564 ( .A(KEYINPUT96), .B(KEYINPUT30), .ZN(n728) );
  XNOR2_X1 U565 ( .A(n729), .B(n728), .ZN(n730) );
  INV_X1 U566 ( .A(KEYINPUT29), .ZN(n723) );
  AND2_X1 U567 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U568 ( .A1(n594), .A2(G68), .ZN(n595) );
  NAND2_X1 U569 ( .A1(n517), .A2(n939), .ZN(n778) );
  INV_X1 U570 ( .A(KEYINPUT100), .ZN(n780) );
  NOR2_X1 U571 ( .A1(n821), .A2(n515), .ZN(n805) );
  INV_X1 U572 ( .A(KEYINPUT68), .ZN(n540) );
  AND2_X1 U573 ( .A1(n806), .A2(n805), .ZN(n817) );
  INV_X1 U574 ( .A(KEYINPUT75), .ZN(n606) );
  XNOR2_X1 U575 ( .A(n541), .B(n540), .ZN(n594) );
  XNOR2_X1 U576 ( .A(n521), .B(KEYINPUT23), .ZN(n522) );
  NOR2_X1 U577 ( .A1(G543), .A2(n545), .ZN(n546) );
  AND2_X1 U578 ( .A1(n526), .A2(G2104), .ZN(n874) );
  NOR2_X1 U579 ( .A1(G651), .A2(n542), .ZN(n663) );
  NOR2_X1 U580 ( .A1(n528), .A2(n516), .ZN(n529) );
  AND2_X1 U581 ( .A1(n530), .A2(n529), .ZN(G160) );
  XNOR2_X2 U582 ( .A(n519), .B(n518), .ZN(n873) );
  NAND2_X1 U583 ( .A1(G137), .A2(n873), .ZN(n520) );
  XOR2_X1 U584 ( .A(KEYINPUT67), .B(n520), .Z(n530) );
  INV_X1 U585 ( .A(G2105), .ZN(n526) );
  NAND2_X1 U586 ( .A1(G101), .A2(n874), .ZN(n523) );
  AND2_X1 U587 ( .A1(G2104), .A2(G2105), .ZN(n869) );
  NAND2_X1 U588 ( .A1(G113), .A2(n869), .ZN(n524) );
  NAND2_X1 U589 ( .A1(n525), .A2(n524), .ZN(n528) );
  NAND2_X1 U590 ( .A1(G125), .A2(n531), .ZN(n527) );
  NAND2_X1 U591 ( .A1(G114), .A2(n869), .ZN(n533) );
  NAND2_X1 U592 ( .A1(G126), .A2(n531), .ZN(n532) );
  AND2_X1 U593 ( .A1(n533), .A2(n532), .ZN(n539) );
  XNOR2_X1 U594 ( .A(n534), .B(KEYINPUT86), .ZN(n536) );
  NAND2_X1 U595 ( .A1(G102), .A2(n874), .ZN(n535) );
  NAND2_X1 U596 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U597 ( .A(n537), .B(KEYINPUT87), .ZN(n538) );
  AND2_X1 U598 ( .A1(n539), .A2(n538), .ZN(G164) );
  XOR2_X1 U599 ( .A(G543), .B(KEYINPUT0), .Z(n542) );
  INV_X1 U600 ( .A(G651), .ZN(n545) );
  OR2_X1 U601 ( .A1(n542), .A2(n545), .ZN(n541) );
  BUF_X1 U602 ( .A(n594), .Z(n659) );
  NAND2_X1 U603 ( .A1(G75), .A2(n659), .ZN(n551) );
  NAND2_X1 U604 ( .A1(G50), .A2(n663), .ZN(n544) );
  NAND2_X1 U605 ( .A1(G88), .A2(n656), .ZN(n543) );
  NAND2_X1 U606 ( .A1(n544), .A2(n543), .ZN(n549) );
  XOR2_X2 U607 ( .A(KEYINPUT1), .B(n546), .Z(n655) );
  NAND2_X1 U608 ( .A1(G62), .A2(n655), .ZN(n547) );
  XNOR2_X1 U609 ( .A(KEYINPUT81), .B(n547), .ZN(n548) );
  NOR2_X1 U610 ( .A1(n549), .A2(n548), .ZN(n550) );
  NAND2_X1 U611 ( .A1(n551), .A2(n550), .ZN(n552) );
  XOR2_X1 U612 ( .A(KEYINPUT82), .B(n552), .Z(G166) );
  INV_X1 U613 ( .A(G166), .ZN(G303) );
  XOR2_X1 U614 ( .A(G2427), .B(G2435), .Z(n554) );
  XNOR2_X1 U615 ( .A(G2454), .B(G2443), .ZN(n553) );
  XNOR2_X1 U616 ( .A(n554), .B(n553), .ZN(n561) );
  XOR2_X1 U617 ( .A(G2451), .B(KEYINPUT103), .Z(n556) );
  XNOR2_X1 U618 ( .A(G2430), .B(G2438), .ZN(n555) );
  XNOR2_X1 U619 ( .A(n556), .B(n555), .ZN(n557) );
  XOR2_X1 U620 ( .A(n557), .B(G2446), .Z(n559) );
  XNOR2_X1 U621 ( .A(G1348), .B(G1341), .ZN(n558) );
  XNOR2_X1 U622 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U623 ( .A(n561), .B(n560), .ZN(n562) );
  AND2_X1 U624 ( .A1(n562), .A2(G14), .ZN(G401) );
  NAND2_X1 U625 ( .A1(G64), .A2(n655), .ZN(n564) );
  NAND2_X1 U626 ( .A1(G52), .A2(n663), .ZN(n563) );
  NAND2_X1 U627 ( .A1(n564), .A2(n563), .ZN(n571) );
  NAND2_X1 U628 ( .A1(G77), .A2(n659), .ZN(n565) );
  XNOR2_X1 U629 ( .A(n565), .B(KEYINPUT70), .ZN(n567) );
  NAND2_X1 U630 ( .A1(G90), .A2(n656), .ZN(n566) );
  NAND2_X1 U631 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U632 ( .A(KEYINPUT9), .B(n568), .ZN(n569) );
  XNOR2_X1 U633 ( .A(KEYINPUT71), .B(n569), .ZN(n570) );
  NOR2_X1 U634 ( .A1(n571), .A2(n570), .ZN(G171) );
  AND2_X1 U635 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U636 ( .A1(G135), .A2(n873), .ZN(n573) );
  NAND2_X1 U637 ( .A1(G111), .A2(n869), .ZN(n572) );
  NAND2_X1 U638 ( .A1(n573), .A2(n572), .ZN(n576) );
  NAND2_X1 U639 ( .A1(n531), .A2(G123), .ZN(n574) );
  XOR2_X1 U640 ( .A(KEYINPUT18), .B(n574), .Z(n575) );
  NOR2_X1 U641 ( .A1(n576), .A2(n575), .ZN(n578) );
  NAND2_X1 U642 ( .A1(n874), .A2(G99), .ZN(n577) );
  NAND2_X1 U643 ( .A1(n578), .A2(n577), .ZN(n1000) );
  XNOR2_X1 U644 ( .A(G2096), .B(n1000), .ZN(n579) );
  OR2_X1 U645 ( .A1(G2100), .A2(n579), .ZN(G156) );
  INV_X1 U646 ( .A(G132), .ZN(G219) );
  INV_X1 U647 ( .A(G82), .ZN(G220) );
  NAND2_X1 U648 ( .A1(G63), .A2(n655), .ZN(n581) );
  NAND2_X1 U649 ( .A1(G51), .A2(n663), .ZN(n580) );
  NAND2_X1 U650 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U651 ( .A(KEYINPUT6), .B(n582), .ZN(n589) );
  NAND2_X1 U652 ( .A1(G89), .A2(n656), .ZN(n583) );
  XNOR2_X1 U653 ( .A(n583), .B(KEYINPUT78), .ZN(n584) );
  XNOR2_X1 U654 ( .A(n584), .B(KEYINPUT4), .ZN(n586) );
  NAND2_X1 U655 ( .A1(G76), .A2(n659), .ZN(n585) );
  NAND2_X1 U656 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U657 ( .A(n587), .B(KEYINPUT5), .Z(n588) );
  NOR2_X1 U658 ( .A1(n589), .A2(n588), .ZN(n590) );
  XOR2_X1 U659 ( .A(KEYINPUT7), .B(n590), .Z(n591) );
  XOR2_X1 U660 ( .A(KEYINPUT79), .B(n591), .Z(G168) );
  XOR2_X1 U661 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U662 ( .A1(G7), .A2(G661), .ZN(n592) );
  XNOR2_X1 U663 ( .A(n592), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U664 ( .A(G223), .ZN(n833) );
  NAND2_X1 U665 ( .A1(n833), .A2(G567), .ZN(n593) );
  XOR2_X1 U666 ( .A(KEYINPUT11), .B(n593), .Z(G234) );
  XNOR2_X1 U667 ( .A(n595), .B(KEYINPUT73), .ZN(n598) );
  NAND2_X1 U668 ( .A1(n656), .A2(G81), .ZN(n596) );
  XOR2_X1 U669 ( .A(KEYINPUT12), .B(n596), .Z(n597) );
  NOR2_X1 U670 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U671 ( .A(n599), .B(KEYINPUT13), .ZN(n602) );
  NAND2_X1 U672 ( .A1(n655), .A2(G56), .ZN(n600) );
  XOR2_X1 U673 ( .A(KEYINPUT14), .B(n600), .Z(n601) );
  NOR2_X1 U674 ( .A1(n602), .A2(n601), .ZN(n603) );
  XNOR2_X1 U675 ( .A(n603), .B(KEYINPUT74), .ZN(n605) );
  NAND2_X1 U676 ( .A1(G43), .A2(n663), .ZN(n604) );
  NAND2_X1 U677 ( .A1(n605), .A2(n604), .ZN(n607) );
  XNOR2_X2 U678 ( .A(n607), .B(n606), .ZN(n699) );
  INV_X1 U679 ( .A(n699), .ZN(n631) );
  NAND2_X1 U680 ( .A1(n631), .A2(G860), .ZN(G153) );
  INV_X1 U681 ( .A(G171), .ZN(G301) );
  NAND2_X1 U682 ( .A1(G79), .A2(n659), .ZN(n614) );
  NAND2_X1 U683 ( .A1(G54), .A2(n663), .ZN(n609) );
  NAND2_X1 U684 ( .A1(G92), .A2(n656), .ZN(n608) );
  NAND2_X1 U685 ( .A1(n609), .A2(n608), .ZN(n612) );
  NAND2_X1 U686 ( .A1(n655), .A2(G66), .ZN(n610) );
  XOR2_X1 U687 ( .A(KEYINPUT76), .B(n610), .Z(n611) );
  NOR2_X1 U688 ( .A1(n612), .A2(n611), .ZN(n613) );
  NAND2_X1 U689 ( .A1(n614), .A2(n613), .ZN(n615) );
  XOR2_X1 U690 ( .A(KEYINPUT15), .B(n615), .Z(n707) );
  INV_X1 U691 ( .A(n707), .ZN(n946) );
  NOR2_X1 U692 ( .A1(n946), .A2(G868), .ZN(n616) );
  XNOR2_X1 U693 ( .A(n616), .B(KEYINPUT77), .ZN(n618) );
  NAND2_X1 U694 ( .A1(G868), .A2(G301), .ZN(n617) );
  NAND2_X1 U695 ( .A1(n618), .A2(n617), .ZN(G284) );
  NAND2_X1 U696 ( .A1(G65), .A2(n655), .ZN(n620) );
  NAND2_X1 U697 ( .A1(G53), .A2(n663), .ZN(n619) );
  NAND2_X1 U698 ( .A1(n620), .A2(n619), .ZN(n624) );
  NAND2_X1 U699 ( .A1(n656), .A2(G91), .ZN(n622) );
  NAND2_X1 U700 ( .A1(G78), .A2(n659), .ZN(n621) );
  NAND2_X1 U701 ( .A1(n622), .A2(n621), .ZN(n623) );
  NOR2_X1 U702 ( .A1(n624), .A2(n623), .ZN(n950) );
  INV_X1 U703 ( .A(n950), .ZN(G299) );
  XOR2_X1 U704 ( .A(KEYINPUT80), .B(G868), .Z(n625) );
  NOR2_X1 U705 ( .A1(G286), .A2(n625), .ZN(n627) );
  NOR2_X1 U706 ( .A1(G868), .A2(G299), .ZN(n626) );
  NOR2_X1 U707 ( .A1(n627), .A2(n626), .ZN(G297) );
  INV_X1 U708 ( .A(G860), .ZN(n635) );
  NAND2_X1 U709 ( .A1(n635), .A2(G559), .ZN(n628) );
  NAND2_X1 U710 ( .A1(n628), .A2(n946), .ZN(n629) );
  XNOR2_X1 U711 ( .A(n629), .B(KEYINPUT16), .ZN(G148) );
  OR2_X1 U712 ( .A1(G559), .A2(n707), .ZN(n630) );
  NAND2_X1 U713 ( .A1(n630), .A2(G868), .ZN(n633) );
  OR2_X1 U714 ( .A1(n631), .A2(G868), .ZN(n632) );
  NAND2_X1 U715 ( .A1(n633), .A2(n632), .ZN(G282) );
  NAND2_X1 U716 ( .A1(G559), .A2(n946), .ZN(n634) );
  XOR2_X1 U717 ( .A(n699), .B(n634), .Z(n672) );
  NAND2_X1 U718 ( .A1(n635), .A2(n672), .ZN(n642) );
  NAND2_X1 U719 ( .A1(G67), .A2(n655), .ZN(n637) );
  NAND2_X1 U720 ( .A1(G55), .A2(n663), .ZN(n636) );
  NAND2_X1 U721 ( .A1(n637), .A2(n636), .ZN(n641) );
  NAND2_X1 U722 ( .A1(n656), .A2(G93), .ZN(n639) );
  NAND2_X1 U723 ( .A1(G80), .A2(n659), .ZN(n638) );
  NAND2_X1 U724 ( .A1(n639), .A2(n638), .ZN(n640) );
  NOR2_X1 U725 ( .A1(n641), .A2(n640), .ZN(n674) );
  XOR2_X1 U726 ( .A(n642), .B(n674), .Z(G145) );
  NAND2_X1 U727 ( .A1(G49), .A2(n663), .ZN(n644) );
  NAND2_X1 U728 ( .A1(G74), .A2(G651), .ZN(n643) );
  NAND2_X1 U729 ( .A1(n644), .A2(n643), .ZN(n645) );
  NOR2_X1 U730 ( .A1(n655), .A2(n645), .ZN(n647) );
  NAND2_X1 U731 ( .A1(n542), .A2(G87), .ZN(n646) );
  NAND2_X1 U732 ( .A1(n647), .A2(n646), .ZN(G288) );
  NAND2_X1 U733 ( .A1(G60), .A2(n655), .ZN(n649) );
  NAND2_X1 U734 ( .A1(G47), .A2(n663), .ZN(n648) );
  NAND2_X1 U735 ( .A1(n649), .A2(n648), .ZN(n650) );
  XNOR2_X1 U736 ( .A(KEYINPUT69), .B(n650), .ZN(n654) );
  NAND2_X1 U737 ( .A1(n659), .A2(G72), .ZN(n652) );
  NAND2_X1 U738 ( .A1(n656), .A2(G85), .ZN(n651) );
  AND2_X1 U739 ( .A1(n652), .A2(n651), .ZN(n653) );
  NAND2_X1 U740 ( .A1(n654), .A2(n653), .ZN(G290) );
  NAND2_X1 U741 ( .A1(G61), .A2(n655), .ZN(n658) );
  NAND2_X1 U742 ( .A1(G86), .A2(n656), .ZN(n657) );
  NAND2_X1 U743 ( .A1(n658), .A2(n657), .ZN(n662) );
  NAND2_X1 U744 ( .A1(n659), .A2(G73), .ZN(n660) );
  XOR2_X1 U745 ( .A(KEYINPUT2), .B(n660), .Z(n661) );
  NOR2_X1 U746 ( .A1(n662), .A2(n661), .ZN(n665) );
  NAND2_X1 U747 ( .A1(n663), .A2(G48), .ZN(n664) );
  NAND2_X1 U748 ( .A1(n665), .A2(n664), .ZN(G305) );
  XNOR2_X1 U749 ( .A(n950), .B(n674), .ZN(n670) );
  XOR2_X1 U750 ( .A(KEYINPUT19), .B(KEYINPUT83), .Z(n666) );
  XNOR2_X1 U751 ( .A(G288), .B(n666), .ZN(n667) );
  XNOR2_X1 U752 ( .A(n667), .B(G290), .ZN(n668) );
  XNOR2_X1 U753 ( .A(n668), .B(G305), .ZN(n669) );
  XNOR2_X1 U754 ( .A(n670), .B(n669), .ZN(n671) );
  XNOR2_X1 U755 ( .A(G303), .B(n671), .ZN(n887) );
  XNOR2_X1 U756 ( .A(n887), .B(n672), .ZN(n673) );
  NAND2_X1 U757 ( .A1(n673), .A2(G868), .ZN(n676) );
  OR2_X1 U758 ( .A1(G868), .A2(n674), .ZN(n675) );
  NAND2_X1 U759 ( .A1(n676), .A2(n675), .ZN(G295) );
  XOR2_X1 U760 ( .A(KEYINPUT84), .B(KEYINPUT20), .Z(n678) );
  NAND2_X1 U761 ( .A1(G2084), .A2(G2078), .ZN(n677) );
  XNOR2_X1 U762 ( .A(n678), .B(n677), .ZN(n679) );
  NAND2_X1 U763 ( .A1(n679), .A2(G2090), .ZN(n680) );
  XOR2_X1 U764 ( .A(KEYINPUT85), .B(n680), .Z(n681) );
  XNOR2_X1 U765 ( .A(KEYINPUT21), .B(n681), .ZN(n682) );
  NAND2_X1 U766 ( .A1(n682), .A2(G2072), .ZN(G158) );
  XOR2_X1 U767 ( .A(KEYINPUT72), .B(G57), .Z(G237) );
  XNOR2_X1 U768 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U769 ( .A1(G108), .A2(G120), .ZN(n683) );
  NOR2_X1 U770 ( .A1(G237), .A2(n683), .ZN(n684) );
  NAND2_X1 U771 ( .A1(G69), .A2(n684), .ZN(n839) );
  NAND2_X1 U772 ( .A1(n839), .A2(G567), .ZN(n689) );
  NOR2_X1 U773 ( .A1(G220), .A2(G219), .ZN(n685) );
  XOR2_X1 U774 ( .A(KEYINPUT22), .B(n685), .Z(n686) );
  NOR2_X1 U775 ( .A1(G218), .A2(n686), .ZN(n687) );
  NAND2_X1 U776 ( .A1(G96), .A2(n687), .ZN(n840) );
  NAND2_X1 U777 ( .A1(n840), .A2(G2106), .ZN(n688) );
  NAND2_X1 U778 ( .A1(n689), .A2(n688), .ZN(n841) );
  NAND2_X1 U779 ( .A1(G483), .A2(G661), .ZN(n690) );
  NOR2_X1 U780 ( .A1(n841), .A2(n690), .ZN(n838) );
  NAND2_X1 U781 ( .A1(n838), .A2(G36), .ZN(G176) );
  NAND2_X1 U782 ( .A1(G160), .A2(G40), .ZN(n784) );
  XNOR2_X1 U783 ( .A(n784), .B(KEYINPUT93), .ZN(n691) );
  NAND2_X1 U784 ( .A1(G8), .A2(n694), .ZN(n776) );
  NOR2_X1 U785 ( .A1(G1966), .A2(n776), .ZN(n738) );
  XNOR2_X1 U786 ( .A(G2078), .B(KEYINPUT25), .ZN(n925) );
  NOR2_X1 U787 ( .A1(n694), .A2(n925), .ZN(n693) );
  INV_X1 U788 ( .A(G1961), .ZN(n963) );
  NOR2_X1 U789 ( .A1(n713), .A2(n963), .ZN(n692) );
  NOR2_X1 U790 ( .A1(n693), .A2(n692), .ZN(n731) );
  NAND2_X1 U791 ( .A1(G171), .A2(n731), .ZN(n726) );
  INV_X1 U792 ( .A(G1996), .ZN(n919) );
  XNOR2_X1 U793 ( .A(n696), .B(n695), .ZN(n698) );
  NAND2_X1 U794 ( .A1(n694), .A2(G1341), .ZN(n697) );
  NAND2_X1 U795 ( .A1(n698), .A2(n697), .ZN(n700) );
  NOR2_X1 U796 ( .A1(n700), .A2(n699), .ZN(n702) );
  INV_X1 U797 ( .A(KEYINPUT64), .ZN(n701) );
  XNOR2_X1 U798 ( .A(n702), .B(n701), .ZN(n708) );
  OR2_X1 U799 ( .A1(n708), .A2(n707), .ZN(n706) );
  NOR2_X1 U800 ( .A1(n713), .A2(G1348), .ZN(n704) );
  NOR2_X1 U801 ( .A1(G2067), .A2(n694), .ZN(n703) );
  NOR2_X1 U802 ( .A1(n704), .A2(n703), .ZN(n705) );
  NAND2_X1 U803 ( .A1(n706), .A2(n705), .ZN(n710) );
  NAND2_X1 U804 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U805 ( .A1(n710), .A2(n709), .ZN(n717) );
  NAND2_X1 U806 ( .A1(G2072), .A2(n713), .ZN(n712) );
  XNOR2_X1 U807 ( .A(KEYINPUT94), .B(KEYINPUT27), .ZN(n711) );
  XNOR2_X1 U808 ( .A(n712), .B(n711), .ZN(n715) );
  INV_X1 U809 ( .A(G1956), .ZN(n949) );
  NOR2_X1 U810 ( .A1(n713), .A2(n949), .ZN(n714) );
  NOR2_X1 U811 ( .A1(n715), .A2(n714), .ZN(n718) );
  NAND2_X1 U812 ( .A1(n950), .A2(n718), .ZN(n716) );
  NAND2_X1 U813 ( .A1(n717), .A2(n716), .ZN(n722) );
  NOR2_X1 U814 ( .A1(n950), .A2(n718), .ZN(n720) );
  XNOR2_X1 U815 ( .A(KEYINPUT95), .B(KEYINPUT28), .ZN(n719) );
  XNOR2_X1 U816 ( .A(n720), .B(n719), .ZN(n721) );
  NAND2_X1 U817 ( .A1(n722), .A2(n721), .ZN(n724) );
  XNOR2_X1 U818 ( .A(n724), .B(n723), .ZN(n725) );
  NAND2_X1 U819 ( .A1(n726), .A2(n725), .ZN(n736) );
  NOR2_X1 U820 ( .A1(G2084), .A2(n694), .ZN(n739) );
  NOR2_X1 U821 ( .A1(n738), .A2(n739), .ZN(n727) );
  NAND2_X1 U822 ( .A1(G8), .A2(n727), .ZN(n729) );
  NOR2_X1 U823 ( .A1(G168), .A2(n730), .ZN(n733) );
  NOR2_X1 U824 ( .A1(G171), .A2(n731), .ZN(n732) );
  NOR2_X1 U825 ( .A1(n733), .A2(n732), .ZN(n734) );
  XOR2_X1 U826 ( .A(KEYINPUT31), .B(n734), .Z(n735) );
  NAND2_X1 U827 ( .A1(n736), .A2(n735), .ZN(n742) );
  INV_X1 U828 ( .A(n742), .ZN(n737) );
  NOR2_X1 U829 ( .A1(n738), .A2(n737), .ZN(n741) );
  NAND2_X1 U830 ( .A1(G8), .A2(n739), .ZN(n740) );
  NAND2_X1 U831 ( .A1(n741), .A2(n740), .ZN(n764) );
  NAND2_X1 U832 ( .A1(n742), .A2(G286), .ZN(n751) );
  INV_X1 U833 ( .A(G8), .ZN(n749) );
  NOR2_X1 U834 ( .A1(G1971), .A2(n776), .ZN(n744) );
  NOR2_X1 U835 ( .A1(G2090), .A2(n694), .ZN(n743) );
  NOR2_X1 U836 ( .A1(n744), .A2(n743), .ZN(n745) );
  XNOR2_X1 U837 ( .A(n745), .B(KEYINPUT97), .ZN(n746) );
  NOR2_X1 U838 ( .A1(G166), .A2(n746), .ZN(n747) );
  XOR2_X1 U839 ( .A(KEYINPUT98), .B(n747), .Z(n748) );
  OR2_X1 U840 ( .A1(n749), .A2(n748), .ZN(n750) );
  XNOR2_X1 U841 ( .A(n752), .B(KEYINPUT32), .ZN(n765) );
  NAND2_X1 U842 ( .A1(n764), .A2(n765), .ZN(n755) );
  NOR2_X1 U843 ( .A1(G303), .A2(G2090), .ZN(n753) );
  NAND2_X1 U844 ( .A1(G8), .A2(n753), .ZN(n754) );
  NAND2_X1 U845 ( .A1(n755), .A2(n754), .ZN(n757) );
  INV_X1 U846 ( .A(KEYINPUT101), .ZN(n756) );
  XNOR2_X1 U847 ( .A(n757), .B(n756), .ZN(n758) );
  NAND2_X1 U848 ( .A1(n758), .A2(n776), .ZN(n762) );
  NOR2_X1 U849 ( .A1(G1981), .A2(G305), .ZN(n759) );
  XOR2_X1 U850 ( .A(n759), .B(KEYINPUT24), .Z(n760) );
  OR2_X1 U851 ( .A1(n776), .A2(n760), .ZN(n761) );
  AND2_X1 U852 ( .A1(n762), .A2(n761), .ZN(n783) );
  INV_X1 U853 ( .A(n776), .ZN(n763) );
  NAND2_X1 U854 ( .A1(G1976), .A2(G288), .ZN(n953) );
  AND2_X1 U855 ( .A1(n763), .A2(n953), .ZN(n767) );
  AND2_X1 U856 ( .A1(n764), .A2(n767), .ZN(n766) );
  AND2_X1 U857 ( .A1(n766), .A2(n765), .ZN(n775) );
  INV_X1 U858 ( .A(n767), .ZN(n771) );
  NOR2_X1 U859 ( .A1(G1976), .A2(G288), .ZN(n952) );
  NOR2_X1 U860 ( .A1(G303), .A2(G1971), .ZN(n768) );
  XOR2_X1 U861 ( .A(n768), .B(KEYINPUT99), .Z(n769) );
  NOR2_X1 U862 ( .A1(n952), .A2(n769), .ZN(n770) );
  OR2_X1 U863 ( .A1(n771), .A2(n770), .ZN(n773) );
  INV_X1 U864 ( .A(KEYINPUT33), .ZN(n772) );
  NAND2_X1 U865 ( .A1(n773), .A2(n772), .ZN(n774) );
  NOR2_X1 U866 ( .A1(n775), .A2(n774), .ZN(n779) );
  NAND2_X1 U867 ( .A1(n952), .A2(KEYINPUT33), .ZN(n777) );
  XOR2_X1 U868 ( .A(G1981), .B(G305), .Z(n939) );
  NOR2_X1 U869 ( .A1(n779), .A2(n778), .ZN(n781) );
  XNOR2_X1 U870 ( .A(n781), .B(n780), .ZN(n782) );
  NAND2_X1 U871 ( .A1(n783), .A2(n782), .ZN(n806) );
  NOR2_X1 U872 ( .A1(n785), .A2(n784), .ZN(n829) );
  XOR2_X1 U873 ( .A(KEYINPUT38), .B(KEYINPUT90), .Z(n787) );
  NAND2_X1 U874 ( .A1(G105), .A2(n874), .ZN(n786) );
  XNOR2_X1 U875 ( .A(n787), .B(n786), .ZN(n792) );
  NAND2_X1 U876 ( .A1(G117), .A2(n869), .ZN(n789) );
  NAND2_X1 U877 ( .A1(G129), .A2(n531), .ZN(n788) );
  NAND2_X1 U878 ( .A1(n789), .A2(n788), .ZN(n790) );
  XOR2_X1 U879 ( .A(KEYINPUT89), .B(n790), .Z(n791) );
  NOR2_X1 U880 ( .A1(n792), .A2(n791), .ZN(n794) );
  NAND2_X1 U881 ( .A1(n873), .A2(G141), .ZN(n793) );
  NAND2_X1 U882 ( .A1(n794), .A2(n793), .ZN(n851) );
  NAND2_X1 U883 ( .A1(G1996), .A2(n851), .ZN(n795) );
  XOR2_X1 U884 ( .A(KEYINPUT91), .B(n795), .Z(n803) );
  NAND2_X1 U885 ( .A1(G131), .A2(n873), .ZN(n797) );
  NAND2_X1 U886 ( .A1(G107), .A2(n869), .ZN(n796) );
  NAND2_X1 U887 ( .A1(n797), .A2(n796), .ZN(n801) );
  NAND2_X1 U888 ( .A1(G95), .A2(n874), .ZN(n799) );
  NAND2_X1 U889 ( .A1(G119), .A2(n531), .ZN(n798) );
  NAND2_X1 U890 ( .A1(n799), .A2(n798), .ZN(n800) );
  OR2_X1 U891 ( .A1(n801), .A2(n800), .ZN(n863) );
  NAND2_X1 U892 ( .A1(G1991), .A2(n863), .ZN(n802) );
  NAND2_X1 U893 ( .A1(n803), .A2(n802), .ZN(n999) );
  NAND2_X1 U894 ( .A1(n829), .A2(n999), .ZN(n804) );
  XOR2_X1 U895 ( .A(KEYINPUT92), .B(n804), .Z(n821) );
  XNOR2_X1 U896 ( .A(G1986), .B(G290), .ZN(n956) );
  XNOR2_X1 U897 ( .A(KEYINPUT34), .B(KEYINPUT88), .ZN(n810) );
  NAND2_X1 U898 ( .A1(G140), .A2(n873), .ZN(n808) );
  NAND2_X1 U899 ( .A1(G104), .A2(n874), .ZN(n807) );
  NAND2_X1 U900 ( .A1(n808), .A2(n807), .ZN(n809) );
  XNOR2_X1 U901 ( .A(n810), .B(n809), .ZN(n815) );
  NAND2_X1 U902 ( .A1(G116), .A2(n869), .ZN(n812) );
  NAND2_X1 U903 ( .A1(G128), .A2(n531), .ZN(n811) );
  NAND2_X1 U904 ( .A1(n812), .A2(n811), .ZN(n813) );
  XOR2_X1 U905 ( .A(KEYINPUT35), .B(n813), .Z(n814) );
  NOR2_X1 U906 ( .A1(n815), .A2(n814), .ZN(n816) );
  XNOR2_X1 U907 ( .A(KEYINPUT36), .B(n816), .ZN(n850) );
  XNOR2_X1 U908 ( .A(KEYINPUT37), .B(G2067), .ZN(n826) );
  NOR2_X1 U909 ( .A1(n850), .A2(n826), .ZN(n996) );
  NAND2_X1 U910 ( .A1(n829), .A2(n996), .ZN(n824) );
  NAND2_X1 U911 ( .A1(n817), .A2(n824), .ZN(n818) );
  XNOR2_X1 U912 ( .A(n818), .B(KEYINPUT102), .ZN(n831) );
  NOR2_X1 U913 ( .A1(G1996), .A2(n851), .ZN(n1013) );
  NOR2_X1 U914 ( .A1(G1991), .A2(n863), .ZN(n1003) );
  NOR2_X1 U915 ( .A1(G1986), .A2(G290), .ZN(n819) );
  NOR2_X1 U916 ( .A1(n1003), .A2(n819), .ZN(n820) );
  NOR2_X1 U917 ( .A1(n821), .A2(n820), .ZN(n822) );
  NOR2_X1 U918 ( .A1(n1013), .A2(n822), .ZN(n823) );
  XNOR2_X1 U919 ( .A(n823), .B(KEYINPUT39), .ZN(n825) );
  NAND2_X1 U920 ( .A1(n825), .A2(n824), .ZN(n827) );
  NAND2_X1 U921 ( .A1(n850), .A2(n826), .ZN(n995) );
  NAND2_X1 U922 ( .A1(n827), .A2(n995), .ZN(n828) );
  NAND2_X1 U923 ( .A1(n829), .A2(n828), .ZN(n830) );
  NAND2_X1 U924 ( .A1(n831), .A2(n830), .ZN(n832) );
  XNOR2_X1 U925 ( .A(n832), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U926 ( .A1(n833), .A2(G2106), .ZN(n834) );
  XNOR2_X1 U927 ( .A(n834), .B(KEYINPUT104), .ZN(G217) );
  AND2_X1 U928 ( .A1(G15), .A2(G2), .ZN(n835) );
  NAND2_X1 U929 ( .A1(G661), .A2(n835), .ZN(G259) );
  NAND2_X1 U930 ( .A1(G3), .A2(G1), .ZN(n836) );
  XOR2_X1 U931 ( .A(KEYINPUT105), .B(n836), .Z(n837) );
  NAND2_X1 U932 ( .A1(n838), .A2(n837), .ZN(G188) );
  INV_X1 U934 ( .A(G120), .ZN(G236) );
  INV_X1 U935 ( .A(G108), .ZN(G238) );
  INV_X1 U936 ( .A(G96), .ZN(G221) );
  INV_X1 U937 ( .A(G69), .ZN(G235) );
  NOR2_X1 U938 ( .A1(n840), .A2(n839), .ZN(G325) );
  INV_X1 U939 ( .A(G325), .ZN(G261) );
  INV_X1 U940 ( .A(n841), .ZN(G319) );
  NAND2_X1 U941 ( .A1(G100), .A2(n874), .ZN(n843) );
  NAND2_X1 U942 ( .A1(G112), .A2(n869), .ZN(n842) );
  NAND2_X1 U943 ( .A1(n843), .A2(n842), .ZN(n849) );
  NAND2_X1 U944 ( .A1(n531), .A2(G124), .ZN(n844) );
  XNOR2_X1 U945 ( .A(n844), .B(KEYINPUT44), .ZN(n846) );
  NAND2_X1 U946 ( .A1(G136), .A2(n873), .ZN(n845) );
  NAND2_X1 U947 ( .A1(n846), .A2(n845), .ZN(n847) );
  XOR2_X1 U948 ( .A(KEYINPUT109), .B(n847), .Z(n848) );
  NOR2_X1 U949 ( .A1(n849), .A2(n848), .ZN(G162) );
  XNOR2_X1 U950 ( .A(G160), .B(n850), .ZN(n852) );
  XNOR2_X1 U951 ( .A(n852), .B(n851), .ZN(n853) );
  XNOR2_X1 U952 ( .A(n1000), .B(n853), .ZN(n862) );
  NAND2_X1 U953 ( .A1(G139), .A2(n873), .ZN(n855) );
  NAND2_X1 U954 ( .A1(G103), .A2(n874), .ZN(n854) );
  NAND2_X1 U955 ( .A1(n855), .A2(n854), .ZN(n860) );
  NAND2_X1 U956 ( .A1(G115), .A2(n869), .ZN(n857) );
  NAND2_X1 U957 ( .A1(G127), .A2(n531), .ZN(n856) );
  NAND2_X1 U958 ( .A1(n857), .A2(n856), .ZN(n858) );
  XOR2_X1 U959 ( .A(KEYINPUT47), .B(n858), .Z(n859) );
  NOR2_X1 U960 ( .A1(n860), .A2(n859), .ZN(n1006) );
  XNOR2_X1 U961 ( .A(n1006), .B(G162), .ZN(n861) );
  XNOR2_X1 U962 ( .A(n862), .B(n861), .ZN(n867) );
  XNOR2_X1 U963 ( .A(KEYINPUT48), .B(KEYINPUT112), .ZN(n865) );
  XNOR2_X1 U964 ( .A(n863), .B(KEYINPUT46), .ZN(n864) );
  XNOR2_X1 U965 ( .A(n865), .B(n864), .ZN(n866) );
  XOR2_X1 U966 ( .A(n867), .B(n866), .Z(n882) );
  NAND2_X1 U967 ( .A1(G130), .A2(n531), .ZN(n868) );
  XNOR2_X1 U968 ( .A(n868), .B(KEYINPUT110), .ZN(n872) );
  NAND2_X1 U969 ( .A1(G118), .A2(n869), .ZN(n870) );
  XOR2_X1 U970 ( .A(KEYINPUT111), .B(n870), .Z(n871) );
  NAND2_X1 U971 ( .A1(n872), .A2(n871), .ZN(n879) );
  NAND2_X1 U972 ( .A1(G142), .A2(n873), .ZN(n876) );
  NAND2_X1 U973 ( .A1(G106), .A2(n874), .ZN(n875) );
  NAND2_X1 U974 ( .A1(n876), .A2(n875), .ZN(n877) );
  XOR2_X1 U975 ( .A(KEYINPUT45), .B(n877), .Z(n878) );
  NOR2_X1 U976 ( .A1(n879), .A2(n878), .ZN(n880) );
  XNOR2_X1 U977 ( .A(G164), .B(n880), .ZN(n881) );
  XNOR2_X1 U978 ( .A(n882), .B(n881), .ZN(n883) );
  NOR2_X1 U979 ( .A1(G37), .A2(n883), .ZN(n884) );
  XOR2_X1 U980 ( .A(KEYINPUT113), .B(n884), .Z(G395) );
  XNOR2_X1 U981 ( .A(n699), .B(G286), .ZN(n886) );
  XNOR2_X1 U982 ( .A(G171), .B(n946), .ZN(n885) );
  XNOR2_X1 U983 ( .A(n886), .B(n885), .ZN(n888) );
  XNOR2_X1 U984 ( .A(n888), .B(n887), .ZN(n889) );
  NOR2_X1 U985 ( .A1(G37), .A2(n889), .ZN(G397) );
  XOR2_X1 U986 ( .A(G1981), .B(G1956), .Z(n891) );
  XNOR2_X1 U987 ( .A(G1966), .B(G1961), .ZN(n890) );
  XNOR2_X1 U988 ( .A(n891), .B(n890), .ZN(n892) );
  XOR2_X1 U989 ( .A(n892), .B(G2474), .Z(n894) );
  XNOR2_X1 U990 ( .A(G1996), .B(G1991), .ZN(n893) );
  XNOR2_X1 U991 ( .A(n894), .B(n893), .ZN(n898) );
  XOR2_X1 U992 ( .A(KEYINPUT41), .B(G1976), .Z(n896) );
  XNOR2_X1 U993 ( .A(G1986), .B(G1971), .ZN(n895) );
  XNOR2_X1 U994 ( .A(n896), .B(n895), .ZN(n897) );
  XNOR2_X1 U995 ( .A(n898), .B(n897), .ZN(G229) );
  XOR2_X1 U996 ( .A(KEYINPUT108), .B(G2678), .Z(n900) );
  XNOR2_X1 U997 ( .A(KEYINPUT43), .B(G2096), .ZN(n899) );
  XNOR2_X1 U998 ( .A(n900), .B(n899), .ZN(n901) );
  XOR2_X1 U999 ( .A(n901), .B(KEYINPUT107), .Z(n903) );
  XNOR2_X1 U1000 ( .A(G2078), .B(G2072), .ZN(n902) );
  XNOR2_X1 U1001 ( .A(n903), .B(n902), .ZN(n907) );
  XOR2_X1 U1002 ( .A(G2100), .B(G2084), .Z(n905) );
  XNOR2_X1 U1003 ( .A(G2067), .B(G2090), .ZN(n904) );
  XNOR2_X1 U1004 ( .A(n905), .B(n904), .ZN(n906) );
  XOR2_X1 U1005 ( .A(n907), .B(n906), .Z(n909) );
  XNOR2_X1 U1006 ( .A(KEYINPUT106), .B(KEYINPUT42), .ZN(n908) );
  XNOR2_X1 U1007 ( .A(n909), .B(n908), .ZN(G227) );
  NOR2_X1 U1008 ( .A1(G395), .A2(G397), .ZN(n910) );
  XNOR2_X1 U1009 ( .A(n910), .B(KEYINPUT114), .ZN(n911) );
  NAND2_X1 U1010 ( .A1(G319), .A2(n911), .ZN(n912) );
  NOR2_X1 U1011 ( .A1(G401), .A2(n912), .ZN(n915) );
  NOR2_X1 U1012 ( .A1(G229), .A2(G227), .ZN(n913) );
  XOR2_X1 U1013 ( .A(KEYINPUT49), .B(n913), .Z(n914) );
  NAND2_X1 U1014 ( .A1(n915), .A2(n914), .ZN(G225) );
  INV_X1 U1015 ( .A(G225), .ZN(G308) );
  XNOR2_X1 U1016 ( .A(G1991), .B(G25), .ZN(n917) );
  XNOR2_X1 U1017 ( .A(G33), .B(G2072), .ZN(n916) );
  NOR2_X1 U1018 ( .A1(n917), .A2(n916), .ZN(n924) );
  XOR2_X1 U1019 ( .A(G2067), .B(G26), .Z(n918) );
  NAND2_X1 U1020 ( .A1(n918), .A2(G28), .ZN(n922) );
  XOR2_X1 U1021 ( .A(G32), .B(n919), .Z(n920) );
  XNOR2_X1 U1022 ( .A(KEYINPUT120), .B(n920), .ZN(n921) );
  NOR2_X1 U1023 ( .A1(n922), .A2(n921), .ZN(n923) );
  NAND2_X1 U1024 ( .A1(n924), .A2(n923), .ZN(n928) );
  XNOR2_X1 U1025 ( .A(G27), .B(n925), .ZN(n926) );
  XNOR2_X1 U1026 ( .A(KEYINPUT119), .B(n926), .ZN(n927) );
  NOR2_X1 U1027 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1028 ( .A(n929), .B(KEYINPUT53), .ZN(n930) );
  XNOR2_X1 U1029 ( .A(n930), .B(KEYINPUT121), .ZN(n933) );
  XOR2_X1 U1030 ( .A(G2084), .B(G34), .Z(n931) );
  XNOR2_X1 U1031 ( .A(KEYINPUT54), .B(n931), .ZN(n932) );
  NAND2_X1 U1032 ( .A1(n933), .A2(n932), .ZN(n935) );
  XNOR2_X1 U1033 ( .A(G35), .B(G2090), .ZN(n934) );
  NOR2_X1 U1034 ( .A1(n935), .A2(n934), .ZN(n936) );
  XOR2_X1 U1035 ( .A(KEYINPUT55), .B(n936), .Z(n937) );
  XNOR2_X1 U1036 ( .A(KEYINPUT122), .B(n937), .ZN(n938) );
  NOR2_X1 U1037 ( .A1(G29), .A2(n938), .ZN(n993) );
  XOR2_X1 U1038 ( .A(G16), .B(KEYINPUT56), .Z(n962) );
  XNOR2_X1 U1039 ( .A(G1966), .B(G168), .ZN(n940) );
  NAND2_X1 U1040 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1041 ( .A(n941), .B(KEYINPUT57), .ZN(n945) );
  XNOR2_X1 U1042 ( .A(G301), .B(G1961), .ZN(n943) );
  XNOR2_X1 U1043 ( .A(n699), .B(G1341), .ZN(n942) );
  NOR2_X1 U1044 ( .A1(n943), .A2(n942), .ZN(n944) );
  NAND2_X1 U1045 ( .A1(n945), .A2(n944), .ZN(n960) );
  XOR2_X1 U1046 ( .A(G1348), .B(n946), .Z(n948) );
  XNOR2_X1 U1047 ( .A(G303), .B(G1971), .ZN(n947) );
  NOR2_X1 U1048 ( .A1(n948), .A2(n947), .ZN(n958) );
  XNOR2_X1 U1049 ( .A(n950), .B(n949), .ZN(n951) );
  NOR2_X1 U1050 ( .A1(n952), .A2(n951), .ZN(n954) );
  NAND2_X1 U1051 ( .A1(n954), .A2(n953), .ZN(n955) );
  NOR2_X1 U1052 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1053 ( .A1(n958), .A2(n957), .ZN(n959) );
  NOR2_X1 U1054 ( .A1(n960), .A2(n959), .ZN(n961) );
  NOR2_X1 U1055 ( .A1(n962), .A2(n961), .ZN(n990) );
  XNOR2_X1 U1056 ( .A(G5), .B(n963), .ZN(n985) );
  XNOR2_X1 U1057 ( .A(KEYINPUT123), .B(G1981), .ZN(n964) );
  XNOR2_X1 U1058 ( .A(n964), .B(G6), .ZN(n970) );
  XOR2_X1 U1059 ( .A(KEYINPUT124), .B(G4), .Z(n966) );
  XNOR2_X1 U1060 ( .A(G1348), .B(KEYINPUT59), .ZN(n965) );
  XNOR2_X1 U1061 ( .A(n966), .B(n965), .ZN(n968) );
  XNOR2_X1 U1062 ( .A(G1341), .B(G19), .ZN(n967) );
  NOR2_X1 U1063 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1064 ( .A1(n970), .A2(n969), .ZN(n972) );
  XNOR2_X1 U1065 ( .A(G20), .B(G1956), .ZN(n971) );
  NOR2_X1 U1066 ( .A1(n972), .A2(n971), .ZN(n973) );
  XOR2_X1 U1067 ( .A(KEYINPUT60), .B(n973), .Z(n975) );
  XNOR2_X1 U1068 ( .A(G1966), .B(G21), .ZN(n974) );
  NOR2_X1 U1069 ( .A1(n975), .A2(n974), .ZN(n976) );
  XNOR2_X1 U1070 ( .A(KEYINPUT125), .B(n976), .ZN(n983) );
  XNOR2_X1 U1071 ( .A(G1971), .B(G22), .ZN(n978) );
  XNOR2_X1 U1072 ( .A(G23), .B(G1976), .ZN(n977) );
  NOR2_X1 U1073 ( .A1(n978), .A2(n977), .ZN(n980) );
  XOR2_X1 U1074 ( .A(G1986), .B(G24), .Z(n979) );
  NAND2_X1 U1075 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1076 ( .A(KEYINPUT58), .B(n981), .ZN(n982) );
  NOR2_X1 U1077 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1078 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1079 ( .A(KEYINPUT61), .B(n986), .ZN(n987) );
  NOR2_X1 U1080 ( .A1(G16), .A2(n987), .ZN(n988) );
  XNOR2_X1 U1081 ( .A(KEYINPUT126), .B(n988), .ZN(n989) );
  NOR2_X1 U1082 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1083 ( .A1(G11), .A2(n991), .ZN(n992) );
  NOR2_X1 U1084 ( .A1(n993), .A2(n992), .ZN(n994) );
  XNOR2_X1 U1085 ( .A(KEYINPUT127), .B(n994), .ZN(n1025) );
  INV_X1 U1086 ( .A(n995), .ZN(n997) );
  NOR2_X1 U1087 ( .A1(n997), .A2(n996), .ZN(n1005) );
  XOR2_X1 U1088 ( .A(G160), .B(G2084), .Z(n998) );
  NOR2_X1 U1089 ( .A1(n999), .A2(n998), .ZN(n1001) );
  NAND2_X1 U1090 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NOR2_X1 U1091 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1092 ( .A1(n1005), .A2(n1004), .ZN(n1018) );
  XNOR2_X1 U1093 ( .A(G2072), .B(n1006), .ZN(n1007) );
  XNOR2_X1 U1094 ( .A(n1007), .B(KEYINPUT115), .ZN(n1009) );
  XOR2_X1 U1095 ( .A(G2078), .B(G164), .Z(n1008) );
  NOR2_X1 U1096 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1097 ( .A(KEYINPUT50), .B(n1010), .ZN(n1011) );
  XNOR2_X1 U1098 ( .A(n1011), .B(KEYINPUT116), .ZN(n1016) );
  XOR2_X1 U1099 ( .A(G2090), .B(G162), .Z(n1012) );
  NOR2_X1 U1100 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XOR2_X1 U1101 ( .A(KEYINPUT51), .B(n1014), .Z(n1015) );
  NAND2_X1 U1102 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NOR2_X1 U1103 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XOR2_X1 U1104 ( .A(KEYINPUT52), .B(n1019), .Z(n1020) );
  NOR2_X1 U1105 ( .A1(KEYINPUT55), .A2(n1020), .ZN(n1021) );
  XNOR2_X1 U1106 ( .A(KEYINPUT117), .B(n1021), .ZN(n1022) );
  NAND2_X1 U1107 ( .A1(n1022), .A2(G29), .ZN(n1023) );
  XOR2_X1 U1108 ( .A(KEYINPUT118), .B(n1023), .Z(n1024) );
  NOR2_X1 U1109 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XNOR2_X1 U1110 ( .A(KEYINPUT62), .B(n1026), .ZN(G311) );
  INV_X1 U1111 ( .A(G311), .ZN(G150) );
endmodule

