//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 0 0 0 0 0 1 0 1 0 1 0 1 1 0 0 0 0 1 0 1 0 0 1 1 1 1 1 0 1 1 1 1 1 1 0 1 1 1 0 0 1 0 0 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n724,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n752, new_n754, new_n755, new_n756,
    new_n757, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n770, new_n771, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n795, new_n796,
    new_n797, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n839, new_n841, new_n842,
    new_n844, new_n845, new_n846, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n896, new_n897, new_n898, new_n899, new_n901, new_n902, new_n903,
    new_n904, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n963, new_n964, new_n965;
  NAND2_X1  g000(.A1(G226gat), .A2(G233gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(G183gat), .A2(G190gat), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  OR2_X1    g003(.A1(G169gat), .A2(G176gat), .ZN(new_n205));
  OR2_X1    g004(.A1(new_n205), .A2(KEYINPUT26), .ZN(new_n206));
  NAND2_X1  g005(.A1(G169gat), .A2(G176gat), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  AOI21_X1  g007(.A(new_n208), .B1(KEYINPUT26), .B2(new_n205), .ZN(new_n209));
  AOI21_X1  g008(.A(new_n204), .B1(new_n206), .B2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(G183gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(KEYINPUT27), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT27), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(G183gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  NOR3_X1   g015(.A1(new_n216), .A2(KEYINPUT28), .A3(G190gat), .ZN(new_n217));
  INV_X1    g016(.A(new_n217), .ZN(new_n218));
  AND3_X1   g017(.A1(new_n213), .A2(new_n215), .A3(KEYINPUT67), .ZN(new_n219));
  AOI21_X1  g018(.A(KEYINPUT67), .B1(new_n213), .B2(new_n215), .ZN(new_n220));
  NOR3_X1   g019(.A1(new_n219), .A2(new_n220), .A3(G190gat), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT28), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n218), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT68), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n211), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT67), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n216), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(G190gat), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n213), .A2(new_n215), .A3(KEYINPUT67), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n227), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  AOI211_X1 g029(.A(new_n224), .B(new_n217), .C1(new_n230), .C2(KEYINPUT28), .ZN(new_n231));
  INV_X1    g030(.A(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT25), .ZN(new_n233));
  XNOR2_X1  g032(.A(new_n205), .B(KEYINPUT23), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(new_n207), .ZN(new_n235));
  AND3_X1   g034(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n236), .B1(new_n212), .B2(new_n228), .ZN(new_n237));
  OR2_X1    g036(.A1(new_n204), .A2(KEYINPUT24), .ZN(new_n238));
  AND2_X1   g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n233), .B1(new_n235), .B2(new_n239), .ZN(new_n240));
  OR2_X1    g039(.A1(new_n207), .A2(KEYINPUT64), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n207), .A2(KEYINPUT64), .ZN(new_n242));
  AND3_X1   g041(.A1(new_n241), .A2(KEYINPUT25), .A3(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT66), .ZN(new_n244));
  XNOR2_X1  g043(.A(KEYINPUT65), .B(KEYINPUT24), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n244), .B1(new_n245), .B2(new_n204), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(new_n237), .ZN(new_n247));
  NOR3_X1   g046(.A1(new_n245), .A2(new_n244), .A3(new_n204), .ZN(new_n248));
  OAI211_X1 g047(.A(new_n234), .B(new_n243), .C1(new_n247), .C2(new_n248), .ZN(new_n249));
  AOI22_X1  g048(.A1(new_n225), .A2(new_n232), .B1(new_n240), .B2(new_n249), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n202), .B1(new_n250), .B2(KEYINPUT29), .ZN(new_n251));
  XNOR2_X1  g050(.A(G197gat), .B(G204gat), .ZN(new_n252));
  NAND2_X1  g051(.A1(G211gat), .A2(G218gat), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n252), .B1(KEYINPUT22), .B2(new_n254), .ZN(new_n255));
  NOR2_X1   g054(.A1(G211gat), .A2(G218gat), .ZN(new_n256));
  NOR3_X1   g055(.A1(new_n254), .A2(new_n256), .A3(KEYINPUT72), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(G197gat), .ZN(new_n259));
  INV_X1    g058(.A(G204gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(G197gat), .A2(G204gat), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT22), .ZN(new_n263));
  AOI22_X1  g062(.A1(new_n261), .A2(new_n262), .B1(new_n263), .B2(new_n253), .ZN(new_n264));
  XNOR2_X1  g063(.A(G211gat), .B(G218gat), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n264), .B1(KEYINPUT72), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n258), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT73), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n258), .A2(KEYINPUT73), .A3(new_n266), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n240), .A2(new_n249), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n217), .B1(new_n230), .B2(KEYINPUT28), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n210), .B1(new_n273), .B2(KEYINPUT68), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n272), .B1(new_n274), .B2(new_n231), .ZN(new_n275));
  INV_X1    g074(.A(new_n202), .ZN(new_n276));
  AND3_X1   g075(.A1(new_n275), .A2(KEYINPUT75), .A3(new_n276), .ZN(new_n277));
  AOI21_X1  g076(.A(KEYINPUT75), .B1(new_n275), .B2(new_n276), .ZN(new_n278));
  OAI211_X1 g077(.A(new_n251), .B(new_n271), .C1(new_n277), .C2(new_n278), .ZN(new_n279));
  AND3_X1   g078(.A1(new_n258), .A2(KEYINPUT73), .A3(new_n266), .ZN(new_n280));
  AOI21_X1  g079(.A(KEYINPUT73), .B1(new_n258), .B2(new_n266), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n250), .A2(new_n202), .ZN(new_n283));
  XOR2_X1   g082(.A(KEYINPUT74), .B(KEYINPUT29), .Z(new_n284));
  AOI21_X1  g083(.A(new_n276), .B1(new_n275), .B2(new_n284), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n282), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(G8gat), .B(G36gat), .ZN(new_n287));
  XNOR2_X1  g086(.A(G64gat), .B(G92gat), .ZN(new_n288));
  XOR2_X1   g087(.A(new_n287), .B(new_n288), .Z(new_n289));
  AND3_X1   g088(.A1(new_n279), .A2(new_n286), .A3(new_n289), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n289), .B1(new_n279), .B2(new_n286), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT30), .ZN(new_n292));
  NOR3_X1   g091(.A1(new_n290), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n279), .A2(new_n286), .ZN(new_n294));
  INV_X1    g093(.A(new_n289), .ZN(new_n295));
  NOR3_X1   g094(.A1(new_n294), .A2(KEYINPUT30), .A3(new_n295), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n293), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  XNOR2_X1  g097(.A(G15gat), .B(G43gat), .ZN(new_n299));
  XNOR2_X1  g098(.A(G71gat), .B(G99gat), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n299), .B(new_n300), .ZN(new_n301));
  OR2_X1    g100(.A1(G113gat), .A2(G120gat), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT70), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT1), .ZN(new_n304));
  NAND2_X1  g103(.A1(G113gat), .A2(G120gat), .ZN(new_n305));
  NAND4_X1  g104(.A1(new_n302), .A2(new_n303), .A3(new_n304), .A4(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(G127gat), .ZN(new_n307));
  INV_X1    g106(.A(G134gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(G127gat), .A2(G134gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT69), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n309), .A2(new_n312), .A3(new_n310), .ZN(new_n313));
  AND2_X1   g112(.A1(G113gat), .A2(G120gat), .ZN(new_n314));
  NOR2_X1   g113(.A1(G113gat), .A2(G120gat), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  AOI21_X1  g115(.A(KEYINPUT1), .B1(new_n313), .B2(new_n316), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n302), .A2(new_n303), .A3(new_n305), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(new_n312), .ZN(new_n319));
  AOI221_X4 g118(.A(KEYINPUT71), .B1(new_n306), .B2(new_n311), .C1(new_n317), .C2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT71), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n313), .A2(new_n316), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n319), .A2(new_n322), .A3(new_n304), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n306), .A2(new_n311), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n321), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n320), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n275), .A2(new_n327), .ZN(new_n328));
  OAI211_X1 g127(.A(new_n326), .B(new_n272), .C1(new_n231), .C2(new_n274), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(G227gat), .A2(G233gat), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT33), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n301), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n328), .A2(new_n329), .A3(new_n331), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(KEYINPUT34), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT34), .ZN(new_n338));
  NAND4_X1  g137(.A1(new_n328), .A2(new_n329), .A3(new_n338), .A4(new_n331), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n335), .A2(new_n340), .ZN(new_n341));
  AOI21_X1  g140(.A(KEYINPUT33), .B1(new_n330), .B2(new_n332), .ZN(new_n342));
  OAI211_X1 g141(.A(new_n337), .B(new_n339), .C1(new_n342), .C2(new_n301), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n333), .A2(KEYINPUT32), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  XNOR2_X1  g145(.A(G78gat), .B(G106gat), .ZN(new_n347));
  XNOR2_X1  g146(.A(new_n347), .B(G50gat), .ZN(new_n348));
  XNOR2_X1  g147(.A(KEYINPUT84), .B(KEYINPUT31), .ZN(new_n349));
  XNOR2_X1  g148(.A(new_n348), .B(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(G155gat), .A2(G162gat), .ZN(new_n351));
  NOR2_X1   g150(.A1(G155gat), .A2(G162gat), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  XNOR2_X1  g152(.A(G141gat), .B(G148gat), .ZN(new_n354));
  XNOR2_X1  g153(.A(KEYINPUT76), .B(KEYINPUT2), .ZN(new_n355));
  OAI211_X1 g154(.A(new_n351), .B(new_n353), .C1(new_n354), .C2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(G148gat), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(KEYINPUT77), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT77), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(G148gat), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n358), .A2(new_n360), .A3(G141gat), .ZN(new_n361));
  INV_X1    g160(.A(G141gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(G148gat), .ZN(new_n363));
  AND2_X1   g162(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT2), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n352), .A2(new_n365), .ZN(new_n366));
  AND2_X1   g165(.A1(new_n366), .A2(new_n351), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n356), .B1(new_n364), .B2(new_n367), .ZN(new_n368));
  AOI21_X1  g167(.A(KEYINPUT29), .B1(new_n258), .B2(new_n266), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n368), .B1(new_n369), .B2(KEYINPUT3), .ZN(new_n370));
  AND2_X1   g169(.A1(G228gat), .A2(G233gat), .ZN(new_n371));
  INV_X1    g170(.A(new_n284), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n353), .A2(new_n351), .ZN(new_n373));
  XOR2_X1   g172(.A(KEYINPUT76), .B(KEYINPUT2), .Z(new_n374));
  NAND2_X1  g173(.A1(new_n357), .A2(G141gat), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n363), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n373), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  AOI22_X1  g176(.A1(new_n361), .A2(new_n363), .B1(new_n351), .B2(new_n366), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT3), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n372), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  OAI211_X1 g180(.A(new_n370), .B(new_n371), .C1(new_n271), .C2(new_n381), .ZN(new_n382));
  OAI211_X1 g181(.A(new_n356), .B(new_n380), .C1(new_n364), .C2(new_n367), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(new_n284), .ZN(new_n384));
  OAI21_X1  g183(.A(KEYINPUT78), .B1(new_n377), .B2(new_n378), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT78), .ZN(new_n386));
  OAI211_X1 g185(.A(new_n356), .B(new_n386), .C1(new_n364), .C2(new_n367), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n255), .A2(new_n265), .ZN(new_n389));
  INV_X1    g188(.A(new_n265), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n284), .B1(new_n390), .B2(new_n264), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n380), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  AOI22_X1  g191(.A1(new_n282), .A2(new_n384), .B1(new_n388), .B2(new_n392), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n382), .B1(new_n393), .B2(new_n371), .ZN(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(G22gat), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n350), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT88), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n394), .A2(KEYINPUT87), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT87), .ZN(new_n400));
  OAI211_X1 g199(.A(new_n382), .B(new_n400), .C1(new_n393), .C2(new_n371), .ZN(new_n401));
  AND4_X1   g200(.A1(new_n398), .A2(new_n399), .A3(G22gat), .A4(new_n401), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n396), .B1(new_n394), .B2(KEYINPUT87), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n398), .B1(new_n403), .B2(new_n401), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n397), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n395), .A2(new_n396), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n394), .A2(G22gat), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n406), .A2(KEYINPUT86), .A3(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT86), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n394), .A2(new_n409), .A3(G22gat), .ZN(new_n410));
  XOR2_X1   g209(.A(new_n350), .B(KEYINPUT85), .Z(new_n411));
  AND2_X1   g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n408), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n405), .A2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(new_n345), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n341), .A2(new_n415), .A3(new_n343), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n346), .A2(new_n414), .A3(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  XNOR2_X1  g217(.A(G1gat), .B(G29gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n419), .B(KEYINPUT0), .ZN(new_n420));
  XNOR2_X1  g219(.A(G57gat), .B(G85gat), .ZN(new_n421));
  XOR2_X1   g220(.A(new_n420), .B(new_n421), .Z(new_n422));
  INV_X1    g221(.A(KEYINPUT4), .ZN(new_n423));
  AND2_X1   g222(.A1(new_n385), .A2(new_n387), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n326), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(KEYINPUT83), .ZN(new_n426));
  NOR3_X1   g225(.A1(new_n388), .A2(new_n320), .A3(new_n325), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT83), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n427), .A2(new_n428), .A3(new_n423), .ZN(new_n429));
  AND2_X1   g228(.A1(new_n323), .A2(new_n324), .ZN(new_n430));
  OAI21_X1  g229(.A(KEYINPUT4), .B1(new_n430), .B2(new_n368), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n426), .A2(new_n429), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n368), .A2(KEYINPUT3), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n433), .A2(new_n430), .A3(new_n383), .ZN(new_n434));
  NAND2_X1  g233(.A1(G225gat), .A2(G233gat), .ZN(new_n435));
  AND2_X1   g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  XOR2_X1   g235(.A(KEYINPUT81), .B(KEYINPUT5), .Z(new_n437));
  NAND3_X1  g236(.A1(new_n432), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n423), .B1(new_n326), .B2(new_n424), .ZN(new_n439));
  AND2_X1   g238(.A1(G127gat), .A2(G134gat), .ZN(new_n440));
  NOR2_X1   g239(.A1(G127gat), .A2(G134gat), .ZN(new_n441));
  NOR3_X1   g240(.A1(new_n440), .A2(new_n441), .A3(KEYINPUT69), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n302), .A2(new_n305), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n304), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  AOI21_X1  g243(.A(KEYINPUT69), .B1(new_n316), .B2(new_n303), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n324), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n446), .A2(new_n423), .A3(new_n379), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(KEYINPUT79), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT79), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n446), .A2(new_n379), .A3(new_n449), .A4(new_n423), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n436), .B1(new_n439), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(KEYINPUT80), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT80), .ZN(new_n454));
  OAI211_X1 g253(.A(new_n436), .B(new_n454), .C1(new_n439), .C2(new_n451), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  XNOR2_X1  g255(.A(new_n446), .B(new_n379), .ZN(new_n457));
  INV_X1    g256(.A(new_n435), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n437), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  AOI21_X1  g258(.A(KEYINPUT82), .B1(new_n456), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT82), .ZN(new_n461));
  INV_X1    g260(.A(new_n459), .ZN(new_n462));
  AOI211_X1 g261(.A(new_n461), .B(new_n462), .C1(new_n453), .C2(new_n455), .ZN(new_n463));
  OAI211_X1 g262(.A(new_n422), .B(new_n438), .C1(new_n460), .C2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT6), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n448), .B(new_n450), .C1(new_n427), .C2(new_n423), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n454), .B1(new_n467), .B2(new_n436), .ZN(new_n468));
  INV_X1    g267(.A(new_n455), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n459), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(new_n461), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n456), .A2(KEYINPUT82), .A3(new_n459), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n422), .B1(new_n473), .B2(new_n438), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n466), .A2(new_n474), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n438), .B1(new_n460), .B2(new_n463), .ZN(new_n476));
  INV_X1    g275(.A(new_n422), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n476), .A2(KEYINPUT6), .A3(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  OAI211_X1 g278(.A(new_n298), .B(new_n418), .C1(new_n475), .C2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(KEYINPUT35), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n476), .A2(new_n477), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n482), .A2(new_n465), .A3(new_n464), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(new_n478), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT35), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n485), .B1(new_n293), .B2(new_n296), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n417), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(KEYINPUT89), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT89), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n484), .A2(new_n487), .A3(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n481), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n484), .A2(new_n298), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n399), .A2(G22gat), .A3(new_n401), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(KEYINPUT88), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n403), .A2(new_n398), .A3(new_n401), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AOI22_X1  g296(.A1(new_n497), .A2(new_n397), .B1(new_n408), .B2(new_n412), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n493), .A2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT38), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n294), .A2(new_n295), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n295), .A2(KEYINPUT37), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n294), .A2(KEYINPUT37), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n500), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n295), .B1(new_n294), .B2(KEYINPUT37), .ZN(new_n506));
  OAI211_X1 g305(.A(new_n251), .B(new_n282), .C1(new_n277), .C2(new_n278), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n271), .B1(new_n283), .B2(new_n285), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n507), .A2(KEYINPUT37), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(new_n500), .ZN(new_n510));
  OAI22_X1  g309(.A1(new_n506), .A2(new_n510), .B1(new_n294), .B2(new_n295), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n505), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n512), .A2(new_n483), .A3(new_n478), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n432), .A2(new_n434), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(new_n458), .ZN(new_n515));
  OR2_X1    g314(.A1(new_n457), .A2(new_n458), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n515), .A2(KEYINPUT39), .A3(new_n516), .ZN(new_n517));
  OAI211_X1 g316(.A(new_n517), .B(new_n422), .C1(KEYINPUT39), .C2(new_n515), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT40), .ZN(new_n519));
  OR2_X1    g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n518), .A2(new_n519), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n520), .A2(new_n482), .A3(new_n297), .A4(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n513), .A2(new_n522), .A3(new_n414), .ZN(new_n523));
  INV_X1    g322(.A(new_n416), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n415), .B1(new_n341), .B2(new_n343), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n526), .B(KEYINPUT36), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n499), .A2(new_n523), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n492), .A2(new_n528), .ZN(new_n529));
  OAI21_X1  g328(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  NOR3_X1   g330(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n532));
  INV_X1    g331(.A(G29gat), .ZN(new_n533));
  INV_X1    g332(.A(G36gat), .ZN(new_n534));
  OAI22_X1  g333(.A1(new_n531), .A2(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  AND2_X1   g334(.A1(G43gat), .A2(G50gat), .ZN(new_n536));
  NOR2_X1   g335(.A1(G43gat), .A2(G50gat), .ZN(new_n537));
  OAI21_X1  g336(.A(KEYINPUT15), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n535), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT91), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT15), .ZN(new_n542));
  AOI22_X1  g341(.A1(new_n541), .A2(new_n542), .B1(G43gat), .B2(G50gat), .ZN(new_n543));
  XNOR2_X1  g342(.A(KEYINPUT92), .B(G50gat), .ZN(new_n544));
  OAI221_X1 g343(.A(new_n543), .B1(new_n541), .B2(new_n542), .C1(new_n544), .C2(G43gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n545), .B(KEYINPUT93), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n538), .B1(new_n533), .B2(new_n534), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n532), .A2(KEYINPUT94), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n548), .A2(new_n531), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n532), .A2(KEYINPUT94), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n547), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n546), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(KEYINPUT95), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n552), .A2(KEYINPUT95), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n540), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT17), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(G15gat), .B(G22gat), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT16), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n559), .B1(new_n560), .B2(G1gat), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n561), .B1(G1gat), .B2(new_n559), .ZN(new_n562));
  INV_X1    g361(.A(G8gat), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n562), .B(new_n563), .ZN(new_n564));
  OAI211_X1 g363(.A(KEYINPUT17), .B(new_n540), .C1(new_n554), .C2(new_n555), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n558), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(G229gat), .A2(G233gat), .ZN(new_n567));
  OR2_X1    g366(.A1(new_n552), .A2(KEYINPUT95), .ZN(new_n568));
  AOI22_X1  g367(.A1(new_n568), .A2(new_n553), .B1(new_n535), .B2(new_n539), .ZN(new_n569));
  OR2_X1    g368(.A1(new_n569), .A2(new_n564), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n566), .A2(new_n567), .A3(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT18), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND4_X1  g372(.A1(new_n566), .A2(KEYINPUT18), .A3(new_n567), .A4(new_n570), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n569), .B(new_n564), .ZN(new_n575));
  XOR2_X1   g374(.A(new_n567), .B(KEYINPUT13), .Z(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(G113gat), .B(G141gat), .ZN(new_n578));
  XNOR2_X1  g377(.A(KEYINPUT90), .B(G197gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(KEYINPUT11), .B(G169gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n580), .B(new_n581), .ZN(new_n582));
  XOR2_X1   g381(.A(new_n582), .B(KEYINPUT12), .Z(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  NAND4_X1  g383(.A1(new_n573), .A2(new_n574), .A3(new_n577), .A4(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  AOI22_X1  g385(.A1(new_n571), .A2(new_n572), .B1(new_n575), .B2(new_n576), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n584), .B1(new_n587), .B2(new_n574), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  AND2_X1   g389(.A1(G232gat), .A2(G233gat), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n591), .A2(KEYINPUT41), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT100), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n593), .A2(KEYINPUT7), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT7), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n595), .A2(KEYINPUT100), .ZN(new_n596));
  NAND4_X1  g395(.A1(new_n594), .A2(new_n596), .A3(G85gat), .A4(G92gat), .ZN(new_n597));
  INV_X1    g396(.A(G85gat), .ZN(new_n598));
  INV_X1    g397(.A(G92gat), .ZN(new_n599));
  OAI211_X1 g398(.A(KEYINPUT100), .B(new_n595), .C1(new_n598), .C2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(G99gat), .A2(G106gat), .ZN(new_n601));
  AOI22_X1  g400(.A1(KEYINPUT8), .A2(new_n601), .B1(new_n598), .B2(new_n599), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n597), .A2(new_n600), .A3(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(G99gat), .B(G106gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(KEYINPUT101), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n592), .B1(new_n569), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(KEYINPUT102), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT102), .ZN(new_n610));
  OAI211_X1 g409(.A(new_n610), .B(new_n592), .C1(new_n569), .C2(new_n607), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n558), .A2(new_n565), .A3(new_n607), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n609), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(G190gat), .B(G218gat), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT103), .ZN(new_n615));
  OR2_X1    g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n614), .A2(new_n615), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n591), .A2(KEYINPUT41), .ZN(new_n618));
  XOR2_X1   g417(.A(new_n617), .B(new_n618), .Z(new_n619));
  XOR2_X1   g418(.A(G134gat), .B(G162gat), .Z(new_n620));
  XOR2_X1   g419(.A(new_n619), .B(new_n620), .Z(new_n621));
  NAND3_X1  g420(.A1(new_n613), .A2(new_n616), .A3(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n621), .B1(new_n613), .B2(new_n616), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT9), .ZN(new_n626));
  INV_X1    g425(.A(G64gat), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n627), .A2(G57gat), .ZN(new_n628));
  INV_X1    g427(.A(G57gat), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n629), .A2(G64gat), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n626), .B1(new_n628), .B2(new_n630), .ZN(new_n631));
  OAI21_X1  g430(.A(KEYINPUT96), .B1(G71gat), .B2(G78gat), .ZN(new_n632));
  INV_X1    g431(.A(G71gat), .ZN(new_n633));
  INV_X1    g432(.A(G78gat), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n632), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NOR3_X1   g434(.A1(KEYINPUT96), .A2(G71gat), .A3(G78gat), .ZN(new_n636));
  OR3_X1    g435(.A1(new_n631), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n633), .A2(new_n634), .A3(KEYINPUT9), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n638), .B1(new_n633), .B2(new_n634), .ZN(new_n639));
  NAND4_X1  g438(.A1(KEYINPUT97), .A2(KEYINPUT98), .A3(G57gat), .A4(G64gat), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT98), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n627), .B1(new_n641), .B2(new_n629), .ZN(new_n642));
  OR2_X1    g441(.A1(KEYINPUT97), .A2(G57gat), .ZN(new_n643));
  NAND4_X1  g442(.A1(new_n639), .A2(new_n640), .A3(new_n642), .A4(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n637), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT21), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(G231gat), .A2(G233gat), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(G127gat), .B(G155gat), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(KEYINPUT99), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n649), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(G183gat), .B(G211gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n652), .B(new_n653), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n564), .B1(new_n646), .B2(new_n645), .ZN(new_n655));
  XOR2_X1   g454(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n656));
  XNOR2_X1  g455(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XOR2_X1   g456(.A(new_n654), .B(new_n657), .Z(new_n658));
  NOR2_X1   g457(.A1(new_n625), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n605), .B(new_n645), .ZN(new_n660));
  NAND2_X1  g459(.A1(G230gat), .A2(G233gat), .ZN(new_n661));
  OR2_X1    g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(KEYINPUT104), .ZN(new_n663));
  INV_X1    g462(.A(new_n645), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n606), .A2(KEYINPUT10), .A3(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT10), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n660), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n668), .A2(new_n661), .ZN(new_n669));
  XNOR2_X1  g468(.A(G120gat), .B(G148gat), .ZN(new_n670));
  XNOR2_X1  g469(.A(G176gat), .B(G204gat), .ZN(new_n671));
  XOR2_X1   g470(.A(new_n670), .B(new_n671), .Z(new_n672));
  NAND3_X1  g471(.A1(new_n663), .A2(new_n669), .A3(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n663), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n669), .A2(KEYINPUT105), .ZN(new_n675));
  INV_X1    g474(.A(new_n661), .ZN(new_n676));
  AOI211_X1 g475(.A(KEYINPUT105), .B(new_n676), .C1(new_n665), .C2(new_n667), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n674), .B1(new_n675), .B2(new_n678), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n673), .B1(new_n679), .B2(new_n672), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  NAND4_X1  g480(.A1(new_n529), .A2(new_n590), .A3(new_n659), .A4(new_n681), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n682), .A2(new_n484), .ZN(new_n683));
  XOR2_X1   g482(.A(new_n683), .B(G1gat), .Z(G1324gat));
  NOR2_X1   g483(.A1(new_n682), .A2(new_n298), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n685), .A2(new_n563), .ZN(new_n686));
  XOR2_X1   g485(.A(new_n686), .B(KEYINPUT106), .Z(new_n687));
  XOR2_X1   g486(.A(KEYINPUT16), .B(G8gat), .Z(new_n688));
  NAND2_X1  g487(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(KEYINPUT42), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n687), .A2(new_n690), .ZN(G1325gat));
  XNOR2_X1  g490(.A(new_n527), .B(KEYINPUT107), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  OAI21_X1  g492(.A(G15gat), .B1(new_n682), .B2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n526), .ZN(new_n695));
  OR2_X1    g494(.A1(new_n695), .A2(G15gat), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n694), .B1(new_n682), .B2(new_n696), .ZN(G1326gat));
  NOR2_X1   g496(.A1(new_n682), .A2(new_n414), .ZN(new_n698));
  XOR2_X1   g497(.A(KEYINPUT43), .B(G22gat), .Z(new_n699));
  XNOR2_X1  g498(.A(new_n698), .B(new_n699), .ZN(G1327gat));
  INV_X1    g499(.A(new_n625), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n701), .B1(new_n492), .B2(new_n528), .ZN(new_n702));
  INV_X1    g501(.A(new_n658), .ZN(new_n703));
  NOR3_X1   g502(.A1(new_n589), .A2(new_n703), .A3(new_n680), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  NOR3_X1   g504(.A1(new_n705), .A2(G29gat), .A3(new_n484), .ZN(new_n706));
  XNOR2_X1  g505(.A(KEYINPUT108), .B(KEYINPUT45), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n706), .B(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT109), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n709), .B1(new_n623), .B2(new_n624), .ZN(new_n710));
  INV_X1    g509(.A(new_n624), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n711), .A2(KEYINPUT109), .A3(new_n622), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT44), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n529), .A2(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n717), .B1(new_n702), .B2(new_n714), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(new_n704), .ZN(new_n719));
  OAI21_X1  g518(.A(KEYINPUT110), .B1(new_n719), .B2(new_n484), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(G29gat), .ZN(new_n721));
  NOR3_X1   g520(.A1(new_n719), .A2(KEYINPUT110), .A3(new_n484), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n708), .B1(new_n721), .B2(new_n722), .ZN(G1328gat));
  NOR3_X1   g522(.A1(new_n705), .A2(G36gat), .A3(new_n298), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n724), .B(KEYINPUT46), .ZN(new_n725));
  OAI21_X1  g524(.A(G36gat), .B1(new_n719), .B2(new_n298), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(G1329gat));
  OAI21_X1  g526(.A(G43gat), .B1(new_n719), .B2(new_n527), .ZN(new_n728));
  INV_X1    g527(.A(new_n705), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n695), .A2(G43gat), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n728), .A2(KEYINPUT47), .A3(new_n731), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n718), .A2(new_n692), .A3(new_n704), .ZN(new_n733));
  AOI22_X1  g532(.A1(new_n733), .A2(G43gat), .B1(new_n729), .B2(new_n730), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n732), .B1(new_n734), .B2(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g534(.A(new_n714), .B1(new_n529), .B2(new_n625), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n715), .B1(new_n492), .B2(new_n528), .ZN(new_n737));
  OAI211_X1 g536(.A(new_n498), .B(new_n704), .C1(new_n736), .C2(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(new_n544), .ZN(new_n739));
  NOR3_X1   g538(.A1(new_n705), .A2(new_n414), .A3(new_n544), .ZN(new_n740));
  INV_X1    g539(.A(new_n740), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n739), .A2(KEYINPUT48), .A3(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT112), .ZN(new_n743));
  AND3_X1   g542(.A1(new_n738), .A2(new_n743), .A3(new_n544), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n743), .B1(new_n738), .B2(new_n544), .ZN(new_n745));
  NOR3_X1   g544(.A1(new_n744), .A2(new_n745), .A3(new_n740), .ZN(new_n746));
  XOR2_X1   g545(.A(KEYINPUT111), .B(KEYINPUT48), .Z(new_n747));
  OAI21_X1  g546(.A(new_n742), .B1(new_n746), .B2(new_n747), .ZN(G1331gat));
  AND3_X1   g547(.A1(new_n529), .A2(new_n589), .A3(new_n659), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(new_n680), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n750), .A2(new_n484), .ZN(new_n751));
  XOR2_X1   g550(.A(KEYINPUT97), .B(G57gat), .Z(new_n752));
  XNOR2_X1  g551(.A(new_n751), .B(new_n752), .ZN(G1332gat));
  NOR2_X1   g552(.A1(new_n750), .A2(new_n298), .ZN(new_n754));
  NOR2_X1   g553(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n755));
  AND2_X1   g554(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n754), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n757), .B1(new_n754), .B2(new_n755), .ZN(G1333gat));
  NOR2_X1   g557(.A1(new_n695), .A2(new_n681), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n749), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(KEYINPUT113), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT113), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n749), .A2(new_n762), .A3(new_n759), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n761), .A2(new_n633), .A3(new_n763), .ZN(new_n764));
  NAND4_X1  g563(.A1(new_n749), .A2(G71gat), .A3(new_n680), .A4(new_n692), .ZN(new_n765));
  XNOR2_X1  g564(.A(KEYINPUT114), .B(KEYINPUT50), .ZN(new_n766));
  AND3_X1   g565(.A1(new_n764), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n766), .B1(new_n764), .B2(new_n765), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n767), .A2(new_n768), .ZN(G1334gat));
  NOR2_X1   g568(.A1(new_n750), .A2(new_n414), .ZN(new_n770));
  XNOR2_X1  g569(.A(KEYINPUT115), .B(G78gat), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n770), .B(new_n771), .ZN(G1335gat));
  NOR2_X1   g571(.A1(new_n590), .A2(new_n703), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT51), .ZN(new_n774));
  AND2_X1   g573(.A1(new_n774), .A2(KEYINPUT116), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n774), .A2(KEYINPUT116), .ZN(new_n776));
  OAI211_X1 g575(.A(new_n702), .B(new_n773), .C1(new_n775), .C2(new_n776), .ZN(new_n777));
  AND2_X1   g576(.A1(new_n702), .A2(new_n773), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n777), .B1(new_n778), .B2(new_n776), .ZN(new_n779));
  INV_X1    g578(.A(new_n484), .ZN(new_n780));
  NAND4_X1  g579(.A1(new_n779), .A2(new_n598), .A3(new_n780), .A4(new_n680), .ZN(new_n781));
  NOR3_X1   g580(.A1(new_n590), .A2(new_n703), .A3(new_n681), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n718), .A2(new_n780), .A3(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n781), .B1(new_n784), .B2(new_n598), .ZN(G1336gat));
  NOR3_X1   g584(.A1(new_n681), .A2(new_n298), .A3(G92gat), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT117), .ZN(new_n787));
  AOI22_X1  g586(.A1(new_n779), .A2(new_n786), .B1(new_n787), .B2(KEYINPUT52), .ZN(new_n788));
  OR2_X1    g587(.A1(new_n787), .A2(KEYINPUT52), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n718), .A2(new_n782), .ZN(new_n790));
  OAI21_X1  g589(.A(G92gat), .B1(new_n790), .B2(new_n298), .ZN(new_n791));
  AND3_X1   g590(.A1(new_n788), .A2(new_n789), .A3(new_n791), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n789), .B1(new_n788), .B2(new_n791), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n792), .A2(new_n793), .ZN(G1337gat));
  OAI21_X1  g593(.A(G99gat), .B1(new_n790), .B2(new_n693), .ZN(new_n795));
  INV_X1    g594(.A(G99gat), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n779), .A2(new_n796), .A3(new_n759), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n795), .A2(new_n797), .ZN(G1338gat));
  OAI21_X1  g597(.A(G106gat), .B1(new_n790), .B2(new_n414), .ZN(new_n799));
  NOR3_X1   g598(.A1(new_n681), .A2(G106gat), .A3(new_n414), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n779), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(KEYINPUT53), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT53), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n799), .A2(new_n804), .A3(new_n801), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n803), .A2(new_n805), .ZN(G1339gat));
  NAND3_X1  g605(.A1(new_n659), .A2(new_n589), .A3(new_n681), .ZN(new_n807));
  INV_X1    g606(.A(new_n807), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n575), .A2(new_n576), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n567), .B1(new_n566), .B2(new_n570), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n582), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n585), .A2(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT55), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n676), .B1(new_n665), .B2(new_n667), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT105), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n816), .A2(new_n677), .A3(KEYINPUT54), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n665), .A2(new_n676), .A3(new_n667), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n669), .A2(KEYINPUT54), .A3(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(new_n672), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n813), .B1(new_n817), .B2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT54), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n678), .A2(new_n675), .A3(new_n823), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n824), .A2(KEYINPUT55), .A3(new_n820), .A4(new_n819), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n822), .A2(new_n825), .A3(new_n673), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n812), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n713), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n573), .A2(new_n574), .A3(new_n577), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(new_n583), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n826), .B1(new_n830), .B2(new_n585), .ZN(new_n831));
  AND3_X1   g630(.A1(new_n680), .A2(new_n585), .A3(new_n811), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n828), .B1(new_n833), .B2(new_n713), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n808), .B1(new_n834), .B2(new_n658), .ZN(new_n835));
  NOR4_X1   g634(.A1(new_n835), .A2(new_n484), .A3(new_n297), .A4(new_n417), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(new_n590), .ZN(new_n837));
  XNOR2_X1  g636(.A(new_n837), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g637(.A1(new_n836), .A2(new_n680), .ZN(new_n839));
  XNOR2_X1  g638(.A(new_n839), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g639(.A1(new_n836), .A2(new_n703), .ZN(new_n841));
  XOR2_X1   g640(.A(KEYINPUT118), .B(G127gat), .Z(new_n842));
  XNOR2_X1  g641(.A(new_n841), .B(new_n842), .ZN(G1342gat));
  INV_X1    g642(.A(KEYINPUT56), .ZN(new_n844));
  OAI211_X1 g643(.A(new_n836), .B(new_n625), .C1(new_n844), .C2(new_n308), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n308), .ZN(new_n846));
  XNOR2_X1  g645(.A(new_n845), .B(new_n846), .ZN(G1343gat));
  OR2_X1    g646(.A1(KEYINPUT121), .A2(KEYINPUT58), .ZN(new_n848));
  NAND2_X1  g647(.A1(KEYINPUT121), .A2(KEYINPUT58), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n484), .A2(new_n297), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(new_n527), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT57), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n414), .A2(new_n852), .ZN(new_n853));
  OAI21_X1  g652(.A(KEYINPUT119), .B1(new_n831), .B2(new_n832), .ZN(new_n854));
  AND3_X1   g653(.A1(new_n822), .A2(new_n825), .A3(new_n673), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n855), .B1(new_n586), .B2(new_n588), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT119), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n680), .A2(new_n585), .A3(new_n811), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n856), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n854), .A2(new_n859), .A3(new_n701), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n703), .B1(new_n860), .B2(new_n828), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n853), .B1(new_n861), .B2(new_n808), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n852), .B1(new_n835), .B2(new_n414), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n851), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n362), .B1(new_n864), .B2(new_n590), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n713), .B1(new_n856), .B2(new_n858), .ZN(new_n866));
  AND2_X1   g665(.A1(new_n713), .A2(new_n827), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n658), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(new_n807), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n869), .A2(new_n498), .A3(new_n693), .ZN(new_n870));
  INV_X1    g669(.A(new_n850), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n590), .A2(new_n362), .ZN(new_n872));
  XNOR2_X1  g671(.A(new_n872), .B(KEYINPUT120), .ZN(new_n873));
  NOR3_X1   g672(.A1(new_n870), .A2(new_n871), .A3(new_n873), .ZN(new_n874));
  OAI211_X1 g673(.A(new_n848), .B(new_n849), .C1(new_n865), .C2(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n862), .A2(new_n863), .ZN(new_n876));
  INV_X1    g675(.A(new_n851), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n876), .A2(new_n590), .A3(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(G141gat), .ZN(new_n879));
  INV_X1    g678(.A(new_n874), .ZN(new_n880));
  NAND4_X1  g679(.A1(new_n879), .A2(KEYINPUT121), .A3(KEYINPUT58), .A4(new_n880), .ZN(new_n881));
  AND2_X1   g680(.A1(new_n875), .A2(new_n881), .ZN(G1344gat));
  INV_X1    g681(.A(KEYINPUT59), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n864), .A2(new_n883), .A3(new_n680), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n870), .A2(new_n871), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n883), .B1(new_n885), .B2(new_n680), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n358), .A2(new_n360), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n827), .A2(new_n625), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n703), .B1(new_n860), .B2(new_n888), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n498), .B1(new_n889), .B2(new_n808), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(new_n852), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n869), .A2(new_n853), .ZN(new_n892));
  AOI211_X1 g691(.A(new_n681), .B(new_n851), .C1(new_n891), .C2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n894));
  OAI221_X1 g693(.A(new_n884), .B1(new_n886), .B2(new_n887), .C1(new_n893), .C2(new_n894), .ZN(G1345gat));
  INV_X1    g694(.A(new_n864), .ZN(new_n896));
  OAI21_X1  g695(.A(G155gat), .B1(new_n896), .B2(new_n658), .ZN(new_n897));
  INV_X1    g696(.A(G155gat), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n885), .A2(new_n898), .A3(new_n703), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n897), .A2(new_n899), .ZN(G1346gat));
  INV_X1    g699(.A(new_n713), .ZN(new_n901));
  OAI21_X1  g700(.A(G162gat), .B1(new_n896), .B2(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(G162gat), .ZN(new_n903));
  NAND4_X1  g702(.A1(new_n780), .A2(new_n903), .A3(new_n298), .A4(new_n625), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n902), .B1(new_n870), .B2(new_n904), .ZN(G1347gat));
  NOR2_X1   g704(.A1(new_n298), .A2(new_n417), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n869), .A2(new_n484), .A3(new_n906), .ZN(new_n907));
  INV_X1    g706(.A(new_n907), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(new_n590), .ZN(new_n909));
  XNOR2_X1  g708(.A(new_n909), .B(G169gat), .ZN(G1348gat));
  AOI21_X1  g709(.A(G176gat), .B1(new_n908), .B2(new_n680), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n835), .A2(new_n780), .ZN(new_n912));
  AND4_X1   g711(.A1(G176gat), .A2(new_n759), .A3(new_n414), .A4(new_n297), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n911), .B1(new_n912), .B2(new_n913), .ZN(G1349gat));
  INV_X1    g713(.A(KEYINPUT122), .ZN(new_n915));
  OAI22_X1  g714(.A1(new_n907), .A2(new_n658), .B1(new_n915), .B2(new_n212), .ZN(new_n916));
  AOI22_X1  g715(.A1(new_n227), .A2(new_n229), .B1(new_n915), .B2(G183gat), .ZN(new_n917));
  NAND4_X1  g716(.A1(new_n912), .A2(new_n703), .A3(new_n906), .A4(new_n917), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  XOR2_X1   g718(.A(KEYINPUT123), .B(KEYINPUT60), .Z(new_n920));
  NAND2_X1  g719(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT124), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n919), .A2(KEYINPUT124), .A3(new_n920), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT60), .ZN(new_n925));
  OAI211_X1 g724(.A(new_n923), .B(new_n924), .C1(new_n925), .C2(new_n919), .ZN(G1350gat));
  NAND3_X1  g725(.A1(new_n908), .A2(new_n228), .A3(new_n713), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n912), .A2(new_n625), .A3(new_n906), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT61), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n928), .A2(new_n929), .A3(G190gat), .ZN(new_n930));
  INV_X1    g729(.A(new_n930), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n929), .B1(new_n928), .B2(G190gat), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n927), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n933), .A2(KEYINPUT125), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT125), .ZN(new_n935));
  OAI211_X1 g734(.A(new_n935), .B(new_n927), .C1(new_n931), .C2(new_n932), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n934), .A2(new_n936), .ZN(G1351gat));
  NOR3_X1   g736(.A1(new_n692), .A2(new_n414), .A3(new_n298), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n912), .A2(new_n938), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT126), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n939), .B(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(new_n590), .ZN(new_n942));
  NOR3_X1   g741(.A1(new_n692), .A2(new_n780), .A3(new_n298), .ZN(new_n943));
  INV_X1    g742(.A(new_n943), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n944), .B1(new_n891), .B2(new_n892), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n589), .A2(new_n259), .ZN(new_n946));
  AOI22_X1  g745(.A1(new_n942), .A2(new_n259), .B1(new_n945), .B2(new_n946), .ZN(G1352gat));
  INV_X1    g746(.A(KEYINPUT127), .ZN(new_n948));
  AOI211_X1 g747(.A(G204gat), .B(new_n681), .C1(new_n948), .C2(KEYINPUT62), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n912), .A2(new_n938), .A3(new_n949), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n948), .A2(KEYINPUT62), .ZN(new_n951));
  XNOR2_X1  g750(.A(new_n950), .B(new_n951), .ZN(new_n952));
  AND2_X1   g751(.A1(new_n945), .A2(new_n680), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n952), .B1(new_n953), .B2(new_n260), .ZN(G1353gat));
  INV_X1    g753(.A(G211gat), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n941), .A2(new_n955), .A3(new_n703), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT63), .ZN(new_n957));
  AOI211_X1 g756(.A(new_n957), .B(new_n955), .C1(new_n945), .C2(new_n703), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n891), .A2(new_n892), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n959), .A2(new_n703), .A3(new_n943), .ZN(new_n960));
  AOI21_X1  g759(.A(KEYINPUT63), .B1(new_n960), .B2(G211gat), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n956), .B1(new_n958), .B2(new_n961), .ZN(G1354gat));
  INV_X1    g761(.A(G218gat), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n941), .A2(new_n963), .A3(new_n713), .ZN(new_n964));
  AND2_X1   g763(.A1(new_n945), .A2(new_n625), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n964), .B1(new_n963), .B2(new_n965), .ZN(G1355gat));
endmodule


