

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778;

  NOR2_X1 U370 ( .A1(n453), .A2(n404), .ZN(n599) );
  NAND2_X1 U371 ( .A1(n703), .A2(n702), .ZN(n699) );
  BUF_X1 U372 ( .A(G146), .Z(n349) );
  XNOR2_X1 U373 ( .A(n536), .B(n435), .ZN(n369) );
  XNOR2_X1 U374 ( .A(n495), .B(G125), .ZN(n544) );
  XNOR2_X2 U375 ( .A(n386), .B(n387), .ZN(n661) );
  NAND2_X2 U376 ( .A1(n446), .A2(n443), .ZN(n620) );
  NAND2_X2 U377 ( .A1(n420), .A2(n419), .ZN(n442) );
  XNOR2_X2 U378 ( .A(n583), .B(n584), .ZN(n703) );
  XNOR2_X2 U379 ( .A(n350), .B(n654), .ZN(n725) );
  NAND2_X1 U380 ( .A1(n403), .A2(n506), .ZN(n350) );
  NAND2_X1 U381 ( .A1(n618), .A2(n686), .ZN(n598) );
  INV_X1 U382 ( .A(G953), .ZN(n765) );
  XNOR2_X2 U383 ( .A(n418), .B(G143), .ZN(n536) );
  XNOR2_X2 U384 ( .A(n414), .B(KEYINPUT22), .ZN(n648) );
  INV_X1 U385 ( .A(n628), .ZN(n649) );
  INV_X1 U386 ( .A(G472), .ZN(n563) );
  INV_X1 U387 ( .A(G469), .ZN(n509) );
  AND2_X1 U388 ( .A1(n422), .A2(n421), .ZN(n420) );
  AND2_X1 U389 ( .A1(n448), .A2(n447), .ZN(n446) );
  AND2_X1 U390 ( .A1(n488), .A2(n431), .ZN(n430) );
  NAND2_X1 U391 ( .A1(n432), .A2(n352), .ZN(n488) );
  NAND2_X1 U392 ( .A1(n383), .A2(n379), .ZN(n606) );
  XNOR2_X1 U393 ( .A(n482), .B(n478), .ZN(n368) );
  XOR2_X1 U394 ( .A(G113), .B(G104), .Z(n541) );
  NAND2_X1 U395 ( .A1(n460), .A2(n461), .ZN(n367) );
  XNOR2_X2 U396 ( .A(n391), .B(n390), .ZN(n695) );
  XOR2_X1 U397 ( .A(G101), .B(KEYINPUT66), .Z(n558) );
  XNOR2_X1 U398 ( .A(n369), .B(n433), .ZN(n762) );
  XNOR2_X1 U399 ( .A(n562), .B(n434), .ZN(n433) );
  XNOR2_X1 U400 ( .A(n512), .B(G137), .ZN(n434) );
  INV_X1 U401 ( .A(KEYINPUT4), .ZN(n512) );
  XNOR2_X1 U402 ( .A(n558), .B(n535), .ZN(n568) );
  INV_X1 U403 ( .A(G110), .ZN(n535) );
  XNOR2_X1 U404 ( .A(n500), .B(G475), .ZN(n499) );
  INV_X1 U405 ( .A(KEYINPUT13), .ZN(n500) );
  INV_X1 U406 ( .A(KEYINPUT19), .ZN(n597) );
  NAND2_X1 U407 ( .A1(n607), .A2(n606), .ZN(n629) );
  AND2_X1 U408 ( .A1(n492), .A2(n773), .ZN(n440) );
  AND2_X1 U409 ( .A1(n604), .A2(n600), .ZN(n492) );
  INV_X1 U410 ( .A(KEYINPUT70), .ZN(n493) );
  XNOR2_X1 U411 ( .A(n497), .B(KEYINPUT83), .ZN(n644) );
  NOR2_X1 U412 ( .A1(G953), .A2(G237), .ZN(n555) );
  XNOR2_X1 U413 ( .A(n558), .B(n560), .ZN(n389) );
  XOR2_X1 U414 ( .A(KEYINPUT5), .B(KEYINPUT73), .Z(n560) );
  XOR2_X1 U415 ( .A(KEYINPUT72), .B(G113), .Z(n557) );
  AND2_X1 U416 ( .A1(n657), .A2(n505), .ZN(n476) );
  NAND2_X1 U417 ( .A1(n504), .A2(n473), .ZN(n472) );
  NAND2_X1 U418 ( .A1(KEYINPUT64), .A2(KEYINPUT2), .ZN(n473) );
  XNOR2_X1 U419 ( .A(n540), .B(KEYINPUT90), .ZN(n486) );
  AND2_X1 U420 ( .A1(n727), .A2(n726), .ZN(n460) );
  INV_X1 U421 ( .A(KEYINPUT39), .ZN(n444) );
  NAND2_X1 U422 ( .A1(n608), .A2(KEYINPUT39), .ZN(n447) );
  INV_X1 U423 ( .A(KEYINPUT33), .ZN(n390) );
  XNOR2_X1 U424 ( .A(n480), .B(n479), .ZN(n754) );
  XNOR2_X1 U425 ( .A(n541), .B(KEYINPUT16), .ZN(n479) );
  INV_X1 U426 ( .A(n542), .ZN(n481) );
  XNOR2_X1 U427 ( .A(n530), .B(n374), .ZN(n580) );
  INV_X1 U428 ( .A(KEYINPUT84), .ZN(n374) );
  XNOR2_X1 U429 ( .A(n578), .B(n463), .ZN(n462) );
  INV_X1 U430 ( .A(KEYINPUT23), .ZN(n463) );
  XNOR2_X1 U431 ( .A(G128), .B(KEYINPUT24), .ZN(n578) );
  XNOR2_X1 U432 ( .A(n494), .B(n522), .ZN(n761) );
  XOR2_X1 U433 ( .A(KEYINPUT68), .B(KEYINPUT10), .Z(n522) );
  XNOR2_X1 U434 ( .A(n544), .B(G140), .ZN(n494) );
  XNOR2_X1 U435 ( .A(G116), .B(KEYINPUT7), .ZN(n531) );
  XOR2_X1 U436 ( .A(KEYINPUT9), .B(KEYINPUT102), .Z(n532) );
  NAND2_X1 U437 ( .A1(n580), .A2(G217), .ZN(n373) );
  XNOR2_X1 U438 ( .A(n570), .B(n459), .ZN(n511) );
  XNOR2_X1 U439 ( .A(n354), .B(n569), .ZN(n459) );
  XNOR2_X1 U440 ( .A(n595), .B(n416), .ZN(n596) );
  INV_X1 U441 ( .A(KEYINPUT28), .ZN(n416) );
  AND2_X1 U442 ( .A1(n594), .A2(n632), .ZN(n595) );
  AND2_X1 U443 ( .A1(n613), .A2(n377), .ZN(n376) );
  NOR2_X1 U444 ( .A1(n641), .A2(n359), .ZN(n423) );
  INV_X1 U445 ( .A(KEYINPUT76), .ZN(n370) );
  BUF_X1 U446 ( .A(n698), .Z(n464) );
  NAND2_X1 U447 ( .A1(n467), .A2(n465), .ZN(n585) );
  XNOR2_X1 U448 ( .A(n567), .B(n456), .ZN(n467) );
  AND2_X1 U449 ( .A1(n385), .A2(n384), .ZN(n383) );
  NAND2_X1 U450 ( .A1(n499), .A2(G902), .ZN(n384) );
  XNOR2_X1 U451 ( .A(n534), .B(n501), .ZN(n607) );
  XNOR2_X1 U452 ( .A(n502), .B(KEYINPUT104), .ZN(n501) );
  INV_X1 U453 ( .A(G478), .ZN(n502) );
  NAND2_X1 U454 ( .A1(n429), .A2(n491), .ZN(n490) );
  NAND2_X1 U455 ( .A1(n627), .A2(n357), .ZN(n491) );
  OR2_X1 U456 ( .A1(n619), .A2(n676), .ZN(n497) );
  NOR2_X1 U457 ( .A1(n397), .A2(n396), .ZN(n395) );
  NAND2_X1 U458 ( .A1(n775), .A2(KEYINPUT44), .ZN(n396) );
  XNOR2_X1 U459 ( .A(n513), .B(G131), .ZN(n562) );
  INV_X1 U460 ( .A(KEYINPUT69), .ZN(n513) );
  NAND2_X1 U461 ( .A1(G234), .A2(G237), .ZN(n548) );
  XNOR2_X1 U462 ( .A(n415), .B(n436), .ZN(n727) );
  INV_X1 U463 ( .A(KEYINPUT48), .ZN(n436) );
  AND2_X1 U464 ( .A1(n441), .A2(n440), .ZN(n439) );
  INV_X1 U465 ( .A(G146), .ZN(n495) );
  XOR2_X1 U466 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n524) );
  XNOR2_X1 U467 ( .A(G143), .B(G122), .ZN(n523) );
  XNOR2_X1 U468 ( .A(KEYINPUT98), .B(KEYINPUT101), .ZN(n518) );
  XOR2_X1 U469 ( .A(KEYINPUT100), .B(KEYINPUT99), .Z(n519) );
  NOR2_X1 U470 ( .A1(G902), .A2(G237), .ZN(n545) );
  INV_X1 U471 ( .A(KEYINPUT30), .ZN(n456) );
  INV_X1 U472 ( .A(n590), .ZN(n466) );
  NAND2_X1 U473 ( .A1(n382), .A2(n381), .ZN(n380) );
  INV_X1 U474 ( .A(G902), .ZN(n381) );
  BUF_X1 U475 ( .A(n589), .Z(n706) );
  XNOR2_X1 U476 ( .A(n388), .B(n561), .ZN(n387) );
  XNOR2_X1 U477 ( .A(n389), .B(n559), .ZN(n388) );
  INV_X1 U478 ( .A(KEYINPUT45), .ZN(n654) );
  NAND2_X1 U479 ( .A1(n474), .A2(n472), .ZN(n471) );
  NAND2_X1 U480 ( .A1(n656), .A2(KEYINPUT64), .ZN(n474) );
  XNOR2_X1 U481 ( .A(n568), .B(n539), .ZN(n483) );
  AND2_X1 U482 ( .A1(n367), .A2(n405), .ZN(n724) );
  INV_X1 U483 ( .A(KEYINPUT85), .ZN(n405) );
  NAND2_X1 U484 ( .A1(n445), .A2(n356), .ZN(n443) );
  BUF_X1 U485 ( .A(n626), .Z(n404) );
  AND2_X1 U486 ( .A1(n630), .A2(n702), .ZN(n431) );
  XNOR2_X1 U487 ( .A(n577), .B(n462), .ZN(n579) );
  XNOR2_X1 U488 ( .A(n372), .B(n371), .ZN(n740) );
  XNOR2_X1 U489 ( .A(n373), .B(n514), .ZN(n372) );
  INV_X1 U490 ( .A(KEYINPUT122), .ZN(n457) );
  XNOR2_X1 U491 ( .A(n376), .B(n592), .ZN(n375) );
  NAND2_X1 U492 ( .A1(n424), .A2(n423), .ZN(n419) );
  INV_X1 U493 ( .A(n678), .ZN(n676) );
  NOR2_X1 U494 ( .A1(n605), .A2(n629), .ZN(n586) );
  AND2_X1 U495 ( .A1(n607), .A2(n498), .ZN(n672) );
  INV_X1 U496 ( .A(n606), .ZN(n498) );
  NAND2_X1 U497 ( .A1(n378), .A2(n606), .ZN(n678) );
  INV_X1 U498 ( .A(n607), .ZN(n378) );
  INV_X1 U499 ( .A(KEYINPUT60), .ZN(n449) );
  INV_X1 U500 ( .A(KEYINPUT124), .ZN(n407) );
  INV_X1 U501 ( .A(KEYINPUT56), .ZN(n409) );
  XNOR2_X1 U502 ( .A(KEYINPUT53), .B(KEYINPUT123), .ZN(n468) );
  XNOR2_X1 U503 ( .A(n634), .B(G119), .ZN(G21) );
  AND2_X1 U504 ( .A1(n641), .A2(n359), .ZN(n351) );
  NOR2_X1 U505 ( .A1(n627), .A2(n357), .ZN(n352) );
  AND2_X1 U506 ( .A1(G210), .A2(n566), .ZN(n353) );
  XNOR2_X1 U507 ( .A(n706), .B(KEYINPUT6), .ZN(n628) );
  XNOR2_X1 U508 ( .A(G104), .B(G140), .ZN(n354) );
  XOR2_X1 U509 ( .A(n629), .B(n370), .Z(n355) );
  AND2_X1 U510 ( .A1(n687), .A2(n444), .ZN(n356) );
  XOR2_X1 U511 ( .A(KEYINPUT0), .B(KEYINPUT65), .Z(n357) );
  XNOR2_X1 U512 ( .A(KEYINPUT78), .B(KEYINPUT32), .ZN(n358) );
  XOR2_X1 U513 ( .A(KEYINPUT34), .B(KEYINPUT77), .Z(n359) );
  XNOR2_X1 U514 ( .A(n737), .B(KEYINPUT59), .ZN(n360) );
  XOR2_X1 U515 ( .A(n735), .B(n734), .Z(n361) );
  XNOR2_X1 U516 ( .A(n659), .B(n658), .ZN(n362) );
  XOR2_X1 U517 ( .A(n661), .B(KEYINPUT62), .Z(n363) );
  INV_X1 U518 ( .A(n656), .ZN(n504) );
  XNOR2_X1 U519 ( .A(G902), .B(KEYINPUT15), .ZN(n656) );
  XOR2_X1 U520 ( .A(KEYINPUT86), .B(KEYINPUT46), .Z(n364) );
  AND2_X1 U521 ( .A1(n504), .A2(KEYINPUT64), .ZN(n365) );
  INV_X1 U522 ( .A(n746), .ZN(n451) );
  XOR2_X1 U523 ( .A(n663), .B(KEYINPUT63), .Z(n366) );
  NAND2_X1 U524 ( .A1(n367), .A2(n476), .ZN(n475) );
  INV_X1 U525 ( .A(n367), .ZN(n723) );
  NAND2_X1 U526 ( .A1(n368), .A2(n656), .ZN(n425) );
  XNOR2_X1 U527 ( .A(n368), .B(KEYINPUT82), .ZN(n658) );
  XNOR2_X1 U528 ( .A(n369), .B(n542), .ZN(n371) );
  NOR2_X1 U529 ( .A1(n375), .A2(n464), .ZN(n593) );
  INV_X1 U530 ( .A(n598), .ZN(n377) );
  OR2_X1 U531 ( .A1(n737), .A2(n380), .ZN(n379) );
  INV_X1 U532 ( .A(n499), .ZN(n382) );
  NAND2_X1 U533 ( .A1(n737), .A2(n499), .ZN(n385) );
  XNOR2_X1 U534 ( .A(n511), .B(n386), .ZN(n735) );
  XNOR2_X2 U535 ( .A(n762), .B(n349), .ZN(n386) );
  INV_X1 U536 ( .A(n393), .ZN(n640) );
  NAND2_X1 U537 ( .A1(n392), .A2(n649), .ZN(n391) );
  XNOR2_X1 U538 ( .A(n393), .B(KEYINPUT109), .ZN(n392) );
  OR2_X2 U539 ( .A1(n698), .A2(n699), .ZN(n393) );
  NAND2_X1 U540 ( .A1(n399), .A2(n394), .ZN(n403) );
  NAND2_X1 U541 ( .A1(n398), .A2(n395), .ZN(n394) );
  INV_X1 U542 ( .A(n634), .ZN(n397) );
  INV_X1 U543 ( .A(n774), .ZN(n398) );
  AND2_X1 U544 ( .A1(n402), .A2(n400), .ZN(n399) );
  NAND2_X1 U545 ( .A1(n401), .A2(n508), .ZN(n400) );
  NAND2_X1 U546 ( .A1(n634), .A2(n775), .ZN(n401) );
  NAND2_X1 U547 ( .A1(n774), .A2(n508), .ZN(n402) );
  NAND2_X1 U548 ( .A1(n428), .A2(n631), .ZN(n426) );
  XNOR2_X1 U549 ( .A(n406), .B(n366), .ZN(G57) );
  NAND2_X1 U550 ( .A1(n412), .A2(n451), .ZN(n406) );
  XNOR2_X1 U551 ( .A(n408), .B(n407), .ZN(G54) );
  NAND2_X1 U552 ( .A1(n413), .A2(n451), .ZN(n408) );
  XNOR2_X1 U553 ( .A(n410), .B(n409), .ZN(G51) );
  NAND2_X1 U554 ( .A1(n411), .A2(n451), .ZN(n410) );
  XNOR2_X1 U555 ( .A(n438), .B(n364), .ZN(n437) );
  NAND2_X1 U556 ( .A1(n437), .A2(n439), .ZN(n415) );
  XNOR2_X1 U557 ( .A(n660), .B(n362), .ZN(n411) );
  XNOR2_X1 U558 ( .A(n662), .B(n363), .ZN(n412) );
  XNOR2_X1 U559 ( .A(n736), .B(n361), .ZN(n413) );
  NAND2_X1 U560 ( .A1(n430), .A2(n489), .ZN(n414) );
  INV_X1 U561 ( .A(n778), .ZN(n507) );
  XNOR2_X1 U562 ( .A(n484), .B(n483), .ZN(n482) );
  INV_X1 U563 ( .A(n490), .ZN(n489) );
  NOR2_X1 U564 ( .A1(n417), .A2(n647), .ZN(n636) );
  XNOR2_X1 U565 ( .A(n417), .B(KEYINPUT1), .ZN(n698) );
  OR2_X1 U566 ( .A1(n596), .A2(n417), .ZN(n453) );
  XNOR2_X2 U567 ( .A(n510), .B(n509), .ZN(n417) );
  XNOR2_X2 U568 ( .A(G128), .B(KEYINPUT80), .ZN(n418) );
  NOR2_X1 U569 ( .A1(n351), .A2(n355), .ZN(n421) );
  NAND2_X1 U570 ( .A1(n695), .A2(n359), .ZN(n422) );
  INV_X1 U571 ( .A(n695), .ZN(n424) );
  XNOR2_X2 U572 ( .A(n425), .B(n353), .ZN(n618) );
  XNOR2_X2 U573 ( .A(n426), .B(n358), .ZN(n634) );
  XNOR2_X2 U574 ( .A(n427), .B(KEYINPUT108), .ZN(n775) );
  NAND2_X1 U575 ( .A1(n428), .A2(n633), .ZN(n427) );
  NOR2_X2 U576 ( .A1(n648), .A2(n703), .ZN(n428) );
  NAND2_X1 U577 ( .A1(n626), .A2(n357), .ZN(n429) );
  INV_X1 U578 ( .A(n626), .ZN(n432) );
  INV_X1 U579 ( .A(G134), .ZN(n435) );
  NAND2_X1 U580 ( .A1(n776), .A2(n777), .ZN(n438) );
  XNOR2_X1 U581 ( .A(n603), .B(n493), .ZN(n441) );
  XNOR2_X2 U582 ( .A(n442), .B(KEYINPUT35), .ZN(n774) );
  INV_X1 U583 ( .A(n605), .ZN(n445) );
  NAND2_X1 U584 ( .A1(n605), .A2(KEYINPUT39), .ZN(n448) );
  NAND2_X1 U585 ( .A1(n620), .A2(n676), .ZN(n454) );
  NAND2_X2 U586 ( .A1(n470), .A2(n469), .ZN(n477) );
  XNOR2_X1 U587 ( .A(n450), .B(n449), .ZN(G60) );
  NAND2_X1 U588 ( .A1(n452), .A2(n451), .ZN(n450) );
  XNOR2_X1 U589 ( .A(n738), .B(n360), .ZN(n452) );
  NAND2_X1 U590 ( .A1(n731), .A2(n732), .ZN(n458) );
  NAND2_X1 U591 ( .A1(n723), .A2(KEYINPUT2), .ZN(n503) );
  XNOR2_X1 U592 ( .A(n458), .B(n457), .ZN(n733) );
  NOR2_X1 U593 ( .A1(n646), .A2(n507), .ZN(n506) );
  OR2_X2 U594 ( .A1(n735), .A2(G902), .ZN(n510) );
  INV_X2 U595 ( .A(n671), .ZN(n601) );
  INV_X1 U596 ( .A(n453), .ZN(n610) );
  XNOR2_X2 U597 ( .A(n454), .B(KEYINPUT40), .ZN(n776) );
  XNOR2_X1 U598 ( .A(n455), .B(n468), .ZN(G75) );
  NAND2_X1 U599 ( .A1(n733), .A2(n765), .ZN(n455) );
  INV_X1 U600 ( .A(n725), .ZN(n461) );
  NOR2_X1 U601 ( .A1(G902), .A2(n744), .ZN(n583) );
  AND2_X1 U602 ( .A1(n636), .A2(n466), .ZN(n465) );
  NAND2_X1 U603 ( .A1(n723), .A2(n365), .ZN(n469) );
  AND2_X2 U604 ( .A1(n475), .A2(n471), .ZN(n470) );
  AND2_X4 U605 ( .A1(n477), .A2(n503), .ZN(n742) );
  INV_X1 U606 ( .A(n754), .ZN(n478) );
  XNOR2_X1 U607 ( .A(n559), .B(n481), .ZN(n480) );
  XNOR2_X1 U608 ( .A(n485), .B(n515), .ZN(n484) );
  XNOR2_X1 U609 ( .A(n536), .B(n486), .ZN(n485) );
  NAND2_X1 U610 ( .A1(n489), .A2(n488), .ZN(n641) );
  NOR2_X1 U611 ( .A1(n490), .A2(n487), .ZN(n635) );
  NAND2_X1 U612 ( .A1(n488), .A2(n702), .ZN(n487) );
  XNOR2_X2 U613 ( .A(n598), .B(n597), .ZN(n626) );
  INV_X1 U614 ( .A(n497), .ZN(n692) );
  NAND2_X1 U615 ( .A1(n496), .A2(n601), .ZN(n602) );
  INV_X1 U616 ( .A(n644), .ZN(n496) );
  INV_X1 U617 ( .A(KEYINPUT2), .ZN(n505) );
  INV_X1 U618 ( .A(KEYINPUT44), .ZN(n508) );
  NAND2_X1 U619 ( .A1(n742), .A2(G210), .ZN(n660) );
  XNOR2_X2 U620 ( .A(n585), .B(KEYINPUT74), .ZN(n605) );
  XNOR2_X1 U621 ( .A(n533), .B(KEYINPUT103), .ZN(n514) );
  XOR2_X1 U622 ( .A(KEYINPUT4), .B(n544), .Z(n515) );
  NOR2_X1 U623 ( .A1(G952), .A2(n765), .ZN(n746) );
  XOR2_X1 U624 ( .A(n562), .B(n541), .Z(n517) );
  NAND2_X1 U625 ( .A1(G214), .A2(n555), .ZN(n516) );
  XNOR2_X1 U626 ( .A(n517), .B(n516), .ZN(n521) );
  XNOR2_X1 U627 ( .A(n519), .B(n518), .ZN(n520) );
  XOR2_X1 U628 ( .A(n521), .B(n520), .Z(n527) );
  XNOR2_X1 U629 ( .A(n524), .B(n523), .ZN(n525) );
  XNOR2_X1 U630 ( .A(n761), .B(n525), .ZN(n526) );
  XNOR2_X1 U631 ( .A(n527), .B(n526), .ZN(n737) );
  XOR2_X1 U632 ( .A(KEYINPUT8), .B(KEYINPUT67), .Z(n529) );
  NAND2_X1 U633 ( .A1(G234), .A2(n765), .ZN(n528) );
  XNOR2_X1 U634 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U635 ( .A(n532), .B(n531), .ZN(n533) );
  XOR2_X1 U636 ( .A(G107), .B(G122), .Z(n542) );
  NOR2_X1 U637 ( .A1(G902), .A2(n740), .ZN(n534) );
  XOR2_X1 U638 ( .A(KEYINPUT105), .B(n672), .Z(n619) );
  NAND2_X1 U639 ( .A1(n692), .A2(KEYINPUT47), .ZN(n587) );
  XOR2_X1 U640 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n538) );
  NAND2_X1 U641 ( .A1(G224), .A2(n765), .ZN(n537) );
  XNOR2_X1 U642 ( .A(n538), .B(n537), .ZN(n539) );
  INV_X1 U643 ( .A(KEYINPUT89), .ZN(n540) );
  XNOR2_X1 U644 ( .A(G119), .B(G116), .ZN(n543) );
  XNOR2_X1 U645 ( .A(n543), .B(KEYINPUT3), .ZN(n559) );
  XNOR2_X1 U646 ( .A(n545), .B(KEYINPUT71), .ZN(n566) );
  NAND2_X1 U647 ( .A1(G234), .A2(n656), .ZN(n546) );
  XNOR2_X1 U648 ( .A(KEYINPUT20), .B(n546), .ZN(n571) );
  NAND2_X1 U649 ( .A1(n571), .A2(G221), .ZN(n547) );
  XOR2_X1 U650 ( .A(KEYINPUT21), .B(n547), .Z(n702) );
  XOR2_X1 U651 ( .A(KEYINPUT14), .B(KEYINPUT91), .Z(n549) );
  XNOR2_X1 U652 ( .A(n549), .B(n548), .ZN(n551) );
  NAND2_X1 U653 ( .A1(n551), .A2(G952), .ZN(n550) );
  XOR2_X1 U654 ( .A(KEYINPUT92), .B(n550), .Z(n718) );
  NAND2_X1 U655 ( .A1(n765), .A2(n718), .ZN(n622) );
  NAND2_X1 U656 ( .A1(G902), .A2(n551), .ZN(n623) );
  NOR2_X1 U657 ( .A1(G900), .A2(n623), .ZN(n552) );
  NAND2_X1 U658 ( .A1(G953), .A2(n552), .ZN(n553) );
  NAND2_X1 U659 ( .A1(n622), .A2(n553), .ZN(n554) );
  NAND2_X1 U660 ( .A1(n702), .A2(n554), .ZN(n590) );
  NAND2_X1 U661 ( .A1(n555), .A2(G210), .ZN(n556) );
  XNOR2_X1 U662 ( .A(n557), .B(n556), .ZN(n561) );
  NOR2_X2 U663 ( .A1(G902), .A2(n661), .ZN(n564) );
  XNOR2_X2 U664 ( .A(n564), .B(n563), .ZN(n589) );
  INV_X1 U665 ( .A(KEYINPUT107), .ZN(n565) );
  XNOR2_X2 U666 ( .A(n589), .B(n565), .ZN(n632) );
  NAND2_X1 U667 ( .A1(G214), .A2(n566), .ZN(n686) );
  NAND2_X1 U668 ( .A1(n632), .A2(n686), .ZN(n567) );
  XOR2_X1 U669 ( .A(G107), .B(n568), .Z(n570) );
  NAND2_X1 U670 ( .A1(G227), .A2(n765), .ZN(n569) );
  XOR2_X1 U671 ( .A(KEYINPUT95), .B(KEYINPUT94), .Z(n573) );
  NAND2_X1 U672 ( .A1(n571), .A2(G217), .ZN(n572) );
  XNOR2_X1 U673 ( .A(n573), .B(n572), .ZN(n574) );
  XNOR2_X1 U674 ( .A(KEYINPUT25), .B(n574), .ZN(n584) );
  XOR2_X1 U675 ( .A(KEYINPUT75), .B(G110), .Z(n576) );
  XNOR2_X1 U676 ( .A(G137), .B(G119), .ZN(n575) );
  XNOR2_X1 U677 ( .A(n576), .B(n575), .ZN(n577) );
  XOR2_X1 U678 ( .A(n761), .B(n579), .Z(n582) );
  NAND2_X1 U679 ( .A1(G221), .A2(n580), .ZN(n581) );
  XNOR2_X1 U680 ( .A(n582), .B(n581), .ZN(n744) );
  INV_X1 U681 ( .A(n703), .ZN(n647) );
  NAND2_X1 U682 ( .A1(n618), .A2(n586), .ZN(n675) );
  NAND2_X1 U683 ( .A1(n587), .A2(n675), .ZN(n588) );
  XNOR2_X1 U684 ( .A(n588), .B(KEYINPUT81), .ZN(n604) );
  NOR2_X1 U685 ( .A1(n703), .A2(n590), .ZN(n594) );
  NAND2_X1 U686 ( .A1(n594), .A2(n676), .ZN(n591) );
  NOR2_X1 U687 ( .A1(n628), .A2(n591), .ZN(n613) );
  XOR2_X1 U688 ( .A(KEYINPUT112), .B(KEYINPUT36), .Z(n592) );
  XNOR2_X1 U689 ( .A(KEYINPUT113), .B(n593), .ZN(n773) );
  XNOR2_X1 U690 ( .A(n599), .B(KEYINPUT79), .ZN(n671) );
  NAND2_X1 U691 ( .A1(KEYINPUT47), .A2(n671), .ZN(n600) );
  NOR2_X1 U692 ( .A1(KEYINPUT47), .A2(n602), .ZN(n603) );
  XNOR2_X1 U693 ( .A(KEYINPUT38), .B(n618), .ZN(n608) );
  XOR2_X1 U694 ( .A(KEYINPUT111), .B(KEYINPUT42), .Z(n612) );
  NOR2_X1 U695 ( .A1(n607), .A2(n606), .ZN(n630) );
  INV_X1 U696 ( .A(n630), .ZN(n690) );
  INV_X1 U697 ( .A(n608), .ZN(n687) );
  NAND2_X1 U698 ( .A1(n687), .A2(n686), .ZN(n691) );
  NOR2_X1 U699 ( .A1(n690), .A2(n691), .ZN(n609) );
  XOR2_X1 U700 ( .A(KEYINPUT41), .B(n609), .Z(n712) );
  NAND2_X1 U701 ( .A1(n712), .A2(n610), .ZN(n611) );
  XNOR2_X1 U702 ( .A(n612), .B(n611), .ZN(n777) );
  INV_X1 U703 ( .A(n464), .ZN(n650) );
  NAND2_X1 U704 ( .A1(n613), .A2(n686), .ZN(n614) );
  NOR2_X1 U705 ( .A1(n650), .A2(n614), .ZN(n616) );
  XNOR2_X1 U706 ( .A(KEYINPUT110), .B(KEYINPUT43), .ZN(n615) );
  XNOR2_X1 U707 ( .A(n616), .B(n615), .ZN(n617) );
  NOR2_X1 U708 ( .A1(n618), .A2(n617), .ZN(n685) );
  NAND2_X1 U709 ( .A1(n620), .A2(n619), .ZN(n684) );
  INV_X1 U710 ( .A(n684), .ZN(n621) );
  NOR2_X1 U711 ( .A1(n685), .A2(n621), .ZN(n726) );
  INV_X1 U712 ( .A(n622), .ZN(n625) );
  XNOR2_X1 U713 ( .A(G898), .B(KEYINPUT93), .ZN(n751) );
  NAND2_X1 U714 ( .A1(G953), .A2(n751), .ZN(n757) );
  NOR2_X1 U715 ( .A1(n623), .A2(n757), .ZN(n624) );
  NOR2_X1 U716 ( .A1(n625), .A2(n624), .ZN(n627) );
  NOR2_X1 U717 ( .A1(n649), .A2(n464), .ZN(n631) );
  NOR2_X1 U718 ( .A1(n650), .A2(n632), .ZN(n633) );
  INV_X1 U719 ( .A(n706), .ZN(n637) );
  AND2_X1 U720 ( .A1(n637), .A2(n636), .ZN(n638) );
  NAND2_X1 U721 ( .A1(n635), .A2(n638), .ZN(n639) );
  XNOR2_X1 U722 ( .A(KEYINPUT96), .B(n639), .ZN(n666) );
  NAND2_X1 U723 ( .A1(n706), .A2(n640), .ZN(n709) );
  NOR2_X1 U724 ( .A1(n709), .A2(n641), .ZN(n642) );
  XNOR2_X1 U725 ( .A(n642), .B(KEYINPUT31), .ZN(n681) );
  NAND2_X1 U726 ( .A1(n666), .A2(n681), .ZN(n643) );
  XNOR2_X1 U727 ( .A(KEYINPUT97), .B(n643), .ZN(n645) );
  NOR2_X1 U728 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U729 ( .A1(n648), .A2(n647), .ZN(n652) );
  NOR2_X1 U730 ( .A1(n650), .A2(n649), .ZN(n651) );
  NAND2_X1 U731 ( .A1(n652), .A2(n651), .ZN(n653) );
  XNOR2_X1 U732 ( .A(KEYINPUT106), .B(n653), .ZN(n778) );
  INV_X1 U733 ( .A(KEYINPUT64), .ZN(n657) );
  XOR2_X1 U734 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n659) );
  NAND2_X1 U735 ( .A1(n742), .A2(G472), .ZN(n662) );
  XNOR2_X1 U736 ( .A(KEYINPUT87), .B(KEYINPUT88), .ZN(n663) );
  NOR2_X1 U737 ( .A1(n666), .A2(n678), .ZN(n664) );
  XOR2_X1 U738 ( .A(KEYINPUT114), .B(n664), .Z(n665) );
  XNOR2_X1 U739 ( .A(G104), .B(n665), .ZN(G6) );
  INV_X1 U740 ( .A(n672), .ZN(n682) );
  NOR2_X1 U741 ( .A1(n682), .A2(n666), .ZN(n670) );
  XOR2_X1 U742 ( .A(KEYINPUT27), .B(KEYINPUT115), .Z(n668) );
  XNOR2_X1 U743 ( .A(G107), .B(KEYINPUT26), .ZN(n667) );
  XNOR2_X1 U744 ( .A(n668), .B(n667), .ZN(n669) );
  XNOR2_X1 U745 ( .A(n670), .B(n669), .ZN(G9) );
  XOR2_X1 U746 ( .A(G128), .B(KEYINPUT29), .Z(n674) );
  NAND2_X1 U747 ( .A1(n601), .A2(n672), .ZN(n673) );
  XNOR2_X1 U748 ( .A(n674), .B(n673), .ZN(G30) );
  XNOR2_X1 U749 ( .A(n675), .B(G143), .ZN(G45) );
  NAND2_X1 U750 ( .A1(n601), .A2(n676), .ZN(n677) );
  XNOR2_X1 U751 ( .A(n677), .B(n349), .ZN(G48) );
  NOR2_X1 U752 ( .A1(n678), .A2(n681), .ZN(n679) );
  XOR2_X1 U753 ( .A(KEYINPUT116), .B(n679), .Z(n680) );
  XNOR2_X1 U754 ( .A(G113), .B(n680), .ZN(G15) );
  NOR2_X1 U755 ( .A1(n682), .A2(n681), .ZN(n683) );
  XOR2_X1 U756 ( .A(G116), .B(n683), .Z(G18) );
  XNOR2_X1 U757 ( .A(G134), .B(n684), .ZN(G36) );
  XOR2_X1 U758 ( .A(G140), .B(n685), .Z(G42) );
  NAND2_X1 U759 ( .A1(n424), .A2(n712), .ZN(n721) );
  XNOR2_X1 U760 ( .A(KEYINPUT52), .B(KEYINPUT120), .ZN(n717) );
  NOR2_X1 U761 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U762 ( .A(n688), .B(KEYINPUT118), .ZN(n689) );
  NOR2_X1 U763 ( .A1(n690), .A2(n689), .ZN(n694) );
  NOR2_X1 U764 ( .A1(n692), .A2(n691), .ZN(n693) );
  NOR2_X1 U765 ( .A1(n694), .A2(n693), .ZN(n696) );
  NOR2_X1 U766 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U767 ( .A(n697), .B(KEYINPUT119), .ZN(n715) );
  NAND2_X1 U768 ( .A1(n699), .A2(n464), .ZN(n700) );
  XOR2_X1 U769 ( .A(KEYINPUT50), .B(n700), .Z(n701) );
  XNOR2_X1 U770 ( .A(n701), .B(KEYINPUT117), .ZN(n708) );
  NOR2_X1 U771 ( .A1(n703), .A2(n702), .ZN(n704) );
  XOR2_X1 U772 ( .A(KEYINPUT49), .B(n704), .Z(n705) );
  NOR2_X1 U773 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U774 ( .A1(n708), .A2(n707), .ZN(n710) );
  NAND2_X1 U775 ( .A1(n710), .A2(n709), .ZN(n711) );
  XOR2_X1 U776 ( .A(KEYINPUT51), .B(n711), .Z(n713) );
  NAND2_X1 U777 ( .A1(n713), .A2(n712), .ZN(n714) );
  NAND2_X1 U778 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U779 ( .A(n717), .B(n716), .ZN(n719) );
  NAND2_X1 U780 ( .A1(n719), .A2(n718), .ZN(n720) );
  NAND2_X1 U781 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U782 ( .A(n722), .B(KEYINPUT121), .ZN(n732) );
  XNOR2_X1 U783 ( .A(n724), .B(KEYINPUT2), .ZN(n730) );
  AND2_X1 U784 ( .A1(n727), .A2(n726), .ZN(n763) );
  OR2_X1 U785 ( .A1(n725), .A2(n763), .ZN(n728) );
  NAND2_X1 U786 ( .A1(KEYINPUT85), .A2(n728), .ZN(n729) );
  NAND2_X1 U787 ( .A1(n730), .A2(n729), .ZN(n731) );
  NAND2_X1 U788 ( .A1(n742), .A2(G469), .ZN(n736) );
  XOR2_X1 U789 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n734) );
  NAND2_X1 U790 ( .A1(n742), .A2(G475), .ZN(n738) );
  NAND2_X1 U791 ( .A1(G478), .A2(n742), .ZN(n739) );
  XNOR2_X1 U792 ( .A(n740), .B(n739), .ZN(n741) );
  NOR2_X1 U793 ( .A1(n746), .A2(n741), .ZN(G63) );
  NAND2_X1 U794 ( .A1(G217), .A2(n742), .ZN(n743) );
  XNOR2_X1 U795 ( .A(n744), .B(n743), .ZN(n745) );
  NOR2_X1 U796 ( .A1(n746), .A2(n745), .ZN(G66) );
  XOR2_X1 U797 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n748) );
  NAND2_X1 U798 ( .A1(G224), .A2(G953), .ZN(n747) );
  XNOR2_X1 U799 ( .A(n748), .B(n747), .ZN(n749) );
  XOR2_X1 U800 ( .A(KEYINPUT125), .B(n749), .Z(n750) );
  NOR2_X1 U801 ( .A1(n751), .A2(n750), .ZN(n753) );
  NOR2_X1 U802 ( .A1(G953), .A2(n725), .ZN(n752) );
  NOR2_X1 U803 ( .A1(n753), .A2(n752), .ZN(n759) );
  XNOR2_X1 U804 ( .A(n754), .B(G101), .ZN(n755) );
  XNOR2_X1 U805 ( .A(n755), .B(G110), .ZN(n756) );
  NAND2_X1 U806 ( .A1(n757), .A2(n756), .ZN(n758) );
  XOR2_X1 U807 ( .A(n759), .B(n758), .Z(n760) );
  XNOR2_X1 U808 ( .A(KEYINPUT127), .B(n760), .ZN(G69) );
  XOR2_X1 U809 ( .A(n761), .B(n762), .Z(n767) );
  INV_X1 U810 ( .A(n767), .ZN(n764) );
  XNOR2_X1 U811 ( .A(n764), .B(n763), .ZN(n766) );
  NAND2_X1 U812 ( .A1(n766), .A2(n765), .ZN(n771) );
  XNOR2_X1 U813 ( .A(G227), .B(n767), .ZN(n768) );
  NAND2_X1 U814 ( .A1(n768), .A2(G900), .ZN(n769) );
  NAND2_X1 U815 ( .A1(n769), .A2(G953), .ZN(n770) );
  NAND2_X1 U816 ( .A1(n771), .A2(n770), .ZN(G72) );
  XOR2_X1 U817 ( .A(G125), .B(KEYINPUT37), .Z(n772) );
  XNOR2_X1 U818 ( .A(n773), .B(n772), .ZN(G27) );
  XOR2_X1 U819 ( .A(n774), .B(G122), .Z(G24) );
  XNOR2_X1 U820 ( .A(n775), .B(G110), .ZN(G12) );
  XNOR2_X1 U821 ( .A(n776), .B(G131), .ZN(G33) );
  XNOR2_X1 U822 ( .A(G137), .B(n777), .ZN(G39) );
  XNOR2_X1 U823 ( .A(G101), .B(n778), .ZN(G3) );
endmodule

