//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 0 0 1 0 0 1 0 0 0 1 0 0 0 0 1 1 1 1 1 0 1 0 0 1 1 1 0 1 0 0 0 0 0 1 1 0 1 0 1 1 1 1 1 1 0 1 0 1 1 1 1 0 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:30 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n757, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n784, new_n785, new_n786, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n855,
    new_n856, new_n857, new_n859, new_n860, new_n861, new_n862, new_n864,
    new_n865, new_n866, new_n867, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n914, new_n915, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n924, new_n925, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n955, new_n956, new_n957, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n966, new_n967;
  XNOR2_X1  g000(.A(G197gat), .B(G204gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT22), .ZN(new_n203));
  INV_X1    g002(.A(G211gat), .ZN(new_n204));
  INV_X1    g003(.A(G218gat), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n203), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n202), .A2(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G211gat), .B(G218gat), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n208), .A2(new_n202), .A3(new_n206), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT72), .ZN(new_n214));
  INV_X1    g013(.A(G169gat), .ZN(new_n215));
  INV_X1    g014(.A(G176gat), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NOR2_X1   g016(.A1(G169gat), .A2(G176gat), .ZN(new_n218));
  NOR3_X1   g017(.A1(new_n217), .A2(KEYINPUT26), .A3(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(KEYINPUT26), .ZN(new_n220));
  NAND2_X1  g019(.A1(G183gat), .A2(G190gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n219), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT64), .ZN(new_n224));
  INV_X1    g023(.A(G183gat), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n224), .B1(new_n225), .B2(KEYINPUT27), .ZN(new_n226));
  AOI21_X1  g025(.A(G190gat), .B1(new_n225), .B2(KEYINPUT27), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT27), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n228), .A2(KEYINPUT64), .A3(G183gat), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n226), .A2(new_n227), .A3(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT28), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n230), .A2(KEYINPUT65), .A3(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n228), .A2(G183gat), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n227), .A2(KEYINPUT28), .A3(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(KEYINPUT66), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT66), .ZN(new_n236));
  NAND4_X1  g035(.A1(new_n227), .A2(new_n236), .A3(KEYINPUT28), .A4(new_n233), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n232), .A2(new_n235), .A3(new_n237), .ZN(new_n238));
  AOI21_X1  g037(.A(KEYINPUT65), .B1(new_n230), .B2(new_n231), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n223), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT23), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n218), .B(new_n241), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n221), .A2(KEYINPUT24), .ZN(new_n243));
  NOR2_X1   g042(.A1(new_n243), .A2(new_n217), .ZN(new_n244));
  OR2_X1    g043(.A1(G183gat), .A2(G190gat), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n245), .A2(KEYINPUT24), .A3(new_n221), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n242), .A2(new_n244), .A3(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT25), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n242), .A2(new_n244), .A3(KEYINPUT25), .A4(new_n246), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  AOI21_X1  g050(.A(KEYINPUT29), .B1(new_n240), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(G226gat), .A2(G233gat), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n214), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n230), .A2(new_n231), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT65), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n258), .A2(new_n232), .A3(new_n235), .A4(new_n237), .ZN(new_n259));
  AOI22_X1  g058(.A1(new_n259), .A2(new_n223), .B1(new_n249), .B2(new_n250), .ZN(new_n260));
  OAI211_X1 g059(.A(KEYINPUT72), .B(new_n253), .C1(new_n260), .C2(KEYINPUT29), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n213), .B1(new_n255), .B2(new_n261), .ZN(new_n262));
  AND3_X1   g061(.A1(new_n240), .A2(KEYINPUT71), .A3(new_n251), .ZN(new_n263));
  AOI21_X1  g062(.A(KEYINPUT71), .B1(new_n240), .B2(new_n251), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  AOI21_X1  g064(.A(KEYINPUT73), .B1(new_n265), .B2(new_n254), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT73), .ZN(new_n267));
  NOR4_X1   g066(.A1(new_n263), .A2(new_n264), .A3(new_n267), .A4(new_n253), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n262), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(G8gat), .B(G36gat), .ZN(new_n270));
  XNOR2_X1  g069(.A(G64gat), .B(G92gat), .ZN(new_n271));
  XOR2_X1   g070(.A(new_n270), .B(new_n271), .Z(new_n272));
  NAND2_X1  g071(.A1(new_n240), .A2(new_n251), .ZN(new_n273));
  INV_X1    g072(.A(new_n264), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n260), .A2(KEYINPUT71), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  OR2_X1    g075(.A1(new_n254), .A2(KEYINPUT29), .ZN(new_n277));
  OAI221_X1 g076(.A(new_n213), .B1(new_n273), .B2(new_n253), .C1(new_n276), .C2(new_n277), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n269), .A2(new_n272), .A3(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT74), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT30), .ZN(new_n281));
  AND3_X1   g080(.A1(new_n279), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n280), .B1(new_n279), .B2(new_n281), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(G127gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(G134gat), .ZN(new_n286));
  INV_X1    g085(.A(G134gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(G127gat), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n286), .A2(new_n288), .A3(KEYINPUT67), .ZN(new_n289));
  INV_X1    g088(.A(G113gat), .ZN(new_n290));
  INV_X1    g089(.A(G120gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT1), .ZN(new_n293));
  NAND2_X1  g092(.A1(G113gat), .A2(G120gat), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n292), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  OAI211_X1 g094(.A(new_n289), .B(new_n295), .C1(KEYINPUT67), .C2(new_n286), .ZN(new_n296));
  AND2_X1   g095(.A1(G113gat), .A2(G120gat), .ZN(new_n297));
  NOR2_X1   g096(.A1(G113gat), .A2(G120gat), .ZN(new_n298));
  OAI21_X1  g097(.A(KEYINPUT68), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT68), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n292), .A2(new_n300), .A3(new_n294), .ZN(new_n301));
  XNOR2_X1  g100(.A(G127gat), .B(G134gat), .ZN(new_n302));
  NAND4_X1  g101(.A1(new_n299), .A2(new_n301), .A3(new_n293), .A4(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT77), .ZN(new_n304));
  AND3_X1   g103(.A1(new_n296), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n304), .B1(new_n296), .B2(new_n303), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(G141gat), .ZN(new_n308));
  OAI21_X1  g107(.A(KEYINPUT75), .B1(new_n308), .B2(G148gat), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT75), .ZN(new_n310));
  INV_X1    g109(.A(G148gat), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n310), .A2(new_n311), .A3(G141gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n308), .A2(G148gat), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n309), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(G155gat), .A2(G162gat), .ZN(new_n315));
  INV_X1    g114(.A(G155gat), .ZN(new_n316));
  INV_X1    g115(.A(G162gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n315), .B1(new_n318), .B2(KEYINPUT2), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n314), .A2(new_n319), .ZN(new_n320));
  XNOR2_X1  g119(.A(G141gat), .B(G148gat), .ZN(new_n321));
  OAI211_X1 g120(.A(new_n315), .B(new_n318), .C1(new_n321), .C2(KEYINPUT2), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(KEYINPUT76), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT76), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n320), .A2(new_n322), .A3(new_n325), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n324), .A2(KEYINPUT3), .A3(new_n326), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n323), .A2(KEYINPUT3), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n307), .A2(new_n327), .A3(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT4), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n296), .A2(new_n303), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n331), .B1(new_n332), .B2(new_n323), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT2), .ZN(new_n334));
  INV_X1    g133(.A(new_n313), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n308), .A2(G148gat), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n334), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  AND2_X1   g136(.A1(new_n318), .A2(new_n315), .ZN(new_n338));
  AOI22_X1  g137(.A1(new_n337), .A2(new_n338), .B1(new_n314), .B2(new_n319), .ZN(new_n339));
  NAND4_X1  g138(.A1(new_n339), .A2(KEYINPUT4), .A3(new_n296), .A4(new_n303), .ZN(new_n340));
  AND2_X1   g139(.A1(new_n333), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(G225gat), .A2(G233gat), .ZN(new_n342));
  XOR2_X1   g141(.A(new_n342), .B(KEYINPUT78), .Z(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  NAND4_X1  g143(.A1(new_n330), .A2(KEYINPUT5), .A3(new_n341), .A4(new_n344), .ZN(new_n345));
  AND3_X1   g144(.A1(new_n330), .A2(new_n344), .A3(new_n341), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT5), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n332), .A2(KEYINPUT77), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n296), .A2(new_n303), .A3(new_n304), .ZN(new_n349));
  NAND4_X1  g148(.A1(new_n348), .A2(new_n324), .A3(new_n326), .A4(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n332), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(new_n339), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n347), .B1(new_n353), .B2(new_n343), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n345), .B1(new_n346), .B2(new_n354), .ZN(new_n355));
  XOR2_X1   g154(.A(G1gat), .B(G29gat), .Z(new_n356));
  XNOR2_X1  g155(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n357));
  XNOR2_X1  g156(.A(new_n356), .B(new_n357), .ZN(new_n358));
  XNOR2_X1  g157(.A(G57gat), .B(G85gat), .ZN(new_n359));
  XNOR2_X1  g158(.A(new_n358), .B(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n355), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT6), .ZN(new_n363));
  OAI211_X1 g162(.A(new_n360), .B(new_n345), .C1(new_n346), .C2(new_n354), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n362), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  OR3_X1    g164(.A1(new_n355), .A2(new_n363), .A3(new_n361), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n269), .A2(new_n278), .ZN(new_n368));
  INV_X1    g167(.A(new_n272), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND4_X1  g169(.A1(new_n269), .A2(KEYINPUT30), .A3(new_n272), .A4(new_n278), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n367), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  OAI21_X1  g171(.A(KEYINPUT80), .B1(new_n284), .B2(new_n372), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n213), .B1(new_n328), .B2(KEYINPUT29), .ZN(new_n374));
  NAND2_X1  g173(.A1(G228gat), .A2(G233gat), .ZN(new_n375));
  AOI21_X1  g174(.A(KEYINPUT29), .B1(new_n210), .B2(new_n211), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n323), .B1(new_n376), .B2(KEYINPUT3), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n374), .A2(new_n375), .A3(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  OAI211_X1 g178(.A(new_n324), .B(new_n326), .C1(KEYINPUT3), .C2(new_n376), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n375), .B1(new_n374), .B2(new_n380), .ZN(new_n381));
  OAI21_X1  g180(.A(G22gat), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(G22gat), .ZN(new_n383));
  AND2_X1   g182(.A1(new_n374), .A2(new_n380), .ZN(new_n384));
  OAI211_X1 g183(.A(new_n378), .B(new_n383), .C1(new_n384), .C2(new_n375), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n382), .A2(new_n385), .A3(KEYINPUT83), .ZN(new_n386));
  XOR2_X1   g185(.A(G78gat), .B(G106gat), .Z(new_n387));
  XNOR2_X1  g186(.A(KEYINPUT81), .B(KEYINPUT31), .ZN(new_n388));
  XNOR2_X1  g187(.A(new_n387), .B(new_n388), .ZN(new_n389));
  XOR2_X1   g188(.A(KEYINPUT82), .B(G50gat), .Z(new_n390));
  XOR2_X1   g189(.A(new_n389), .B(new_n390), .Z(new_n391));
  AND3_X1   g190(.A1(new_n386), .A2(KEYINPUT84), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n386), .A2(KEYINPUT84), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT84), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n382), .A2(new_n385), .A3(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n391), .ZN(new_n396));
  AND2_X1   g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n392), .B1(new_n393), .B2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n279), .A2(new_n281), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(KEYINPUT74), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n279), .A2(new_n280), .A3(new_n281), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  AND3_X1   g202(.A1(new_n367), .A2(new_n370), .A3(new_n371), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT80), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n403), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n373), .A2(new_n399), .A3(new_n406), .ZN(new_n407));
  AND2_X1   g206(.A1(G227gat), .A2(G233gat), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n273), .A2(new_n351), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n240), .A2(new_n332), .A3(new_n251), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n408), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT34), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(KEYINPUT70), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT70), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n411), .A2(new_n415), .A3(new_n412), .ZN(new_n416));
  OR2_X1    g215(.A1(new_n411), .A2(new_n412), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n414), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT32), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n409), .A2(new_n408), .A3(new_n410), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT69), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND4_X1  g221(.A1(new_n409), .A2(KEYINPUT69), .A3(new_n408), .A4(new_n410), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n419), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(KEYINPUT33), .B1(new_n422), .B2(new_n423), .ZN(new_n425));
  XOR2_X1   g224(.A(G15gat), .B(G43gat), .Z(new_n426));
  XNOR2_X1  g225(.A(G71gat), .B(G99gat), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n426), .B(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  NOR3_X1   g228(.A1(new_n424), .A2(new_n425), .A3(new_n429), .ZN(new_n430));
  AOI221_X4 g229(.A(new_n419), .B1(KEYINPUT33), .B2(new_n428), .C1(new_n422), .C2(new_n423), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n418), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n424), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n422), .A2(new_n423), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT33), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n433), .A2(new_n436), .A3(new_n428), .ZN(new_n437));
  INV_X1    g236(.A(new_n431), .ZN(new_n438));
  INV_X1    g237(.A(new_n418), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n437), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n432), .A2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT36), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n432), .A2(KEYINPUT36), .A3(new_n440), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n407), .A2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(new_n368), .ZN(new_n447));
  XOR2_X1   g246(.A(KEYINPUT85), .B(KEYINPUT37), .Z(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(new_n369), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT37), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n447), .A2(new_n451), .ZN(new_n452));
  OAI21_X1  g251(.A(KEYINPUT38), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n279), .A2(new_n365), .A3(new_n366), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n272), .B1(new_n447), .B2(new_n448), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n276), .A2(new_n277), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n456), .B1(new_n260), .B2(new_n254), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n451), .B1(new_n457), .B2(new_n212), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n212), .B1(new_n255), .B2(new_n261), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n459), .B1(new_n266), .B2(new_n268), .ZN(new_n460));
  AOI21_X1  g259(.A(KEYINPUT38), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n454), .B1(new_n455), .B2(new_n461), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n399), .B1(new_n453), .B2(new_n462), .ZN(new_n463));
  AND2_X1   g262(.A1(new_n370), .A2(new_n371), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n403), .A2(new_n464), .ZN(new_n465));
  AND2_X1   g264(.A1(new_n330), .A2(new_n341), .ZN(new_n466));
  OR3_X1    g265(.A1(new_n466), .A2(KEYINPUT39), .A3(new_n344), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n466), .A2(new_n344), .ZN(new_n468));
  OAI21_X1  g267(.A(KEYINPUT39), .B1(new_n353), .B2(new_n343), .ZN(new_n469));
  OAI211_X1 g268(.A(new_n467), .B(new_n361), .C1(new_n468), .C2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT40), .ZN(new_n471));
  OR2_X1    g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n470), .A2(new_n471), .ZN(new_n473));
  NAND4_X1  g272(.A1(new_n465), .A2(new_n364), .A3(new_n472), .A4(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n463), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(KEYINPUT86), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT86), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n463), .A2(new_n474), .A3(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n446), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  NOR3_X1   g278(.A1(new_n284), .A2(KEYINPUT80), .A3(new_n372), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n405), .B1(new_n403), .B2(new_n404), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n432), .A2(new_n398), .A3(new_n440), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT88), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND4_X1  g284(.A1(new_n432), .A2(new_n398), .A3(new_n440), .A4(KEYINPUT88), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  OAI21_X1  g286(.A(KEYINPUT35), .B1(new_n482), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(KEYINPUT89), .ZN(new_n489));
  OAI211_X1 g288(.A(new_n485), .B(new_n486), .C1(new_n480), .C2(new_n481), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT89), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n490), .A2(new_n491), .A3(KEYINPUT35), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT87), .ZN(new_n494));
  XNOR2_X1  g293(.A(new_n441), .B(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(new_n398), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  NOR3_X1   g296(.A1(new_n284), .A2(KEYINPUT35), .A3(new_n372), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n479), .B1(new_n493), .B2(new_n499), .ZN(new_n500));
  XNOR2_X1  g299(.A(G15gat), .B(G22gat), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT16), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n501), .B1(new_n502), .B2(G1gat), .ZN(new_n503));
  OAI211_X1 g302(.A(new_n503), .B(KEYINPUT92), .C1(G1gat), .C2(new_n501), .ZN(new_n504));
  XNOR2_X1  g303(.A(new_n504), .B(G8gat), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT14), .ZN(new_n506));
  INV_X1    g305(.A(G29gat), .ZN(new_n507));
  INV_X1    g306(.A(G36gat), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n506), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  OAI21_X1  g308(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n510));
  AOI22_X1  g309(.A1(new_n509), .A2(new_n510), .B1(G29gat), .B2(G36gat), .ZN(new_n511));
  XNOR2_X1  g310(.A(G43gat), .B(G50gat), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(KEYINPUT15), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n514), .B(KEYINPUT90), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT91), .ZN(new_n516));
  AND2_X1   g315(.A1(new_n509), .A2(new_n516), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n509), .A2(new_n516), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n510), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  OR2_X1    g318(.A1(new_n512), .A2(KEYINPUT15), .ZN(new_n520));
  NAND2_X1  g319(.A1(G29gat), .A2(G36gat), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n519), .A2(new_n520), .A3(new_n513), .A4(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n515), .A2(new_n522), .ZN(new_n523));
  NOR2_X1   g322(.A1(KEYINPUT93), .A2(KEYINPUT17), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(KEYINPUT93), .A2(KEYINPUT17), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n523), .A2(KEYINPUT93), .A3(KEYINPUT17), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n505), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(G229gat), .A2(G233gat), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  AND2_X1   g330(.A1(new_n523), .A2(new_n505), .ZN(new_n532));
  NOR3_X1   g331(.A1(new_n529), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  OR2_X1    g332(.A1(new_n533), .A2(KEYINPUT18), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(KEYINPUT18), .ZN(new_n535));
  XOR2_X1   g334(.A(new_n530), .B(KEYINPUT13), .Z(new_n536));
  NOR2_X1   g335(.A1(new_n523), .A2(new_n505), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n536), .B1(new_n532), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n534), .A2(new_n535), .A3(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(G113gat), .B(G141gat), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n540), .B(G197gat), .ZN(new_n541));
  XNOR2_X1  g340(.A(KEYINPUT11), .B(G169gat), .ZN(new_n542));
  XOR2_X1   g341(.A(new_n541), .B(new_n542), .Z(new_n543));
  XOR2_X1   g342(.A(new_n543), .B(KEYINPUT12), .Z(new_n544));
  NAND2_X1  g343(.A1(new_n539), .A2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(new_n544), .ZN(new_n546));
  NAND4_X1  g345(.A1(new_n534), .A2(new_n546), .A3(new_n535), .A4(new_n538), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n500), .A2(new_n549), .ZN(new_n550));
  XNOR2_X1  g349(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n551), .B(new_n316), .ZN(new_n552));
  XNOR2_X1  g351(.A(G183gat), .B(G211gat), .ZN(new_n553));
  XOR2_X1   g352(.A(new_n552), .B(new_n553), .Z(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  NOR2_X1   g354(.A1(G71gat), .A2(G78gat), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT94), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n556), .B(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(G64gat), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n559), .A2(G57gat), .ZN(new_n560));
  INV_X1    g359(.A(G57gat), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n561), .A2(G64gat), .ZN(new_n562));
  OAI21_X1  g361(.A(KEYINPUT9), .B1(new_n560), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(G71gat), .A2(G78gat), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n558), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT95), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n565), .B(new_n566), .ZN(new_n567));
  OR2_X1    g366(.A1(new_n562), .A2(KEYINPUT96), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n562), .A2(KEYINPUT96), .ZN(new_n569));
  OAI211_X1 g368(.A(new_n568), .B(new_n569), .C1(G57gat), .C2(new_n559), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n556), .A2(KEYINPUT9), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(new_n564), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n567), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n575), .A2(KEYINPUT21), .ZN(new_n576));
  NAND2_X1  g375(.A1(G231gat), .A2(G233gat), .ZN(new_n577));
  XOR2_X1   g376(.A(new_n576), .B(new_n577), .Z(new_n578));
  XNOR2_X1  g377(.A(new_n578), .B(new_n285), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n505), .B1(new_n575), .B2(KEYINPUT21), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n578), .B(G127gat), .ZN(new_n582));
  INV_X1    g381(.A(new_n580), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n555), .B1(new_n581), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n579), .A2(new_n580), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n582), .A2(new_n583), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n586), .A2(new_n587), .A3(new_n554), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n527), .A2(new_n528), .ZN(new_n590));
  NAND2_X1  g389(.A1(G85gat), .A2(G92gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n591), .B(KEYINPUT7), .ZN(new_n592));
  NAND2_X1  g391(.A1(G99gat), .A2(G106gat), .ZN(new_n593));
  INV_X1    g392(.A(G85gat), .ZN(new_n594));
  INV_X1    g393(.A(G92gat), .ZN(new_n595));
  AOI22_X1  g394(.A1(KEYINPUT8), .A2(new_n593), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n592), .A2(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(G99gat), .B(G106gat), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n597), .B(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n590), .A2(new_n600), .ZN(new_n601));
  AND2_X1   g400(.A1(G232gat), .A2(G233gat), .ZN(new_n602));
  AOI22_X1  g401(.A1(new_n523), .A2(new_n599), .B1(KEYINPUT41), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  XOR2_X1   g403(.A(G190gat), .B(G218gat), .Z(new_n605));
  AND2_X1   g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n604), .A2(new_n605), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n602), .A2(KEYINPUT41), .ZN(new_n609));
  XNOR2_X1  g408(.A(G134gat), .B(G162gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  OR2_X1    g410(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n608), .A2(new_n611), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n589), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(G230gat), .A2(G233gat), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n575), .A2(new_n599), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n574), .A2(new_n600), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n616), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  XOR2_X1   g418(.A(new_n619), .B(KEYINPUT98), .Z(new_n620));
  NOR2_X1   g419(.A1(new_n574), .A2(new_n600), .ZN(new_n621));
  AND3_X1   g420(.A1(new_n621), .A2(KEYINPUT97), .A3(KEYINPUT10), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT10), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n617), .A2(new_n623), .A3(new_n618), .ZN(new_n624));
  AOI21_X1  g423(.A(KEYINPUT97), .B1(new_n621), .B2(KEYINPUT10), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n622), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n626), .A2(new_n616), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n627), .A2(KEYINPUT102), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT102), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n626), .A2(new_n629), .A3(new_n616), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n620), .B1(new_n628), .B2(new_n630), .ZN(new_n631));
  XOR2_X1   g430(.A(G176gat), .B(G204gat), .Z(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(KEYINPUT101), .ZN(new_n633));
  XNOR2_X1  g432(.A(G120gat), .B(G148gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(KEYINPUT99), .B(KEYINPUT100), .ZN(new_n636));
  XOR2_X1   g435(.A(new_n635), .B(new_n636), .Z(new_n637));
  NOR2_X1   g436(.A1(new_n631), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n627), .ZN(new_n639));
  INV_X1    g438(.A(new_n637), .ZN(new_n640));
  NOR3_X1   g439(.A1(new_n639), .A2(new_n620), .A3(new_n640), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n638), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n615), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n550), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n645), .A2(new_n367), .ZN(new_n646));
  XOR2_X1   g445(.A(KEYINPUT103), .B(G1gat), .Z(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(G1324gat));
  NAND3_X1  g447(.A1(new_n550), .A2(new_n465), .A3(new_n644), .ZN(new_n649));
  AND2_X1   g448(.A1(new_n649), .A2(G8gat), .ZN(new_n650));
  XNOR2_X1  g449(.A(KEYINPUT16), .B(G8gat), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  OAI21_X1  g451(.A(KEYINPUT42), .B1(new_n650), .B2(new_n652), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n653), .B1(KEYINPUT42), .B2(new_n652), .ZN(G1325gat));
  NOR2_X1   g453(.A1(new_n445), .A2(KEYINPUT104), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT104), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n656), .B1(new_n443), .B2(new_n444), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  OAI21_X1  g457(.A(G15gat), .B1(new_n645), .B2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(G15gat), .ZN(new_n660));
  NAND4_X1  g459(.A1(new_n550), .A2(new_n660), .A3(new_n495), .A4(new_n644), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n659), .A2(new_n661), .ZN(G1326gat));
  NOR2_X1   g461(.A1(new_n645), .A2(new_n398), .ZN(new_n663));
  XOR2_X1   g462(.A(KEYINPUT43), .B(G22gat), .Z(new_n664));
  XNOR2_X1  g463(.A(new_n663), .B(new_n664), .ZN(G1327gat));
  INV_X1    g464(.A(new_n367), .ZN(new_n666));
  NOR3_X1   g465(.A1(new_n589), .A2(new_n643), .A3(new_n614), .ZN(new_n667));
  AND4_X1   g466(.A1(new_n507), .A2(new_n550), .A3(new_n666), .A4(new_n667), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(KEYINPUT105), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n669), .A2(KEYINPUT45), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT105), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n668), .B(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT45), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  OAI21_X1  g473(.A(KEYINPUT44), .B1(new_n500), .B2(new_n614), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT108), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT35), .ZN(new_n677));
  AND2_X1   g476(.A1(new_n485), .A2(new_n486), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n373), .A2(new_n406), .ZN(new_n679));
  AOI211_X1 g478(.A(KEYINPUT89), .B(new_n677), .C1(new_n678), .C2(new_n679), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n491), .B1(new_n490), .B2(KEYINPUT35), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n499), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n478), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n477), .B1(new_n463), .B2(new_n474), .ZN(new_n684));
  OAI211_X1 g483(.A(new_n658), .B(new_n407), .C1(new_n683), .C2(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n614), .A2(KEYINPUT44), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n676), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n687), .ZN(new_n689));
  AOI211_X1 g488(.A(KEYINPUT108), .B(new_n689), .C1(new_n682), .C2(new_n685), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n675), .B1(new_n688), .B2(new_n690), .ZN(new_n691));
  OR2_X1    g490(.A1(new_n643), .A2(KEYINPUT107), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n643), .A2(KEYINPUT107), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n589), .B(KEYINPUT106), .ZN(new_n696));
  AND3_X1   g495(.A1(new_n695), .A2(new_n548), .A3(new_n696), .ZN(new_n697));
  AND2_X1   g496(.A1(new_n691), .A2(new_n697), .ZN(new_n698));
  AND2_X1   g497(.A1(new_n698), .A2(new_n666), .ZN(new_n699));
  OAI211_X1 g498(.A(new_n670), .B(new_n674), .C1(new_n507), .C2(new_n699), .ZN(G1328gat));
  NAND2_X1  g499(.A1(new_n550), .A2(new_n667), .ZN(new_n701));
  INV_X1    g500(.A(new_n465), .ZN(new_n702));
  NOR3_X1   g501(.A1(new_n701), .A2(G36gat), .A3(new_n702), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(KEYINPUT46), .ZN(new_n704));
  AND2_X1   g503(.A1(new_n698), .A2(new_n465), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n704), .B1(new_n508), .B2(new_n705), .ZN(G1329gat));
  INV_X1    g505(.A(G43gat), .ZN(new_n707));
  NAND4_X1  g506(.A1(new_n550), .A2(new_n707), .A3(new_n495), .A4(new_n667), .ZN(new_n708));
  INV_X1    g507(.A(new_n658), .ZN(new_n709));
  AND2_X1   g508(.A1(new_n698), .A2(new_n709), .ZN(new_n710));
  OAI211_X1 g509(.A(KEYINPUT47), .B(new_n708), .C1(new_n710), .C2(new_n707), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT47), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n707), .B1(new_n698), .B2(new_n709), .ZN(new_n713));
  INV_X1    g512(.A(new_n708), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n712), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n711), .A2(new_n715), .ZN(G1330gat));
  INV_X1    g515(.A(G50gat), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n399), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n701), .A2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT48), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n721), .B1(new_n719), .B2(KEYINPUT109), .ZN(new_n722));
  AND2_X1   g521(.A1(new_n698), .A2(new_n399), .ZN(new_n723));
  OAI211_X1 g522(.A(new_n720), .B(new_n722), .C1(new_n723), .C2(new_n717), .ZN(new_n724));
  INV_X1    g523(.A(new_n722), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n717), .B1(new_n698), .B2(new_n399), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n725), .B1(new_n726), .B2(new_n719), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n724), .A2(new_n727), .ZN(G1331gat));
  NAND3_X1  g527(.A1(new_n589), .A2(new_n549), .A3(new_n614), .ZN(new_n729));
  INV_X1    g528(.A(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n694), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(KEYINPUT110), .ZN(new_n732));
  INV_X1    g531(.A(new_n686), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(KEYINPUT111), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(new_n666), .ZN(new_n736));
  XNOR2_X1  g535(.A(KEYINPUT112), .B(G57gat), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n736), .B(new_n737), .ZN(G1332gat));
  INV_X1    g537(.A(KEYINPUT111), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n734), .B(new_n739), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n740), .A2(new_n702), .ZN(new_n741));
  NOR2_X1   g540(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n742));
  AND2_X1   g541(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n741), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n744), .B1(new_n741), .B2(new_n742), .ZN(G1333gat));
  INV_X1    g544(.A(KEYINPUT50), .ZN(new_n746));
  INV_X1    g545(.A(new_n495), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n747), .A2(G71gat), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n735), .A2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(G71gat), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n751), .B1(new_n735), .B2(new_n709), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n746), .B1(new_n750), .B2(new_n752), .ZN(new_n753));
  OAI21_X1  g552(.A(G71gat), .B1(new_n740), .B2(new_n658), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n754), .A2(KEYINPUT50), .A3(new_n749), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n753), .A2(new_n755), .ZN(G1334gat));
  NAND2_X1  g555(.A1(new_n735), .A2(new_n399), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g557(.A1(new_n589), .A2(new_n548), .A3(new_n642), .ZN(new_n759));
  AND2_X1   g558(.A1(new_n691), .A2(new_n759), .ZN(new_n760));
  AND2_X1   g559(.A1(new_n760), .A2(new_n666), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT51), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n589), .A2(new_n548), .ZN(new_n763));
  AND2_X1   g562(.A1(new_n612), .A2(new_n613), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n762), .B1(new_n733), .B2(new_n765), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n686), .A2(KEYINPUT51), .A3(new_n764), .A4(new_n763), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n642), .B1(new_n768), .B2(KEYINPUT113), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n769), .B1(KEYINPUT113), .B2(new_n768), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n666), .A2(new_n594), .ZN(new_n771));
  OAI22_X1  g570(.A1(new_n761), .A2(new_n594), .B1(new_n770), .B2(new_n771), .ZN(G1336gat));
  INV_X1    g571(.A(KEYINPUT115), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n691), .A2(new_n465), .A3(new_n759), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n773), .B1(new_n774), .B2(G92gat), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n694), .A2(new_n595), .A3(new_n465), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(KEYINPUT114), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n777), .B1(new_n766), .B2(new_n767), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n778), .B1(new_n774), .B2(G92gat), .ZN(new_n779));
  NOR3_X1   g578(.A1(new_n775), .A2(new_n779), .A3(KEYINPUT52), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT52), .ZN(new_n781));
  AOI221_X4 g580(.A(new_n778), .B1(new_n773), .B2(new_n781), .C1(new_n774), .C2(G92gat), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n780), .A2(new_n782), .ZN(G1337gat));
  NAND2_X1  g582(.A1(new_n760), .A2(new_n709), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(G99gat), .ZN(new_n785));
  OR2_X1    g584(.A1(new_n747), .A2(G99gat), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n785), .B1(new_n770), .B2(new_n786), .ZN(G1338gat));
  INV_X1    g586(.A(G106gat), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n694), .A2(new_n788), .A3(new_n399), .ZN(new_n789));
  INV_X1    g588(.A(new_n789), .ZN(new_n790));
  AOI21_X1  g589(.A(KEYINPUT53), .B1(new_n768), .B2(new_n790), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n691), .A2(new_n399), .A3(new_n759), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT117), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(G106gat), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n792), .A2(new_n793), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n791), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  AND2_X1   g596(.A1(new_n792), .A2(G106gat), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n789), .B(KEYINPUT116), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n799), .B1(new_n766), .B2(new_n767), .ZN(new_n800));
  OAI21_X1  g599(.A(KEYINPUT53), .B1(new_n798), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n797), .A2(new_n801), .ZN(G1339gat));
  NAND2_X1  g601(.A1(new_n702), .A2(new_n666), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT54), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n628), .A2(new_n630), .A3(new_n804), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n804), .B1(new_n626), .B2(new_n616), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT119), .ZN(new_n807));
  INV_X1    g606(.A(new_n616), .ZN(new_n808));
  AND2_X1   g607(.A1(new_n624), .A2(new_n625), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n808), .B1(new_n809), .B2(new_n622), .ZN(new_n810));
  AND3_X1   g609(.A1(new_n806), .A2(new_n807), .A3(new_n810), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n807), .B1(new_n806), .B2(new_n810), .ZN(new_n812));
  OAI211_X1 g611(.A(new_n640), .B(new_n805), .C1(new_n811), .C2(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT55), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n641), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(new_n812), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n806), .A2(new_n810), .A3(new_n807), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n818), .A2(KEYINPUT55), .A3(new_n640), .A4(new_n805), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n815), .A2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT120), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n815), .A2(KEYINPUT120), .A3(new_n819), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n822), .A2(new_n548), .A3(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(new_n543), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n531), .B1(new_n529), .B2(new_n532), .ZN(new_n826));
  OR2_X1    g625(.A1(new_n826), .A2(KEYINPUT121), .ZN(new_n827));
  NOR3_X1   g626(.A1(new_n532), .A2(new_n537), .A3(new_n536), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n828), .B1(new_n826), .B2(KEYINPUT121), .ZN(new_n829));
  AND2_X1   g628(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  OAI221_X1 g629(.A(new_n547), .B1(new_n825), .B2(new_n830), .C1(new_n638), .C2(new_n641), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n764), .B1(new_n824), .B2(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT122), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n830), .A2(new_n825), .ZN(new_n834));
  INV_X1    g633(.A(new_n547), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n833), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  OAI211_X1 g635(.A(new_n547), .B(KEYINPUT122), .C1(new_n830), .C2(new_n825), .ZN(new_n837));
  AND3_X1   g636(.A1(new_n764), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n822), .A2(new_n838), .A3(new_n823), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n696), .B1(new_n832), .B2(new_n840), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n764), .B1(new_n588), .B2(new_n585), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT118), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n842), .A2(new_n549), .A3(new_n642), .A4(new_n843), .ZN(new_n844));
  OAI21_X1  g643(.A(KEYINPUT118), .B1(new_n729), .B2(new_n643), .ZN(new_n845));
  AND2_X1   g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n803), .B1(new_n841), .B2(new_n847), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n848), .A2(new_n678), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n849), .A2(new_n290), .A3(new_n548), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n848), .A2(new_n548), .A3(new_n497), .ZN(new_n851));
  AND3_X1   g650(.A1(new_n851), .A2(KEYINPUT123), .A3(G113gat), .ZN(new_n852));
  AOI21_X1  g651(.A(KEYINPUT123), .B1(new_n851), .B2(G113gat), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n850), .B1(new_n852), .B2(new_n853), .ZN(G1340gat));
  AOI21_X1  g653(.A(G120gat), .B1(new_n849), .B2(new_n643), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n848), .A2(new_n497), .ZN(new_n856));
  NOR3_X1   g655(.A1(new_n856), .A2(new_n291), .A3(new_n695), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n855), .A2(new_n857), .ZN(G1341gat));
  NAND3_X1  g657(.A1(new_n849), .A2(new_n285), .A3(new_n589), .ZN(new_n859));
  OAI21_X1  g658(.A(G127gat), .B1(new_n856), .B2(new_n696), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT124), .ZN(new_n862));
  XNOR2_X1  g661(.A(new_n861), .B(new_n862), .ZN(G1342gat));
  NAND3_X1  g662(.A1(new_n849), .A2(new_n287), .A3(new_n764), .ZN(new_n864));
  OR2_X1    g663(.A1(new_n864), .A2(KEYINPUT56), .ZN(new_n865));
  OAI21_X1  g664(.A(G134gat), .B1(new_n856), .B2(new_n614), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n864), .A2(KEYINPUT56), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(G1343gat));
  NOR2_X1   g667(.A1(new_n709), .A2(new_n803), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n841), .A2(new_n847), .ZN(new_n870));
  AOI21_X1  g669(.A(KEYINPUT57), .B1(new_n870), .B2(new_n399), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT57), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n398), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n815), .A2(new_n548), .A3(new_n819), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(new_n831), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(new_n614), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n589), .B1(new_n839), .B2(new_n876), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n873), .B1(new_n877), .B2(new_n846), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT125), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  OAI211_X1 g679(.A(KEYINPUT125), .B(new_n873), .C1(new_n877), .C2(new_n846), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  OAI211_X1 g681(.A(new_n548), .B(new_n869), .C1(new_n871), .C2(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(G141gat), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n709), .A2(new_n398), .ZN(new_n885));
  AND2_X1   g684(.A1(new_n848), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n886), .A2(new_n308), .A3(new_n548), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(KEYINPUT58), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT58), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n884), .A2(new_n890), .A3(new_n887), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n889), .A2(new_n891), .ZN(G1344gat));
  NAND3_X1  g691(.A1(new_n886), .A2(new_n311), .A3(new_n643), .ZN(new_n893));
  XNOR2_X1  g692(.A(new_n893), .B(KEYINPUT126), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT59), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n895), .A2(G148gat), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n869), .B1(new_n871), .B2(new_n882), .ZN(new_n897));
  INV_X1    g696(.A(new_n897), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n896), .B1(new_n898), .B2(new_n643), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n803), .A2(new_n642), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n838), .A2(new_n819), .A3(new_n815), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n589), .B1(new_n876), .B2(new_n901), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n729), .A2(new_n643), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n399), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  AND2_X1   g703(.A1(new_n904), .A2(new_n872), .ZN(new_n905));
  INV_X1    g704(.A(new_n873), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n906), .B1(new_n841), .B2(new_n847), .ZN(new_n907));
  OAI211_X1 g706(.A(new_n658), .B(new_n900), .C1(new_n905), .C2(new_n907), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n895), .B1(new_n908), .B2(G148gat), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n894), .B1(new_n899), .B2(new_n909), .ZN(G1345gat));
  OAI21_X1  g709(.A(G155gat), .B1(new_n897), .B2(new_n696), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n886), .A2(new_n316), .A3(new_n589), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(G1346gat));
  AOI21_X1  g712(.A(G162gat), .B1(new_n886), .B2(new_n764), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n614), .A2(new_n317), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n914), .B1(new_n898), .B2(new_n915), .ZN(G1347gat));
  NOR2_X1   g715(.A1(new_n702), .A2(new_n666), .ZN(new_n917));
  AND2_X1   g716(.A1(new_n870), .A2(new_n917), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n918), .A2(new_n678), .ZN(new_n919));
  AOI21_X1  g718(.A(G169gat), .B1(new_n919), .B2(new_n548), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n918), .A2(new_n497), .ZN(new_n921));
  NOR3_X1   g720(.A1(new_n921), .A2(new_n215), .A3(new_n549), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n920), .A2(new_n922), .ZN(G1348gat));
  NAND3_X1  g722(.A1(new_n919), .A2(new_n216), .A3(new_n643), .ZN(new_n924));
  OAI21_X1  g723(.A(G176gat), .B1(new_n921), .B2(new_n695), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(G1349gat));
  NAND2_X1  g725(.A1(new_n225), .A2(KEYINPUT27), .ZN(new_n927));
  AND3_X1   g726(.A1(new_n589), .A2(new_n233), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n919), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g728(.A(G183gat), .B1(new_n921), .B2(new_n696), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(KEYINPUT60), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT60), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n929), .A2(new_n930), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n932), .A2(new_n934), .ZN(G1350gat));
  INV_X1    g734(.A(KEYINPUT127), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n918), .A2(new_n497), .A3(new_n764), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n936), .B1(new_n937), .B2(G190gat), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT61), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n614), .A2(G190gat), .ZN(new_n940));
  AOI22_X1  g739(.A1(new_n938), .A2(new_n939), .B1(new_n919), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n937), .A2(G190gat), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n942), .A2(KEYINPUT127), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n943), .A2(KEYINPUT61), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n942), .A2(KEYINPUT127), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n941), .B1(new_n944), .B2(new_n945), .ZN(G1351gat));
  NAND2_X1  g745(.A1(new_n918), .A2(new_n885), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n947), .A2(new_n549), .ZN(new_n948));
  OAI211_X1 g747(.A(new_n658), .B(new_n917), .C1(new_n905), .C2(new_n907), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n548), .A2(G197gat), .ZN(new_n950));
  OAI22_X1  g749(.A1(new_n948), .A2(G197gat), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  INV_X1    g750(.A(new_n951), .ZN(G1352gat));
  NOR3_X1   g751(.A1(new_n947), .A2(G204gat), .A3(new_n642), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT62), .ZN(new_n954));
  OR2_X1    g753(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n953), .A2(new_n954), .ZN(new_n956));
  OAI21_X1  g755(.A(G204gat), .B1(new_n949), .B2(new_n695), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n955), .A2(new_n956), .A3(new_n957), .ZN(G1353gat));
  INV_X1    g757(.A(new_n589), .ZN(new_n959));
  OR2_X1    g758(.A1(new_n949), .A2(new_n959), .ZN(new_n960));
  AOI21_X1  g759(.A(KEYINPUT63), .B1(new_n960), .B2(G211gat), .ZN(new_n961));
  OAI211_X1 g760(.A(KEYINPUT63), .B(G211gat), .C1(new_n949), .C2(new_n959), .ZN(new_n962));
  INV_X1    g761(.A(new_n962), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n589), .A2(new_n204), .ZN(new_n964));
  OAI22_X1  g763(.A1(new_n961), .A2(new_n963), .B1(new_n947), .B2(new_n964), .ZN(G1354gat));
  OAI21_X1  g764(.A(G218gat), .B1(new_n949), .B2(new_n614), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n764), .A2(new_n205), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n966), .B1(new_n947), .B2(new_n967), .ZN(G1355gat));
endmodule


