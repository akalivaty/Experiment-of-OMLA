//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 1 0 1 1 0 1 1 0 0 0 1 1 0 0 0 1 0 1 1 1 1 1 1 0 0 0 1 0 0 1 1 0 0 1 0 1 1 0 1 0 1 1 1 0 1 1 0 1 1 0 1 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:30 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n703,
    new_n704, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n748, new_n749, new_n750,
    new_n752, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n856, new_n857, new_n859, new_n860, new_n861, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n917, new_n918, new_n920, new_n921, new_n922, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n936, new_n937, new_n938, new_n939, new_n940, new_n942,
    new_n943, new_n944, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n956, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n981,
    new_n982;
  OR2_X1    g000(.A1(KEYINPUT69), .A2(KEYINPUT1), .ZN(new_n202));
  XNOR2_X1  g001(.A(G127gat), .B(G134gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(G113gat), .B(G120gat), .ZN(new_n204));
  OAI211_X1 g003(.A(new_n202), .B(new_n203), .C1(new_n204), .C2(KEYINPUT1), .ZN(new_n205));
  INV_X1    g004(.A(G120gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(G113gat), .ZN(new_n207));
  INV_X1    g006(.A(G113gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(G120gat), .ZN(new_n209));
  AOI21_X1  g008(.A(KEYINPUT1), .B1(new_n207), .B2(new_n209), .ZN(new_n210));
  AND2_X1   g009(.A1(G127gat), .A2(G134gat), .ZN(new_n211));
  NOR2_X1   g010(.A1(G127gat), .A2(G134gat), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n202), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n210), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n205), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT25), .ZN(new_n217));
  OAI21_X1  g016(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(G183gat), .A2(G190gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND3_X1  g019(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(G169gat), .A2(G176gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(KEYINPUT23), .ZN(new_n224));
  INV_X1    g023(.A(G169gat), .ZN(new_n225));
  INV_X1    g024(.A(G176gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n224), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n222), .A2(new_n228), .ZN(new_n229));
  NOR2_X1   g028(.A1(G169gat), .A2(G176gat), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT65), .ZN(new_n231));
  AND3_X1   g030(.A1(new_n230), .A2(new_n231), .A3(KEYINPUT23), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n231), .B1(new_n230), .B2(KEYINPUT23), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n217), .B1(new_n229), .B2(new_n234), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n225), .A2(new_n226), .A3(KEYINPUT23), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n228), .A2(KEYINPUT25), .A3(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n221), .A2(KEYINPUT66), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT66), .ZN(new_n239));
  NAND4_X1  g038(.A1(new_n239), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n240));
  AOI22_X1  g039(.A1(new_n238), .A2(new_n240), .B1(new_n219), .B2(new_n218), .ZN(new_n241));
  OR2_X1    g040(.A1(new_n237), .A2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT67), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n235), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  AOI22_X1  g043(.A1(new_n220), .A2(new_n221), .B1(new_n227), .B2(new_n224), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n236), .A2(KEYINPUT65), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n230), .A2(new_n231), .A3(KEYINPUT23), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  AOI21_X1  g047(.A(KEYINPUT25), .B1(new_n245), .B2(new_n248), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n237), .A2(new_n241), .ZN(new_n250));
  OAI21_X1  g049(.A(KEYINPUT67), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n244), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT26), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n227), .A2(new_n253), .A3(new_n223), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n230), .A2(KEYINPUT26), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n254), .A2(new_n255), .A3(new_n219), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(G183gat), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(KEYINPUT27), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT27), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(G183gat), .ZN(new_n261));
  AND3_X1   g060(.A1(new_n259), .A2(new_n261), .A3(KEYINPUT68), .ZN(new_n262));
  AOI21_X1  g061(.A(KEYINPUT68), .B1(new_n259), .B2(new_n261), .ZN(new_n263));
  INV_X1    g062(.A(G190gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(KEYINPUT28), .ZN(new_n265));
  NOR3_X1   g064(.A1(new_n262), .A2(new_n263), .A3(new_n265), .ZN(new_n266));
  XNOR2_X1  g065(.A(KEYINPUT27), .B(G183gat), .ZN(new_n267));
  AOI21_X1  g066(.A(KEYINPUT28), .B1(new_n267), .B2(new_n264), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n257), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n216), .B1(new_n252), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n259), .A2(new_n261), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT68), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n267), .A2(KEYINPUT68), .ZN(new_n274));
  NAND4_X1  g073(.A1(new_n273), .A2(new_n274), .A3(KEYINPUT28), .A4(new_n264), .ZN(new_n275));
  INV_X1    g074(.A(new_n268), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n256), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  AOI211_X1 g076(.A(new_n215), .B(new_n277), .C1(new_n244), .C2(new_n251), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n270), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(G227gat), .A2(G233gat), .ZN(new_n280));
  XOR2_X1   g079(.A(new_n280), .B(KEYINPUT64), .Z(new_n281));
  OAI21_X1  g080(.A(KEYINPUT34), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n243), .B1(new_n235), .B2(new_n242), .ZN(new_n283));
  NOR3_X1   g082(.A1(new_n249), .A2(new_n250), .A3(KEYINPUT67), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n269), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(new_n215), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n277), .B1(new_n244), .B2(new_n251), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(new_n216), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT34), .ZN(new_n290));
  INV_X1    g089(.A(new_n281), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n289), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  AOI21_X1  g091(.A(KEYINPUT33), .B1(new_n279), .B2(new_n281), .ZN(new_n293));
  XNOR2_X1  g092(.A(G15gat), .B(G43gat), .ZN(new_n294));
  XNOR2_X1  g093(.A(G71gat), .B(G99gat), .ZN(new_n295));
  XNOR2_X1  g094(.A(new_n294), .B(new_n295), .ZN(new_n296));
  OAI211_X1 g095(.A(new_n282), .B(new_n292), .C1(new_n293), .C2(new_n296), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n286), .A2(new_n281), .A3(new_n288), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT33), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n296), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n290), .B1(new_n289), .B2(new_n291), .ZN(new_n301));
  AOI211_X1 g100(.A(KEYINPUT34), .B(new_n281), .C1(new_n286), .C2(new_n288), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n300), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n297), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n298), .A2(KEYINPUT32), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(G22gat), .ZN(new_n307));
  AND2_X1   g106(.A1(G228gat), .A2(G233gat), .ZN(new_n308));
  XNOR2_X1  g107(.A(G211gat), .B(G218gat), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(G197gat), .B(G204gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(G211gat), .A2(G218gat), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT70), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT22), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n312), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n311), .A2(new_n315), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n313), .B1(new_n312), .B2(new_n314), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n310), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n317), .ZN(new_n319));
  NAND4_X1  g118(.A1(new_n319), .A2(new_n309), .A3(new_n311), .A4(new_n315), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT29), .ZN(new_n322));
  AOI21_X1  g121(.A(KEYINPUT3), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(G155gat), .A2(G162gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(KEYINPUT73), .ZN(new_n325));
  XNOR2_X1  g124(.A(G141gat), .B(G148gat), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT2), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n327), .B1(G155gat), .B2(G162gat), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n325), .B1(new_n326), .B2(new_n328), .ZN(new_n329));
  XNOR2_X1  g128(.A(G155gat), .B(G162gat), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n324), .A2(KEYINPUT2), .ZN(new_n333));
  INV_X1    g132(.A(G141gat), .ZN(new_n334));
  INV_X1    g133(.A(G148gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(G141gat), .A2(G148gat), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n333), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n338), .A2(new_n330), .A3(new_n325), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n332), .A2(new_n339), .ZN(new_n340));
  OR2_X1    g139(.A1(new_n323), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n321), .ZN(new_n342));
  XOR2_X1   g141(.A(KEYINPUT74), .B(KEYINPUT3), .Z(new_n343));
  AOI21_X1  g142(.A(KEYINPUT29), .B1(new_n340), .B2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT81), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n342), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  AND3_X1   g145(.A1(new_n338), .A2(new_n330), .A3(new_n325), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n330), .B1(new_n338), .B2(new_n325), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n343), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(new_n322), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n350), .A2(KEYINPUT81), .ZN(new_n351));
  OAI211_X1 g150(.A(new_n308), .B(new_n341), .C1(new_n346), .C2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(new_n308), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT80), .ZN(new_n354));
  OAI211_X1 g153(.A(new_n354), .B(new_n310), .C1(new_n316), .C2(new_n317), .ZN(new_n355));
  OAI211_X1 g154(.A(new_n322), .B(new_n355), .C1(new_n321), .C2(new_n354), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n340), .B1(new_n356), .B2(new_n343), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n344), .A2(new_n321), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n353), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n307), .B1(new_n352), .B2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n352), .A2(new_n359), .A3(new_n307), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  XNOR2_X1  g162(.A(KEYINPUT79), .B(KEYINPUT31), .ZN(new_n364));
  INV_X1    g163(.A(G50gat), .ZN(new_n365));
  XNOR2_X1  g164(.A(new_n364), .B(new_n365), .ZN(new_n366));
  XOR2_X1   g165(.A(G78gat), .B(G106gat), .Z(new_n367));
  XNOR2_X1  g166(.A(new_n366), .B(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT82), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n368), .B1(new_n360), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n363), .A2(new_n370), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n361), .A2(new_n369), .A3(new_n362), .A4(new_n368), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n305), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n297), .A2(new_n303), .A3(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n306), .A2(new_n373), .A3(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(G226gat), .A2(G233gat), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n285), .A2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT71), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n235), .A2(new_n242), .ZN(new_n382));
  AOI21_X1  g181(.A(KEYINPUT29), .B1(new_n382), .B2(new_n269), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n381), .B1(new_n383), .B2(new_n379), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n249), .A2(new_n250), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n385), .A2(new_n277), .ZN(new_n386));
  OAI211_X1 g185(.A(KEYINPUT71), .B(new_n378), .C1(new_n386), .C2(KEYINPUT29), .ZN(new_n387));
  NAND4_X1  g186(.A1(new_n380), .A2(new_n384), .A3(new_n387), .A4(new_n321), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n382), .A2(new_n269), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n379), .A2(KEYINPUT29), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  OAI221_X1 g190(.A(new_n342), .B1(new_n378), .B2(new_n389), .C1(new_n287), .C2(new_n391), .ZN(new_n392));
  XNOR2_X1  g191(.A(G8gat), .B(G36gat), .ZN(new_n393));
  XNOR2_X1  g192(.A(G64gat), .B(G92gat), .ZN(new_n394));
  XOR2_X1   g193(.A(new_n393), .B(new_n394), .Z(new_n395));
  NAND3_X1  g194(.A1(new_n388), .A2(new_n392), .A3(new_n395), .ZN(new_n396));
  XOR2_X1   g195(.A(KEYINPUT72), .B(KEYINPUT30), .Z(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(G225gat), .A2(G233gat), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n347), .A2(new_n348), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n215), .B1(new_n401), .B2(KEYINPUT3), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n400), .B1(new_n402), .B2(new_n349), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n215), .B1(new_n347), .B2(new_n348), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(KEYINPUT4), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT77), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT4), .ZN(new_n407));
  OAI211_X1 g206(.A(new_n215), .B(new_n407), .C1(new_n348), .C2(new_n347), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n405), .A2(new_n406), .A3(new_n408), .ZN(new_n409));
  XOR2_X1   g208(.A(KEYINPUT75), .B(KEYINPUT5), .Z(new_n410));
  INV_X1    g209(.A(new_n408), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(KEYINPUT77), .ZN(new_n412));
  NAND4_X1  g211(.A1(new_n403), .A2(new_n409), .A3(new_n410), .A4(new_n412), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n332), .A2(new_n339), .A3(new_n214), .A4(new_n205), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n404), .A2(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n410), .B1(new_n415), .B2(new_n400), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n407), .B1(new_n340), .B2(new_n215), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n411), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n332), .A2(new_n339), .A3(KEYINPUT3), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n349), .A2(new_n419), .A3(new_n216), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(new_n399), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n416), .B1(new_n418), .B2(new_n421), .ZN(new_n422));
  XOR2_X1   g221(.A(G1gat), .B(G29gat), .Z(new_n423));
  XNOR2_X1  g222(.A(G57gat), .B(G85gat), .ZN(new_n424));
  XNOR2_X1  g223(.A(new_n423), .B(new_n424), .ZN(new_n425));
  XNOR2_X1  g224(.A(KEYINPUT76), .B(KEYINPUT0), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n425), .B(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n413), .A2(new_n422), .A3(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT6), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n428), .B1(new_n413), .B2(new_n422), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  AOI211_X1 g232(.A(new_n430), .B(new_n428), .C1(new_n413), .C2(new_n422), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n398), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n388), .A2(new_n392), .ZN(new_n436));
  INV_X1    g235(.A(new_n395), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n388), .A2(KEYINPUT30), .A3(new_n392), .A4(new_n395), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NOR3_X1   g239(.A1(new_n435), .A2(KEYINPUT35), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n377), .A2(new_n441), .ZN(new_n442));
  OAI21_X1  g241(.A(KEYINPUT78), .B1(new_n435), .B2(new_n440), .ZN(new_n443));
  INV_X1    g242(.A(new_n440), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT78), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n413), .A2(new_n422), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(new_n427), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n447), .A2(new_n430), .A3(new_n429), .ZN(new_n448));
  INV_X1    g247(.A(new_n434), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n444), .A2(new_n445), .A3(new_n450), .A4(new_n398), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n376), .B1(new_n443), .B2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT35), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n442), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  AND3_X1   g253(.A1(new_n448), .A2(new_n449), .A3(new_n396), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT37), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n395), .A2(new_n456), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n457), .B1(new_n436), .B2(new_n437), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT38), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n380), .A2(new_n384), .A3(new_n387), .A4(new_n342), .ZN(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  OAI22_X1  g260(.A1(new_n287), .A2(new_n391), .B1(new_n378), .B2(new_n389), .ZN(new_n462));
  OAI21_X1  g261(.A(KEYINPUT37), .B1(new_n462), .B2(new_n342), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n459), .B1(new_n461), .B2(new_n463), .ZN(new_n464));
  OAI21_X1  g263(.A(KEYINPUT83), .B1(new_n458), .B2(new_n464), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n456), .B1(new_n388), .B2(new_n392), .ZN(new_n466));
  OAI21_X1  g265(.A(KEYINPUT38), .B1(new_n458), .B2(new_n466), .ZN(new_n467));
  AOI22_X1  g266(.A1(new_n285), .A2(new_n390), .B1(new_n386), .B2(new_n379), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n456), .B1(new_n468), .B2(new_n321), .ZN(new_n469));
  AOI21_X1  g268(.A(KEYINPUT38), .B1(new_n469), .B2(new_n460), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT83), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n395), .B1(new_n388), .B2(new_n392), .ZN(new_n472));
  OAI211_X1 g271(.A(new_n470), .B(new_n471), .C1(new_n472), .C2(new_n457), .ZN(new_n473));
  NAND4_X1  g272(.A1(new_n455), .A2(new_n465), .A3(new_n467), .A4(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT40), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n409), .A2(new_n412), .A3(new_n420), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT39), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n476), .A2(new_n477), .A3(new_n400), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(new_n428), .ZN(new_n479));
  OAI21_X1  g278(.A(KEYINPUT39), .B1(new_n415), .B2(new_n400), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n480), .B1(new_n476), .B2(new_n400), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n475), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n476), .A2(new_n400), .ZN(new_n483));
  INV_X1    g282(.A(new_n480), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND4_X1  g284(.A1(new_n485), .A2(KEYINPUT40), .A3(new_n428), .A4(new_n478), .ZN(new_n486));
  AND3_X1   g285(.A1(new_n482), .A2(new_n447), .A3(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n398), .A2(new_n438), .A3(new_n439), .ZN(new_n488));
  AOI22_X1  g287(.A1(new_n487), .A2(new_n488), .B1(new_n371), .B2(new_n372), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n474), .A2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(new_n373), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n443), .A2(new_n491), .A3(new_n451), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT36), .ZN(new_n494));
  AND3_X1   g293(.A1(new_n297), .A2(new_n303), .A3(new_n374), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n374), .B1(new_n297), .B2(new_n303), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n306), .A2(KEYINPUT36), .A3(new_n375), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(new_n499), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n454), .B1(new_n493), .B2(new_n500), .ZN(new_n501));
  XNOR2_X1  g300(.A(G113gat), .B(G141gat), .ZN(new_n502));
  XNOR2_X1  g301(.A(KEYINPUT84), .B(KEYINPUT11), .ZN(new_n503));
  XNOR2_X1  g302(.A(new_n502), .B(new_n503), .ZN(new_n504));
  XOR2_X1   g303(.A(G169gat), .B(G197gat), .Z(new_n505));
  XNOR2_X1  g304(.A(new_n504), .B(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n506), .B(KEYINPUT12), .ZN(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  XNOR2_X1  g307(.A(G15gat), .B(G22gat), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT85), .ZN(new_n510));
  INV_X1    g309(.A(G1gat), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n509), .A2(new_n510), .A3(KEYINPUT16), .A4(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT16), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n509), .A2(new_n514), .ZN(new_n515));
  AOI22_X1  g314(.A1(new_n515), .A2(new_n511), .B1(new_n510), .B2(new_n509), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT86), .ZN(new_n517));
  INV_X1    g316(.A(G8gat), .ZN(new_n518));
  OAI22_X1  g317(.A1(new_n513), .A2(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n515), .A2(new_n511), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n509), .A2(new_n510), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(KEYINPUT86), .B(G8gat), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n522), .A2(new_n512), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n519), .A2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  XOR2_X1   g325(.A(G43gat), .B(G50gat), .Z(new_n527));
  INV_X1    g326(.A(G36gat), .ZN(new_n528));
  AND2_X1   g327(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n529));
  NOR2_X1   g328(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(G29gat), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n532), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n527), .B1(new_n534), .B2(KEYINPUT15), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n535), .B1(KEYINPUT15), .B2(new_n534), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n534), .A2(KEYINPUT15), .A3(new_n527), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n538), .A2(KEYINPUT17), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT17), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n540), .B1(new_n536), .B2(new_n537), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n526), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT87), .ZN(new_n543));
  AND3_X1   g342(.A1(new_n519), .A2(new_n543), .A3(new_n524), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n543), .B1(new_n519), .B2(new_n524), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n538), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(G229gat), .A2(G233gat), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n542), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT18), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n548), .A2(KEYINPUT88), .A3(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(new_n544), .ZN(new_n551));
  INV_X1    g350(.A(new_n538), .ZN(new_n552));
  INV_X1    g351(.A(new_n545), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(new_n546), .ZN(new_n555));
  XNOR2_X1  g354(.A(KEYINPUT89), .B(KEYINPUT13), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n556), .B(new_n547), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n550), .A2(new_n559), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n549), .B1(new_n548), .B2(KEYINPUT88), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n508), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n561), .ZN(new_n563));
  NAND4_X1  g362(.A1(new_n563), .A2(new_n559), .A3(new_n550), .A4(new_n507), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(G85gat), .A2(G92gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n566), .B(KEYINPUT7), .ZN(new_n567));
  NAND2_X1  g366(.A1(G99gat), .A2(G106gat), .ZN(new_n568));
  INV_X1    g367(.A(G85gat), .ZN(new_n569));
  INV_X1    g368(.A(G92gat), .ZN(new_n570));
  AOI22_X1  g369(.A1(KEYINPUT8), .A2(new_n568), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n567), .A2(new_n571), .ZN(new_n572));
  XOR2_X1   g371(.A(G99gat), .B(G106gat), .Z(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n573), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n575), .A2(new_n567), .A3(new_n571), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n577), .B1(new_n539), .B2(new_n541), .ZN(new_n578));
  XOR2_X1   g377(.A(G190gat), .B(G218gat), .Z(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n577), .ZN(new_n581));
  AND2_X1   g380(.A1(G232gat), .A2(G233gat), .ZN(new_n582));
  AOI22_X1  g381(.A1(new_n538), .A2(new_n581), .B1(KEYINPUT41), .B2(new_n582), .ZN(new_n583));
  AND3_X1   g382(.A1(new_n578), .A2(new_n580), .A3(new_n583), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n580), .B1(new_n578), .B2(new_n583), .ZN(new_n585));
  XOR2_X1   g384(.A(G134gat), .B(G162gat), .Z(new_n586));
  NOR2_X1   g385(.A1(new_n582), .A2(KEYINPUT41), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  XOR2_X1   g387(.A(KEYINPUT91), .B(KEYINPUT92), .Z(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  OR3_X1    g390(.A1(new_n584), .A2(new_n585), .A3(new_n591), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n591), .B1(new_n584), .B2(new_n585), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  XOR2_X1   g393(.A(G57gat), .B(G64gat), .Z(new_n595));
  NAND2_X1  g394(.A1(G71gat), .A2(G78gat), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT9), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(G71gat), .B(G78gat), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n595), .A2(new_n600), .A3(new_n598), .ZN(new_n603));
  AND3_X1   g402(.A1(new_n602), .A2(KEYINPUT90), .A3(new_n603), .ZN(new_n604));
  AOI21_X1  g403(.A(KEYINPUT90), .B1(new_n602), .B2(new_n603), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT21), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(G231gat), .A2(G233gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(G127gat), .ZN(new_n611));
  OR2_X1    g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n610), .A2(new_n611), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n551), .A2(new_n553), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n606), .A2(new_n607), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  OR2_X1    g416(.A1(new_n614), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n614), .A2(new_n617), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n621));
  INV_X1    g420(.A(G155gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(G183gat), .B(G211gat), .ZN(new_n624));
  XOR2_X1   g423(.A(new_n623), .B(new_n624), .Z(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n620), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n618), .A2(new_n619), .A3(new_n625), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n594), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(G230gat), .A2(G233gat), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n577), .B1(new_n604), .B2(new_n605), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n602), .A2(new_n603), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n581), .A2(new_n632), .ZN(new_n633));
  AOI21_X1  g432(.A(KEYINPUT10), .B1(new_n631), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n581), .A2(KEYINPUT10), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n635), .A2(new_n606), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n630), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(G120gat), .B(G148gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(G176gat), .B(G204gat), .ZN(new_n639));
  XOR2_X1   g438(.A(new_n638), .B(new_n639), .Z(new_n640));
  NAND2_X1  g439(.A1(new_n631), .A2(new_n633), .ZN(new_n641));
  OAI211_X1 g440(.A(new_n637), .B(new_n640), .C1(new_n630), .C2(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n641), .A2(new_n630), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT93), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n637), .A2(new_n644), .ZN(new_n645));
  OAI211_X1 g444(.A(KEYINPUT93), .B(new_n630), .C1(new_n634), .C2(new_n636), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n643), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n642), .B1(new_n647), .B2(new_n640), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NAND4_X1  g448(.A1(new_n501), .A2(new_n565), .A3(new_n629), .A4(new_n649), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n650), .A2(new_n450), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(new_n511), .ZN(G1324gat));
  INV_X1    g451(.A(new_n650), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n518), .B1(new_n653), .B2(new_n488), .ZN(new_n654));
  INV_X1    g453(.A(new_n488), .ZN(new_n655));
  XNOR2_X1  g454(.A(KEYINPUT16), .B(G8gat), .ZN(new_n656));
  NOR3_X1   g455(.A1(new_n650), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  OAI21_X1  g456(.A(KEYINPUT42), .B1(new_n654), .B2(new_n657), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n658), .B1(KEYINPUT42), .B2(new_n657), .ZN(G1325gat));
  INV_X1    g458(.A(KEYINPUT94), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n497), .A2(new_n498), .A3(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n660), .B1(new_n497), .B2(new_n498), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  OAI21_X1  g463(.A(G15gat), .B1(new_n650), .B2(new_n664), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n495), .A2(new_n496), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  OR2_X1    g466(.A1(new_n667), .A2(G15gat), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n665), .B1(new_n650), .B2(new_n668), .ZN(G1326gat));
  NOR2_X1   g468(.A1(new_n650), .A2(new_n373), .ZN(new_n670));
  XOR2_X1   g469(.A(KEYINPUT43), .B(G22gat), .Z(new_n671));
  XNOR2_X1  g470(.A(new_n670), .B(new_n671), .ZN(G1327gat));
  NAND2_X1  g471(.A1(new_n501), .A2(new_n594), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n627), .A2(new_n628), .ZN(new_n675));
  INV_X1    g474(.A(new_n565), .ZN(new_n676));
  NOR3_X1   g475(.A1(new_n675), .A2(new_n676), .A3(new_n648), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n450), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n679), .A2(new_n532), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n681), .B(KEYINPUT45), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT95), .ZN(new_n683));
  NOR3_X1   g482(.A1(new_n662), .A2(new_n493), .A3(new_n663), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n443), .A2(new_n451), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n377), .A2(new_n685), .ZN(new_n686));
  AOI22_X1  g485(.A1(new_n686), .A2(KEYINPUT35), .B1(new_n377), .B2(new_n441), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n683), .B1(new_n684), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n499), .A2(KEYINPUT94), .ZN(new_n689));
  NAND4_X1  g488(.A1(new_n689), .A2(new_n492), .A3(new_n490), .A4(new_n661), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n690), .A2(new_n454), .A3(KEYINPUT95), .ZN(new_n691));
  INV_X1    g490(.A(new_n594), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n692), .A2(KEYINPUT44), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n688), .A2(new_n691), .A3(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(KEYINPUT96), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n673), .A2(KEYINPUT44), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT96), .ZN(new_n697));
  NAND4_X1  g496(.A1(new_n688), .A2(new_n697), .A3(new_n691), .A4(new_n693), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n695), .A2(new_n696), .A3(new_n698), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n699), .A2(new_n680), .A3(new_n677), .ZN(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n682), .B1(new_n532), .B2(new_n701), .ZN(G1328gat));
  NOR3_X1   g501(.A1(new_n678), .A2(G36gat), .A3(new_n655), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(KEYINPUT46), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n699), .A2(new_n677), .ZN(new_n705));
  OAI21_X1  g504(.A(G36gat), .B1(new_n705), .B2(new_n655), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n704), .A2(new_n706), .ZN(G1329gat));
  INV_X1    g506(.A(KEYINPUT47), .ZN(new_n708));
  INV_X1    g507(.A(new_n664), .ZN(new_n709));
  AND3_X1   g508(.A1(new_n690), .A2(KEYINPUT95), .A3(new_n454), .ZN(new_n710));
  AOI21_X1  g509(.A(KEYINPUT95), .B1(new_n690), .B2(new_n454), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n697), .B1(new_n712), .B2(new_n693), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n698), .A2(new_n696), .ZN(new_n714));
  OAI211_X1 g513(.A(new_n709), .B(new_n677), .C1(new_n713), .C2(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(KEYINPUT97), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT97), .ZN(new_n717));
  NAND4_X1  g516(.A1(new_n699), .A2(new_n717), .A3(new_n709), .A4(new_n677), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n716), .A2(new_n718), .A3(G43gat), .ZN(new_n719));
  NOR3_X1   g518(.A1(new_n678), .A2(G43gat), .A3(new_n667), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n708), .B1(new_n719), .B2(new_n721), .ZN(new_n722));
  AOI211_X1 g521(.A(KEYINPUT47), .B(new_n720), .C1(new_n715), .C2(G43gat), .ZN(new_n723));
  OAI21_X1  g522(.A(KEYINPUT98), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(new_n723), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT98), .ZN(new_n726));
  INV_X1    g525(.A(G43gat), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n727), .B1(new_n715), .B2(KEYINPUT97), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n720), .B1(new_n728), .B2(new_n718), .ZN(new_n729));
  OAI211_X1 g528(.A(new_n725), .B(new_n726), .C1(new_n729), .C2(new_n708), .ZN(new_n730));
  AND2_X1   g529(.A1(new_n724), .A2(new_n730), .ZN(G1330gat));
  OAI21_X1  g530(.A(G50gat), .B1(new_n705), .B2(new_n373), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n679), .A2(new_n365), .A3(new_n491), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT99), .ZN(new_n735));
  AOI21_X1  g534(.A(KEYINPUT48), .B1(new_n733), .B2(new_n735), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n734), .B(new_n736), .ZN(G1331gat));
  NAND4_X1  g536(.A1(new_n712), .A2(new_n676), .A3(new_n629), .A4(new_n648), .ZN(new_n738));
  INV_X1    g537(.A(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(new_n680), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g540(.A(new_n655), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n742));
  XOR2_X1   g541(.A(new_n742), .B(KEYINPUT100), .Z(new_n743));
  NAND2_X1  g542(.A1(new_n739), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(KEYINPUT101), .ZN(new_n745));
  NOR2_X1   g544(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n745), .B(new_n746), .ZN(G1333gat));
  OAI21_X1  g546(.A(G71gat), .B1(new_n738), .B2(new_n664), .ZN(new_n748));
  OR2_X1    g547(.A1(new_n667), .A2(G71gat), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n748), .B1(new_n738), .B2(new_n749), .ZN(new_n750));
  XOR2_X1   g549(.A(new_n750), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g550(.A1(new_n739), .A2(new_n491), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g552(.A1(new_n684), .A2(new_n687), .ZN(new_n754));
  INV_X1    g553(.A(new_n675), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n755), .A2(new_n676), .A3(new_n594), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(KEYINPUT51), .ZN(new_n758));
  INV_X1    g557(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n759), .A2(new_n649), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n760), .A2(new_n569), .A3(new_n680), .ZN(new_n761));
  NOR3_X1   g560(.A1(new_n675), .A2(new_n565), .A3(new_n649), .ZN(new_n762));
  AND2_X1   g561(.A1(new_n699), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(new_n680), .ZN(new_n764));
  INV_X1    g563(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n761), .B1(new_n765), .B2(new_n569), .ZN(G1336gat));
  OAI211_X1 g565(.A(new_n488), .B(new_n762), .C1(new_n713), .C2(new_n714), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(G92gat), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT52), .ZN(new_n769));
  NOR3_X1   g568(.A1(new_n649), .A2(new_n655), .A3(G92gat), .ZN(new_n770));
  INV_X1    g569(.A(new_n770), .ZN(new_n771));
  OAI211_X1 g570(.A(new_n768), .B(new_n769), .C1(new_n759), .C2(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT102), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n757), .B1(new_n773), .B2(KEYINPUT51), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n773), .A2(KEYINPUT51), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n775), .B1(new_n754), .B2(new_n756), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n771), .B1(new_n774), .B2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n768), .A2(new_n778), .ZN(new_n779));
  AOI21_X1  g578(.A(KEYINPUT103), .B1(new_n779), .B2(KEYINPUT52), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n777), .B1(new_n767), .B2(G92gat), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT103), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n781), .A2(new_n782), .A3(new_n769), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n772), .B1(new_n780), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(KEYINPUT104), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT104), .ZN(new_n786));
  OAI211_X1 g585(.A(new_n786), .B(new_n772), .C1(new_n780), .C2(new_n783), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n785), .A2(new_n787), .ZN(G1337gat));
  INV_X1    g587(.A(G99gat), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n760), .A2(new_n789), .A3(new_n666), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n763), .A2(new_n709), .ZN(new_n791));
  INV_X1    g590(.A(new_n791), .ZN(new_n792));
  OAI21_X1  g591(.A(G99gat), .B1(new_n792), .B2(KEYINPUT105), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT105), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n791), .A2(new_n794), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n790), .B1(new_n793), .B2(new_n795), .ZN(G1338gat));
  NAND2_X1  g595(.A1(new_n763), .A2(new_n491), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(G106gat), .ZN(new_n798));
  NOR3_X1   g597(.A1(new_n373), .A2(new_n649), .A3(G106gat), .ZN(new_n799));
  AOI21_X1  g598(.A(KEYINPUT53), .B1(new_n758), .B2(new_n799), .ZN(new_n800));
  AND3_X1   g599(.A1(new_n798), .A2(KEYINPUT106), .A3(new_n800), .ZN(new_n801));
  AOI21_X1  g600(.A(KEYINPUT106), .B1(new_n798), .B2(new_n800), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n774), .A2(new_n776), .ZN(new_n803));
  AOI22_X1  g602(.A1(new_n797), .A2(G106gat), .B1(new_n803), .B2(new_n799), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT53), .ZN(new_n805));
  OAI22_X1  g604(.A1(new_n801), .A2(new_n802), .B1(new_n804), .B2(new_n805), .ZN(G1339gat));
  NAND3_X1  g605(.A1(new_n629), .A2(new_n676), .A3(new_n649), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT54), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT10), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n641), .A2(new_n809), .ZN(new_n810));
  OR2_X1    g609(.A1(new_n635), .A2(new_n606), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n808), .B1(new_n812), .B2(new_n630), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT107), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n634), .A2(new_n636), .ZN(new_n815));
  INV_X1    g614(.A(new_n630), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n814), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NOR4_X1   g616(.A1(new_n634), .A2(new_n636), .A3(KEYINPUT107), .A4(new_n630), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n813), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(new_n640), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n645), .A2(new_n808), .A3(new_n646), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n819), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT55), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n819), .A2(KEYINPUT55), .A3(new_n820), .A4(new_n821), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n565), .A2(new_n824), .A3(new_n642), .A4(new_n825), .ZN(new_n826));
  AND3_X1   g625(.A1(new_n554), .A2(new_n546), .A3(new_n557), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n547), .B1(new_n542), .B2(new_n546), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n506), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(KEYINPUT108), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT108), .ZN(new_n831));
  OAI211_X1 g630(.A(new_n831), .B(new_n506), .C1(new_n827), .C2(new_n828), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n648), .A2(new_n564), .A3(new_n830), .A4(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n594), .B1(new_n826), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n824), .A2(new_n594), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n825), .A2(new_n642), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n564), .A2(new_n830), .A3(new_n832), .ZN(new_n837));
  NOR3_X1   g636(.A1(new_n835), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n834), .A2(new_n838), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n807), .B1(new_n839), .B2(new_n675), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT109), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  OAI211_X1 g641(.A(new_n807), .B(KEYINPUT109), .C1(new_n839), .C2(new_n675), .ZN(new_n843));
  AND2_X1   g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  AND2_X1   g643(.A1(new_n844), .A2(new_n373), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n488), .A2(new_n450), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n845), .A2(new_n666), .A3(new_n846), .ZN(new_n847));
  NOR3_X1   g646(.A1(new_n847), .A2(new_n208), .A3(new_n676), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n844), .A2(new_n680), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(new_n377), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n850), .A2(new_n488), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(new_n565), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n848), .B1(new_n852), .B2(new_n208), .ZN(G1340gat));
  NAND2_X1  g652(.A1(new_n648), .A2(new_n206), .ZN(new_n854));
  XOR2_X1   g653(.A(new_n854), .B(KEYINPUT110), .Z(new_n855));
  NAND2_X1  g654(.A1(new_n851), .A2(new_n855), .ZN(new_n856));
  OAI21_X1  g655(.A(G120gat), .B1(new_n847), .B2(new_n649), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(G1341gat));
  NOR3_X1   g657(.A1(new_n847), .A2(new_n611), .A3(new_n755), .ZN(new_n859));
  XNOR2_X1  g658(.A(new_n859), .B(KEYINPUT111), .ZN(new_n860));
  AOI21_X1  g659(.A(G127gat), .B1(new_n851), .B2(new_n675), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n860), .A2(new_n861), .ZN(G1342gat));
  NAND2_X1  g661(.A1(new_n655), .A2(new_n594), .ZN(new_n863));
  XNOR2_X1  g662(.A(new_n863), .B(KEYINPUT112), .ZN(new_n864));
  INV_X1    g663(.A(G134gat), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  OAI22_X1  g665(.A1(new_n850), .A2(new_n866), .B1(KEYINPUT114), .B2(KEYINPUT56), .ZN(new_n867));
  NAND2_X1  g666(.A1(KEYINPUT114), .A2(KEYINPUT56), .ZN(new_n868));
  XOR2_X1   g667(.A(new_n867), .B(new_n868), .Z(new_n869));
  OAI21_X1  g668(.A(G134gat), .B1(new_n847), .B2(new_n692), .ZN(new_n870));
  XNOR2_X1  g669(.A(new_n870), .B(KEYINPUT113), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n869), .A2(new_n871), .ZN(G1343gat));
  NAND2_X1  g671(.A1(new_n664), .A2(new_n846), .ZN(new_n873));
  INV_X1    g672(.A(new_n873), .ZN(new_n874));
  XNOR2_X1  g673(.A(KEYINPUT115), .B(KEYINPUT55), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n822), .A2(new_n875), .ZN(new_n876));
  NAND4_X1  g675(.A1(new_n565), .A2(new_n876), .A3(new_n642), .A4(new_n825), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n594), .B1(new_n877), .B2(new_n833), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n755), .B1(new_n878), .B2(new_n838), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(new_n807), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT57), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n373), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  XNOR2_X1  g682(.A(new_n883), .B(KEYINPUT116), .ZN(new_n884));
  INV_X1    g683(.A(new_n884), .ZN(new_n885));
  AOI21_X1  g684(.A(KEYINPUT57), .B1(new_n844), .B2(new_n491), .ZN(new_n886));
  OAI211_X1 g685(.A(new_n565), .B(new_n874), .C1(new_n885), .C2(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT119), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n334), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n889), .B1(new_n888), .B2(new_n887), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT58), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n709), .A2(new_n373), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n849), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n565), .A2(new_n334), .ZN(new_n894));
  XOR2_X1   g693(.A(new_n894), .B(KEYINPUT117), .Z(new_n895));
  NAND3_X1  g694(.A1(new_n893), .A2(new_n655), .A3(new_n895), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n890), .A2(new_n891), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n887), .A2(G141gat), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(new_n896), .ZN(new_n899));
  AND3_X1   g698(.A1(new_n899), .A2(KEYINPUT118), .A3(KEYINPUT58), .ZN(new_n900));
  AOI21_X1  g699(.A(KEYINPUT118), .B1(new_n899), .B2(KEYINPUT58), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n897), .B1(new_n900), .B2(new_n901), .ZN(G1344gat));
  NAND4_X1  g701(.A1(new_n893), .A2(new_n335), .A3(new_n655), .A4(new_n648), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n880), .A2(new_n491), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT120), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n904), .A2(new_n905), .A3(new_n881), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n373), .B1(new_n879), .B2(new_n807), .ZN(new_n907));
  OAI21_X1  g706(.A(KEYINPUT120), .B1(new_n907), .B2(KEYINPUT57), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n842), .A2(new_n843), .A3(new_n882), .ZN(new_n910));
  AOI211_X1 g709(.A(new_n649), .B(new_n873), .C1(new_n909), .C2(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n912));
  INV_X1    g711(.A(new_n886), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n873), .B1(new_n913), .B2(new_n884), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n335), .B1(new_n914), .B2(new_n648), .ZN(new_n915));
  OAI221_X1 g714(.A(new_n903), .B1(new_n911), .B2(new_n912), .C1(new_n915), .C2(KEYINPUT59), .ZN(G1345gat));
  NAND4_X1  g715(.A1(new_n893), .A2(new_n622), .A3(new_n655), .A4(new_n675), .ZN(new_n917));
  AND2_X1   g716(.A1(new_n914), .A2(new_n675), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n917), .B1(new_n918), .B2(new_n622), .ZN(G1346gat));
  INV_X1    g718(.A(G162gat), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n893), .A2(new_n920), .A3(new_n864), .ZN(new_n921));
  AND2_X1   g720(.A1(new_n914), .A2(new_n594), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n921), .B1(new_n922), .B2(new_n920), .ZN(G1347gat));
  NOR2_X1   g722(.A1(new_n655), .A2(new_n680), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n844), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(new_n377), .ZN(new_n926));
  INV_X1    g725(.A(new_n926), .ZN(new_n927));
  AOI21_X1  g726(.A(G169gat), .B1(new_n927), .B2(new_n565), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n845), .A2(new_n666), .A3(new_n924), .ZN(new_n929));
  NOR3_X1   g728(.A1(new_n929), .A2(new_n225), .A3(new_n676), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n928), .A2(new_n930), .ZN(G1348gat));
  OAI21_X1  g730(.A(G176gat), .B1(new_n929), .B2(new_n649), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n648), .A2(new_n226), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n932), .B1(new_n926), .B2(new_n933), .ZN(new_n934));
  XNOR2_X1  g733(.A(new_n934), .B(KEYINPUT121), .ZN(G1349gat));
  NAND4_X1  g734(.A1(new_n927), .A2(new_n273), .A3(new_n274), .A4(new_n675), .ZN(new_n936));
  OAI21_X1  g735(.A(G183gat), .B1(new_n929), .B2(new_n755), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT60), .ZN(new_n938));
  AOI22_X1  g737(.A1(new_n936), .A2(new_n937), .B1(KEYINPUT122), .B2(new_n938), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n938), .A2(KEYINPUT122), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n939), .B(new_n940), .ZN(G1350gat));
  OAI21_X1  g740(.A(G190gat), .B1(new_n929), .B2(new_n692), .ZN(new_n942));
  XNOR2_X1  g741(.A(new_n942), .B(KEYINPUT61), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n927), .A2(new_n264), .A3(new_n594), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(G1351gat));
  NAND2_X1  g744(.A1(new_n925), .A2(new_n892), .ZN(new_n946));
  NOR3_X1   g745(.A1(new_n946), .A2(G197gat), .A3(new_n676), .ZN(new_n947));
  XOR2_X1   g746(.A(new_n947), .B(KEYINPUT123), .Z(new_n948));
  NAND2_X1  g747(.A1(new_n664), .A2(new_n924), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n949), .B1(new_n909), .B2(new_n910), .ZN(new_n950));
  INV_X1    g749(.A(new_n950), .ZN(new_n951));
  OAI21_X1  g750(.A(G197gat), .B1(new_n951), .B2(new_n676), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n948), .A2(new_n952), .ZN(G1352gat));
  NOR3_X1   g752(.A1(new_n946), .A2(G204gat), .A3(new_n649), .ZN(new_n954));
  XNOR2_X1  g753(.A(new_n954), .B(KEYINPUT62), .ZN(new_n955));
  OAI21_X1  g754(.A(G204gat), .B1(new_n951), .B2(new_n649), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n955), .A2(new_n956), .ZN(G1353gat));
  INV_X1    g756(.A(KEYINPUT125), .ZN(new_n958));
  INV_X1    g757(.A(G211gat), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n959), .B1(new_n950), .B2(new_n675), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n958), .B1(new_n960), .B2(KEYINPUT63), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n905), .B1(new_n904), .B2(new_n881), .ZN(new_n962));
  NOR3_X1   g761(.A1(new_n907), .A2(KEYINPUT120), .A3(KEYINPUT57), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n910), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  INV_X1    g763(.A(new_n949), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n964), .A2(new_n675), .A3(new_n965), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n966), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n967), .A2(KEYINPUT124), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT63), .ZN(new_n969));
  AOI211_X1 g768(.A(new_n755), .B(new_n949), .C1(new_n909), .C2(new_n910), .ZN(new_n970));
  OAI211_X1 g769(.A(KEYINPUT125), .B(new_n969), .C1(new_n970), .C2(new_n959), .ZN(new_n971));
  INV_X1    g770(.A(KEYINPUT124), .ZN(new_n972));
  NAND4_X1  g771(.A1(new_n966), .A2(new_n972), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n973));
  NAND4_X1  g772(.A1(new_n961), .A2(new_n968), .A3(new_n971), .A4(new_n973), .ZN(new_n974));
  NAND4_X1  g773(.A1(new_n925), .A2(new_n959), .A3(new_n675), .A4(new_n892), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n976), .A2(KEYINPUT126), .ZN(new_n977));
  INV_X1    g776(.A(KEYINPUT126), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n974), .A2(new_n978), .A3(new_n975), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n977), .A2(new_n979), .ZN(G1354gat));
  OAI21_X1  g779(.A(G218gat), .B1(new_n951), .B2(new_n692), .ZN(new_n981));
  OR2_X1    g780(.A1(new_n692), .A2(G218gat), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n981), .B1(new_n946), .B2(new_n982), .ZN(G1355gat));
endmodule


