//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 0 1 1 0 0 1 0 0 1 0 0 1 0 0 0 1 0 0 0 0 1 0 0 0 0 0 1 0 1 0 1 1 1 1 1 0 1 1 1 1 0 0 0 0 0 0 0 1 1 0 0 1 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n636, new_n637,
    new_n638, new_n640, new_n641, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n669, new_n670, new_n671, new_n673, new_n674, new_n675, new_n677,
    new_n678, new_n679, new_n680, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n811, new_n812, new_n814,
    new_n815, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n893, new_n894, new_n895,
    new_n896, new_n898, new_n899, new_n900, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n914, new_n915, new_n916, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n935, new_n936, new_n937,
    new_n938, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n948, new_n949, new_n950, new_n951;
  XNOR2_X1  g000(.A(G43gat), .B(G50gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT87), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(KEYINPUT15), .ZN(new_n205));
  NAND2_X1  g004(.A1(G29gat), .A2(G36gat), .ZN(new_n206));
  OAI21_X1  g005(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  NOR3_X1   g007(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n206), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n205), .A2(new_n210), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n202), .A2(KEYINPUT15), .ZN(new_n212));
  AOI21_X1  g011(.A(new_n212), .B1(new_n204), .B2(KEYINPUT15), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n211), .B1(new_n213), .B2(new_n210), .ZN(new_n214));
  XOR2_X1   g013(.A(new_n214), .B(KEYINPUT17), .Z(new_n215));
  INV_X1    g014(.A(KEYINPUT16), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n216), .A2(G1gat), .ZN(new_n217));
  XNOR2_X1  g016(.A(G15gat), .B(G22gat), .ZN(new_n218));
  MUX2_X1   g017(.A(G1gat), .B(new_n217), .S(new_n218), .Z(new_n219));
  XNOR2_X1  g018(.A(new_n219), .B(G8gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n215), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(G229gat), .A2(G233gat), .ZN(new_n222));
  OR2_X1    g021(.A1(new_n214), .A2(new_n220), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT18), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND4_X1  g025(.A1(new_n221), .A2(KEYINPUT18), .A3(new_n222), .A4(new_n223), .ZN(new_n227));
  XNOR2_X1  g026(.A(new_n214), .B(new_n220), .ZN(new_n228));
  XOR2_X1   g027(.A(new_n222), .B(KEYINPUT13), .Z(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n226), .A2(new_n227), .A3(new_n230), .ZN(new_n231));
  XNOR2_X1  g030(.A(G113gat), .B(G141gat), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n232), .B(KEYINPUT11), .ZN(new_n233));
  INV_X1    g032(.A(G169gat), .ZN(new_n234));
  XNOR2_X1  g033(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(new_n235), .B(G197gat), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n236), .B(KEYINPUT12), .ZN(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n231), .A2(new_n238), .ZN(new_n239));
  NAND4_X1  g038(.A1(new_n226), .A2(new_n227), .A3(new_n230), .A4(new_n237), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(KEYINPUT77), .B(KEYINPUT6), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(G120gat), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(G113gat), .ZN(new_n246));
  INV_X1    g045(.A(G113gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(G120gat), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n246), .A2(new_n248), .A3(KEYINPUT68), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT1), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  AOI21_X1  g050(.A(KEYINPUT68), .B1(new_n246), .B2(new_n248), .ZN(new_n252));
  INV_X1    g051(.A(G127gat), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n253), .A2(G134gat), .ZN(new_n254));
  INV_X1    g053(.A(G134gat), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n255), .A2(G127gat), .ZN(new_n256));
  OAI22_X1  g055(.A1(new_n251), .A2(new_n252), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT75), .ZN(new_n258));
  INV_X1    g057(.A(G148gat), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n258), .A2(new_n259), .A3(G141gat), .ZN(new_n260));
  INV_X1    g059(.A(G141gat), .ZN(new_n261));
  AOI21_X1  g060(.A(KEYINPUT75), .B1(new_n261), .B2(G148gat), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n261), .A2(G148gat), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n260), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NOR2_X1   g063(.A1(G155gat), .A2(G162gat), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT2), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  AND2_X1   g066(.A1(G155gat), .A2(G162gat), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n259), .A2(G141gat), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n266), .B1(new_n263), .B2(new_n271), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n268), .A2(new_n265), .ZN(new_n273));
  AOI22_X1  g072(.A1(new_n264), .A2(new_n270), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT69), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n275), .A2(new_n245), .A3(G113gat), .ZN(new_n276));
  AOI21_X1  g075(.A(KEYINPUT69), .B1(new_n247), .B2(G120gat), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n247), .A2(G120gat), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n276), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(G127gat), .B(G134gat), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT70), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  OAI21_X1  g081(.A(KEYINPUT70), .B1(new_n254), .B2(new_n256), .ZN(new_n283));
  NAND4_X1  g082(.A1(new_n279), .A2(new_n282), .A3(new_n283), .A4(new_n250), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n257), .A2(new_n274), .A3(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT4), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n257), .A2(new_n284), .ZN(new_n288));
  XNOR2_X1  g087(.A(G141gat), .B(G148gat), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n273), .B1(new_n289), .B2(KEYINPUT2), .ZN(new_n290));
  XNOR2_X1  g089(.A(KEYINPUT76), .B(KEYINPUT3), .ZN(new_n291));
  NOR3_X1   g090(.A1(new_n261), .A2(KEYINPUT75), .A3(G148gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n259), .A2(G141gat), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n258), .B1(new_n259), .B2(G141gat), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n292), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n268), .B1(new_n266), .B2(new_n265), .ZN(new_n296));
  OAI211_X1 g095(.A(new_n290), .B(new_n291), .C1(new_n295), .C2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n294), .A2(new_n293), .ZN(new_n298));
  AOI22_X1  g097(.A1(new_n298), .A2(new_n260), .B1(new_n269), .B2(new_n267), .ZN(new_n299));
  XNOR2_X1  g098(.A(G155gat), .B(G162gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n261), .A2(G148gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n293), .A2(new_n301), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n300), .B1(new_n266), .B2(new_n302), .ZN(new_n303));
  OAI21_X1  g102(.A(KEYINPUT3), .B1(new_n299), .B2(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n288), .A2(new_n297), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(G225gat), .A2(G233gat), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n257), .A2(new_n274), .A3(KEYINPUT4), .A4(new_n284), .ZN(new_n307));
  NAND4_X1  g106(.A1(new_n287), .A2(new_n305), .A3(new_n306), .A4(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT5), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(new_n306), .ZN(new_n312));
  INV_X1    g111(.A(new_n285), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n274), .B1(new_n257), .B2(new_n284), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n312), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n309), .B1(new_n308), .B2(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(G1gat), .B(G29gat), .ZN(new_n317));
  XNOR2_X1  g116(.A(new_n317), .B(KEYINPUT0), .ZN(new_n318));
  XNOR2_X1  g117(.A(G57gat), .B(G85gat), .ZN(new_n319));
  XNOR2_X1  g118(.A(new_n318), .B(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  NOR3_X1   g120(.A1(new_n311), .A2(new_n316), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n308), .A2(new_n315), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(KEYINPUT5), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n320), .B1(new_n324), .B2(new_n310), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n244), .B1(new_n322), .B2(new_n325), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n324), .A2(new_n320), .A3(new_n310), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(new_n243), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(G183gat), .A2(G190gat), .ZN(new_n330));
  AOI21_X1  g129(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n331));
  INV_X1    g130(.A(G176gat), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n331), .B1(new_n234), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n234), .A2(new_n332), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n334), .A2(KEYINPUT26), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n330), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  XOR2_X1   g135(.A(KEYINPUT67), .B(KEYINPUT28), .Z(new_n337));
  XNOR2_X1  g136(.A(KEYINPUT27), .B(G183gat), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT66), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT27), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n339), .B1(new_n341), .B2(G183gat), .ZN(new_n342));
  INV_X1    g141(.A(G190gat), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n337), .B1(new_n340), .B2(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n338), .A2(KEYINPUT28), .A3(new_n343), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n336), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT25), .ZN(new_n348));
  NAND3_X1  g147(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT64), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND4_X1  g150(.A1(KEYINPUT64), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n352));
  OAI21_X1  g151(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n353));
  AOI22_X1  g152(.A1(new_n351), .A2(new_n352), .B1(new_n330), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(KEYINPUT65), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT23), .ZN(new_n357));
  NOR3_X1   g156(.A1(new_n357), .A2(G169gat), .A3(G176gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(G169gat), .A2(G176gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(KEYINPUT23), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n358), .B1(new_n334), .B2(new_n360), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n361), .B1(new_n354), .B2(KEYINPUT65), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n348), .B1(new_n356), .B2(new_n362), .ZN(new_n363));
  AND2_X1   g162(.A1(new_n361), .A2(KEYINPUT25), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n353), .A2(new_n330), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(new_n349), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n347), .B1(new_n363), .B2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(G226gat), .ZN(new_n369));
  INV_X1    g168(.A(G233gat), .ZN(new_n370));
  OAI22_X1  g169(.A1(new_n368), .A2(KEYINPUT29), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n369), .A2(new_n370), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n351), .A2(new_n352), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(new_n365), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT65), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n376), .A2(new_n355), .A3(new_n361), .ZN(new_n377));
  AOI22_X1  g176(.A1(new_n377), .A2(new_n348), .B1(new_n366), .B2(new_n364), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n372), .B1(new_n378), .B2(new_n347), .ZN(new_n379));
  NAND2_X1  g178(.A1(G211gat), .A2(G218gat), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT22), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(G204gat), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(G197gat), .ZN(new_n384));
  INV_X1    g183(.A(G197gat), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(G204gat), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n382), .A2(new_n384), .A3(new_n386), .ZN(new_n387));
  XOR2_X1   g186(.A(G211gat), .B(G218gat), .Z(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  XNOR2_X1  g188(.A(G211gat), .B(G218gat), .ZN(new_n390));
  XNOR2_X1  g189(.A(G197gat), .B(G204gat), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n390), .A2(new_n391), .A3(new_n382), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n389), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n371), .A2(new_n379), .A3(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT74), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND4_X1  g195(.A1(new_n371), .A2(new_n379), .A3(KEYINPUT74), .A4(new_n393), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n371), .A2(new_n379), .ZN(new_n398));
  INV_X1    g197(.A(new_n393), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n396), .A2(new_n397), .A3(new_n400), .ZN(new_n401));
  XNOR2_X1  g200(.A(G8gat), .B(G36gat), .ZN(new_n402));
  XNOR2_X1  g201(.A(G64gat), .B(G92gat), .ZN(new_n403));
  XNOR2_X1  g202(.A(new_n402), .B(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(new_n404), .ZN(new_n406));
  NAND4_X1  g205(.A1(new_n396), .A2(new_n400), .A3(new_n397), .A4(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n405), .A2(KEYINPUT30), .A3(new_n407), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n393), .B1(new_n371), .B2(new_n379), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n409), .B1(new_n395), .B2(new_n394), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT30), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n410), .A2(new_n411), .A3(new_n397), .A4(new_n406), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n329), .B1(new_n408), .B2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(G22gat), .ZN(new_n414));
  NAND2_X1  g213(.A1(G228gat), .A2(G233gat), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT29), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n387), .A2(new_n388), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n390), .B1(new_n382), .B2(new_n391), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n416), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n274), .B1(new_n419), .B2(new_n291), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n393), .B1(new_n297), .B2(new_n416), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n415), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT80), .ZN(new_n423));
  AND3_X1   g222(.A1(new_n297), .A2(new_n423), .A3(new_n416), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n423), .B1(new_n297), .B2(new_n416), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n399), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n304), .A2(G228gat), .A3(G233gat), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n419), .A2(new_n274), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  AOI22_X1  g228(.A1(KEYINPUT79), .A2(new_n422), .B1(new_n426), .B2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT79), .ZN(new_n431));
  OAI211_X1 g230(.A(new_n431), .B(new_n415), .C1(new_n420), .C2(new_n421), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n414), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n422), .A2(KEYINPUT79), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n426), .A2(new_n429), .ZN(new_n435));
  AND4_X1   g234(.A1(new_n414), .A2(new_n434), .A3(new_n435), .A4(new_n432), .ZN(new_n436));
  NOR3_X1   g235(.A1(new_n433), .A2(new_n436), .A3(KEYINPUT81), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT81), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n434), .A2(new_n435), .A3(new_n432), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(G22gat), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n430), .A2(new_n414), .A3(new_n432), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n439), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  XOR2_X1   g242(.A(G78gat), .B(G106gat), .Z(new_n444));
  XNOR2_X1  g243(.A(new_n444), .B(KEYINPUT78), .ZN(new_n445));
  XOR2_X1   g244(.A(KEYINPUT31), .B(G50gat), .Z(new_n446));
  XNOR2_X1  g245(.A(new_n445), .B(new_n446), .ZN(new_n447));
  NOR3_X1   g246(.A1(new_n443), .A2(KEYINPUT82), .A3(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT82), .ZN(new_n449));
  OAI21_X1  g248(.A(KEYINPUT81), .B1(new_n433), .B2(new_n436), .ZN(new_n450));
  INV_X1    g249(.A(new_n447), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n449), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n438), .B1(new_n448), .B2(new_n452), .ZN(new_n453));
  OAI21_X1  g252(.A(KEYINPUT82), .B1(new_n443), .B2(new_n447), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n450), .A2(new_n449), .A3(new_n451), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n454), .A2(new_n455), .A3(new_n437), .ZN(new_n456));
  INV_X1    g255(.A(new_n288), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n457), .B1(new_n378), .B2(new_n347), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n368), .A2(new_n288), .ZN(new_n459));
  AND2_X1   g258(.A1(G227gat), .A2(G233gat), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n458), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(KEYINPUT32), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT33), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  XOR2_X1   g263(.A(G15gat), .B(G43gat), .Z(new_n465));
  XNOR2_X1  g264(.A(G71gat), .B(G99gat), .ZN(new_n466));
  XNOR2_X1  g265(.A(new_n465), .B(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n462), .A2(new_n464), .A3(new_n467), .ZN(new_n468));
  XOR2_X1   g267(.A(new_n467), .B(KEYINPUT71), .Z(new_n469));
  OAI211_X1 g268(.A(new_n461), .B(KEYINPUT32), .C1(new_n463), .C2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT72), .ZN(new_n472));
  AND2_X1   g271(.A1(new_n458), .A2(new_n459), .ZN(new_n473));
  OAI211_X1 g272(.A(new_n472), .B(KEYINPUT34), .C1(new_n473), .C2(new_n460), .ZN(new_n474));
  AOI211_X1 g273(.A(KEYINPUT34), .B(new_n460), .C1(new_n458), .C2(new_n459), .ZN(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n460), .B1(new_n458), .B2(new_n459), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT34), .ZN(new_n478));
  OAI21_X1  g277(.A(KEYINPUT72), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n474), .A2(new_n476), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n471), .A2(new_n480), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n477), .A2(new_n478), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n475), .B1(new_n482), .B2(new_n472), .ZN(new_n483));
  NAND4_X1  g282(.A1(new_n483), .A2(new_n479), .A3(new_n470), .A4(new_n468), .ZN(new_n484));
  AND2_X1   g283(.A1(new_n481), .A2(new_n484), .ZN(new_n485));
  NAND4_X1  g284(.A1(new_n413), .A2(new_n453), .A3(new_n456), .A4(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(KEYINPUT35), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(KEYINPUT86), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT86), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n486), .A2(new_n489), .A3(KEYINPUT35), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n407), .A2(KEYINPUT30), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n406), .B1(new_n410), .B2(new_n397), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n412), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(KEYINPUT83), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT35), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT83), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n408), .A2(new_n496), .A3(new_n412), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n494), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(new_n329), .ZN(new_n499));
  NAND4_X1  g298(.A1(new_n453), .A2(new_n485), .A3(new_n499), .A4(new_n456), .ZN(new_n500));
  OR2_X1    g299(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n488), .A2(new_n490), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n494), .A2(new_n497), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n287), .A2(new_n305), .A3(new_n307), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(new_n312), .ZN(new_n505));
  OR2_X1    g304(.A1(new_n313), .A2(new_n314), .ZN(new_n506));
  OAI211_X1 g305(.A(new_n505), .B(KEYINPUT39), .C1(new_n312), .C2(new_n506), .ZN(new_n507));
  OAI211_X1 g306(.A(new_n507), .B(new_n321), .C1(KEYINPUT39), .C2(new_n505), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT40), .ZN(new_n509));
  AND2_X1   g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n508), .A2(new_n509), .ZN(new_n511));
  NOR3_X1   g310(.A1(new_n510), .A2(new_n511), .A3(new_n322), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n503), .A2(new_n512), .ZN(new_n513));
  AND2_X1   g312(.A1(new_n453), .A2(new_n456), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT84), .ZN(new_n515));
  AND2_X1   g314(.A1(new_n400), .A2(new_n394), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT37), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n517), .B1(new_n400), .B2(new_n394), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(KEYINPUT84), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n410), .A2(new_n517), .A3(new_n397), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n406), .A2(KEYINPUT38), .ZN(new_n522));
  NAND4_X1  g321(.A1(new_n518), .A2(new_n520), .A3(new_n521), .A4(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(KEYINPUT85), .ZN(new_n524));
  AOI211_X1 g323(.A(KEYINPUT38), .B(new_n406), .C1(new_n519), .C2(KEYINPUT84), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT85), .ZN(new_n526));
  NAND4_X1  g325(.A1(new_n525), .A2(new_n526), .A3(new_n518), .A4(new_n521), .ZN(new_n527));
  AND2_X1   g326(.A1(new_n329), .A2(new_n407), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n521), .A2(new_n404), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n517), .B1(new_n410), .B2(new_n397), .ZN(new_n530));
  OAI21_X1  g329(.A(KEYINPUT38), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND4_X1  g330(.A1(new_n524), .A2(new_n527), .A3(new_n528), .A4(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n513), .A2(new_n514), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n481), .A2(new_n484), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT73), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n534), .A2(new_n535), .A3(KEYINPUT36), .ZN(new_n536));
  XNOR2_X1  g335(.A(KEYINPUT73), .B(KEYINPUT36), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n481), .A2(new_n484), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n453), .A2(new_n456), .ZN(new_n540));
  INV_X1    g339(.A(new_n413), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n533), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n242), .B1(new_n502), .B2(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(G57gat), .B(G64gat), .ZN(new_n545));
  AOI21_X1  g344(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n546));
  OR2_X1    g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  XOR2_X1   g346(.A(G71gat), .B(G78gat), .Z(new_n548));
  OR2_X1    g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n547), .A2(new_n548), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT21), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(G231gat), .A2(G233gat), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n553), .B(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(G127gat), .B(G155gat), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n555), .B(new_n556), .ZN(new_n557));
  XOR2_X1   g356(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n558));
  XNOR2_X1  g357(.A(new_n557), .B(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n551), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(KEYINPUT21), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(new_n220), .ZN(new_n562));
  XOR2_X1   g361(.A(new_n559), .B(new_n562), .Z(new_n563));
  XOR2_X1   g362(.A(G183gat), .B(G211gat), .Z(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n559), .B(new_n562), .ZN(new_n566));
  INV_X1    g365(.A(new_n564), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  AOI21_X1  g369(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n571), .B(KEYINPUT88), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n572), .B(KEYINPUT89), .ZN(new_n573));
  XNOR2_X1  g372(.A(G134gat), .B(G162gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n574), .B(KEYINPUT90), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n573), .B(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n577));
  NAND3_X1  g376(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT7), .ZN(new_n579));
  NAND2_X1  g378(.A1(G85gat), .A2(G92gat), .ZN(new_n580));
  NAND2_X1  g379(.A1(G99gat), .A2(G106gat), .ZN(new_n581));
  AOI22_X1  g380(.A1(new_n579), .A2(new_n580), .B1(new_n581), .B2(KEYINPUT8), .ZN(new_n582));
  XOR2_X1   g381(.A(KEYINPUT91), .B(G85gat), .Z(new_n583));
  OAI211_X1 g382(.A(new_n578), .B(new_n582), .C1(new_n583), .C2(G92gat), .ZN(new_n584));
  XOR2_X1   g383(.A(G99gat), .B(G106gat), .Z(new_n585));
  AND2_X1   g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(KEYINPUT92), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT92), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  OR2_X1    g389(.A1(new_n584), .A2(new_n585), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n588), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n577), .B1(new_n592), .B2(new_n214), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n593), .B1(new_n215), .B2(new_n592), .ZN(new_n594));
  XNOR2_X1  g393(.A(G190gat), .B(G218gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(KEYINPUT93), .ZN(new_n596));
  OR2_X1    g395(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n576), .B1(new_n597), .B2(KEYINPUT94), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n594), .A2(new_n596), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  OAI211_X1 g400(.A(new_n597), .B(new_n599), .C1(KEYINPUT94), .C2(new_n576), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(G230gat), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n604), .A2(new_n370), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n592), .A2(new_n551), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT10), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n560), .A2(new_n587), .A3(new_n591), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  OR3_X1    g408(.A1(new_n592), .A2(new_n607), .A3(new_n551), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n605), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n606), .A2(new_n608), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n613), .A2(new_n605), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(G120gat), .B(G148gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(G176gat), .B(G204gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n616), .B(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n615), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n618), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n612), .A2(new_n614), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  NOR3_X1   g421(.A1(new_n570), .A2(new_n603), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n544), .A2(new_n623), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n624), .A2(new_n499), .ZN(new_n625));
  XOR2_X1   g424(.A(new_n625), .B(G1gat), .Z(G1324gat));
  INV_X1    g425(.A(new_n503), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  XOR2_X1   g427(.A(KEYINPUT16), .B(G8gat), .Z(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT42), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(KEYINPUT95), .ZN(new_n633));
  INV_X1    g432(.A(G8gat), .ZN(new_n634));
  OAI221_X1 g433(.A(new_n633), .B1(new_n631), .B2(new_n630), .C1(new_n634), .C2(new_n628), .ZN(G1325gat));
  INV_X1    g434(.A(new_n539), .ZN(new_n636));
  OAI21_X1  g435(.A(G15gat), .B1(new_n624), .B2(new_n636), .ZN(new_n637));
  OR2_X1    g436(.A1(new_n534), .A2(G15gat), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n637), .B1(new_n624), .B2(new_n638), .ZN(G1326gat));
  NOR2_X1   g438(.A1(new_n624), .A2(new_n514), .ZN(new_n640));
  XOR2_X1   g439(.A(KEYINPUT43), .B(G22gat), .Z(new_n641));
  XNOR2_X1  g440(.A(new_n640), .B(new_n641), .ZN(G1327gat));
  AND3_X1   g441(.A1(new_n486), .A2(new_n489), .A3(KEYINPUT35), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n489), .B1(new_n486), .B2(KEYINPUT35), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n498), .A2(new_n500), .ZN(new_n645));
  NOR3_X1   g444(.A1(new_n643), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  OAI211_X1 g445(.A(new_n538), .B(new_n536), .C1(new_n514), .C2(new_n413), .ZN(new_n647));
  AND2_X1   g446(.A1(new_n532), .A2(new_n514), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n647), .B1(new_n648), .B2(new_n513), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n603), .B1(new_n646), .B2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT97), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n650), .A2(new_n651), .A3(KEYINPUT44), .ZN(new_n652));
  INV_X1    g451(.A(new_n603), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n653), .B1(new_n502), .B2(new_n543), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT44), .ZN(new_n655));
  OAI21_X1  g454(.A(KEYINPUT97), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  AOI22_X1  g455(.A1(new_n652), .A2(new_n656), .B1(new_n655), .B2(new_n654), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n569), .B(KEYINPUT96), .ZN(new_n658));
  INV_X1    g457(.A(new_n622), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n658), .A2(new_n241), .A3(new_n659), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  OAI21_X1  g461(.A(G29gat), .B1(new_n662), .B2(new_n499), .ZN(new_n663));
  NOR3_X1   g462(.A1(new_n569), .A2(new_n653), .A3(new_n622), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n544), .A2(new_n664), .ZN(new_n665));
  NOR3_X1   g464(.A1(new_n665), .A2(G29gat), .A3(new_n499), .ZN(new_n666));
  XOR2_X1   g465(.A(new_n666), .B(KEYINPUT45), .Z(new_n667));
  NAND2_X1  g466(.A1(new_n663), .A2(new_n667), .ZN(G1328gat));
  OAI21_X1  g467(.A(G36gat), .B1(new_n662), .B2(new_n627), .ZN(new_n669));
  NOR3_X1   g468(.A1(new_n665), .A2(G36gat), .A3(new_n627), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(KEYINPUT46), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n669), .A2(new_n671), .ZN(G1329gat));
  NAND3_X1  g471(.A1(new_n661), .A2(G43gat), .A3(new_n539), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n665), .A2(new_n534), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n673), .B1(G43gat), .B2(new_n674), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g475(.A(new_n665), .ZN(new_n677));
  AOI21_X1  g476(.A(G50gat), .B1(new_n677), .B2(new_n540), .ZN(new_n678));
  AND2_X1   g477(.A1(new_n540), .A2(G50gat), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n678), .B1(new_n661), .B2(new_n679), .ZN(new_n680));
  XOR2_X1   g479(.A(new_n680), .B(KEYINPUT48), .Z(G1331gat));
  NAND3_X1  g480(.A1(new_n569), .A2(new_n242), .A3(new_n653), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n682), .A2(new_n659), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n502), .A2(new_n543), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n686), .A2(new_n329), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g487(.A(new_n685), .B(KEYINPUT98), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n627), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g490(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n692));
  XOR2_X1   g491(.A(new_n692), .B(KEYINPUT99), .Z(new_n693));
  XNOR2_X1  g492(.A(new_n691), .B(new_n693), .ZN(G1333gat));
  AND3_X1   g493(.A1(new_n689), .A2(G71gat), .A3(new_n539), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(KEYINPUT100), .ZN(new_n696));
  AOI21_X1  g495(.A(G71gat), .B1(new_n686), .B2(new_n485), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT100), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n696), .B1(new_n695), .B2(new_n699), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g500(.A1(new_n689), .A2(new_n540), .ZN(new_n702));
  XNOR2_X1  g501(.A(KEYINPUT101), .B(G78gat), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n702), .B(new_n703), .ZN(G1335gat));
  NOR2_X1   g503(.A1(new_n569), .A2(new_n241), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(new_n622), .ZN(new_n706));
  OAI21_X1  g505(.A(KEYINPUT102), .B1(new_n657), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n654), .A2(new_n655), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n651), .B1(new_n650), .B2(KEYINPUT44), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n654), .A2(KEYINPUT97), .A3(new_n655), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n708), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT102), .ZN(new_n712));
  INV_X1    g511(.A(new_n706), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n711), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n707), .A2(new_n714), .A3(new_n329), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(new_n583), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n684), .A2(new_n603), .A3(new_n705), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT51), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n717), .B(new_n718), .ZN(new_n719));
  NOR3_X1   g518(.A1(new_n659), .A2(new_n499), .A3(new_n583), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n716), .A2(new_n721), .ZN(G1336gat));
  NOR3_X1   g521(.A1(new_n627), .A2(new_n659), .A3(G92gat), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n719), .A2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT52), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(G92gat), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n711), .A2(new_n503), .A3(new_n713), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n727), .B1(new_n728), .B2(KEYINPUT104), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT104), .ZN(new_n730));
  NAND4_X1  g529(.A1(new_n711), .A2(new_n730), .A3(new_n503), .A4(new_n713), .ZN(new_n731));
  AOI211_X1 g530(.A(KEYINPUT105), .B(new_n726), .C1(new_n729), .C2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT105), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n728), .A2(KEYINPUT104), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n734), .A2(G92gat), .A3(new_n731), .ZN(new_n735));
  INV_X1    g534(.A(new_n726), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n733), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT103), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n724), .A2(new_n738), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n719), .A2(KEYINPUT103), .A3(new_n723), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n707), .A2(new_n714), .A3(new_n503), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n741), .B1(G92gat), .B2(new_n742), .ZN(new_n743));
  OAI22_X1  g542(.A1(new_n732), .A2(new_n737), .B1(new_n725), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(KEYINPUT106), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT106), .ZN(new_n746));
  OAI221_X1 g545(.A(new_n746), .B1(new_n743), .B2(new_n725), .C1(new_n732), .C2(new_n737), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n745), .A2(new_n747), .ZN(G1337gat));
  NOR3_X1   g547(.A1(new_n659), .A2(G99gat), .A3(new_n534), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(KEYINPUT108), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n719), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n707), .A2(new_n714), .A3(new_n539), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT107), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(G99gat), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n752), .A2(new_n753), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n751), .B1(new_n755), .B2(new_n756), .ZN(G1338gat));
  INV_X1    g556(.A(G106gat), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n719), .A2(new_n758), .A3(new_n540), .A4(new_n622), .ZN(new_n759));
  AND3_X1   g558(.A1(new_n707), .A2(new_n714), .A3(new_n540), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n759), .B1(new_n760), .B2(new_n758), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(KEYINPUT53), .ZN(new_n762));
  OR2_X1    g561(.A1(new_n762), .A2(KEYINPUT109), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(KEYINPUT109), .ZN(new_n764));
  XNOR2_X1  g563(.A(KEYINPUT110), .B(KEYINPUT53), .ZN(new_n765));
  NOR3_X1   g564(.A1(new_n657), .A2(new_n514), .A3(new_n706), .ZN(new_n766));
  OAI211_X1 g565(.A(new_n759), .B(new_n765), .C1(new_n766), .C2(new_n758), .ZN(new_n767));
  XOR2_X1   g566(.A(new_n767), .B(KEYINPUT111), .Z(new_n768));
  NAND3_X1  g567(.A1(new_n763), .A2(new_n764), .A3(new_n768), .ZN(G1339gat));
  AOI21_X1  g568(.A(new_n222), .B1(new_n221), .B2(new_n223), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n228), .A2(new_n229), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n236), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n240), .A2(new_n772), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n773), .B1(new_n602), .B2(new_n601), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n609), .A2(new_n610), .A3(new_n605), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n612), .A2(KEYINPUT54), .A3(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT54), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n620), .B1(new_n611), .B2(new_n777), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n776), .A2(KEYINPUT55), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(new_n621), .ZN(new_n780));
  INV_X1    g579(.A(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n776), .A2(new_n778), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT55), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n774), .A2(new_n781), .A3(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(KEYINPUT112), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT112), .ZN(new_n787));
  NAND4_X1  g586(.A1(new_n774), .A2(new_n787), .A3(new_n781), .A4(new_n784), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n659), .A2(new_n773), .ZN(new_n790));
  INV_X1    g589(.A(new_n790), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n781), .A2(new_n241), .A3(new_n784), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n603), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  OAI21_X1  g592(.A(KEYINPUT113), .B1(new_n789), .B2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(new_n793), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT113), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n795), .A2(new_n796), .A3(new_n786), .A4(new_n788), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n794), .A2(new_n658), .A3(new_n797), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n682), .A2(new_n622), .ZN(new_n799));
  INV_X1    g598(.A(new_n799), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n540), .B1(new_n798), .B2(new_n800), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n534), .A2(new_n499), .ZN(new_n802));
  AND2_X1   g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(new_n627), .ZN(new_n804));
  XNOR2_X1  g603(.A(new_n804), .B(KEYINPUT115), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n805), .A2(new_n247), .A3(new_n241), .ZN(new_n806));
  XOR2_X1   g605(.A(new_n801), .B(KEYINPUT114), .Z(new_n807));
  NAND3_X1  g606(.A1(new_n807), .A2(new_n627), .A3(new_n802), .ZN(new_n808));
  OAI21_X1  g607(.A(G113gat), .B1(new_n808), .B2(new_n242), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n806), .A2(new_n809), .ZN(G1340gat));
  NAND3_X1  g609(.A1(new_n805), .A2(new_n245), .A3(new_n622), .ZN(new_n811));
  OAI21_X1  g610(.A(G120gat), .B1(new_n808), .B2(new_n659), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(G1341gat));
  OAI21_X1  g612(.A(G127gat), .B1(new_n808), .B2(new_n658), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n569), .A2(new_n253), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n814), .B1(new_n804), .B2(new_n815), .ZN(G1342gat));
  NOR2_X1   g615(.A1(new_n653), .A2(new_n503), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n803), .A2(new_n255), .A3(new_n817), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n818), .A2(KEYINPUT56), .ZN(new_n819));
  XOR2_X1   g618(.A(new_n819), .B(KEYINPUT116), .Z(new_n820));
  OAI21_X1  g619(.A(G134gat), .B1(new_n808), .B2(new_n653), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n818), .A2(KEYINPUT56), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n820), .A2(new_n821), .A3(new_n822), .ZN(G1343gat));
  AOI21_X1  g622(.A(new_n514), .B1(new_n798), .B2(new_n800), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT57), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n539), .A2(new_n499), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(new_n627), .ZN(new_n828));
  INV_X1    g627(.A(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n826), .A2(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT117), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n782), .A2(new_n831), .A3(new_n783), .ZN(new_n832));
  INV_X1    g631(.A(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n831), .B1(new_n782), .B2(new_n783), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n781), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT118), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  OAI211_X1 g636(.A(KEYINPUT118), .B(new_n781), .C1(new_n833), .C2(new_n834), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n837), .A2(new_n241), .A3(new_n838), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n603), .B1(new_n839), .B2(new_n791), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n570), .B1(new_n840), .B2(new_n789), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(new_n800), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n825), .B1(new_n842), .B2(new_n540), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n830), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(new_n241), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(G141gat), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n824), .A2(new_n827), .ZN(new_n847));
  XNOR2_X1  g646(.A(new_n847), .B(KEYINPUT119), .ZN(new_n848));
  NAND4_X1  g647(.A1(new_n848), .A2(new_n261), .A3(new_n241), .A4(new_n627), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT58), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n846), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  NOR4_X1   g650(.A1(new_n847), .A2(G141gat), .A3(new_n242), .A4(new_n503), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n852), .B1(new_n845), .B2(G141gat), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n851), .B1(new_n850), .B2(new_n853), .ZN(G1344gat));
  XNOR2_X1  g653(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n798), .A2(new_n800), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n856), .A2(KEYINPUT57), .A3(new_n540), .ZN(new_n857));
  INV_X1    g656(.A(new_n785), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n570), .B1(new_n840), .B2(new_n858), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n514), .B1(new_n859), .B2(new_n800), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n857), .B1(KEYINPUT57), .B2(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT121), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n861), .A2(new_n862), .A3(new_n622), .A4(new_n829), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(G148gat), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n838), .A2(new_n241), .ZN(new_n865));
  INV_X1    g664(.A(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n790), .B1(new_n866), .B2(new_n837), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n785), .B1(new_n867), .B2(new_n603), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n799), .B1(new_n868), .B2(new_n570), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n825), .B1(new_n869), .B2(new_n514), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n659), .B1(new_n870), .B2(new_n857), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n862), .B1(new_n871), .B2(new_n829), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n855), .B1(new_n864), .B2(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT59), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(G148gat), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n875), .B1(new_n844), .B2(new_n622), .ZN(new_n876));
  INV_X1    g675(.A(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n873), .A2(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT122), .ZN(new_n879));
  INV_X1    g678(.A(new_n848), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n880), .A2(new_n503), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n881), .A2(new_n259), .A3(new_n622), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n878), .A2(new_n879), .A3(new_n882), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n860), .A2(KEYINPUT57), .ZN(new_n884));
  AOI211_X1 g683(.A(new_n825), .B(new_n514), .C1(new_n798), .C2(new_n800), .ZN(new_n885));
  OAI211_X1 g684(.A(new_n622), .B(new_n829), .C1(new_n884), .C2(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(KEYINPUT121), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n887), .A2(G148gat), .A3(new_n863), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n876), .B1(new_n888), .B2(new_n855), .ZN(new_n889));
  NOR4_X1   g688(.A1(new_n880), .A2(G148gat), .A3(new_n503), .A4(new_n659), .ZN(new_n890));
  OAI21_X1  g689(.A(KEYINPUT122), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n883), .A2(new_n891), .ZN(G1345gat));
  INV_X1    g691(.A(G155gat), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n881), .A2(new_n893), .A3(new_n569), .ZN(new_n894));
  INV_X1    g693(.A(new_n844), .ZN(new_n895));
  OAI21_X1  g694(.A(G155gat), .B1(new_n895), .B2(new_n658), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n894), .A2(new_n896), .ZN(G1346gat));
  OAI21_X1  g696(.A(G162gat), .B1(new_n895), .B2(new_n653), .ZN(new_n898));
  INV_X1    g697(.A(G162gat), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n848), .A2(new_n899), .A3(new_n817), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n898), .A2(new_n900), .ZN(G1347gat));
  NAND3_X1  g700(.A1(new_n503), .A2(new_n499), .A3(new_n485), .ZN(new_n902));
  XOR2_X1   g701(.A(new_n902), .B(KEYINPUT124), .Z(new_n903));
  NAND2_X1  g702(.A1(new_n807), .A2(new_n903), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n904), .A2(new_n234), .A3(new_n242), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n627), .A2(new_n500), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n856), .A2(new_n906), .ZN(new_n907));
  XNOR2_X1  g706(.A(new_n907), .B(KEYINPUT123), .ZN(new_n908));
  AOI21_X1  g707(.A(G169gat), .B1(new_n908), .B2(new_n241), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n905), .A2(new_n909), .ZN(G1348gat));
  OAI21_X1  g709(.A(G176gat), .B1(new_n904), .B2(new_n659), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n908), .A2(new_n332), .A3(new_n622), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(G1349gat));
  OAI21_X1  g712(.A(G183gat), .B1(new_n904), .B2(new_n658), .ZN(new_n914));
  NAND4_X1  g713(.A1(new_n856), .A2(new_n338), .A3(new_n569), .A4(new_n906), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g715(.A(new_n916), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g716(.A1(new_n807), .A2(new_n603), .A3(new_n903), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(G190gat), .ZN(new_n919));
  OAI21_X1  g718(.A(KEYINPUT125), .B1(new_n919), .B2(KEYINPUT61), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT125), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT61), .ZN(new_n922));
  NAND4_X1  g721(.A1(new_n918), .A2(new_n921), .A3(new_n922), .A4(G190gat), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n919), .A2(KEYINPUT61), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n920), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n908), .A2(new_n343), .A3(new_n603), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(new_n926), .ZN(G1351gat));
  NOR3_X1   g726(.A1(new_n627), .A2(new_n539), .A3(new_n329), .ZN(new_n928));
  AND2_X1   g727(.A1(new_n824), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g728(.A(G197gat), .B1(new_n929), .B2(new_n241), .ZN(new_n930));
  XNOR2_X1  g729(.A(new_n928), .B(KEYINPUT126), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n931), .B1(new_n870), .B2(new_n857), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n242), .A2(new_n385), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n930), .B1(new_n932), .B2(new_n933), .ZN(G1352gat));
  NAND3_X1  g733(.A1(new_n929), .A2(new_n383), .A3(new_n622), .ZN(new_n935));
  XOR2_X1   g734(.A(new_n935), .B(KEYINPUT62), .Z(new_n936));
  INV_X1    g735(.A(new_n871), .ZN(new_n937));
  OAI21_X1  g736(.A(G204gat), .B1(new_n937), .B2(new_n931), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n936), .A2(new_n938), .ZN(G1353gat));
  NAND2_X1  g738(.A1(new_n932), .A2(new_n569), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(G211gat), .ZN(new_n941));
  OR2_X1    g740(.A1(new_n941), .A2(KEYINPUT63), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(KEYINPUT63), .ZN(new_n943));
  INV_X1    g742(.A(G211gat), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n929), .A2(new_n944), .A3(new_n569), .ZN(new_n945));
  XNOR2_X1  g744(.A(new_n945), .B(KEYINPUT127), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n942), .A2(new_n943), .A3(new_n946), .ZN(G1354gat));
  INV_X1    g746(.A(G218gat), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n929), .A2(new_n948), .A3(new_n603), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n932), .A2(new_n603), .ZN(new_n950));
  INV_X1    g749(.A(new_n950), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n949), .B1(new_n951), .B2(new_n948), .ZN(G1355gat));
endmodule


