//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 1 0 1 1 1 1 1 1 0 0 1 1 0 1 0 1 1 1 1 0 1 0 1 1 0 0 0 1 0 1 1 0 0 0 0 1 0 0 0 0 1 1 1 1 1 0 1 1 0 0 0 0 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:35 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1290, new_n1291,
    new_n1292, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1361, new_n1362, new_n1363, new_n1364, new_n1365,
    new_n1366, new_n1367;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  OAI21_X1  g0009(.A(G50), .B1(G58), .B2(G68), .ZN(new_n210));
  XOR2_X1   g0010(.A(new_n210), .B(KEYINPUT64), .Z(new_n211));
  NAND4_X1  g0011(.A1(new_n211), .A2(G1), .A3(G13), .A4(G20), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n213));
  INV_X1    g0013(.A(G68), .ZN(new_n214));
  INV_X1    g0014(.A(G238), .ZN(new_n215));
  INV_X1    g0015(.A(G87), .ZN(new_n216));
  INV_X1    g0016(.A(G250), .ZN(new_n217));
  OAI221_X1 g0017(.A(new_n213), .B1(new_n214), .B2(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n219));
  INV_X1    g0019(.A(G58), .ZN(new_n220));
  INV_X1    g0020(.A(G232), .ZN(new_n221));
  INV_X1    g0021(.A(G97), .ZN(new_n222));
  INV_X1    g0022(.A(G257), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n206), .B1(new_n218), .B2(new_n224), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n209), .B(new_n212), .C1(KEYINPUT1), .C2(new_n225), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(new_n221), .ZN(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT2), .B(G226), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(G264), .B(G270), .Z(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n231), .B(new_n234), .Z(G358));
  XNOR2_X1  g0035(.A(G50), .B(G68), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G58), .B(G77), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n236), .B(new_n237), .Z(new_n238));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XNOR2_X1  g0039(.A(G107), .B(G116), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G351));
  NAND2_X1  g0042(.A1(G33), .A2(G41), .ZN(new_n243));
  NAND3_X1  g0043(.A1(new_n243), .A2(G1), .A3(G13), .ZN(new_n244));
  OR2_X1    g0044(.A1(KEYINPUT3), .A2(G33), .ZN(new_n245));
  NAND2_X1  g0045(.A1(KEYINPUT3), .A2(G33), .ZN(new_n246));
  AOI21_X1  g0046(.A(G1698), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(G222), .ZN(new_n248));
  XNOR2_X1  g0048(.A(KEYINPUT3), .B(G33), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n249), .A2(G223), .A3(G1698), .ZN(new_n250));
  AND2_X1   g0050(.A1(KEYINPUT3), .A2(G33), .ZN(new_n251));
  NOR2_X1   g0051(.A1(KEYINPUT3), .A2(G33), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G77), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n248), .A2(new_n250), .A3(new_n254), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n244), .B1(new_n255), .B2(KEYINPUT67), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n256), .B1(KEYINPUT67), .B2(new_n255), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT66), .ZN(new_n258));
  NAND2_X1  g0058(.A1(G1), .A2(G13), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n259), .B1(G33), .B2(G41), .ZN(new_n260));
  INV_X1    g0060(.A(G41), .ZN(new_n261));
  INV_X1    g0061(.A(G45), .ZN(new_n262));
  AOI21_X1  g0062(.A(G1), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n258), .B1(new_n260), .B2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G1), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n265), .B1(G41), .B2(G45), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n244), .A2(KEYINPUT66), .A3(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n264), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n263), .A2(new_n244), .A3(G274), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT65), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND4_X1  g0071(.A1(new_n263), .A2(new_n244), .A3(KEYINPUT65), .A4(G274), .ZN(new_n272));
  AOI22_X1  g0072(.A1(new_n268), .A2(G226), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n257), .A2(new_n273), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n274), .A2(G179), .ZN(new_n275));
  XNOR2_X1  g0075(.A(new_n275), .B(KEYINPUT70), .ZN(new_n276));
  XNOR2_X1  g0076(.A(KEYINPUT8), .B(G58), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(KEYINPUT68), .ZN(new_n278));
  OR3_X1    g0078(.A1(new_n220), .A2(KEYINPUT68), .A3(KEYINPUT8), .ZN(new_n279));
  AND2_X1   g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G33), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n281), .A2(G20), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n203), .A2(KEYINPUT69), .A3(G20), .ZN(new_n284));
  NOR2_X1   g0084(.A1(G20), .A2(G33), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G150), .ZN(new_n286));
  INV_X1    g0086(.A(G20), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n287), .B1(new_n201), .B2(new_n202), .ZN(new_n288));
  OR2_X1    g0088(.A1(new_n288), .A2(KEYINPUT69), .ZN(new_n289));
  NAND4_X1  g0089(.A1(new_n283), .A2(new_n284), .A3(new_n286), .A4(new_n289), .ZN(new_n290));
  NAND3_X1  g0090(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(new_n259), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n265), .A2(G13), .A3(G20), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n294), .A2(G50), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n292), .B1(new_n265), .B2(G20), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n295), .B1(new_n296), .B2(G50), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n293), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G169), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n299), .B1(new_n300), .B2(new_n274), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n276), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n274), .A2(G200), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT74), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n274), .A2(KEYINPUT74), .A3(G200), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT9), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n298), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n257), .A2(G190), .A3(new_n273), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n293), .A2(KEYINPUT9), .A3(new_n297), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n309), .A2(KEYINPUT73), .A3(new_n310), .A4(new_n311), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n307), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT10), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NOR3_X1   g0115(.A1(new_n307), .A2(new_n312), .A3(KEYINPUT10), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n302), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT16), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n245), .A2(new_n287), .A3(new_n246), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT7), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND4_X1  g0121(.A1(new_n245), .A2(KEYINPUT7), .A3(new_n287), .A4(new_n246), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n214), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n220), .A2(new_n214), .ZN(new_n324));
  OAI21_X1  g0124(.A(G20), .B1(new_n324), .B2(new_n201), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n285), .A2(G159), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n318), .B1(new_n323), .B2(new_n327), .ZN(new_n328));
  AOI21_X1  g0128(.A(KEYINPUT7), .B1(new_n253), .B2(new_n287), .ZN(new_n329));
  INV_X1    g0129(.A(new_n322), .ZN(new_n330));
  OAI21_X1  g0130(.A(G68), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n327), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n331), .A2(KEYINPUT16), .A3(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n328), .A2(new_n333), .A3(new_n292), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT78), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n328), .A2(new_n333), .A3(KEYINPUT78), .A4(new_n292), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(G200), .ZN(new_n339));
  AND3_X1   g0139(.A1(new_n244), .A2(G232), .A3(new_n266), .ZN(new_n340));
  NAND2_X1  g0140(.A1(G33), .A2(G87), .ZN(new_n341));
  INV_X1    g0141(.A(G226), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(G1698), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n343), .B1(G223), .B2(G1698), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n341), .B1(new_n344), .B2(new_n253), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n340), .B1(new_n345), .B2(new_n260), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT79), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n271), .A2(new_n272), .ZN(new_n348));
  AND3_X1   g0148(.A1(new_n346), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n347), .B1(new_n346), .B2(new_n348), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n339), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n346), .A2(new_n348), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(G190), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n351), .A2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(new_n280), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(new_n294), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n358), .B1(new_n357), .B2(new_n296), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n338), .A2(new_n356), .A3(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT17), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n338), .A2(new_n359), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT18), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n300), .B1(new_n349), .B2(new_n350), .ZN(new_n365));
  INV_X1    g0165(.A(G179), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n353), .A2(new_n366), .ZN(new_n367));
  AND2_X1   g0167(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n363), .A2(new_n364), .A3(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n359), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n370), .B1(new_n336), .B2(new_n337), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n365), .B1(G179), .B2(new_n352), .ZN(new_n372));
  OAI21_X1  g0172(.A(KEYINPUT18), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n371), .A2(KEYINPUT17), .A3(new_n356), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n362), .A2(new_n369), .A3(new_n373), .A4(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n268), .A2(G238), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(new_n348), .ZN(new_n377));
  INV_X1    g0177(.A(G1698), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n342), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n221), .A2(G1698), .ZN(new_n380));
  OAI211_X1 g0180(.A(new_n379), .B(new_n380), .C1(new_n251), .C2(new_n252), .ZN(new_n381));
  NAND2_X1  g0181(.A1(G33), .A2(G97), .ZN(new_n382));
  AND3_X1   g0182(.A1(new_n381), .A2(KEYINPUT75), .A3(new_n382), .ZN(new_n383));
  AOI21_X1  g0183(.A(KEYINPUT75), .B1(new_n381), .B2(new_n382), .ZN(new_n384));
  NOR3_X1   g0184(.A1(new_n383), .A2(new_n384), .A3(new_n244), .ZN(new_n385));
  OAI21_X1  g0185(.A(KEYINPUT13), .B1(new_n377), .B2(new_n385), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n384), .A2(new_n244), .ZN(new_n387));
  INV_X1    g0187(.A(new_n383), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT13), .ZN(new_n390));
  AOI22_X1  g0190(.A1(new_n268), .A2(G238), .B1(new_n271), .B2(new_n272), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n389), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n386), .A2(new_n392), .ZN(new_n393));
  OAI21_X1  g0193(.A(KEYINPUT76), .B1(new_n393), .B2(new_n354), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT76), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n386), .A2(new_n392), .A3(new_n395), .A4(G190), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  NOR3_X1   g0197(.A1(new_n377), .A2(new_n385), .A3(KEYINPUT13), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n390), .B1(new_n389), .B2(new_n391), .ZN(new_n399));
  OAI21_X1  g0199(.A(G200), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n296), .A2(G68), .ZN(new_n401));
  XOR2_X1   g0201(.A(new_n401), .B(KEYINPUT77), .Z(new_n402));
  NAND2_X1  g0202(.A1(new_n282), .A2(G77), .ZN(new_n403));
  INV_X1    g0203(.A(new_n285), .ZN(new_n404));
  OAI221_X1 g0204(.A(new_n403), .B1(new_n287), .B2(G68), .C1(new_n202), .C2(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n405), .A2(KEYINPUT11), .A3(new_n292), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n292), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT11), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(new_n294), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(new_n214), .ZN(new_n411));
  XNOR2_X1  g0211(.A(new_n411), .B(KEYINPUT12), .ZN(new_n412));
  AND4_X1   g0212(.A1(new_n402), .A2(new_n406), .A3(new_n409), .A4(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n400), .A2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n397), .A2(new_n415), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n402), .A2(new_n409), .A3(new_n412), .A4(new_n406), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT14), .ZN(new_n418));
  OAI211_X1 g0218(.A(new_n418), .B(G169), .C1(new_n398), .C2(new_n399), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n386), .A2(G179), .A3(new_n392), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n418), .B1(new_n393), .B2(G169), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n417), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n296), .A2(G77), .ZN(new_n424));
  INV_X1    g0224(.A(G77), .ZN(new_n425));
  OAI22_X1  g0225(.A1(new_n277), .A2(new_n404), .B1(new_n287), .B2(new_n425), .ZN(new_n426));
  XNOR2_X1  g0226(.A(KEYINPUT15), .B(G87), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT71), .ZN(new_n428));
  XNOR2_X1  g0228(.A(new_n427), .B(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n426), .B1(new_n429), .B2(new_n282), .ZN(new_n430));
  INV_X1    g0230(.A(new_n292), .ZN(new_n431));
  OAI221_X1 g0231(.A(new_n424), .B1(G77), .B2(new_n294), .C1(new_n430), .C2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n247), .A2(G232), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n249), .A2(G238), .A3(G1698), .ZN(new_n434));
  INV_X1    g0234(.A(G107), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n433), .B(new_n434), .C1(new_n435), .C2(new_n249), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(new_n260), .ZN(new_n437));
  AOI22_X1  g0237(.A1(new_n268), .A2(G244), .B1(new_n271), .B2(new_n272), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(new_n300), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n437), .A2(new_n438), .A3(new_n366), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n432), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n339), .B1(new_n437), .B2(new_n438), .ZN(new_n443));
  OR3_X1    g0243(.A1(new_n432), .A2(KEYINPUT72), .A3(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n437), .A2(new_n438), .A3(G190), .ZN(new_n445));
  OAI21_X1  g0245(.A(KEYINPUT72), .B1(new_n432), .B2(new_n443), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n444), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n416), .A2(new_n423), .A3(new_n442), .A4(new_n447), .ZN(new_n448));
  NOR3_X1   g0248(.A1(new_n317), .A2(new_n375), .A3(new_n448), .ZN(new_n449));
  OAI211_X1 g0249(.A(G244), .B(new_n378), .C1(new_n251), .C2(new_n252), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT4), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n249), .A2(KEYINPUT4), .A3(G244), .A4(new_n378), .ZN(new_n453));
  NAND2_X1  g0253(.A1(G33), .A2(G283), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n249), .A2(G250), .A3(G1698), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n452), .A2(new_n453), .A3(new_n454), .A4(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(new_n260), .ZN(new_n457));
  OR2_X1    g0257(.A1(KEYINPUT5), .A2(G41), .ZN(new_n458));
  NAND2_X1  g0258(.A1(KEYINPUT5), .A2(G41), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n265), .A2(G45), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n460), .A2(G274), .A3(new_n244), .A4(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n244), .A2(new_n458), .A3(new_n459), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n244), .A2(new_n461), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n223), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n457), .A2(G179), .A3(new_n463), .A4(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(new_n463), .ZN(new_n469));
  AOI211_X1 g0269(.A(new_n469), .B(new_n466), .C1(new_n456), .C2(new_n260), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n468), .B1(new_n470), .B2(new_n300), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n285), .A2(G77), .ZN(new_n472));
  AND3_X1   g0272(.A1(new_n435), .A2(KEYINPUT6), .A3(G97), .ZN(new_n473));
  XNOR2_X1  g0273(.A(G97), .B(G107), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT6), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n473), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n472), .B1(new_n476), .B2(new_n287), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n435), .B1(new_n321), .B2(new_n322), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n292), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n294), .A2(G97), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n265), .A2(G33), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n431), .A2(new_n294), .A3(new_n482), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n481), .B1(new_n483), .B2(new_n222), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n479), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n471), .A2(new_n486), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n287), .B(G87), .C1(new_n251), .C2(new_n252), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(KEYINPUT22), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT22), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n249), .A2(new_n490), .A3(new_n287), .A4(G87), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT23), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n493), .B1(new_n287), .B2(G107), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n435), .A2(KEYINPUT23), .A3(G20), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(G116), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n281), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(new_n287), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n496), .A2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n492), .A2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT83), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT24), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n502), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n500), .B1(new_n489), .B2(new_n491), .ZN(new_n506));
  OAI21_X1  g0306(.A(KEYINPUT24), .B1(new_n506), .B2(KEYINPUT83), .ZN(new_n507));
  AND3_X1   g0307(.A1(new_n492), .A2(KEYINPUT83), .A3(new_n501), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n505), .B(new_n292), .C1(new_n507), .C2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT25), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n510), .B1(new_n294), .B2(G107), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  NOR3_X1   g0312(.A1(new_n294), .A2(new_n510), .A3(G107), .ZN(new_n513));
  OAI22_X1  g0313(.A1(new_n483), .A2(new_n435), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(new_n514), .ZN(new_n515));
  AOI22_X1  g0315(.A1(new_n247), .A2(G250), .B1(G33), .B2(G294), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n249), .A2(G257), .A3(G1698), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n244), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  AND2_X1   g0318(.A1(KEYINPUT5), .A2(G41), .ZN(new_n519));
  NOR2_X1   g0319(.A1(KEYINPUT5), .A2(G41), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  OAI211_X1 g0321(.A(G264), .B(new_n244), .C1(new_n521), .C2(new_n461), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(new_n463), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n339), .B1(new_n518), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n249), .A2(G250), .A3(new_n378), .ZN(new_n525));
  INV_X1    g0325(.A(G294), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n517), .B(new_n525), .C1(new_n281), .C2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(new_n260), .ZN(new_n528));
  INV_X1    g0328(.A(new_n523), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n528), .A2(new_n354), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n524), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n509), .A2(new_n515), .A3(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n466), .B1(new_n456), .B2(new_n260), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n533), .A2(G190), .A3(new_n463), .ZN(new_n534));
  OAI21_X1  g0334(.A(G107), .B1(new_n329), .B2(new_n330), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n474), .A2(new_n475), .ZN(new_n536));
  INV_X1    g0336(.A(new_n473), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(G20), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n535), .A2(new_n539), .A3(new_n472), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n484), .B1(new_n540), .B2(new_n292), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n534), .B(new_n541), .C1(new_n339), .C2(new_n470), .ZN(new_n542));
  AND3_X1   g0342(.A1(new_n487), .A2(new_n532), .A3(new_n542), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n300), .B1(new_n518), .B2(new_n523), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n528), .A2(new_n366), .A3(new_n529), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n546), .B1(new_n509), .B2(new_n515), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n410), .A2(new_n497), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n431), .A2(G116), .A3(new_n294), .A4(new_n482), .ZN(new_n549));
  AOI22_X1  g0349(.A1(new_n291), .A2(new_n259), .B1(G20), .B2(new_n497), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n454), .B(new_n287), .C1(G33), .C2(new_n222), .ZN(new_n551));
  AND3_X1   g0351(.A1(new_n550), .A2(KEYINPUT20), .A3(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(KEYINPUT20), .B1(new_n550), .B2(new_n551), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n548), .B(new_n549), .C1(new_n552), .C2(new_n553), .ZN(new_n554));
  OAI211_X1 g0354(.A(G264), .B(G1698), .C1(new_n251), .C2(new_n252), .ZN(new_n555));
  OAI211_X1 g0355(.A(G257), .B(new_n378), .C1(new_n251), .C2(new_n252), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n245), .A2(G303), .A3(new_n246), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n555), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(new_n260), .ZN(new_n559));
  INV_X1    g0359(.A(new_n559), .ZN(new_n560));
  OAI211_X1 g0360(.A(G270), .B(new_n244), .C1(new_n521), .C2(new_n461), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n463), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n554), .B(G169), .C1(new_n560), .C2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT21), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  AND2_X1   g0365(.A1(new_n561), .A2(new_n463), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n554), .A2(G179), .A3(new_n559), .A4(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n559), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n568), .A2(KEYINPUT21), .A3(G169), .A4(new_n554), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n565), .A2(new_n567), .A3(new_n569), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n547), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n215), .A2(new_n378), .ZN(new_n572));
  INV_X1    g0372(.A(G244), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(G1698), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n572), .B(new_n574), .C1(new_n251), .C2(new_n252), .ZN(new_n575));
  INV_X1    g0375(.A(new_n498), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT80), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n575), .A2(KEYINPUT80), .A3(new_n576), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n579), .A2(new_n260), .A3(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n462), .A2(new_n244), .A3(G274), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n582), .B1(new_n465), .B2(new_n217), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n339), .B1(new_n581), .B2(new_n584), .ZN(new_n585));
  XOR2_X1   g0385(.A(KEYINPUT15), .B(G87), .Z(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(new_n428), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n427), .A2(KEYINPUT71), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(new_n410), .ZN(new_n590));
  OR2_X1    g0390(.A1(new_n483), .A2(new_n216), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n287), .B(G68), .C1(new_n251), .C2(new_n252), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n287), .A2(G33), .A3(G97), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT19), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(KEYINPUT81), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT81), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(KEYINPUT19), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n593), .A2(new_n595), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n592), .A2(new_n598), .ZN(new_n599));
  XNOR2_X1  g0399(.A(KEYINPUT81), .B(KEYINPUT19), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n287), .B1(new_n600), .B2(new_n382), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n216), .A2(new_n222), .A3(new_n435), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n599), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n590), .B(new_n591), .C1(new_n603), .C2(new_n431), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n585), .A2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT82), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n581), .A2(new_n606), .A3(G190), .A4(new_n584), .ZN(new_n607));
  INV_X1    g0407(.A(new_n607), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n244), .B1(new_n577), .B2(new_n578), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n583), .B1(new_n609), .B2(new_n580), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n606), .B1(new_n610), .B2(G190), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n605), .B1(new_n608), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n581), .A2(new_n584), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(new_n300), .ZN(new_n614));
  OAI221_X1 g0414(.A(new_n590), .B1(new_n589), .B2(new_n483), .C1(new_n603), .C2(new_n431), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n610), .A2(new_n366), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n560), .A2(new_n562), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n554), .B1(new_n618), .B2(G190), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n619), .B1(new_n339), .B2(new_n618), .ZN(new_n620));
  AND3_X1   g0420(.A1(new_n612), .A2(new_n617), .A3(new_n620), .ZN(new_n621));
  AND4_X1   g0421(.A1(new_n449), .A2(new_n543), .A3(new_n571), .A4(new_n621), .ZN(G372));
  AND3_X1   g0422(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n623));
  NOR2_X1   g0423(.A1(G238), .A2(G1698), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n624), .B1(new_n573), .B2(G1698), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n498), .B1(new_n625), .B2(new_n249), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n260), .B1(new_n626), .B2(KEYINPUT80), .ZN(new_n627));
  AND3_X1   g0427(.A1(new_n575), .A2(KEYINPUT80), .A3(new_n576), .ZN(new_n628));
  OAI211_X1 g0428(.A(G190), .B(new_n584), .C1(new_n627), .C2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(KEYINPUT82), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(new_n607), .ZN(new_n631));
  AOI21_X1  g0431(.A(KEYINPUT80), .B1(new_n575), .B2(new_n576), .ZN(new_n632));
  NOR3_X1   g0432(.A1(new_n628), .A2(new_n632), .A3(new_n244), .ZN(new_n633));
  OAI21_X1  g0433(.A(G200), .B1(new_n633), .B2(new_n583), .ZN(new_n634));
  INV_X1    g0434(.A(new_n599), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n382), .B1(new_n595), .B2(new_n597), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n602), .B1(new_n636), .B2(G20), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n431), .B1(new_n635), .B2(new_n637), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n294), .B1(new_n587), .B2(new_n588), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n483), .A2(new_n216), .ZN(new_n640));
  NOR3_X1   g0440(.A1(new_n638), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT84), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n634), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  OAI21_X1  g0443(.A(KEYINPUT84), .B1(new_n585), .B2(new_n604), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n631), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(new_n617), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n487), .A2(new_n532), .A3(new_n542), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT85), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n569), .A2(new_n567), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n300), .B1(new_n566), .B2(new_n559), .ZN(new_n651));
  AOI21_X1  g0451(.A(KEYINPUT21), .B1(new_n651), .B2(new_n554), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n649), .B1(new_n650), .B2(new_n652), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n565), .A2(KEYINPUT85), .A3(new_n567), .A4(new_n569), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n547), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n623), .B1(new_n648), .B2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT26), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT86), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n471), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n457), .A2(new_n463), .A3(new_n467), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(G169), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n663), .A2(KEYINPUT86), .A3(new_n468), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n661), .A2(new_n486), .A3(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n659), .B1(new_n646), .B2(new_n665), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n541), .B1(new_n663), .B2(new_n468), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n612), .A2(new_n667), .A3(KEYINPUT26), .A4(new_n617), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n658), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n449), .A2(new_n670), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n414), .B1(new_n396), .B2(new_n394), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n423), .B1(new_n672), .B2(new_n442), .ZN(new_n673));
  AND2_X1   g0473(.A1(new_n362), .A2(new_n374), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n675), .A2(new_n373), .A3(new_n369), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n315), .A2(new_n316), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n671), .A2(new_n302), .A3(new_n679), .ZN(G369));
  NAND3_X1  g0480(.A1(new_n265), .A2(new_n287), .A3(G13), .ZN(new_n681));
  OR2_X1    g0481(.A1(new_n681), .A2(KEYINPUT27), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(KEYINPUT27), .ZN(new_n683));
  AND3_X1   g0483(.A1(new_n682), .A2(G213), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g0484(.A(KEYINPUT87), .B(G343), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  XOR2_X1   g0486(.A(new_n686), .B(KEYINPUT88), .Z(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(new_n554), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n650), .A2(new_n652), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n689), .A2(new_n690), .A3(new_n620), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n691), .B1(new_n655), .B2(new_n689), .ZN(new_n692));
  XNOR2_X1  g0492(.A(new_n692), .B(KEYINPUT89), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(G330), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n656), .A2(new_n532), .ZN(new_n696));
  AND2_X1   g0496(.A1(new_n505), .A2(new_n292), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n502), .A2(new_n503), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n506), .A2(KEYINPUT83), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n698), .A2(KEYINPUT24), .A3(new_n699), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n514), .B1(new_n697), .B2(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n701), .A2(new_n687), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n696), .A2(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n656), .A2(new_n687), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n695), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n570), .A2(new_n687), .ZN(new_n708));
  NOR3_X1   g0508(.A1(new_n696), .A2(new_n702), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n547), .A2(new_n687), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n707), .A2(new_n712), .ZN(new_n713));
  XOR2_X1   g0513(.A(new_n713), .B(KEYINPUT90), .Z(G399));
  INV_X1    g0514(.A(new_n207), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n715), .A2(G41), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n602), .A2(G116), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n717), .A2(G1), .A3(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n211), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n719), .B1(new_n720), .B2(new_n717), .ZN(new_n721));
  XNOR2_X1  g0521(.A(new_n721), .B(KEYINPUT28), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n612), .A2(new_n667), .A3(new_n617), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(new_n659), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n541), .B1(new_n471), .B2(new_n660), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n725), .A2(new_n645), .A3(new_n617), .A4(new_n664), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n724), .B1(new_n726), .B2(new_n659), .ZN(new_n727));
  OAI211_X1 g0527(.A(new_n690), .B(KEYINPUT91), .C1(new_n701), .C2(new_n546), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n635), .A2(new_n637), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n639), .B1(new_n729), .B2(new_n292), .ZN(new_n730));
  OAI211_X1 g0530(.A(new_n730), .B(new_n591), .C1(new_n610), .C2(new_n339), .ZN(new_n731));
  AOI22_X1  g0531(.A1(new_n731), .A2(KEYINPUT84), .B1(new_n630), .B2(new_n607), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n623), .B1(new_n732), .B2(new_n643), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT91), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n734), .B1(new_n547), .B2(new_n570), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n543), .A2(new_n728), .A3(new_n733), .A4(new_n735), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n727), .A2(new_n617), .A3(new_n736), .ZN(new_n737));
  AND3_X1   g0537(.A1(new_n737), .A2(KEYINPUT92), .A3(new_n687), .ZN(new_n738));
  AOI21_X1  g0538(.A(KEYINPUT92), .B1(new_n737), .B2(new_n687), .ZN(new_n739));
  OAI21_X1  g0539(.A(KEYINPUT29), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n688), .B1(new_n658), .B2(new_n669), .ZN(new_n741));
  OR2_X1    g0541(.A1(new_n741), .A2(KEYINPUT29), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n621), .A2(new_n543), .A3(new_n571), .A4(new_n687), .ZN(new_n743));
  NOR3_X1   g0543(.A1(new_n560), .A2(new_n366), .A3(new_n562), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n518), .A2(new_n523), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n744), .A2(new_n533), .A3(new_n745), .A4(new_n610), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT30), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n528), .A2(new_n529), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n613), .A2(new_n749), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n750), .A2(KEYINPUT30), .A3(new_n533), .A4(new_n744), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n745), .A2(new_n610), .ZN(new_n752));
  NAND4_X1  g0552(.A1(new_n752), .A2(new_n366), .A3(new_n662), .A4(new_n568), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n748), .A2(new_n751), .A3(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(new_n688), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT31), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n754), .A2(KEYINPUT31), .A3(new_n688), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n743), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  AOI22_X1  g0559(.A1(new_n740), .A2(new_n742), .B1(G330), .B2(new_n759), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n722), .B1(new_n760), .B2(G1), .ZN(G364));
  INV_X1    g0561(.A(G13), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(G20), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n265), .B1(new_n763), .B2(G45), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n716), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n249), .A2(new_n207), .ZN(new_n767));
  INV_X1    g0567(.A(G355), .ZN(new_n768));
  OAI22_X1  g0568(.A1(new_n767), .A2(new_n768), .B1(G116), .B2(new_n207), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n715), .A2(new_n249), .ZN(new_n770));
  XNOR2_X1  g0570(.A(new_n770), .B(KEYINPUT93), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n771), .B1(new_n262), .B2(new_n211), .ZN(new_n772));
  OR2_X1    g0572(.A1(new_n238), .A2(new_n262), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n769), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(G13), .A2(G33), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(G20), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n259), .B1(G20), .B2(new_n300), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n766), .B1(new_n774), .B2(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n287), .A2(G179), .ZN(new_n782));
  NOR2_X1   g0582(.A1(G190), .A2(G200), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(G159), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n782), .A2(new_n354), .A3(G200), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  AOI22_X1  g0588(.A1(new_n786), .A2(KEYINPUT32), .B1(G107), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(G20), .A2(G179), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(G200), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(new_n354), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n354), .A2(G200), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n287), .B1(new_n795), .B2(new_n366), .ZN(new_n796));
  OAI221_X1 g0596(.A(new_n789), .B1(new_n202), .B2(new_n794), .C1(new_n222), .C2(new_n796), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n782), .A2(G190), .A3(G200), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(new_n216), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n792), .A2(G190), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  OAI221_X1 g0602(.A(new_n800), .B1(new_n786), .B2(KEYINPUT32), .C1(new_n214), .C2(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n791), .A2(new_n783), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n795), .A2(new_n791), .ZN(new_n805));
  OAI221_X1 g0605(.A(new_n249), .B1(new_n804), .B2(new_n425), .C1(new_n220), .C2(new_n805), .ZN(new_n806));
  OR3_X1    g0606(.A1(new_n797), .A2(new_n803), .A3(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(G322), .ZN(new_n808));
  INV_X1    g0608(.A(G329), .ZN(new_n809));
  OAI22_X1  g0609(.A1(new_n805), .A2(new_n808), .B1(new_n784), .B2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n804), .ZN(new_n811));
  AOI211_X1 g0611(.A(new_n249), .B(new_n810), .C1(G311), .C2(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n793), .A2(G326), .ZN(new_n813));
  XNOR2_X1  g0613(.A(KEYINPUT33), .B(G317), .ZN(new_n814));
  INV_X1    g0614(.A(new_n798), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n801), .A2(new_n814), .B1(new_n815), .B2(G303), .ZN(new_n816));
  INV_X1    g0616(.A(new_n796), .ZN(new_n817));
  AOI22_X1  g0617(.A1(G294), .A2(new_n817), .B1(new_n788), .B2(G283), .ZN(new_n818));
  NAND4_X1  g0618(.A1(new_n812), .A2(new_n813), .A3(new_n816), .A4(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n807), .A2(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n781), .B1(new_n778), .B2(new_n820), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n777), .B(KEYINPUT94), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n821), .B1(new_n693), .B2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n766), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n694), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n693), .A2(G330), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n823), .B1(new_n825), .B2(new_n826), .ZN(G396));
  NOR2_X1   g0627(.A1(new_n688), .A2(new_n442), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n688), .A2(new_n432), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n447), .A2(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n828), .B1(new_n830), .B2(new_n442), .ZN(new_n831));
  XNOR2_X1  g0631(.A(new_n741), .B(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n759), .A2(G330), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n766), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n834), .B1(new_n833), .B2(new_n832), .ZN(new_n835));
  INV_X1    g0635(.A(new_n805), .ZN(new_n836));
  AOI22_X1  g0636(.A1(G143), .A2(new_n836), .B1(new_n811), .B2(G159), .ZN(new_n837));
  INV_X1    g0637(.A(G150), .ZN(new_n838));
  INV_X1    g0638(.A(G137), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n837), .B1(new_n802), .B2(new_n838), .C1(new_n839), .C2(new_n794), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT34), .ZN(new_n841));
  AND2_X1   g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n840), .A2(new_n841), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n788), .A2(G68), .ZN(new_n844));
  INV_X1    g0644(.A(G132), .ZN(new_n845));
  OAI211_X1 g0645(.A(new_n844), .B(new_n249), .C1(new_n845), .C2(new_n784), .ZN(new_n846));
  OAI22_X1  g0646(.A1(new_n796), .A2(new_n220), .B1(new_n798), .B2(new_n202), .ZN(new_n847));
  NOR4_X1   g0647(.A1(new_n842), .A2(new_n843), .A3(new_n846), .A4(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(G303), .ZN(new_n849));
  OAI22_X1  g0649(.A1(new_n794), .A2(new_n849), .B1(new_n435), .B2(new_n798), .ZN(new_n850));
  XOR2_X1   g0650(.A(KEYINPUT95), .B(G283), .Z(new_n851));
  AOI22_X1  g0651(.A1(G97), .A2(new_n817), .B1(new_n801), .B2(new_n851), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n249), .B1(new_n836), .B2(G294), .ZN(new_n853));
  AOI22_X1  g0653(.A1(G311), .A2(new_n785), .B1(new_n811), .B2(G116), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n852), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  AOI211_X1 g0655(.A(new_n850), .B(new_n855), .C1(G87), .C2(new_n788), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n778), .B1(new_n848), .B2(new_n856), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n778), .A2(new_n775), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n824), .B1(new_n425), .B2(new_n858), .ZN(new_n859));
  OAI211_X1 g0659(.A(new_n857), .B(new_n859), .C1(new_n831), .C2(new_n776), .ZN(new_n860));
  AND2_X1   g0660(.A1(new_n835), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(G384));
  NOR2_X1   g0662(.A1(new_n763), .A2(new_n265), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n679), .A2(new_n302), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n740), .A2(new_n449), .A3(new_n742), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(KEYINPUT98), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT98), .ZN(new_n867));
  NAND4_X1  g0667(.A1(new_n740), .A2(new_n449), .A3(new_n867), .A4(new_n742), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n864), .B1(new_n866), .B2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT39), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n334), .A2(new_n359), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(new_n684), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(KEYINPUT97), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT97), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n871), .A2(new_n874), .A3(new_n684), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n375), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n871), .A2(new_n365), .A3(new_n367), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n360), .A2(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(KEYINPUT37), .B1(new_n879), .B2(new_n876), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n363), .A2(new_n368), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n363), .A2(new_n684), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT37), .ZN(new_n883));
  NAND4_X1  g0683(.A1(new_n881), .A2(new_n882), .A3(new_n883), .A4(new_n360), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n880), .A2(new_n884), .ZN(new_n885));
  AND3_X1   g0685(.A1(new_n877), .A2(new_n885), .A3(KEYINPUT38), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n360), .B1(new_n372), .B2(new_n371), .ZN(new_n887));
  INV_X1    g0687(.A(new_n684), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n371), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(KEYINPUT37), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(new_n884), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n375), .A2(new_n889), .ZN(new_n892));
  AOI21_X1  g0692(.A(KEYINPUT38), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n870), .B1(new_n886), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n877), .A2(new_n885), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT38), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n877), .A2(new_n885), .A3(KEYINPUT38), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n897), .A2(KEYINPUT39), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n393), .A2(G169), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(KEYINPUT14), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n901), .A2(new_n420), .A3(new_n419), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n902), .A2(new_n417), .A3(new_n687), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n894), .A2(new_n899), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n684), .B1(new_n369), .B2(new_n373), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n897), .A2(new_n898), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n688), .A2(new_n417), .ZN(new_n908));
  AND3_X1   g0708(.A1(new_n416), .A2(new_n423), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n908), .B1(new_n416), .B2(new_n423), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(new_n668), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n912), .B1(new_n659), .B2(new_n726), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n486), .B1(G200), .B2(new_n662), .ZN(new_n914));
  AOI22_X1  g0714(.A1(new_n914), .A2(new_n534), .B1(new_n471), .B2(new_n486), .ZN(new_n915));
  NAND4_X1  g0715(.A1(new_n915), .A2(new_n532), .A3(new_n617), .A4(new_n645), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n547), .B1(new_n653), .B2(new_n654), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n617), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  OAI211_X1 g0718(.A(new_n687), .B(new_n831), .C1(new_n913), .C2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(new_n828), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n911), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n906), .B1(new_n907), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n905), .A2(new_n922), .ZN(new_n923));
  XOR2_X1   g0723(.A(new_n869), .B(new_n923), .Z(new_n924));
  NOR2_X1   g0724(.A1(new_n886), .A2(new_n893), .ZN(new_n925));
  OAI211_X1 g0725(.A(new_n417), .B(new_n688), .C1(new_n672), .C2(new_n902), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n416), .A2(new_n423), .A3(new_n908), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT99), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n758), .A2(new_n929), .ZN(new_n930));
  NAND4_X1  g0730(.A1(new_n754), .A2(KEYINPUT99), .A3(KEYINPUT31), .A4(new_n688), .ZN(new_n931));
  NAND4_X1  g0731(.A1(new_n930), .A2(new_n743), .A3(new_n757), .A4(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n928), .A2(new_n932), .A3(new_n831), .ZN(new_n933));
  OAI21_X1  g0733(.A(KEYINPUT40), .B1(new_n925), .B2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT40), .ZN(new_n935));
  AND3_X1   g0735(.A1(new_n928), .A2(new_n932), .A3(new_n831), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n907), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n934), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n938), .A2(new_n449), .A3(new_n932), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n449), .A2(new_n932), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n934), .A2(new_n940), .A3(new_n937), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n939), .A2(G330), .A3(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n863), .B1(new_n924), .B2(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n943), .B1(new_n924), .B2(new_n942), .ZN(new_n944));
  NOR3_X1   g0744(.A1(new_n259), .A2(new_n287), .A3(new_n497), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n538), .B(KEYINPUT96), .ZN(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT35), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n945), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n949), .B1(new_n948), .B2(new_n947), .ZN(new_n950));
  XOR2_X1   g0750(.A(new_n950), .B(KEYINPUT36), .Z(new_n951));
  NOR3_X1   g0751(.A1(new_n720), .A2(new_n425), .A3(new_n324), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n214), .A2(G50), .ZN(new_n953));
  OAI211_X1 g0753(.A(G1), .B(new_n762), .C1(new_n952), .C2(new_n953), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n944), .A2(new_n951), .A3(new_n954), .ZN(G367));
  NOR2_X1   g0755(.A1(new_n687), .A2(new_n641), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n956), .B(KEYINPUT100), .ZN(new_n957));
  OR3_X1    g0757(.A1(new_n957), .A2(KEYINPUT101), .A3(new_n617), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n733), .ZN(new_n959));
  OAI21_X1  g0759(.A(KEYINPUT101), .B1(new_n957), .B2(new_n617), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n958), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  AND2_X1   g0761(.A1(new_n961), .A2(KEYINPUT43), .ZN(new_n962));
  XOR2_X1   g0762(.A(KEYINPUT102), .B(KEYINPUT43), .Z(new_n963));
  NOR2_X1   g0763(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n915), .B1(new_n541), .B2(new_n687), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n725), .A2(new_n664), .A3(new_n688), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n709), .A2(new_n968), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n969), .B(KEYINPUT42), .ZN(new_n970));
  INV_X1    g0770(.A(new_n968), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n487), .B1(new_n971), .B2(new_n656), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n970), .B1(new_n687), .B2(new_n972), .ZN(new_n973));
  MUX2_X1   g0773(.A(new_n965), .B(new_n964), .S(new_n973), .Z(new_n974));
  NOR2_X1   g0774(.A1(new_n707), .A2(new_n971), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n974), .B(new_n975), .ZN(new_n976));
  XOR2_X1   g0776(.A(new_n716), .B(KEYINPUT41), .Z(new_n977));
  AOI21_X1  g0777(.A(new_n709), .B1(new_n705), .B2(new_n708), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n694), .B(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n712), .A2(new_n968), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(KEYINPUT103), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT103), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n712), .A2(new_n982), .A3(new_n968), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT45), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n712), .A2(new_n968), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT44), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n981), .A2(new_n983), .A3(KEYINPUT45), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n986), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n990), .A2(KEYINPUT104), .A3(new_n707), .ZN(new_n991));
  INV_X1    g0791(.A(new_n991), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n707), .B1(new_n990), .B2(KEYINPUT104), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n979), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n977), .B1(new_n994), .B2(new_n760), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n976), .B1(new_n995), .B2(new_n765), .ZN(new_n996));
  OR2_X1    g0796(.A1(new_n961), .A2(new_n822), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n771), .A2(new_n234), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n779), .B1(new_n589), .B2(new_n207), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n766), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(G159), .ZN(new_n1001));
  OAI22_X1  g0801(.A1(new_n802), .A2(new_n1001), .B1(new_n787), .B2(new_n425), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n1002), .B1(G58), .B2(new_n815), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n805), .A2(new_n838), .B1(new_n804), .B2(new_n202), .ZN(new_n1004));
  AOI211_X1 g0804(.A(new_n253), .B(new_n1004), .C1(G137), .C2(new_n785), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(G68), .A2(new_n817), .B1(new_n793), .B2(G143), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n1003), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(KEYINPUT105), .B(G311), .ZN(new_n1008));
  OAI22_X1  g0808(.A1(new_n794), .A2(new_n1008), .B1(new_n849), .B2(new_n805), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n1009), .ZN(new_n1010));
  OR2_X1    g0810(.A1(new_n1010), .A2(KEYINPUT106), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1010), .A2(KEYINPUT106), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n787), .A2(new_n222), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n796), .A2(new_n435), .ZN(new_n1014));
  AOI211_X1 g0814(.A(new_n1013), .B(new_n1014), .C1(G294), .C2(new_n801), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1011), .A2(new_n1012), .A3(new_n1015), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n815), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n249), .B1(new_n785), .B2(G317), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT46), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1019), .B1(new_n798), .B2(new_n497), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n811), .A2(new_n851), .ZN(new_n1021));
  NAND4_X1  g0821(.A1(new_n1017), .A2(new_n1018), .A3(new_n1020), .A4(new_n1021), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1007), .B1(new_n1016), .B2(new_n1022), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT47), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1000), .B1(new_n1024), .B2(new_n778), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n997), .A2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n996), .A2(new_n1026), .ZN(G387));
  OR2_X1    g0827(.A1(new_n706), .A2(new_n822), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n767), .A2(new_n718), .B1(G107), .B2(new_n207), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n231), .A2(G45), .ZN(new_n1030));
  XOR2_X1   g0830(.A(new_n1030), .B(KEYINPUT107), .Z(new_n1031));
  XOR2_X1   g0831(.A(KEYINPUT108), .B(KEYINPUT50), .Z(new_n1032));
  NOR3_X1   g0832(.A1(new_n1032), .A2(G50), .A3(new_n277), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n262), .B1(new_n214), .B2(new_n425), .ZN(new_n1034));
  NOR4_X1   g0834(.A1(new_n1033), .A2(G116), .A3(new_n602), .A4(new_n1034), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1032), .B1(G50), .B2(new_n277), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n771), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1029), .B1(new_n1031), .B2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n766), .B1(new_n1038), .B2(new_n780), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(G317), .A2(new_n836), .B1(new_n811), .B2(G303), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n1040), .B1(new_n802), .B2(new_n1008), .C1(new_n808), .C2(new_n794), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT48), .ZN(new_n1042));
  OR2_X1    g0842(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n817), .A2(new_n851), .B1(new_n815), .B2(G294), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1043), .A2(new_n1044), .A3(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT49), .ZN(new_n1047));
  OR2_X1    g0847(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n787), .A2(new_n497), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n249), .B(new_n1050), .C1(G326), .C2(new_n785), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1048), .A2(new_n1049), .A3(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1013), .B1(G159), .B2(new_n793), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(new_n425), .B2(new_n798), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n805), .A2(new_n202), .B1(new_n784), .B2(new_n838), .ZN(new_n1055));
  AOI211_X1 g0855(.A(new_n253), .B(new_n1055), .C1(G68), .C2(new_n811), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n429), .A2(new_n817), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n1056), .B(new_n1057), .C1(new_n357), .C2(new_n802), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1052), .B1(new_n1054), .B2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1039), .B1(new_n1059), .B2(new_n778), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT109), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n979), .A2(new_n765), .B1(new_n1028), .B2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n760), .A2(new_n979), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n716), .B(KEYINPUT110), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n760), .A2(new_n979), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1062), .B1(new_n1065), .B2(new_n1066), .ZN(G393));
  NAND2_X1  g0867(.A1(new_n990), .A2(KEYINPUT104), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n707), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n1063), .ZN(new_n1071));
  NAND4_X1  g0871(.A1(new_n1070), .A2(new_n991), .A3(new_n1071), .A4(new_n1064), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n971), .A2(new_n777), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n796), .A2(new_n425), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n802), .A2(new_n202), .B1(new_n787), .B2(new_n216), .ZN(new_n1075));
  AOI211_X1 g0875(.A(new_n1074), .B(new_n1075), .C1(G68), .C2(new_n815), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n793), .A2(G150), .B1(new_n836), .B2(G159), .ZN(new_n1077));
  XOR2_X1   g0877(.A(new_n1077), .B(KEYINPUT51), .Z(new_n1078));
  OR2_X1    g0878(.A1(new_n804), .A2(new_n277), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n253), .B1(new_n785), .B2(G143), .ZN(new_n1080));
  NAND4_X1  g0880(.A1(new_n1076), .A2(new_n1078), .A3(new_n1079), .A4(new_n1080), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n793), .A2(G317), .B1(new_n836), .B2(G311), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1082), .B(KEYINPUT52), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n253), .B1(new_n784), .B2(new_n808), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1084), .B1(G294), .B2(new_n811), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(G116), .A2(new_n817), .B1(new_n801), .B2(G303), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n815), .A2(new_n851), .B1(new_n788), .B2(G107), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1085), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1081), .B1(new_n1083), .B2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(new_n778), .ZN(new_n1090));
  OAI221_X1 g0890(.A(new_n779), .B1(new_n222), .B2(new_n207), .C1(new_n771), .C2(new_n241), .ZN(new_n1091));
  NAND4_X1  g0891(.A1(new_n1073), .A2(new_n766), .A3(new_n1090), .A4(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1072), .A2(new_n1092), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n990), .B(new_n1069), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1094), .B1(new_n764), .B2(new_n1065), .ZN(new_n1095));
  OR2_X1    g0895(.A1(new_n1093), .A2(new_n1095), .ZN(G390));
  INV_X1    g0896(.A(KEYINPUT116), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n928), .A2(new_n831), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n932), .A2(G330), .ZN(new_n1099));
  OR2_X1    g0899(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n894), .A2(new_n899), .ZN(new_n1102));
  INV_X1    g0902(.A(KEYINPUT111), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1103), .B1(new_n921), .B2(new_n904), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n828), .B1(new_n741), .B2(new_n831), .ZN(new_n1105));
  OAI211_X1 g0905(.A(KEYINPUT111), .B(new_n903), .C1(new_n1105), .C2(new_n911), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1102), .A2(new_n1104), .A3(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n830), .A2(new_n442), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1109), .B1(new_n738), .B2(new_n739), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n911), .B1(new_n1110), .B2(new_n920), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n884), .A2(new_n890), .B1(new_n375), .B2(new_n889), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n898), .B1(new_n1112), .B2(KEYINPUT38), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1113), .A2(new_n903), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n1111), .A2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1101), .B1(new_n1108), .B2(new_n1115), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n928), .A2(G330), .A3(new_n759), .A4(new_n831), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n1107), .B(new_n1117), .C1(new_n1111), .C2(new_n1114), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1116), .A2(new_n765), .A3(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n858), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n766), .B1(new_n280), .B2(new_n1120), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n805), .A2(new_n497), .B1(new_n784), .B2(new_n526), .ZN(new_n1122));
  AOI211_X1 g0922(.A(new_n249), .B(new_n1122), .C1(G97), .C2(new_n811), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1123), .A2(new_n800), .A3(new_n844), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1074), .B1(G283), .B2(new_n793), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1125), .B1(new_n435), .B2(new_n802), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(KEYINPUT54), .B(G143), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n801), .A2(G137), .B1(new_n811), .B2(new_n1128), .ZN(new_n1129));
  XOR2_X1   g0929(.A(new_n1129), .B(KEYINPUT113), .Z(new_n1130));
  NOR2_X1   g0930(.A1(new_n798), .A2(new_n838), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(new_n1131), .B(KEYINPUT53), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n249), .B1(new_n805), .B2(new_n845), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1133), .B1(G125), .B2(new_n785), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n788), .A2(G50), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(G159), .A2(new_n817), .B1(new_n793), .B2(G128), .ZN(new_n1136));
  NAND4_X1  g0936(.A1(new_n1132), .A2(new_n1134), .A3(new_n1135), .A4(new_n1136), .ZN(new_n1137));
  OAI22_X1  g0937(.A1(new_n1124), .A2(new_n1126), .B1(new_n1130), .B2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1121), .B1(new_n1138), .B2(new_n778), .ZN(new_n1139));
  XOR2_X1   g0939(.A(new_n1139), .B(KEYINPUT114), .Z(new_n1140));
  INV_X1    g0940(.A(new_n1102), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1140), .B1(new_n1141), .B2(new_n776), .ZN(new_n1142));
  AND3_X1   g0942(.A1(new_n1119), .A2(KEYINPUT115), .A3(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(KEYINPUT115), .B1(new_n1119), .B2(new_n1142), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n903), .B1(new_n1105), .B2(new_n911), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n1146), .A2(new_n1103), .B1(new_n894), .B2(new_n899), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1109), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n737), .A2(new_n687), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT92), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n737), .A2(KEYINPUT92), .A3(new_n687), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1148), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n928), .B1(new_n1153), .B2(new_n828), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1114), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(new_n1147), .A2(new_n1106), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1118), .B1(new_n1156), .B2(new_n1100), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n449), .A2(G330), .A3(new_n932), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1105), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n833), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n928), .B1(new_n1160), .B2(new_n831), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1159), .B1(new_n1101), .B2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n831), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n911), .B1(new_n1099), .B2(new_n1163), .ZN(new_n1164));
  NAND4_X1  g0964(.A1(new_n1110), .A2(new_n920), .A3(new_n1117), .A4(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1162), .A2(new_n1165), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n869), .A2(new_n1158), .A3(new_n1166), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1064), .B1(new_n1157), .B2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1116), .A2(KEYINPUT112), .A3(new_n1118), .ZN(new_n1169));
  INV_X1    g0969(.A(KEYINPUT112), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1158), .ZN(new_n1171));
  AOI211_X1 g0971(.A(new_n864), .B(new_n1171), .C1(new_n866), .C2(new_n868), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n1157), .A2(new_n1170), .B1(new_n1172), .B2(new_n1166), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1168), .B1(new_n1169), .B2(new_n1173), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1097), .B1(new_n1145), .B2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1119), .A2(new_n1142), .ZN(new_n1176));
  INV_X1    g0976(.A(KEYINPUT115), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1119), .A2(KEYINPUT115), .A3(new_n1142), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1168), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1157), .A2(new_n1170), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1182), .A2(new_n1169), .A3(new_n1167), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1181), .A2(new_n1183), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1180), .A2(new_n1184), .A3(KEYINPUT116), .ZN(new_n1185));
  AND2_X1   g0985(.A1(new_n1175), .A2(new_n1185), .ZN(G378));
  NOR2_X1   g0986(.A1(new_n299), .A2(new_n888), .ZN(new_n1187));
  AND2_X1   g0987(.A1(new_n317), .A2(new_n1187), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n317), .A2(new_n1187), .ZN(new_n1189));
  OAI21_X1  g0989(.A(KEYINPUT120), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  OR2_X1    g0990(.A1(new_n317), .A2(new_n1187), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n317), .A2(new_n1187), .ZN(new_n1192));
  INV_X1    g0992(.A(KEYINPUT120), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1191), .A2(new_n1192), .A3(new_n1193), .ZN(new_n1194));
  XOR2_X1   g0994(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1195));
  AND3_X1   g0995(.A1(new_n1190), .A2(new_n1194), .A3(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1195), .B1(new_n1190), .B2(new_n1194), .ZN(new_n1197));
  NOR3_X1   g0997(.A1(new_n1196), .A2(new_n1197), .A3(new_n776), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n766), .B1(new_n1120), .B2(G50), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n253), .A2(new_n261), .ZN(new_n1200));
  OAI211_X1 g1000(.A(new_n1200), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1201));
  XNOR2_X1  g1001(.A(new_n1201), .B(KEYINPUT117), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n794), .A2(new_n497), .B1(new_n787), .B2(new_n220), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(G97), .B2(new_n801), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n429), .A2(new_n811), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n805), .A2(new_n435), .ZN(new_n1206));
  AOI211_X1 g1006(.A(new_n1200), .B(new_n1206), .C1(G283), .C2(new_n785), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(G68), .A2(new_n817), .B1(new_n815), .B2(G77), .ZN(new_n1208));
  NAND4_X1  g1008(.A1(new_n1204), .A2(new_n1205), .A3(new_n1207), .A4(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT58), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1202), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  XOR2_X1   g1011(.A(new_n1211), .B(KEYINPUT118), .Z(new_n1212));
  AOI211_X1 g1012(.A(G33), .B(G41), .C1(new_n785), .C2(G124), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1213), .B1(new_n1001), .B2(new_n787), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n801), .A2(G132), .B1(new_n811), .B2(G137), .ZN(new_n1215));
  XOR2_X1   g1015(.A(new_n1215), .B(KEYINPUT119), .Z(new_n1216));
  AOI22_X1  g1016(.A1(new_n817), .A2(G150), .B1(new_n836), .B2(G128), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(new_n793), .A2(G125), .B1(new_n815), .B2(new_n1128), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1216), .A2(new_n1217), .A3(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1214), .B1(new_n1219), .B2(KEYINPUT59), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1220), .B1(KEYINPUT59), .B2(new_n1219), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n1212), .B(new_n1221), .C1(new_n1210), .C2(new_n1209), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1199), .B1(new_n1222), .B2(new_n778), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n1198), .A2(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT121), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  OAI21_X1  g1027(.A(KEYINPUT121), .B1(new_n1198), .B2(new_n1224), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n923), .A2(new_n938), .A3(G330), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n935), .B1(new_n1113), .B2(new_n936), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n928), .A2(new_n932), .A3(new_n935), .A4(new_n831), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1233), .B1(new_n898), .B2(new_n897), .ZN(new_n1234));
  OAI21_X1  g1034(.A(G330), .B1(new_n1232), .B2(new_n1234), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1235), .A2(new_n905), .A3(new_n922), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1230), .A2(new_n1231), .A3(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1230), .B1(new_n1231), .B2(new_n1236), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n765), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1229), .A2(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1166), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1172), .B1(new_n1157), .B2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1231), .A2(new_n1236), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1230), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(new_n1237), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1243), .A2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT57), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1064), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1249), .B1(new_n1246), .B2(new_n1237), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1251), .B1(new_n1252), .B2(new_n1243), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1241), .B1(new_n1250), .B2(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(G375));
  NAND2_X1  g1055(.A1(new_n869), .A2(new_n1158), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1256), .A2(new_n1242), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n977), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1257), .A2(new_n1258), .A3(new_n1167), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n911), .A2(new_n775), .ZN(new_n1260));
  XNOR2_X1  g1060(.A(new_n1260), .B(KEYINPUT122), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n778), .ZN(new_n1262));
  OAI22_X1  g1062(.A1(new_n794), .A2(new_n845), .B1(new_n202), .B2(new_n796), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1263), .B1(G159), .B2(new_n815), .ZN(new_n1264));
  OAI22_X1  g1064(.A1(new_n805), .A2(new_n839), .B1(new_n804), .B2(new_n838), .ZN(new_n1265));
  AOI211_X1 g1065(.A(new_n253), .B(new_n1265), .C1(G128), .C2(new_n785), .ZN(new_n1266));
  AOI22_X1  g1066(.A1(new_n801), .A2(new_n1128), .B1(new_n788), .B2(G58), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1264), .A2(new_n1266), .A3(new_n1267), .ZN(new_n1268));
  OAI22_X1  g1068(.A1(new_n794), .A2(new_n526), .B1(new_n787), .B2(new_n425), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1269), .B1(G116), .B2(new_n801), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n804), .A2(new_n435), .ZN(new_n1271));
  AOI211_X1 g1071(.A(new_n249), .B(new_n1271), .C1(G283), .C2(new_n836), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1270), .A2(new_n1057), .A3(new_n1272), .ZN(new_n1273));
  OAI22_X1  g1073(.A1(new_n798), .A2(new_n222), .B1(new_n784), .B2(new_n849), .ZN(new_n1274));
  XNOR2_X1  g1074(.A(new_n1274), .B(KEYINPUT123), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1268), .B1(new_n1273), .B2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT124), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1262), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1278), .B1(new_n1277), .B2(new_n1276), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n824), .B1(new_n214), .B2(new_n858), .ZN(new_n1280));
  AND2_X1   g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  AOI22_X1  g1081(.A1(new_n1166), .A2(new_n765), .B1(new_n1261), .B2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1259), .A2(new_n1282), .ZN(G381));
  NOR2_X1   g1083(.A1(new_n1145), .A2(new_n1174), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1284), .ZN(new_n1285));
  NOR2_X1   g1085(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(new_n861), .ZN(new_n1287));
  OR4_X1    g1087(.A1(G396), .A2(G387), .A3(G393), .A4(new_n1287), .ZN(new_n1288));
  OR4_X1    g1088(.A1(new_n1285), .A2(new_n1288), .A3(G375), .A4(G381), .ZN(G407));
  INV_X1    g1089(.A(G213), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n685), .A2(new_n1290), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1254), .A2(new_n1284), .A3(new_n1291), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(G407), .A2(G213), .A3(new_n1292), .ZN(G409));
  INV_X1    g1093(.A(new_n975), .ZN(new_n1294));
  XNOR2_X1  g1094(.A(new_n974), .B(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n979), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1296), .B1(new_n1070), .B2(new_n991), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n760), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1258), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1295), .B1(new_n1299), .B2(new_n764), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1026), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1286), .B1(new_n1300), .B2(new_n1301), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n996), .A2(G390), .A3(new_n1026), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT125), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1306));
  XOR2_X1   g1106(.A(G393), .B(G396), .Z(new_n1307));
  NAND2_X1  g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1307), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1304), .A2(new_n1305), .A3(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1308), .A2(new_n1310), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1175), .A2(new_n1254), .A3(new_n1185), .ZN(new_n1312));
  OAI221_X1 g1112(.A(new_n1240), .B1(new_n1198), .B2(new_n1224), .C1(new_n1248), .C2(new_n977), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1313), .A2(new_n1284), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1312), .A2(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1291), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1317));
  AOI21_X1  g1117(.A(KEYINPUT60), .B1(new_n1256), .B2(new_n1242), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1167), .A2(new_n1064), .ZN(new_n1319));
  NOR2_X1   g1119(.A1(new_n1318), .A2(new_n1319), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1256), .A2(KEYINPUT60), .A3(new_n1242), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1322), .A2(G384), .A3(new_n1282), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1323), .ZN(new_n1324));
  AOI21_X1  g1124(.A(G384), .B1(new_n1322), .B2(new_n1282), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1291), .A2(G2897), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1326), .ZN(new_n1327));
  NOR3_X1   g1127(.A1(new_n1324), .A2(new_n1325), .A3(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1321), .ZN(new_n1329));
  NOR3_X1   g1129(.A1(new_n1329), .A2(new_n1318), .A3(new_n1319), .ZN(new_n1330));
  INV_X1    g1130(.A(new_n1282), .ZN(new_n1331));
  OAI21_X1  g1131(.A(new_n861), .B1(new_n1330), .B2(new_n1331), .ZN(new_n1332));
  AOI21_X1  g1132(.A(new_n1326), .B1(new_n1332), .B2(new_n1323), .ZN(new_n1333));
  NOR2_X1   g1133(.A1(new_n1328), .A2(new_n1333), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1317), .A2(new_n1334), .ZN(new_n1335));
  INV_X1    g1135(.A(KEYINPUT61), .ZN(new_n1336));
  AOI21_X1  g1136(.A(KEYINPUT126), .B1(new_n1335), .B2(new_n1336), .ZN(new_n1337));
  NOR2_X1   g1137(.A1(new_n1324), .A2(new_n1325), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1315), .A2(new_n1316), .A3(new_n1338), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1339), .A2(KEYINPUT62), .ZN(new_n1340));
  AOI21_X1  g1140(.A(new_n1291), .B1(new_n1312), .B2(new_n1314), .ZN(new_n1341));
  INV_X1    g1141(.A(KEYINPUT62), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1341), .A2(new_n1342), .A3(new_n1338), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1340), .A2(new_n1343), .ZN(new_n1344));
  OAI21_X1  g1144(.A(new_n1311), .B1(new_n1337), .B2(new_n1344), .ZN(new_n1345));
  AOI21_X1  g1145(.A(new_n1309), .B1(new_n1304), .B2(new_n1305), .ZN(new_n1346));
  AOI211_X1 g1146(.A(KEYINPUT125), .B(new_n1307), .C1(new_n1302), .C2(new_n1303), .ZN(new_n1347));
  NOR2_X1   g1147(.A1(new_n1346), .A2(new_n1347), .ZN(new_n1348));
  AND3_X1   g1148(.A1(new_n1341), .A2(KEYINPUT63), .A3(new_n1338), .ZN(new_n1349));
  AOI21_X1  g1149(.A(KEYINPUT63), .B1(new_n1341), .B2(new_n1338), .ZN(new_n1350));
  OAI21_X1  g1150(.A(new_n1348), .B1(new_n1349), .B2(new_n1350), .ZN(new_n1351));
  INV_X1    g1151(.A(KEYINPUT126), .ZN(new_n1352));
  OAI21_X1  g1152(.A(new_n1352), .B1(new_n1346), .B2(new_n1347), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1338), .A2(new_n1326), .ZN(new_n1354));
  INV_X1    g1154(.A(new_n1333), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1354), .A2(new_n1355), .ZN(new_n1356));
  OAI211_X1 g1156(.A(new_n1353), .B(new_n1336), .C1(new_n1356), .C2(new_n1341), .ZN(new_n1357));
  INV_X1    g1157(.A(new_n1357), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1351), .A2(new_n1358), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1345), .A2(new_n1359), .ZN(G405));
  NAND3_X1  g1160(.A1(new_n1311), .A2(KEYINPUT127), .A3(new_n1338), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1338), .A2(KEYINPUT127), .ZN(new_n1362));
  NAND2_X1  g1162(.A1(new_n1348), .A2(new_n1362), .ZN(new_n1363));
  NAND2_X1  g1163(.A1(new_n1361), .A2(new_n1363), .ZN(new_n1364));
  NOR2_X1   g1164(.A1(new_n1338), .A2(KEYINPUT127), .ZN(new_n1365));
  NAND2_X1  g1165(.A1(G375), .A2(new_n1284), .ZN(new_n1366));
  AOI21_X1  g1166(.A(new_n1365), .B1(new_n1312), .B2(new_n1366), .ZN(new_n1367));
  XNOR2_X1  g1167(.A(new_n1364), .B(new_n1367), .ZN(G402));
endmodule


