

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710;

  NOR2_X1 U366 ( .A1(n709), .A2(n704), .ZN(n565) );
  XNOR2_X1 U367 ( .A(G146), .B(G125), .ZN(n447) );
  XNOR2_X2 U368 ( .A(n461), .B(KEYINPUT4), .ZN(n694) );
  XNOR2_X2 U369 ( .A(n474), .B(n678), .ZN(n399) );
  XNOR2_X2 U370 ( .A(n694), .B(G101), .ZN(n474) );
  XNOR2_X1 U371 ( .A(n447), .B(KEYINPUT10), .ZN(n487) );
  XNOR2_X1 U372 ( .A(n677), .B(n434), .ZN(n471) );
  INV_X1 U373 ( .A(KEYINPUT72), .ZN(n434) );
  NAND2_X1 U374 ( .A1(n384), .A2(n566), .ZN(n506) );
  XNOR2_X1 U375 ( .A(n518), .B(n385), .ZN(n384) );
  INV_X1 U376 ( .A(KEYINPUT100), .ZN(n385) );
  XNOR2_X1 U377 ( .A(KEYINPUT13), .B(G475), .ZN(n397) );
  OR2_X1 U378 ( .A1(n669), .A2(G902), .ZN(n398) );
  INV_X1 U379 ( .A(n575), .ZN(n396) );
  INV_X1 U380 ( .A(n559), .ZN(n624) );
  XOR2_X1 U381 ( .A(G137), .B(G140), .Z(n488) );
  XNOR2_X1 U382 ( .A(n426), .B(n427), .ZN(n415) );
  XOR2_X1 U383 ( .A(KEYINPUT17), .B(KEYINPUT85), .Z(n427) );
  XOR2_X1 U384 ( .A(KEYINPUT79), .B(KEYINPUT18), .Z(n425) );
  INV_X1 U385 ( .A(n598), .ZN(n407) );
  XNOR2_X1 U386 ( .A(n410), .B(n409), .ZN(n408) );
  INV_X1 U387 ( .A(KEYINPUT44), .ZN(n409) );
  AND2_X1 U388 ( .A1(n706), .A2(n708), .ZN(n513) );
  INV_X1 U389 ( .A(KEYINPUT48), .ZN(n401) );
  AND2_X1 U390 ( .A1(n618), .A2(n574), .ZN(n402) );
  NAND2_X1 U391 ( .A1(n624), .A2(n623), .ZN(n627) );
  XNOR2_X1 U392 ( .A(n577), .B(KEYINPUT38), .ZN(n559) );
  XNOR2_X1 U393 ( .A(n535), .B(KEYINPUT1), .ZN(n642) );
  XOR2_X1 U394 ( .A(KEYINPUT16), .B(G122), .Z(n676) );
  XOR2_X1 U395 ( .A(KEYINPUT24), .B(G110), .Z(n490) );
  XNOR2_X1 U396 ( .A(n487), .B(n377), .ZN(n692) );
  INV_X1 U397 ( .A(n488), .ZN(n377) );
  XNOR2_X1 U398 ( .A(G134), .B(G107), .ZN(n457) );
  XNOR2_X1 U399 ( .A(G116), .B(G122), .ZN(n458) );
  XOR2_X1 U400 ( .A(KEYINPUT94), .B(KEYINPUT93), .Z(n459) );
  XNOR2_X1 U401 ( .A(n456), .B(n487), .ZN(n669) );
  XNOR2_X1 U402 ( .A(n388), .B(n472), .ZN(n665) );
  NAND2_X1 U403 ( .A1(G234), .A2(G237), .ZN(n441) );
  INV_X1 U404 ( .A(n552), .ZN(n577) );
  NOR2_X1 U405 ( .A1(n372), .A2(n439), .ZN(n395) );
  XNOR2_X1 U406 ( .A(n568), .B(KEYINPUT102), .ZN(n575) );
  AND2_X1 U407 ( .A1(n566), .A2(n567), .ZN(n391) );
  OR2_X1 U408 ( .A1(n594), .A2(G902), .ZN(n380) );
  INV_X1 U409 ( .A(KEYINPUT98), .ZN(n374) );
  XNOR2_X1 U410 ( .A(n639), .B(n486), .ZN(n566) );
  XNOR2_X1 U411 ( .A(KEYINPUT97), .B(KEYINPUT6), .ZN(n486) );
  XNOR2_X1 U412 ( .A(n498), .B(n497), .ZN(n636) );
  XNOR2_X1 U413 ( .A(n496), .B(n495), .ZN(n497) );
  INV_X1 U414 ( .A(KEYINPUT25), .ZN(n495) );
  XNOR2_X1 U415 ( .A(n379), .B(n564), .ZN(n709) );
  XNOR2_X1 U416 ( .A(G146), .B(G137), .ZN(n476) );
  NOR2_X1 U417 ( .A1(G953), .A2(G237), .ZN(n479) );
  XNOR2_X1 U418 ( .A(n471), .B(n473), .ZN(n389) );
  NAND2_X1 U419 ( .A1(n642), .A2(n641), .ZN(n518) );
  OR2_X1 U420 ( .A1(n665), .A2(G902), .ZN(n373) );
  XNOR2_X1 U421 ( .A(n414), .B(n412), .ZN(n411) );
  XNOR2_X1 U422 ( .A(n424), .B(n413), .ZN(n412) );
  XNOR2_X1 U423 ( .A(n471), .B(n415), .ZN(n414) );
  AND2_X1 U424 ( .A1(n583), .A2(n581), .ZN(n699) );
  NAND2_X1 U425 ( .A1(n408), .A2(n406), .ZN(n387) );
  AND2_X1 U426 ( .A1(n525), .A2(n407), .ZN(n406) );
  XNOR2_X1 U427 ( .A(n404), .B(n403), .ZN(n656) );
  XNOR2_X1 U428 ( .A(n553), .B(KEYINPUT106), .ZN(n403) );
  NOR2_X1 U429 ( .A1(n627), .A2(n626), .ZN(n404) );
  INV_X1 U430 ( .A(KEYINPUT39), .ZN(n562) );
  NOR2_X1 U431 ( .A1(n561), .A2(n560), .ZN(n563) );
  XNOR2_X1 U432 ( .A(n569), .B(KEYINPUT19), .ZN(n537) );
  INV_X1 U433 ( .A(KEYINPUT64), .ZN(n405) );
  XNOR2_X1 U434 ( .A(n376), .B(n375), .ZN(n673) );
  XNOR2_X1 U435 ( .A(n491), .B(G128), .ZN(n375) );
  XNOR2_X1 U436 ( .A(n493), .B(n692), .ZN(n376) );
  XNOR2_X1 U437 ( .A(n462), .B(n371), .ZN(n467) );
  XNOR2_X1 U438 ( .A(n463), .B(n344), .ZN(n371) );
  INV_X1 U439 ( .A(G953), .ZN(n685) );
  XNOR2_X1 U440 ( .A(n394), .B(n393), .ZN(n576) );
  XNOR2_X1 U441 ( .A(KEYINPUT43), .B(KEYINPUT103), .ZN(n393) );
  NAND2_X1 U442 ( .A1(n396), .A2(n395), .ZN(n394) );
  XNOR2_X1 U443 ( .A(KEYINPUT36), .B(KEYINPUT110), .ZN(n570) );
  NOR2_X1 U444 ( .A1(n511), .A2(n510), .ZN(n512) );
  XNOR2_X1 U445 ( .A(n504), .B(KEYINPUT32), .ZN(n708) );
  AND2_X1 U446 ( .A1(n502), .A2(n346), .ZN(n503) );
  INV_X1 U447 ( .A(KEYINPUT99), .ZN(n382) );
  XNOR2_X1 U448 ( .A(n392), .B(KEYINPUT95), .ZN(n611) );
  INV_X1 U449 ( .A(KEYINPUT60), .ZN(n358) );
  INV_X1 U450 ( .A(KEYINPUT122), .ZN(n362) );
  BUF_X1 U451 ( .A(n642), .Z(n372) );
  XNOR2_X1 U452 ( .A(KEYINPUT9), .B(KEYINPUT7), .ZN(n344) );
  AND2_X1 U453 ( .A1(n505), .A2(n533), .ZN(n641) );
  AND2_X1 U454 ( .A1(n699), .A2(n580), .ZN(n345) );
  NOR2_X1 U455 ( .A1(n566), .A2(n416), .ZN(n346) );
  XOR2_X1 U456 ( .A(KEYINPUT68), .B(KEYINPUT0), .Z(n347) );
  XOR2_X1 U457 ( .A(KEYINPUT22), .B(KEYINPUT74), .Z(n348) );
  XOR2_X1 U458 ( .A(KEYINPUT65), .B(KEYINPUT45), .Z(n349) );
  XOR2_X1 U459 ( .A(n588), .B(KEYINPUT124), .Z(n350) );
  XOR2_X1 U460 ( .A(n596), .B(n595), .Z(n351) );
  XOR2_X1 U461 ( .A(n669), .B(n418), .Z(n352) );
  XOR2_X1 U462 ( .A(n592), .B(n591), .Z(n353) );
  XOR2_X1 U463 ( .A(n667), .B(n666), .Z(n354) );
  XOR2_X1 U464 ( .A(n420), .B(KEYINPUT67), .Z(n355) );
  XOR2_X1 U465 ( .A(KEYINPUT56), .B(KEYINPUT120), .Z(n356) );
  INV_X1 U466 ( .A(n675), .ZN(n367) );
  XNOR2_X1 U467 ( .A(n383), .B(n382), .ZN(n514) );
  XNOR2_X1 U468 ( .A(n500), .B(n374), .ZN(n370) );
  XNOR2_X1 U469 ( .A(n357), .B(KEYINPUT125), .ZN(G63) );
  NAND2_X1 U470 ( .A1(n366), .A2(n367), .ZN(n357) );
  XNOR2_X1 U471 ( .A(n359), .B(n358), .ZN(G60) );
  NAND2_X1 U472 ( .A1(n364), .A2(n367), .ZN(n359) );
  XNOR2_X1 U473 ( .A(n360), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U474 ( .A1(n365), .A2(n367), .ZN(n360) );
  XNOR2_X1 U475 ( .A(n361), .B(n356), .ZN(G51) );
  NAND2_X1 U476 ( .A1(n369), .A2(n367), .ZN(n361) );
  XNOR2_X1 U477 ( .A(n363), .B(n362), .ZN(G54) );
  NAND2_X1 U478 ( .A1(n368), .A2(n367), .ZN(n363) );
  XNOR2_X1 U479 ( .A(n670), .B(n352), .ZN(n364) );
  XNOR2_X1 U480 ( .A(n597), .B(n351), .ZN(n365) );
  XNOR2_X1 U481 ( .A(n589), .B(n350), .ZN(n366) );
  XNOR2_X1 U482 ( .A(n668), .B(n354), .ZN(n368) );
  XNOR2_X1 U483 ( .A(n593), .B(n353), .ZN(n369) );
  NAND2_X1 U484 ( .A1(n370), .A2(n501), .ZN(n383) );
  NOR2_X2 U485 ( .A1(n586), .A2(n585), .ZN(n390) );
  NAND2_X1 U486 ( .A1(n514), .A2(n513), .ZN(n410) );
  XNOR2_X1 U487 ( .A(n378), .B(n401), .ZN(n583) );
  XNOR2_X1 U488 ( .A(n571), .B(n570), .ZN(n572) );
  NAND2_X1 U489 ( .A1(n517), .A2(n516), .ZN(n392) );
  XNOR2_X1 U490 ( .A(n563), .B(n562), .ZN(n578) );
  XNOR2_X2 U491 ( .A(n373), .B(n475), .ZN(n535) );
  NAND2_X2 U492 ( .A1(n502), .A2(n416), .ZN(n500) );
  NAND2_X1 U493 ( .A1(n573), .A2(n402), .ZN(n378) );
  NAND2_X1 U494 ( .A1(n578), .A2(n611), .ZN(n379) );
  NAND2_X1 U495 ( .A1(n639), .A2(n623), .ZN(n542) );
  XNOR2_X2 U496 ( .A(n380), .B(n485), .ZN(n639) );
  XNOR2_X1 U497 ( .A(n399), .B(n484), .ZN(n594) );
  NAND2_X1 U498 ( .A1(n520), .A2(n470), .ZN(n417) );
  XNOR2_X2 U499 ( .A(n381), .B(n347), .ZN(n520) );
  NAND2_X1 U500 ( .A1(n537), .A2(n443), .ZN(n381) );
  INV_X1 U501 ( .A(n514), .ZN(n707) );
  AND2_X2 U502 ( .A1(n386), .A2(n355), .ZN(n587) );
  NAND2_X1 U503 ( .A1(n686), .A2(n345), .ZN(n386) );
  XNOR2_X2 U504 ( .A(n387), .B(n349), .ZN(n686) );
  XNOR2_X1 U505 ( .A(n474), .B(n389), .ZN(n388) );
  NOR2_X1 U506 ( .A1(n660), .A2(n390), .ZN(n661) );
  NOR2_X4 U507 ( .A1(n587), .A2(n390), .ZN(n671) );
  NAND2_X1 U508 ( .A1(n611), .A2(n391), .ZN(n568) );
  XNOR2_X2 U509 ( .A(n398), .B(n397), .ZN(n515) );
  XNOR2_X1 U510 ( .A(n399), .B(n411), .ZN(n590) );
  XNOR2_X2 U511 ( .A(n400), .B(G143), .ZN(n461) );
  XNOR2_X2 U512 ( .A(G128), .B(KEYINPUT66), .ZN(n400) );
  XNOR2_X2 U513 ( .A(n405), .B(G953), .ZN(n700) );
  XNOR2_X1 U514 ( .A(n425), .B(n447), .ZN(n413) );
  INV_X1 U515 ( .A(n372), .ZN(n416) );
  XNOR2_X2 U516 ( .A(n417), .B(n348), .ZN(n502) );
  XNOR2_X1 U517 ( .A(KEYINPUT123), .B(KEYINPUT59), .ZN(n418) );
  AND2_X1 U518 ( .A1(G227), .A2(n700), .ZN(n419) );
  XNOR2_X1 U519 ( .A(n691), .B(n419), .ZN(n472) );
  AND2_X1 U520 ( .A1(n442), .A2(n530), .ZN(n443) );
  XNOR2_X1 U521 ( .A(n490), .B(n489), .ZN(n491) );
  NOR2_X1 U522 ( .A1(n639), .A2(n533), .ZN(n501) );
  NOR2_X1 U523 ( .A1(n700), .A2(G952), .ZN(n675) );
  XNOR2_X1 U524 ( .A(G902), .B(KEYINPUT15), .ZN(n444) );
  INV_X1 U525 ( .A(n444), .ZN(n580) );
  NAND2_X1 U526 ( .A1(n580), .A2(KEYINPUT2), .ZN(n420) );
  XOR2_X1 U527 ( .A(KEYINPUT71), .B(G119), .Z(n422) );
  XNOR2_X1 U528 ( .A(G116), .B(G113), .ZN(n421) );
  XNOR2_X1 U529 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U530 ( .A(KEYINPUT3), .B(n423), .Z(n678) );
  XNOR2_X1 U531 ( .A(n676), .B(KEYINPUT80), .ZN(n424) );
  NAND2_X1 U532 ( .A1(G224), .A2(n700), .ZN(n426) );
  INV_X1 U533 ( .A(G107), .ZN(n428) );
  NAND2_X1 U534 ( .A1(G104), .A2(n428), .ZN(n431) );
  INV_X1 U535 ( .A(G104), .ZN(n429) );
  NAND2_X1 U536 ( .A1(n429), .A2(G107), .ZN(n430) );
  NAND2_X1 U537 ( .A1(n431), .A2(n430), .ZN(n433) );
  XNOR2_X2 U538 ( .A(G110), .B(KEYINPUT78), .ZN(n432) );
  XNOR2_X2 U539 ( .A(n433), .B(n432), .ZN(n677) );
  OR2_X2 U540 ( .A1(n590), .A2(n580), .ZN(n437) );
  NOR2_X1 U541 ( .A1(G237), .A2(G902), .ZN(n435) );
  XOR2_X1 U542 ( .A(KEYINPUT76), .B(n435), .Z(n438) );
  NAND2_X1 U543 ( .A1(n438), .A2(G210), .ZN(n436) );
  XNOR2_X2 U544 ( .A(n437), .B(n436), .ZN(n552) );
  NAND2_X1 U545 ( .A1(n438), .A2(G214), .ZN(n623) );
  INV_X1 U546 ( .A(n623), .ZN(n439) );
  OR2_X2 U547 ( .A1(n552), .A2(n439), .ZN(n569) );
  NOR2_X1 U548 ( .A1(G898), .A2(n685), .ZN(n681) );
  NAND2_X1 U549 ( .A1(n681), .A2(G902), .ZN(n440) );
  NAND2_X1 U550 ( .A1(G952), .A2(n685), .ZN(n528) );
  NAND2_X1 U551 ( .A1(n440), .A2(n528), .ZN(n442) );
  XNOR2_X1 U552 ( .A(KEYINPUT14), .B(n441), .ZN(n530) );
  INV_X1 U553 ( .A(n530), .ZN(n654) );
  NAND2_X1 U554 ( .A1(n444), .A2(G234), .ZN(n445) );
  XNOR2_X1 U555 ( .A(n445), .B(KEYINPUT20), .ZN(n494) );
  NAND2_X1 U556 ( .A1(G221), .A2(n494), .ZN(n446) );
  XNOR2_X1 U557 ( .A(KEYINPUT21), .B(n446), .ZN(n635) );
  XOR2_X1 U558 ( .A(KEYINPUT88), .B(n635), .Z(n505) );
  XOR2_X1 U559 ( .A(G104), .B(G140), .Z(n449) );
  XNOR2_X1 U560 ( .A(G143), .B(G131), .ZN(n448) );
  XNOR2_X1 U561 ( .A(n449), .B(n448), .ZN(n453) );
  XOR2_X1 U562 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n451) );
  XNOR2_X1 U563 ( .A(G113), .B(G122), .ZN(n450) );
  XNOR2_X1 U564 ( .A(n451), .B(n450), .ZN(n452) );
  XOR2_X1 U565 ( .A(n453), .B(n452), .Z(n455) );
  NAND2_X1 U566 ( .A1(G214), .A2(n479), .ZN(n454) );
  XNOR2_X1 U567 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U568 ( .A(n457), .B(KEYINPUT92), .ZN(n463) );
  XNOR2_X1 U569 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U570 ( .A(n461), .B(n460), .ZN(n462) );
  NAND2_X1 U571 ( .A1(n700), .A2(G234), .ZN(n465) );
  XNOR2_X1 U572 ( .A(KEYINPUT83), .B(KEYINPUT8), .ZN(n464) );
  XNOR2_X1 U573 ( .A(n465), .B(n464), .ZN(n492) );
  NAND2_X1 U574 ( .A1(G217), .A2(n492), .ZN(n466) );
  XNOR2_X1 U575 ( .A(n467), .B(n466), .ZN(n588) );
  NOR2_X1 U576 ( .A1(n588), .A2(G902), .ZN(n468) );
  XNOR2_X1 U577 ( .A(n468), .B(G478), .ZN(n516) );
  NAND2_X1 U578 ( .A1(n515), .A2(n516), .ZN(n626) );
  INV_X1 U579 ( .A(n626), .ZN(n469) );
  AND2_X1 U580 ( .A1(n505), .A2(n469), .ZN(n470) );
  XOR2_X1 U581 ( .A(G131), .B(G134), .Z(n478) );
  XOR2_X1 U582 ( .A(KEYINPUT87), .B(n478), .Z(n691) );
  XNOR2_X1 U583 ( .A(G146), .B(n488), .ZN(n473) );
  XNOR2_X1 U584 ( .A(KEYINPUT70), .B(G469), .ZN(n475) );
  XOR2_X1 U585 ( .A(KEYINPUT5), .B(KEYINPUT89), .Z(n477) );
  XNOR2_X1 U586 ( .A(n477), .B(n476), .ZN(n483) );
  XOR2_X1 U587 ( .A(n478), .B(KEYINPUT77), .Z(n481) );
  NAND2_X1 U588 ( .A1(n479), .A2(G210), .ZN(n480) );
  XNOR2_X1 U589 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U590 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U591 ( .A(G472), .B(KEYINPUT90), .ZN(n485) );
  XOR2_X1 U592 ( .A(G119), .B(KEYINPUT23), .Z(n489) );
  NAND2_X1 U593 ( .A1(n492), .A2(G221), .ZN(n493) );
  NOR2_X1 U594 ( .A1(G902), .A2(n673), .ZN(n498) );
  NAND2_X1 U595 ( .A1(G217), .A2(n494), .ZN(n496) );
  OR2_X1 U596 ( .A1(n566), .A2(n636), .ZN(n499) );
  NOR2_X1 U597 ( .A1(n500), .A2(n499), .ZN(n598) );
  INV_X1 U598 ( .A(n639), .ZN(n521) );
  INV_X1 U599 ( .A(n636), .ZN(n533) );
  NAND2_X1 U600 ( .A1(n503), .A2(n636), .ZN(n504) );
  XNOR2_X1 U601 ( .A(n506), .B(KEYINPUT33), .ZN(n632) );
  NAND2_X1 U602 ( .A1(n632), .A2(n520), .ZN(n508) );
  XOR2_X1 U603 ( .A(KEYINPUT73), .B(KEYINPUT34), .Z(n507) );
  XNOR2_X1 U604 ( .A(n508), .B(n507), .ZN(n511) );
  OR2_X1 U605 ( .A1(n515), .A2(n516), .ZN(n509) );
  XOR2_X1 U606 ( .A(KEYINPUT101), .B(n509), .Z(n545) );
  XOR2_X1 U607 ( .A(KEYINPUT81), .B(n545), .Z(n510) );
  XNOR2_X1 U608 ( .A(n512), .B(KEYINPUT35), .ZN(n706) );
  XNOR2_X1 U609 ( .A(n515), .B(KEYINPUT91), .ZN(n517) );
  NOR2_X1 U610 ( .A1(n517), .A2(n516), .ZN(n613) );
  NOR2_X1 U611 ( .A1(n611), .A2(n613), .ZN(n628) );
  NOR2_X1 U612 ( .A1(n521), .A2(n518), .ZN(n647) );
  NAND2_X1 U613 ( .A1(n647), .A2(n520), .ZN(n519) );
  XNOR2_X1 U614 ( .A(n519), .B(KEYINPUT31), .ZN(n614) );
  NAND2_X1 U615 ( .A1(n641), .A2(n535), .ZN(n541) );
  NAND2_X1 U616 ( .A1(n521), .A2(n520), .ZN(n522) );
  NOR2_X1 U617 ( .A1(n541), .A2(n522), .ZN(n603) );
  NOR2_X1 U618 ( .A1(n614), .A2(n603), .ZN(n523) );
  NOR2_X1 U619 ( .A1(n628), .A2(n523), .ZN(n524) );
  XOR2_X1 U620 ( .A(KEYINPUT96), .B(n524), .Z(n525) );
  NOR2_X1 U621 ( .A1(KEYINPUT47), .A2(KEYINPUT75), .ZN(n540) );
  NOR2_X1 U622 ( .A1(G900), .A2(n700), .ZN(n526) );
  NAND2_X1 U623 ( .A1(G902), .A2(n526), .ZN(n527) );
  NAND2_X1 U624 ( .A1(n528), .A2(n527), .ZN(n529) );
  NAND2_X1 U625 ( .A1(n530), .A2(n529), .ZN(n558) );
  NOR2_X1 U626 ( .A1(n635), .A2(n558), .ZN(n531) );
  XNOR2_X1 U627 ( .A(n531), .B(KEYINPUT69), .ZN(n532) );
  NOR2_X1 U628 ( .A1(n533), .A2(n532), .ZN(n567) );
  AND2_X1 U629 ( .A1(n639), .A2(n567), .ZN(n534) );
  XNOR2_X1 U630 ( .A(n534), .B(KEYINPUT28), .ZN(n536) );
  AND2_X1 U631 ( .A1(n536), .A2(n535), .ZN(n554) );
  AND2_X1 U632 ( .A1(n537), .A2(n554), .ZN(n608) );
  INV_X1 U633 ( .A(n628), .ZN(n538) );
  NAND2_X1 U634 ( .A1(n608), .A2(n538), .ZN(n539) );
  XNOR2_X1 U635 ( .A(n540), .B(n539), .ZN(n551) );
  NAND2_X1 U636 ( .A1(KEYINPUT47), .A2(KEYINPUT75), .ZN(n549) );
  INV_X1 U637 ( .A(n541), .ZN(n544) );
  XOR2_X1 U638 ( .A(KEYINPUT30), .B(n542), .Z(n543) );
  NAND2_X1 U639 ( .A1(n544), .A2(n543), .ZN(n561) );
  NOR2_X1 U640 ( .A1(n558), .A2(n561), .ZN(n547) );
  NOR2_X1 U641 ( .A1(n552), .A2(n545), .ZN(n546) );
  NAND2_X1 U642 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U643 ( .A(KEYINPUT104), .B(n548), .ZN(n710) );
  AND2_X1 U644 ( .A1(n549), .A2(n710), .ZN(n550) );
  AND2_X1 U645 ( .A1(n551), .A2(n550), .ZN(n574) );
  XNOR2_X1 U646 ( .A(KEYINPUT107), .B(KEYINPUT41), .ZN(n553) );
  NAND2_X1 U647 ( .A1(n656), .A2(n554), .ZN(n557) );
  XNOR2_X1 U648 ( .A(KEYINPUT109), .B(KEYINPUT42), .ZN(n555) );
  XNOR2_X1 U649 ( .A(n555), .B(KEYINPUT108), .ZN(n556) );
  XNOR2_X1 U650 ( .A(n557), .B(n556), .ZN(n704) );
  XNOR2_X1 U651 ( .A(KEYINPUT40), .B(KEYINPUT105), .ZN(n564) );
  OR2_X1 U652 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U653 ( .A(n565), .B(KEYINPUT46), .ZN(n573) );
  NOR2_X1 U654 ( .A1(n569), .A2(n575), .ZN(n571) );
  NAND2_X1 U655 ( .A1(n572), .A2(n372), .ZN(n618) );
  NOR2_X1 U656 ( .A1(n577), .A2(n576), .ZN(n621) );
  NAND2_X1 U657 ( .A1(n613), .A2(n578), .ZN(n620) );
  INV_X1 U658 ( .A(n620), .ZN(n579) );
  NOR2_X1 U659 ( .A1(n621), .A2(n579), .ZN(n581) );
  INV_X1 U660 ( .A(n686), .ZN(n586) );
  AND2_X1 U661 ( .A1(n581), .A2(KEYINPUT2), .ZN(n582) );
  NAND2_X1 U662 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U663 ( .A(KEYINPUT84), .B(n584), .ZN(n585) );
  NAND2_X1 U664 ( .A1(n671), .A2(G478), .ZN(n589) );
  XOR2_X1 U665 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n592) );
  XNOR2_X1 U666 ( .A(n590), .B(KEYINPUT82), .ZN(n591) );
  NAND2_X1 U667 ( .A1(n671), .A2(G210), .ZN(n593) );
  NAND2_X1 U668 ( .A1(n671), .A2(G472), .ZN(n597) );
  XNOR2_X1 U669 ( .A(n594), .B(KEYINPUT62), .ZN(n596) );
  XOR2_X1 U670 ( .A(KEYINPUT86), .B(KEYINPUT111), .Z(n595) );
  XOR2_X1 U671 ( .A(G101), .B(n598), .Z(G3) );
  NAND2_X1 U672 ( .A1(n603), .A2(n611), .ZN(n599) );
  XNOR2_X1 U673 ( .A(n599), .B(G104), .ZN(G6) );
  XOR2_X1 U674 ( .A(KEYINPUT27), .B(KEYINPUT113), .Z(n601) );
  XNOR2_X1 U675 ( .A(G107), .B(KEYINPUT26), .ZN(n600) );
  XNOR2_X1 U676 ( .A(n601), .B(n600), .ZN(n602) );
  XOR2_X1 U677 ( .A(KEYINPUT112), .B(n602), .Z(n605) );
  NAND2_X1 U678 ( .A1(n603), .A2(n613), .ZN(n604) );
  XNOR2_X1 U679 ( .A(n605), .B(n604), .ZN(G9) );
  XOR2_X1 U680 ( .A(G128), .B(KEYINPUT29), .Z(n607) );
  NAND2_X1 U681 ( .A1(n608), .A2(n613), .ZN(n606) );
  XNOR2_X1 U682 ( .A(n607), .B(n606), .ZN(G30) );
  NAND2_X1 U683 ( .A1(n608), .A2(n611), .ZN(n609) );
  XNOR2_X1 U684 ( .A(n609), .B(KEYINPUT114), .ZN(n610) );
  XNOR2_X1 U685 ( .A(G146), .B(n610), .ZN(G48) );
  NAND2_X1 U686 ( .A1(n614), .A2(n611), .ZN(n612) );
  XNOR2_X1 U687 ( .A(n612), .B(G113), .ZN(G15) );
  XOR2_X1 U688 ( .A(G116), .B(KEYINPUT115), .Z(n616) );
  NAND2_X1 U689 ( .A1(n614), .A2(n613), .ZN(n615) );
  XNOR2_X1 U690 ( .A(n616), .B(n615), .ZN(G18) );
  XOR2_X1 U691 ( .A(KEYINPUT37), .B(KEYINPUT116), .Z(n617) );
  XNOR2_X1 U692 ( .A(n618), .B(n617), .ZN(n619) );
  XNOR2_X1 U693 ( .A(G125), .B(n619), .ZN(G27) );
  XNOR2_X1 U694 ( .A(G134), .B(n620), .ZN(G36) );
  XNOR2_X1 U695 ( .A(G140), .B(n621), .ZN(n622) );
  XNOR2_X1 U696 ( .A(n622), .B(KEYINPUT117), .ZN(G42) );
  NOR2_X1 U697 ( .A1(n624), .A2(n623), .ZN(n625) );
  NOR2_X1 U698 ( .A1(n626), .A2(n625), .ZN(n630) );
  NOR2_X1 U699 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U700 ( .A1(n630), .A2(n629), .ZN(n631) );
  XNOR2_X1 U701 ( .A(n631), .B(KEYINPUT119), .ZN(n634) );
  BUF_X1 U702 ( .A(n632), .Z(n633) );
  NAND2_X1 U703 ( .A1(n634), .A2(n633), .ZN(n651) );
  AND2_X1 U704 ( .A1(n636), .A2(n635), .ZN(n637) );
  XOR2_X1 U705 ( .A(KEYINPUT49), .B(n637), .Z(n638) );
  NOR2_X1 U706 ( .A1(n639), .A2(n638), .ZN(n640) );
  XOR2_X1 U707 ( .A(KEYINPUT118), .B(n640), .Z(n645) );
  NOR2_X1 U708 ( .A1(n372), .A2(n641), .ZN(n643) );
  XNOR2_X1 U709 ( .A(KEYINPUT50), .B(n643), .ZN(n644) );
  NOR2_X1 U710 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U711 ( .A1(n647), .A2(n646), .ZN(n648) );
  XNOR2_X1 U712 ( .A(n648), .B(KEYINPUT51), .ZN(n649) );
  NAND2_X1 U713 ( .A1(n649), .A2(n656), .ZN(n650) );
  NAND2_X1 U714 ( .A1(n651), .A2(n650), .ZN(n652) );
  XOR2_X1 U715 ( .A(KEYINPUT52), .B(n652), .Z(n653) );
  NOR2_X1 U716 ( .A1(n654), .A2(n653), .ZN(n655) );
  NAND2_X1 U717 ( .A1(G952), .A2(n655), .ZN(n658) );
  NAND2_X1 U718 ( .A1(n633), .A2(n656), .ZN(n657) );
  NAND2_X1 U719 ( .A1(n658), .A2(n657), .ZN(n662) );
  AND2_X1 U720 ( .A1(n686), .A2(n699), .ZN(n659) );
  NOR2_X1 U721 ( .A1(n659), .A2(KEYINPUT2), .ZN(n660) );
  NOR2_X1 U722 ( .A1(n662), .A2(n661), .ZN(n663) );
  NAND2_X1 U723 ( .A1(n685), .A2(n663), .ZN(n664) );
  XOR2_X1 U724 ( .A(KEYINPUT53), .B(n664), .Z(G75) );
  XNOR2_X1 U725 ( .A(KEYINPUT58), .B(KEYINPUT121), .ZN(n667) );
  XNOR2_X1 U726 ( .A(n665), .B(KEYINPUT57), .ZN(n666) );
  NAND2_X1 U727 ( .A1(n671), .A2(G469), .ZN(n668) );
  NAND2_X1 U728 ( .A1(n671), .A2(G475), .ZN(n670) );
  NAND2_X1 U729 ( .A1(G217), .A2(n671), .ZN(n672) );
  XNOR2_X1 U730 ( .A(n673), .B(n672), .ZN(n674) );
  NOR2_X1 U731 ( .A1(n675), .A2(n674), .ZN(G66) );
  XOR2_X1 U732 ( .A(n677), .B(n676), .Z(n680) );
  XNOR2_X1 U733 ( .A(G101), .B(n678), .ZN(n679) );
  XNOR2_X1 U734 ( .A(n680), .B(n679), .ZN(n682) );
  NOR2_X1 U735 ( .A1(n682), .A2(n681), .ZN(n690) );
  NAND2_X1 U736 ( .A1(G953), .A2(G224), .ZN(n683) );
  XNOR2_X1 U737 ( .A(KEYINPUT61), .B(n683), .ZN(n684) );
  NAND2_X1 U738 ( .A1(n684), .A2(G898), .ZN(n688) );
  NAND2_X1 U739 ( .A1(n686), .A2(n685), .ZN(n687) );
  NAND2_X1 U740 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U741 ( .A(n690), .B(n689), .ZN(G69) );
  XNOR2_X1 U742 ( .A(n692), .B(n691), .ZN(n693) );
  XOR2_X1 U743 ( .A(n694), .B(n693), .Z(n698) );
  XOR2_X1 U744 ( .A(KEYINPUT126), .B(n698), .Z(n695) );
  XNOR2_X1 U745 ( .A(G227), .B(n695), .ZN(n696) );
  NAND2_X1 U746 ( .A1(n696), .A2(G900), .ZN(n697) );
  NAND2_X1 U747 ( .A1(n697), .A2(G953), .ZN(n703) );
  XNOR2_X1 U748 ( .A(n699), .B(n698), .ZN(n701) );
  NAND2_X1 U749 ( .A1(n701), .A2(n700), .ZN(n702) );
  NAND2_X1 U750 ( .A1(n703), .A2(n702), .ZN(G72) );
  XNOR2_X1 U751 ( .A(G137), .B(n704), .ZN(n705) );
  XNOR2_X1 U752 ( .A(n705), .B(KEYINPUT127), .ZN(G39) );
  XNOR2_X1 U753 ( .A(n706), .B(G122), .ZN(G24) );
  XOR2_X1 U754 ( .A(n707), .B(G110), .Z(G12) );
  XNOR2_X1 U755 ( .A(G119), .B(n708), .ZN(G21) );
  XOR2_X1 U756 ( .A(n709), .B(G131), .Z(G33) );
  XNOR2_X1 U757 ( .A(G143), .B(n710), .ZN(G45) );
endmodule

