//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 1 1 1 1 1 0 1 0 1 0 0 0 0 0 0 0 0 1 0 1 0 1 0 0 1 0 0 1 0 1 1 1 0 1 0 0 1 0 0 1 0 1 0 0 1 0 0 0 0 1 1 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:14 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1200, new_n1201,
    new_n1202, new_n1203, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1253, new_n1254, new_n1255, new_n1256, new_n1257;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT64), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  INV_X1    g0012(.A(G20), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT65), .ZN(new_n215));
  OAI21_X1  g0015(.A(G50), .B1(G58), .B2(G68), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT66), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n219));
  XOR2_X1   g0019(.A(new_n219), .B(KEYINPUT67), .Z(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n223));
  NAND3_X1  g0023(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n208), .B1(new_n220), .B2(new_n224), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n211), .B1(new_n215), .B2(new_n218), .C1(new_n225), .C2(KEYINPUT1), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XOR2_X1   g0027(.A(G226), .B(G232), .Z(new_n228));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT68), .B(KEYINPUT2), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XOR2_X1   g0036(.A(G68), .B(G77), .Z(new_n237));
  XNOR2_X1  g0037(.A(G50), .B(G58), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G351));
  INV_X1    g0043(.A(KEYINPUT3), .ZN(new_n244));
  NOR2_X1   g0044(.A1(new_n244), .A2(G33), .ZN(new_n245));
  INV_X1    g0045(.A(new_n245), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n244), .A2(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(G1698), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(G222), .ZN(new_n251));
  NAND2_X1  g0051(.A1(G223), .A2(G1698), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n249), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  AOI21_X1  g0053(.A(new_n212), .B1(G33), .B2(G41), .ZN(new_n254));
  OAI211_X1 g0054(.A(new_n253), .B(new_n254), .C1(G77), .C2(new_n249), .ZN(new_n255));
  INV_X1    g0055(.A(G274), .ZN(new_n256));
  INV_X1    g0056(.A(G1), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n257), .B1(G41), .B2(G45), .ZN(new_n258));
  AOI211_X1 g0058(.A(new_n256), .B(new_n254), .C1(KEYINPUT69), .C2(new_n258), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n259), .B1(KEYINPUT69), .B2(new_n258), .ZN(new_n260));
  INV_X1    g0060(.A(G226), .ZN(new_n261));
  INV_X1    g0061(.A(new_n254), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(new_n258), .ZN(new_n263));
  OAI211_X1 g0063(.A(new_n255), .B(new_n260), .C1(new_n261), .C2(new_n263), .ZN(new_n264));
  XNOR2_X1  g0064(.A(new_n264), .B(KEYINPUT70), .ZN(new_n265));
  INV_X1    g0065(.A(G169), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NOR2_X1   g0067(.A1(G20), .A2(G33), .ZN(new_n268));
  AOI22_X1  g0068(.A1(new_n204), .A2(G20), .B1(G150), .B2(new_n268), .ZN(new_n269));
  XNOR2_X1  g0069(.A(KEYINPUT8), .B(G58), .ZN(new_n270));
  XNOR2_X1  g0070(.A(new_n270), .B(KEYINPUT71), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n213), .A2(G33), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n269), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G33), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n212), .B1(new_n208), .B2(new_n274), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n257), .A2(G13), .A3(G20), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(KEYINPUT72), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT72), .ZN(new_n278));
  NAND4_X1  g0078(.A1(new_n278), .A2(new_n257), .A3(G13), .A4(G20), .ZN(new_n279));
  AND2_X1   g0079(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  AOI22_X1  g0080(.A1(new_n273), .A2(new_n275), .B1(new_n201), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n277), .A2(new_n279), .ZN(new_n282));
  INV_X1    g0082(.A(new_n275), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n284), .B1(new_n257), .B2(G20), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n281), .B1(new_n201), .B2(new_n286), .ZN(new_n287));
  OAI211_X1 g0087(.A(new_n267), .B(new_n287), .C1(G179), .C2(new_n265), .ZN(new_n288));
  INV_X1    g0088(.A(G190), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n265), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n290), .B1(G200), .B2(new_n265), .ZN(new_n291));
  XNOR2_X1  g0091(.A(new_n287), .B(KEYINPUT9), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  AND2_X1   g0093(.A1(new_n293), .A2(KEYINPUT10), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n293), .A2(KEYINPUT10), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n288), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G238), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n260), .B1(new_n297), .B2(new_n263), .ZN(new_n298));
  INV_X1    g0098(.A(G232), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(G1698), .ZN(new_n300));
  OAI211_X1 g0100(.A(new_n249), .B(new_n300), .C1(G226), .C2(G1698), .ZN(new_n301));
  NAND2_X1  g0101(.A1(G33), .A2(G97), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n262), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  OR3_X1    g0103(.A1(new_n298), .A2(KEYINPUT13), .A3(new_n303), .ZN(new_n304));
  OAI21_X1  g0104(.A(KEYINPUT13), .B1(new_n298), .B2(new_n303), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(G200), .ZN(new_n307));
  XNOR2_X1  g0107(.A(new_n307), .B(KEYINPUT74), .ZN(new_n308));
  INV_X1    g0108(.A(new_n306), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(G190), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n280), .A2(KEYINPUT12), .A3(new_n203), .ZN(new_n311));
  INV_X1    g0111(.A(new_n268), .ZN(new_n312));
  OAI22_X1  g0112(.A1(new_n312), .A2(new_n201), .B1(new_n213), .B2(G68), .ZN(new_n313));
  INV_X1    g0113(.A(G77), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n272), .A2(new_n314), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n275), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT11), .ZN(new_n317));
  OAI221_X1 g0117(.A(new_n311), .B1(KEYINPUT12), .B2(new_n280), .C1(new_n316), .C2(new_n317), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n203), .B1(new_n286), .B2(KEYINPUT12), .ZN(new_n319));
  AOI211_X1 g0119(.A(new_n318), .B(new_n319), .C1(new_n317), .C2(new_n316), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n310), .A2(new_n320), .ZN(new_n321));
  OR2_X1    g0121(.A1(new_n308), .A2(new_n321), .ZN(new_n322));
  XNOR2_X1  g0122(.A(new_n320), .B(KEYINPUT76), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n306), .A2(G169), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n324), .A2(KEYINPUT75), .A3(KEYINPUT14), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n309), .A2(G179), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n324), .B1(KEYINPUT75), .B2(KEYINPUT14), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n323), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(G238), .A2(G1698), .ZN(new_n330));
  OAI211_X1 g0130(.A(new_n249), .B(new_n330), .C1(new_n299), .C2(G1698), .ZN(new_n331));
  XNOR2_X1  g0131(.A(KEYINPUT73), .B(G107), .ZN(new_n332));
  OAI211_X1 g0132(.A(new_n331), .B(new_n254), .C1(new_n249), .C2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(G244), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n260), .B(new_n333), .C1(new_n334), .C2(new_n263), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(G200), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n336), .B1(new_n289), .B2(new_n335), .ZN(new_n337));
  NAND2_X1  g0137(.A1(G20), .A2(G77), .ZN(new_n338));
  XOR2_X1   g0138(.A(KEYINPUT15), .B(G87), .Z(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  OAI221_X1 g0140(.A(new_n338), .B1(new_n312), .B2(new_n270), .C1(new_n340), .C2(new_n272), .ZN(new_n341));
  AOI22_X1  g0141(.A1(new_n341), .A2(new_n275), .B1(new_n314), .B2(new_n280), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n342), .B1(new_n314), .B2(new_n286), .ZN(new_n343));
  OR2_X1    g0143(.A1(new_n337), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n335), .A2(new_n266), .ZN(new_n345));
  OAI211_X1 g0145(.A(new_n345), .B(new_n343), .C1(G179), .C2(new_n335), .ZN(new_n346));
  NAND4_X1  g0146(.A1(new_n322), .A2(new_n329), .A3(new_n344), .A4(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(G58), .A2(G68), .ZN(new_n348));
  XOR2_X1   g0148(.A(new_n348), .B(KEYINPUT81), .Z(new_n349));
  OAI21_X1  g0149(.A(new_n349), .B1(G58), .B2(G68), .ZN(new_n350));
  AOI22_X1  g0150(.A1(new_n350), .A2(G20), .B1(G159), .B2(new_n268), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT77), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(new_n244), .ZN(new_n353));
  NAND2_X1  g0153(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n353), .A2(G33), .A3(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n245), .B1(new_n355), .B2(KEYINPUT78), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT78), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n353), .A2(new_n357), .A3(G33), .A4(new_n354), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(new_n213), .ZN(new_n360));
  XNOR2_X1  g0160(.A(KEYINPUT79), .B(KEYINPUT7), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n203), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(G20), .B1(new_n356), .B2(new_n358), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT79), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT7), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n364), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(KEYINPUT80), .B1(new_n363), .B2(new_n367), .ZN(new_n368));
  OAI21_X1  g0168(.A(G68), .B1(new_n364), .B2(new_n361), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT80), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n365), .A2(new_n366), .ZN(new_n371));
  AOI211_X1 g0171(.A(G20), .B(new_n371), .C1(new_n356), .C2(new_n358), .ZN(new_n372));
  NOR3_X1   g0172(.A1(new_n369), .A2(new_n370), .A3(new_n372), .ZN(new_n373));
  OAI211_X1 g0173(.A(KEYINPUT16), .B(new_n351), .C1(new_n368), .C2(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(KEYINPUT7), .B1(new_n248), .B2(new_n213), .ZN(new_n375));
  AND2_X1   g0175(.A1(new_n353), .A2(new_n354), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n247), .B1(new_n376), .B2(G33), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n366), .A2(G20), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n375), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n351), .B1(new_n379), .B2(new_n203), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT16), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n374), .A2(new_n382), .A3(new_n275), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n271), .A2(new_n280), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n384), .B1(new_n286), .B2(new_n271), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(G200), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n355), .A2(KEYINPUT78), .ZN(new_n388));
  AND3_X1   g0188(.A1(new_n388), .A2(new_n246), .A3(new_n358), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n261), .A2(G1698), .ZN(new_n390));
  OAI211_X1 g0190(.A(new_n389), .B(new_n390), .C1(G223), .C2(G1698), .ZN(new_n391));
  NAND2_X1  g0191(.A1(G33), .A2(G87), .ZN(new_n392));
  XOR2_X1   g0192(.A(new_n392), .B(KEYINPUT82), .Z(new_n393));
  AOI21_X1  g0193(.A(new_n262), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n260), .B1(new_n299), .B2(new_n263), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n387), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  OR2_X1    g0196(.A1(new_n394), .A2(new_n395), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n396), .B1(new_n397), .B2(G190), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n383), .A2(new_n386), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(KEYINPUT83), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT83), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n383), .A2(new_n398), .A3(new_n401), .A4(new_n386), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n400), .A2(KEYINPUT17), .A3(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n351), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n370), .B1(new_n369), .B2(new_n372), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n360), .A2(new_n362), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n406), .A2(new_n367), .A3(KEYINPUT80), .A4(G68), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n404), .B1(new_n405), .B2(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n283), .B1(new_n408), .B2(KEYINPUT16), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n385), .B1(new_n409), .B2(new_n382), .ZN(new_n410));
  XNOR2_X1  g0210(.A(KEYINPUT84), .B(KEYINPUT17), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n410), .A2(new_n398), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n403), .A2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(G179), .ZN(new_n414));
  NOR3_X1   g0214(.A1(new_n394), .A2(new_n414), .A3(new_n395), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n415), .B1(G169), .B2(new_n397), .ZN(new_n416));
  OAI21_X1  g0216(.A(KEYINPUT18), .B1(new_n410), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n383), .A2(new_n386), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT18), .ZN(new_n419));
  INV_X1    g0219(.A(new_n416), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n418), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n417), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n413), .A2(new_n423), .ZN(new_n424));
  NOR3_X1   g0224(.A1(new_n296), .A2(new_n347), .A3(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(G41), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n257), .B(G45), .C1(new_n426), .C2(KEYINPUT5), .ZN(new_n427));
  AND2_X1   g0227(.A1(new_n426), .A2(KEYINPUT5), .ZN(new_n428));
  OR2_X1    g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  AND2_X1   g0229(.A1(new_n429), .A2(new_n262), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(G264), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n356), .A2(G257), .A3(G1698), .A4(new_n358), .ZN(new_n433));
  NAND2_X1  g0233(.A1(G33), .A2(G294), .ZN(new_n434));
  AND2_X1   g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(G250), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n436), .A2(G1698), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n388), .A2(new_n246), .A3(new_n358), .A4(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(KEYINPUT93), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT93), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n356), .A2(new_n440), .A3(new_n358), .A4(new_n437), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n435), .A2(new_n442), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n432), .B1(new_n443), .B2(new_n254), .ZN(new_n444));
  NOR3_X1   g0244(.A1(new_n429), .A2(new_n256), .A3(new_n254), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(KEYINPUT94), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n262), .B1(new_n435), .B2(new_n442), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT94), .ZN(new_n449));
  NOR4_X1   g0249(.A1(new_n448), .A2(new_n449), .A3(new_n445), .A4(new_n432), .ZN(new_n450));
  OAI21_X1  g0250(.A(G169), .B1(new_n447), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n433), .A2(new_n434), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n452), .B1(new_n441), .B2(new_n439), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n446), .B(new_n431), .C1(new_n453), .C2(new_n262), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n454), .A2(new_n414), .ZN(new_n455));
  INV_X1    g0255(.A(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n451), .A2(new_n456), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n282), .B(new_n283), .C1(G1), .C2(new_n274), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(G107), .ZN(new_n460));
  OAI21_X1  g0260(.A(KEYINPUT25), .B1(new_n282), .B2(G107), .ZN(new_n461));
  OR3_X1    g0261(.A1(new_n282), .A2(KEYINPUT25), .A3(G107), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n460), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n356), .A2(new_n213), .A3(G87), .A4(new_n358), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(KEYINPUT22), .ZN(new_n466));
  XNOR2_X1  g0266(.A(KEYINPUT90), .B(KEYINPUT22), .ZN(new_n467));
  INV_X1    g0267(.A(G87), .ZN(new_n468));
  NOR4_X1   g0268(.A1(new_n248), .A2(new_n467), .A3(G20), .A4(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n466), .A2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT24), .ZN(new_n472));
  NOR3_X1   g0272(.A1(new_n213), .A2(KEYINPUT23), .A3(G107), .ZN(new_n473));
  XNOR2_X1  g0273(.A(new_n473), .B(KEYINPUT91), .ZN(new_n474));
  OAI21_X1  g0274(.A(KEYINPUT23), .B1(new_n332), .B2(new_n213), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n213), .A2(G33), .A3(G116), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n474), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n471), .A2(new_n472), .A3(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n469), .B1(new_n465), .B2(KEYINPUT22), .ZN(new_n480));
  OAI21_X1  g0280(.A(KEYINPUT24), .B1(new_n480), .B2(new_n477), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  AOI21_X1  g0282(.A(KEYINPUT92), .B1(new_n482), .B2(new_n275), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT92), .ZN(new_n484));
  AOI211_X1 g0284(.A(new_n484), .B(new_n283), .C1(new_n479), .C2(new_n481), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n464), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n457), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n454), .A2(new_n449), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n443), .A2(new_n254), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n489), .A2(KEYINPUT94), .A3(new_n446), .A4(new_n431), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n488), .A2(new_n289), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n454), .A2(new_n387), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n472), .B1(new_n471), .B2(new_n478), .ZN(new_n494));
  NOR3_X1   g0294(.A1(new_n480), .A2(KEYINPUT24), .A3(new_n477), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n275), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(new_n484), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n482), .A2(KEYINPUT92), .A3(new_n275), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n463), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n493), .A2(new_n499), .ZN(new_n500));
  AND2_X1   g0300(.A1(new_n487), .A2(new_n500), .ZN(new_n501));
  NOR2_X1   g0301(.A1(G238), .A2(G1698), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n502), .B1(new_n334), .B2(G1698), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n356), .A2(new_n358), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(G33), .A2(G116), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n262), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n257), .A2(new_n256), .A3(G45), .ZN(new_n507));
  INV_X1    g0307(.A(G45), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n436), .B1(new_n508), .B2(G1), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n262), .A2(new_n507), .A3(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n506), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(G179), .ZN(new_n513));
  OAI21_X1  g0313(.A(G169), .B1(new_n506), .B2(new_n511), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n282), .A2(new_n339), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n356), .A2(new_n213), .A3(G68), .A4(new_n358), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT19), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n213), .B1(new_n302), .B2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(G97), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n468), .A2(new_n519), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n518), .B1(new_n332), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n213), .A2(G33), .A3(G97), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT87), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n522), .A2(new_n523), .A3(new_n517), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n522), .A2(new_n517), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(KEYINPUT87), .ZN(new_n526));
  AND3_X1   g0326(.A1(new_n521), .A2(new_n524), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n516), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n515), .B1(new_n528), .B2(new_n275), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n459), .A2(new_n339), .ZN(new_n530));
  AOI22_X1  g0330(.A1(new_n513), .A2(new_n514), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n283), .B1(new_n516), .B2(new_n527), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n458), .A2(new_n468), .ZN(new_n533));
  NOR3_X1   g0333(.A1(new_n532), .A2(new_n515), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n504), .A2(new_n505), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n254), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n387), .B1(new_n536), .B2(new_n510), .ZN(new_n537));
  NOR3_X1   g0337(.A1(new_n506), .A2(new_n289), .A3(new_n511), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n531), .B1(new_n534), .B2(new_n539), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n280), .A2(G97), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n541), .B1(G97), .B2(new_n458), .ZN(new_n542));
  XNOR2_X1  g0342(.A(new_n542), .B(KEYINPUT85), .ZN(new_n543));
  INV_X1    g0343(.A(G107), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n544), .A2(KEYINPUT6), .A3(G97), .ZN(new_n545));
  XOR2_X1   g0345(.A(G97), .B(G107), .Z(new_n546));
  OAI21_X1  g0346(.A(new_n545), .B1(new_n546), .B2(KEYINPUT6), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n547), .A2(G20), .B1(G77), .B2(new_n268), .ZN(new_n548));
  INV_X1    g0348(.A(new_n332), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n548), .B1(new_n379), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n275), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n543), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n430), .A2(G257), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(new_n446), .ZN(new_n554));
  INV_X1    g0354(.A(new_n554), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n334), .A2(G1698), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n556), .A2(KEYINPUT4), .B1(G250), .B2(G1698), .ZN(new_n557));
  OR2_X1    g0357(.A1(new_n248), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(G33), .A2(G283), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n356), .A2(new_n358), .A3(new_n556), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT4), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(KEYINPUT86), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT86), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n561), .A2(new_n565), .A3(new_n562), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n560), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n414), .B(new_n555), .C1(new_n567), .C2(new_n262), .ZN(new_n568));
  INV_X1    g0368(.A(new_n560), .ZN(new_n569));
  AND3_X1   g0369(.A1(new_n561), .A2(new_n565), .A3(new_n562), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n565), .B1(new_n561), .B2(new_n562), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n569), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n554), .B1(new_n572), .B2(new_n254), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n552), .B(new_n568), .C1(G169), .C2(new_n573), .ZN(new_n574));
  OAI211_X1 g0374(.A(G190), .B(new_n555), .C1(new_n567), .C2(new_n262), .ZN(new_n575));
  OR2_X1    g0375(.A1(new_n542), .A2(KEYINPUT85), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n542), .A2(KEYINPUT85), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n576), .A2(new_n577), .B1(new_n550), .B2(new_n275), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n575), .B(new_n578), .C1(new_n387), .C2(new_n573), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n540), .A2(new_n574), .A3(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n429), .A2(G270), .A3(new_n262), .ZN(new_n581));
  OR2_X1    g0381(.A1(new_n581), .A2(KEYINPUT88), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(KEYINPUT88), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n445), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(G264), .A2(G1698), .ZN(new_n585));
  INV_X1    g0385(.A(G303), .ZN(new_n586));
  OAI22_X1  g0386(.A1(new_n359), .A2(new_n585), .B1(new_n586), .B2(new_n249), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n389), .A2(KEYINPUT89), .A3(G257), .A4(new_n250), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n356), .A2(G257), .A3(new_n250), .A4(new_n358), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT89), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n587), .B1(new_n588), .B2(new_n591), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n584), .B1(new_n592), .B2(new_n262), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(G200), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n559), .B(new_n213), .C1(G33), .C2(new_n519), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n595), .B(new_n275), .C1(new_n213), .C2(G116), .ZN(new_n596));
  XNOR2_X1  g0396(.A(new_n596), .B(KEYINPUT20), .ZN(new_n597));
  INV_X1    g0397(.A(G116), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n597), .B1(new_n598), .B2(new_n280), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n459), .A2(G116), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(new_n601), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n594), .B(new_n602), .C1(new_n289), .C2(new_n593), .ZN(new_n603));
  INV_X1    g0403(.A(new_n603), .ZN(new_n604));
  XNOR2_X1  g0404(.A(new_n581), .B(KEYINPUT88), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(new_n446), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n588), .A2(new_n591), .ZN(new_n607));
  INV_X1    g0407(.A(new_n587), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n606), .B1(new_n609), .B2(new_n254), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n610), .A2(G179), .A3(new_n601), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT21), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n266), .B1(new_n599), .B2(new_n600), .ZN(new_n613));
  AND3_X1   g0413(.A1(new_n593), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n612), .B1(new_n593), .B2(new_n613), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n611), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NOR3_X1   g0416(.A1(new_n580), .A2(new_n604), .A3(new_n616), .ZN(new_n617));
  AND3_X1   g0417(.A1(new_n425), .A2(new_n501), .A3(new_n617), .ZN(G372));
  NOR2_X1   g0418(.A1(new_n308), .A2(new_n321), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n329), .B1(new_n619), .B2(new_n346), .ZN(new_n620));
  AND2_X1   g0420(.A1(new_n620), .A2(new_n413), .ZN(new_n621));
  OAI22_X1  g0421(.A1(new_n621), .A2(new_n422), .B1(new_n294), .B2(new_n295), .ZN(new_n622));
  AND2_X1   g0422(.A1(new_n622), .A2(new_n288), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT26), .ZN(new_n624));
  INV_X1    g0424(.A(new_n533), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n529), .A2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT95), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NOR4_X1   g0428(.A1(new_n532), .A2(new_n627), .A3(new_n533), .A4(new_n515), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n628), .A2(new_n630), .A3(new_n539), .ZN(new_n631));
  INV_X1    g0431(.A(new_n531), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n624), .B1(new_n633), .B2(new_n574), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT96), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n555), .B1(new_n567), .B2(new_n262), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n578), .B1(new_n266), .B2(new_n637), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n540), .A2(new_n638), .A3(KEYINPUT26), .A4(new_n568), .ZN(new_n639));
  OAI211_X1 g0439(.A(KEYINPUT96), .B(new_n624), .C1(new_n633), .C2(new_n574), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n636), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n616), .B1(new_n457), .B2(new_n486), .ZN(new_n642));
  AOI21_X1  g0442(.A(KEYINPUT95), .B1(new_n529), .B2(new_n625), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n643), .A2(new_n629), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n531), .B1(new_n644), .B2(new_n539), .ZN(new_n645));
  AND3_X1   g0445(.A1(new_n645), .A2(new_n574), .A3(new_n579), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n500), .A2(new_n646), .ZN(new_n647));
  OAI211_X1 g0447(.A(new_n641), .B(new_n632), .C1(new_n642), .C2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n425), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n623), .A2(new_n649), .ZN(G369));
  INV_X1    g0450(.A(G13), .ZN(new_n651));
  NOR3_X1   g0451(.A1(new_n651), .A2(G1), .A3(G20), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n653), .A2(KEYINPUT97), .A3(KEYINPUT27), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  AOI21_X1  g0455(.A(KEYINPUT97), .B1(new_n653), .B2(KEYINPUT27), .ZN(new_n656));
  OAI221_X1 g0456(.A(G213), .B1(KEYINPUT27), .B2(new_n653), .C1(new_n655), .C2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(G343), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n501), .B1(new_n499), .B2(new_n660), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n499), .B1(new_n451), .B2(new_n456), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(new_n659), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n616), .A2(new_n601), .A3(new_n659), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT98), .ZN(new_n667));
  OR2_X1    g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n616), .ZN(new_n669));
  OAI211_X1 g0469(.A(new_n669), .B(new_n603), .C1(new_n602), .C2(new_n660), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n666), .A2(new_n667), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n668), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(G330), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n665), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n669), .A2(new_n659), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n501), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n662), .A2(new_n660), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  OR2_X1    g0478(.A1(new_n674), .A2(new_n678), .ZN(G399));
  INV_X1    g0479(.A(new_n209), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n680), .A2(G41), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NOR3_X1   g0482(.A1(new_n332), .A2(G116), .A3(new_n520), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n682), .A2(G1), .A3(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n684), .B1(new_n216), .B2(new_n682), .ZN(new_n685));
  XNOR2_X1  g0485(.A(new_n685), .B(KEYINPUT28), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n617), .A2(new_n487), .A3(new_n500), .A4(new_n660), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n512), .A2(G179), .ZN(new_n688));
  AND2_X1   g0488(.A1(new_n593), .A2(new_n688), .ZN(new_n689));
  AND2_X1   g0489(.A1(new_n637), .A2(new_n454), .ZN(new_n690));
  INV_X1    g0490(.A(new_n513), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n610), .A2(new_n573), .A3(new_n444), .A4(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT30), .ZN(new_n693));
  AOI22_X1  g0493(.A1(new_n689), .A2(new_n690), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NOR3_X1   g0494(.A1(new_n513), .A2(new_n448), .A3(new_n432), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n695), .A2(KEYINPUT30), .A3(new_n610), .A4(new_n573), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n660), .B1(new_n694), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(KEYINPUT31), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n692), .A2(new_n693), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n637), .A2(new_n454), .A3(new_n593), .A4(new_n688), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n699), .A2(new_n696), .A3(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(new_n659), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT31), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n687), .A2(new_n698), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(G330), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n648), .A2(new_n660), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n708), .A2(KEYINPUT29), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT29), .ZN(new_n710));
  INV_X1    g0510(.A(new_n642), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n645), .A2(new_n574), .A3(new_n579), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n712), .B1(new_n499), .B2(new_n493), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n531), .B1(new_n711), .B2(new_n713), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n645), .A2(new_n568), .A3(new_n638), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(KEYINPUT26), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n540), .A2(new_n624), .A3(new_n638), .A4(new_n568), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n714), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n710), .B1(new_n718), .B2(new_n660), .ZN(new_n719));
  NOR3_X1   g0519(.A1(new_n707), .A2(new_n709), .A3(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n686), .B1(new_n720), .B2(G1), .ZN(G364));
  NOR2_X1   g0521(.A1(new_n651), .A2(G20), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n257), .B1(new_n722), .B2(G45), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n681), .A2(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n725), .B1(new_n672), .B2(G330), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n726), .B1(G330), .B2(new_n672), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n212), .B1(G20), .B2(new_n266), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n213), .A2(new_n414), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(G200), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(new_n289), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(G326), .ZN(new_n734));
  INV_X1    g0534(.A(G294), .ZN(new_n735));
  NOR3_X1   g0535(.A1(new_n289), .A2(G179), .A3(G200), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(new_n213), .ZN(new_n737));
  OAI22_X1  g0537(.A1(new_n733), .A2(new_n734), .B1(new_n735), .B2(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n731), .A2(G190), .ZN(new_n739));
  XNOR2_X1  g0539(.A(KEYINPUT33), .B(G317), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n738), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n213), .A2(G179), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n742), .A2(G190), .A3(G200), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n248), .B1(new_n743), .B2(new_n586), .ZN(new_n744));
  XOR2_X1   g0544(.A(new_n744), .B(KEYINPUT100), .Z(new_n745));
  NAND3_X1  g0545(.A1(new_n742), .A2(new_n289), .A3(G200), .ZN(new_n746));
  XOR2_X1   g0546(.A(new_n746), .B(KEYINPUT99), .Z(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(G283), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n730), .A2(G190), .A3(new_n387), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(G190), .A2(G200), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n742), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  AOI22_X1  g0553(.A1(new_n750), .A2(G322), .B1(new_n753), .B2(G329), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n730), .A2(new_n751), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(G311), .ZN(new_n757));
  AND2_X1   g0557(.A1(new_n754), .A2(new_n757), .ZN(new_n758));
  NAND4_X1  g0558(.A1(new_n741), .A2(new_n745), .A3(new_n748), .A4(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n739), .ZN(new_n760));
  OAI22_X1  g0560(.A1(new_n201), .A2(new_n733), .B1(new_n760), .B2(new_n203), .ZN(new_n761));
  OAI22_X1  g0561(.A1(new_n737), .A2(new_n519), .B1(new_n743), .B2(new_n468), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n747), .A2(G107), .ZN(new_n764));
  INV_X1    g0564(.A(G159), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n752), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g0566(.A(new_n766), .B(KEYINPUT32), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n249), .B1(new_n749), .B2(new_n202), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n768), .B1(G77), .B2(new_n756), .ZN(new_n769));
  NAND4_X1  g0569(.A1(new_n763), .A2(new_n764), .A3(new_n767), .A4(new_n769), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n729), .B1(new_n759), .B2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n725), .ZN(new_n772));
  NOR2_X1   g0572(.A1(G13), .A2(G33), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(G20), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(new_n728), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n389), .A2(new_n680), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n217), .A2(new_n508), .ZN(new_n779));
  OAI211_X1 g0579(.A(new_n778), .B(new_n779), .C1(new_n508), .C2(new_n239), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n248), .A2(new_n680), .ZN(new_n781));
  AOI22_X1  g0581(.A1(new_n781), .A2(G355), .B1(new_n598), .B2(new_n680), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n777), .B1(new_n780), .B2(new_n782), .ZN(new_n783));
  NOR3_X1   g0583(.A1(new_n771), .A2(new_n772), .A3(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n775), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n784), .B1(new_n672), .B2(new_n785), .ZN(new_n786));
  AND2_X1   g0586(.A1(new_n727), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(G396));
  NOR2_X1   g0588(.A1(new_n728), .A2(new_n773), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n772), .B1(new_n314), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n346), .A2(new_n659), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n343), .A2(new_n659), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n344), .A2(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n791), .B1(new_n793), .B2(new_n346), .ZN(new_n794));
  INV_X1    g0594(.A(G311), .ZN(new_n795));
  OAI22_X1  g0595(.A1(new_n749), .A2(new_n735), .B1(new_n752), .B2(new_n795), .ZN(new_n796));
  AOI211_X1 g0596(.A(new_n249), .B(new_n796), .C1(G116), .C2(new_n756), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n747), .A2(G87), .ZN(new_n798));
  INV_X1    g0598(.A(new_n737), .ZN(new_n799));
  INV_X1    g0599(.A(new_n743), .ZN(new_n800));
  AOI22_X1  g0600(.A1(new_n799), .A2(G97), .B1(new_n800), .B2(G107), .ZN(new_n801));
  AOI22_X1  g0601(.A1(G283), .A2(new_n739), .B1(new_n732), .B2(G303), .ZN(new_n802));
  NAND4_X1  g0602(.A1(new_n797), .A2(new_n798), .A3(new_n801), .A4(new_n802), .ZN(new_n803));
  AOI22_X1  g0603(.A1(G137), .A2(new_n732), .B1(new_n739), .B2(G150), .ZN(new_n804));
  XOR2_X1   g0604(.A(new_n804), .B(KEYINPUT101), .Z(new_n805));
  INV_X1    g0605(.A(G143), .ZN(new_n806));
  OAI221_X1 g0606(.A(new_n805), .B1(new_n806), .B2(new_n749), .C1(new_n765), .C2(new_n755), .ZN(new_n807));
  XOR2_X1   g0607(.A(new_n807), .B(KEYINPUT34), .Z(new_n808));
  INV_X1    g0608(.A(new_n747), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n809), .A2(new_n203), .ZN(new_n810));
  AOI22_X1  g0610(.A1(new_n799), .A2(G58), .B1(G132), .B2(new_n753), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n811), .B1(new_n201), .B2(new_n743), .ZN(new_n812));
  OR3_X1    g0612(.A1(new_n810), .A2(new_n812), .A3(new_n359), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n803), .B1(new_n808), .B2(new_n813), .ZN(new_n814));
  XOR2_X1   g0614(.A(new_n814), .B(KEYINPUT102), .Z(new_n815));
  OAI221_X1 g0615(.A(new_n790), .B1(new_n774), .B2(new_n794), .C1(new_n815), .C2(new_n729), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n632), .B1(new_n647), .B2(new_n642), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n640), .A2(new_n639), .ZN(new_n818));
  AOI21_X1  g0618(.A(KEYINPUT96), .B1(new_n715), .B2(new_n624), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  OAI211_X1 g0620(.A(new_n660), .B(new_n794), .C1(new_n817), .C2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(KEYINPUT103), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND4_X1  g0623(.A1(new_n648), .A2(KEYINPUT103), .A3(new_n660), .A4(new_n794), .ZN(new_n824));
  INV_X1    g0624(.A(new_n794), .ZN(new_n825));
  AOI22_X1  g0625(.A1(new_n823), .A2(new_n824), .B1(new_n708), .B2(new_n825), .ZN(new_n826));
  AND2_X1   g0626(.A1(new_n826), .A2(new_n707), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n772), .B1(new_n826), .B2(new_n707), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n816), .B1(new_n827), .B2(new_n828), .ZN(G384));
  AND2_X1   g0629(.A1(new_n547), .A2(KEYINPUT35), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n547), .A2(KEYINPUT35), .ZN(new_n831));
  NOR4_X1   g0631(.A1(new_n830), .A2(new_n831), .A3(new_n598), .A4(new_n215), .ZN(new_n832));
  XNOR2_X1  g0632(.A(new_n832), .B(KEYINPUT36), .ZN(new_n833));
  INV_X1    g0633(.A(new_n216), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n349), .A2(G77), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n201), .A2(G68), .ZN(new_n836));
  AOI211_X1 g0636(.A(new_n257), .B(G13), .C1(new_n835), .C2(new_n836), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n833), .A2(new_n837), .ZN(new_n838));
  XOR2_X1   g0638(.A(KEYINPUT105), .B(KEYINPUT38), .Z(new_n839));
  INV_X1    g0639(.A(new_n657), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n418), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n841), .B1(new_n413), .B2(new_n423), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n418), .A2(new_n420), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT37), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n843), .A2(new_n841), .A3(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n400), .A2(new_n402), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n843), .A2(new_n841), .A3(new_n399), .ZN(new_n849));
  AOI22_X1  g0649(.A1(new_n846), .A2(new_n848), .B1(KEYINPUT37), .B2(new_n849), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n839), .B1(new_n842), .B2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT39), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n845), .A2(new_n847), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n374), .A2(new_n275), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n408), .A2(KEYINPUT16), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n386), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n416), .A2(new_n657), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n400), .A2(new_n858), .A3(new_n402), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n859), .A2(KEYINPUT37), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT104), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n859), .A2(KEYINPUT104), .A3(KEYINPUT37), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n853), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n422), .B1(new_n403), .B2(new_n412), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n856), .A2(new_n840), .ZN(new_n866));
  OAI21_X1  g0666(.A(KEYINPUT38), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  OAI211_X1 g0667(.A(new_n851), .B(new_n852), .C1(new_n864), .C2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(KEYINPUT106), .ZN(new_n869));
  AND3_X1   g0669(.A1(new_n859), .A2(KEYINPUT104), .A3(KEYINPUT37), .ZN(new_n870));
  AOI21_X1  g0670(.A(KEYINPUT104), .B1(new_n859), .B2(KEYINPUT37), .ZN(new_n871));
  OAI22_X1  g0671(.A1(new_n870), .A2(new_n871), .B1(new_n847), .B2(new_n845), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n424), .A2(new_n840), .A3(new_n856), .ZN(new_n873));
  AOI21_X1  g0673(.A(KEYINPUT38), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n864), .A2(new_n867), .ZN(new_n875));
  OAI21_X1  g0675(.A(KEYINPUT39), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n872), .A2(KEYINPUT38), .A3(new_n873), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT106), .ZN(new_n878));
  NAND4_X1  g0678(.A1(new_n877), .A2(new_n878), .A3(new_n852), .A4(new_n851), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n869), .A2(new_n876), .A3(new_n879), .ZN(new_n880));
  OR2_X1    g0680(.A1(new_n327), .A2(new_n328), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n881), .A2(new_n323), .A3(new_n660), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n791), .B1(new_n823), .B2(new_n824), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n323), .B(new_n659), .C1(new_n881), .C2(new_n619), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n323), .A2(new_n659), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n322), .A2(new_n329), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n885), .A2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT38), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n865), .A2(new_n866), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n892), .B1(new_n864), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n877), .ZN(new_n895));
  AOI22_X1  g0695(.A1(new_n891), .A2(new_n895), .B1(new_n422), .B2(new_n657), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n884), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n425), .B1(new_n709), .B2(new_n719), .ZN(new_n898));
  AND2_X1   g0698(.A1(new_n623), .A2(new_n898), .ZN(new_n899));
  XOR2_X1   g0699(.A(new_n897), .B(new_n899), .Z(new_n900));
  NAND2_X1  g0700(.A1(new_n687), .A2(new_n698), .ZN(new_n901));
  AOI21_X1  g0701(.A(KEYINPUT31), .B1(new_n702), .B2(KEYINPUT107), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT107), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n697), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(KEYINPUT108), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT108), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n902), .A2(new_n907), .A3(new_n904), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n901), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n889), .A2(new_n794), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n877), .A2(new_n851), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n911), .A2(new_n912), .A3(KEYINPUT40), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(KEYINPUT40), .B1(new_n895), .B2(new_n911), .ZN(new_n915));
  AND2_X1   g0715(.A1(new_n687), .A2(new_n698), .ZN(new_n916));
  AND3_X1   g0716(.A1(new_n902), .A2(new_n907), .A3(new_n904), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n907), .B1(new_n902), .B2(new_n904), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n916), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n425), .A2(new_n919), .ZN(new_n920));
  OR3_X1    g0720(.A1(new_n914), .A2(new_n915), .A3(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n920), .B1(new_n914), .B2(new_n915), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n921), .A2(G330), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n900), .A2(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n924), .B1(new_n257), .B2(new_n722), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n900), .A2(new_n923), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n838), .B1(new_n925), .B2(new_n926), .ZN(G367));
  OAI211_X1 g0727(.A(new_n574), .B(new_n579), .C1(new_n578), .C2(new_n660), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n638), .A2(new_n568), .A3(new_n659), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n501), .A2(new_n675), .A3(new_n930), .ZN(new_n931));
  OR2_X1    g0731(.A1(new_n931), .A2(KEYINPUT42), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n574), .B1(new_n487), .B2(new_n928), .ZN(new_n933));
  AOI22_X1  g0733(.A1(new_n931), .A2(KEYINPUT42), .B1(new_n660), .B2(new_n933), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n644), .A2(new_n660), .ZN(new_n935));
  MUX2_X1   g0735(.A(new_n645), .B(new_n531), .S(new_n935), .Z(new_n936));
  AOI22_X1  g0736(.A1(new_n932), .A2(new_n934), .B1(KEYINPUT43), .B2(new_n936), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n936), .A2(KEYINPUT43), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n937), .B(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n674), .A2(new_n930), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n939), .B(new_n940), .ZN(new_n941));
  XOR2_X1   g0741(.A(new_n681), .B(KEYINPUT41), .Z(new_n942));
  INV_X1    g0742(.A(new_n930), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT109), .ZN(new_n944));
  OAI211_X1 g0744(.A(new_n678), .B(new_n943), .C1(new_n944), .C2(KEYINPUT44), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT110), .ZN(new_n946));
  AND2_X1   g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n945), .A2(new_n946), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n944), .A2(KEYINPUT44), .ZN(new_n949));
  OR3_X1    g0749(.A1(new_n947), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n949), .B1(new_n947), .B2(new_n948), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n678), .A2(new_n943), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n952), .B(KEYINPUT45), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n950), .A2(new_n951), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(new_n674), .ZN(new_n955));
  INV_X1    g0755(.A(new_n720), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n676), .B1(new_n664), .B2(new_n675), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n957), .B(new_n673), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT111), .ZN(new_n959));
  OR3_X1    g0759(.A1(new_n956), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n959), .B1(new_n956), .B2(new_n958), .ZN(new_n961));
  INV_X1    g0761(.A(new_n674), .ZN(new_n962));
  NAND4_X1  g0762(.A1(new_n950), .A2(new_n962), .A3(new_n951), .A4(new_n953), .ZN(new_n963));
  NAND4_X1  g0763(.A1(new_n955), .A2(new_n960), .A3(new_n961), .A4(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n942), .B1(new_n964), .B2(new_n720), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n941), .B1(new_n965), .B2(new_n724), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n776), .B1(new_n209), .B2(new_n340), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n967), .B1(new_n778), .B2(new_n235), .ZN(new_n968));
  OAI22_X1  g0768(.A1(new_n806), .A2(new_n733), .B1(new_n760), .B2(new_n765), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n969), .B1(G68), .B2(new_n799), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n248), .B1(new_n753), .B2(G137), .ZN(new_n971));
  AOI22_X1  g0771(.A1(new_n750), .A2(G150), .B1(new_n756), .B2(G50), .ZN(new_n972));
  INV_X1    g0772(.A(new_n746), .ZN(new_n973));
  AOI22_X1  g0773(.A1(new_n800), .A2(G58), .B1(new_n973), .B2(G77), .ZN(new_n974));
  NAND4_X1  g0774(.A1(new_n970), .A2(new_n971), .A3(new_n972), .A4(new_n974), .ZN(new_n975));
  AOI22_X1  g0775(.A1(new_n750), .A2(G303), .B1(new_n753), .B2(G317), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT46), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n977), .B1(new_n743), .B2(new_n598), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n800), .A2(KEYINPUT46), .A3(G116), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n756), .A2(G283), .ZN(new_n980));
  NAND4_X1  g0780(.A1(new_n976), .A2(new_n978), .A3(new_n979), .A4(new_n980), .ZN(new_n981));
  AOI22_X1  g0781(.A1(new_n332), .A2(new_n799), .B1(new_n739), .B2(G294), .ZN(new_n982));
  AOI22_X1  g0782(.A1(new_n732), .A2(G311), .B1(new_n973), .B2(G97), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n982), .A2(new_n359), .A3(new_n983), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n975), .B1(new_n981), .B2(new_n984), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n985), .B(KEYINPUT47), .ZN(new_n986));
  AOI211_X1 g0786(.A(new_n772), .B(new_n968), .C1(new_n986), .C2(new_n728), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n987), .B1(new_n936), .B2(new_n785), .ZN(new_n988));
  XOR2_X1   g0788(.A(new_n988), .B(KEYINPUT112), .Z(new_n989));
  NAND2_X1  g0789(.A1(new_n966), .A2(new_n989), .ZN(G387));
  NOR2_X1   g0790(.A1(new_n958), .A2(new_n723), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT113), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n665), .A2(new_n775), .ZN(new_n993));
  INV_X1    g0793(.A(new_n781), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n994), .A2(new_n683), .B1(G107), .B2(new_n209), .ZN(new_n995));
  INV_X1    g0795(.A(new_n778), .ZN(new_n996));
  INV_X1    g0796(.A(new_n683), .ZN(new_n997));
  AOI211_X1 g0797(.A(G45), .B(new_n997), .C1(G68), .C2(G77), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n270), .A2(G50), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(KEYINPUT50), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n996), .B1(new_n998), .B2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n232), .A2(G45), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n995), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n725), .B1(new_n1003), .B2(new_n777), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(G68), .A2(new_n756), .B1(new_n753), .B2(G150), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(new_n201), .B2(new_n749), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n271), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1006), .B1(new_n1007), .B2(new_n739), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n743), .A2(new_n314), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n340), .A2(new_n737), .ZN(new_n1010));
  AOI211_X1 g0810(.A(new_n1009), .B(new_n1010), .C1(G159), .C2(new_n732), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n359), .B1(new_n747), .B2(G97), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1008), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(G311), .A2(new_n739), .B1(new_n732), .B2(G322), .ZN(new_n1014));
  OR2_X1    g0814(.A1(new_n1014), .A2(KEYINPUT114), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1014), .A2(KEYINPUT114), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n750), .A2(G317), .B1(new_n756), .B2(G303), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1015), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT48), .ZN(new_n1019));
  OR2_X1    g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g0820(.A(G283), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n737), .A2(new_n1021), .B1(new_n743), .B2(new_n735), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1022), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1020), .A2(KEYINPUT49), .A3(new_n1023), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n746), .A2(new_n598), .B1(new_n752), .B2(new_n734), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n1025), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1024), .A2(new_n359), .A3(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(KEYINPUT49), .B1(new_n1020), .B2(new_n1023), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1013), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1004), .B1(new_n1029), .B2(new_n728), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n992), .B1(new_n993), .B2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n960), .A2(new_n961), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n682), .B1(new_n956), .B2(new_n958), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1031), .A2(new_n1034), .ZN(G393));
  NAND3_X1  g0835(.A1(new_n955), .A2(new_n724), .A3(new_n963), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n776), .B1(new_n519), .B2(new_n209), .C1(new_n996), .C2(new_n242), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1037), .A2(new_n725), .ZN(new_n1038));
  INV_X1    g0838(.A(G150), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n733), .A2(new_n1039), .B1(new_n765), .B2(new_n749), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT51), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n755), .A2(new_n270), .B1(new_n752), .B2(new_n806), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n737), .A2(new_n314), .B1(new_n743), .B2(new_n203), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n1042), .B(new_n1043), .C1(G50), .C2(new_n739), .ZN(new_n1044));
  NAND4_X1  g0844(.A1(new_n1041), .A2(new_n389), .A3(new_n798), .A4(new_n1044), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(G317), .A2(new_n732), .B1(new_n750), .B2(G311), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1046), .B(KEYINPUT115), .ZN(new_n1047));
  XOR2_X1   g0847(.A(new_n1047), .B(KEYINPUT52), .Z(new_n1048));
  OAI21_X1  g0848(.A(new_n248), .B1(new_n755), .B2(new_n735), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1049), .B1(G322), .B2(new_n753), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n800), .A2(G283), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(G116), .A2(new_n799), .B1(new_n739), .B2(G303), .ZN(new_n1052));
  NAND4_X1  g0852(.A1(new_n764), .A2(new_n1050), .A3(new_n1051), .A4(new_n1052), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1045), .B1(new_n1048), .B2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1038), .B1(new_n1054), .B2(new_n728), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1055), .B1(new_n930), .B2(new_n785), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n964), .A2(new_n681), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n955), .A2(new_n963), .B1(new_n961), .B2(new_n960), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1036), .B(new_n1056), .C1(new_n1057), .C2(new_n1058), .ZN(G390));
  AOI21_X1  g0859(.A(new_n825), .B1(new_n886), .B2(new_n888), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n919), .A2(G330), .A3(new_n1060), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n882), .B1(new_n885), .B2(new_n890), .ZN(new_n1062));
  NAND4_X1  g0862(.A1(new_n1062), .A2(new_n879), .A3(new_n876), .A4(new_n869), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n793), .A2(new_n346), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n718), .A2(new_n660), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n791), .ZN(new_n1066));
  AND2_X1   g0866(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n912), .B(new_n882), .C1(new_n1067), .C2(new_n890), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1061), .B1(new_n1063), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n1069), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n425), .A2(new_n919), .A3(G330), .ZN(new_n1071));
  AND3_X1   g0871(.A1(new_n623), .A2(new_n898), .A3(new_n1071), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n890), .B1(new_n706), .B2(new_n825), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n885), .B1(new_n1073), .B2(new_n1061), .ZN(new_n1074));
  NAND4_X1  g0874(.A1(new_n889), .A2(G330), .A3(new_n705), .A4(new_n794), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1075), .A2(new_n1066), .A3(new_n1065), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n919), .A2(G330), .A3(new_n794), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1076), .B1(new_n890), .B2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1072), .B1(new_n1074), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1079), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1063), .A2(new_n1068), .A3(new_n1075), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1070), .A2(new_n1080), .A3(new_n1081), .ZN(new_n1082));
  AND3_X1   g0882(.A1(new_n1063), .A2(new_n1068), .A3(new_n1075), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1079), .B1(new_n1083), .B2(new_n1069), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1082), .A2(new_n1084), .A3(new_n681), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n1083), .A2(new_n1069), .ZN(new_n1086));
  OR2_X1    g0886(.A1(new_n880), .A2(new_n774), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n789), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n725), .B1(new_n1007), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(G132), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(KEYINPUT54), .B(G143), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n749), .A2(new_n1090), .B1(new_n755), .B2(new_n1091), .ZN(new_n1092));
  AOI211_X1 g0892(.A(new_n248), .B(new_n1092), .C1(G125), .C2(new_n753), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n743), .A2(new_n1039), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(new_n1094), .B(KEYINPUT53), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n732), .A2(G128), .B1(new_n973), .B2(G50), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(G159), .A2(new_n799), .B1(new_n739), .B2(G137), .ZN(new_n1097));
  NAND4_X1  g0897(.A1(new_n1093), .A2(new_n1095), .A3(new_n1096), .A4(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n810), .B1(G294), .B2(new_n753), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(new_n1099), .B(KEYINPUT116), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n549), .A2(new_n760), .B1(new_n733), .B2(new_n1021), .ZN(new_n1101));
  OAI221_X1 g0901(.A(new_n248), .B1(new_n755), .B2(new_n519), .C1(new_n598), .C2(new_n749), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n737), .A2(new_n314), .B1(new_n743), .B2(new_n468), .ZN(new_n1103));
  OR3_X1    g0903(.A1(new_n1101), .A2(new_n1102), .A3(new_n1103), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1098), .B1(new_n1100), .B2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1089), .B1(new_n1105), .B2(new_n728), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n1086), .A2(new_n724), .B1(new_n1087), .B2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1085), .A2(new_n1107), .ZN(G378));
  XNOR2_X1  g0908(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1109));
  XOR2_X1   g0909(.A(new_n296), .B(new_n1109), .Z(new_n1110));
  NAND2_X1  g0910(.A1(new_n287), .A2(new_n840), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(new_n1110), .B(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(KEYINPUT118), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n919), .A2(new_n1060), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1114), .B1(new_n877), .B2(new_n894), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n913), .B(G330), .C1(new_n1115), .C2(KEYINPUT40), .ZN(new_n1116));
  AND3_X1   g0916(.A1(new_n884), .A2(new_n1116), .A3(new_n896), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1116), .B1(new_n884), .B2(new_n896), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1113), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1116), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n897), .A2(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1113), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n884), .A2(new_n1116), .A3(new_n896), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1121), .A2(new_n1122), .A3(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1119), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1112), .A2(new_n773), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n725), .B1(new_n1088), .B2(G50), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n389), .A2(G41), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n746), .A2(new_n202), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1009), .B1(G283), .B2(new_n753), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1128), .A2(new_n1130), .A3(new_n1131), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(new_n1132), .B(KEYINPUT117), .ZN(new_n1133));
  OAI22_X1  g0933(.A1(new_n340), .A2(new_n755), .B1(new_n544), .B2(new_n749), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1134), .B1(G68), .B2(new_n799), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(G97), .A2(new_n739), .B1(new_n732), .B2(G116), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1133), .A2(new_n1135), .A3(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(KEYINPUT58), .ZN(new_n1138));
  OR2_X1    g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(G33), .A2(G41), .ZN(new_n1141));
  NOR3_X1   g0941(.A1(new_n1128), .A2(G50), .A3(new_n1141), .ZN(new_n1142));
  AOI22_X1  g0942(.A1(G150), .A2(new_n799), .B1(new_n732), .B2(G125), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n739), .A2(G132), .ZN(new_n1144));
  AND2_X1   g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(new_n750), .A2(G128), .B1(new_n756), .B2(G137), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n1145), .B(new_n1146), .C1(new_n743), .C2(new_n1091), .ZN(new_n1147));
  OR2_X1    g0947(.A1(new_n1147), .A2(KEYINPUT59), .ZN(new_n1148));
  INV_X1    g0948(.A(G124), .ZN(new_n1149));
  OAI221_X1 g0949(.A(new_n1141), .B1(new_n752), .B2(new_n1149), .C1(new_n765), .C2(new_n746), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1150), .B1(new_n1147), .B2(KEYINPUT59), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1142), .B1(new_n1148), .B2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1139), .A2(new_n1140), .A3(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1127), .B1(new_n1153), .B2(new_n728), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n1125), .A2(new_n724), .B1(new_n1126), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT119), .ZN(new_n1157));
  NOR3_X1   g0957(.A1(new_n1083), .A2(new_n1069), .A3(new_n1079), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1072), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1157), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1082), .A2(KEYINPUT119), .A3(new_n1072), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1160), .A2(new_n1125), .A3(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(KEYINPUT57), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n682), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  NAND4_X1  g0964(.A1(new_n1160), .A2(new_n1125), .A3(new_n1161), .A4(KEYINPUT57), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1156), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1166), .ZN(G375));
  OAI21_X1  g0967(.A(new_n724), .B1(new_n1078), .B2(new_n1074), .ZN(new_n1168));
  INV_X1    g0968(.A(KEYINPUT120), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n890), .A2(new_n773), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n725), .B1(new_n1088), .B2(G68), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n598), .A2(new_n760), .B1(new_n733), .B2(new_n735), .ZN(new_n1172));
  AOI211_X1 g0972(.A(new_n1010), .B(new_n1172), .C1(G97), .C2(new_n800), .ZN(new_n1173));
  OAI22_X1  g0973(.A1(new_n549), .A2(new_n755), .B1(new_n749), .B2(new_n1021), .ZN(new_n1174));
  AOI211_X1 g0974(.A(new_n249), .B(new_n1174), .C1(G303), .C2(new_n753), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n1173), .B(new_n1175), .C1(new_n314), .C2(new_n809), .ZN(new_n1176));
  OAI22_X1  g0976(.A1(new_n737), .A2(new_n201), .B1(new_n755), .B2(new_n1039), .ZN(new_n1177));
  XOR2_X1   g0977(.A(new_n1177), .B(KEYINPUT121), .Z(new_n1178));
  OAI22_X1  g0978(.A1(new_n1090), .A2(new_n733), .B1(new_n760), .B2(new_n1091), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1179), .B1(G159), .B2(new_n800), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(new_n750), .A2(G137), .B1(new_n753), .B2(G128), .ZN(new_n1181));
  NAND4_X1  g0981(.A1(new_n1180), .A2(new_n389), .A3(new_n1130), .A4(new_n1181), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1176), .B1(new_n1178), .B2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1171), .B1(new_n1183), .B2(new_n728), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(new_n1168), .A2(new_n1169), .B1(new_n1170), .B2(new_n1184), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1185), .B1(new_n1169), .B2(new_n1168), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n1080), .A2(new_n942), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n1078), .A2(new_n1074), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1159), .A2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1188), .A2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1187), .A2(new_n1191), .ZN(G381));
  NAND3_X1  g0992(.A1(new_n1031), .A2(new_n787), .A3(new_n1034), .ZN(new_n1193));
  OR3_X1    g0993(.A1(G390), .A2(G384), .A3(new_n1193), .ZN(new_n1194));
  NOR3_X1   g0994(.A1(new_n1194), .A2(G387), .A3(G381), .ZN(new_n1195));
  AND3_X1   g0995(.A1(new_n1085), .A2(new_n1107), .A3(KEYINPUT122), .ZN(new_n1196));
  AOI21_X1  g0996(.A(KEYINPUT122), .B1(new_n1085), .B2(new_n1107), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1195), .A2(new_n1166), .A3(new_n1198), .ZN(G407));
  INV_X1    g0999(.A(G213), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n1200), .A2(G343), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1166), .A2(new_n1198), .A3(new_n1201), .ZN(new_n1202));
  XOR2_X1   g1002(.A(new_n1202), .B(KEYINPUT123), .Z(new_n1203));
  NAND3_X1  g1003(.A1(new_n1203), .A2(G213), .A3(G407), .ZN(G409));
  AOI21_X1  g1004(.A(G390), .B1(new_n966), .B2(new_n989), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n966), .A2(new_n989), .A3(G390), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(G393), .A2(G396), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1209), .A2(new_n1193), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1210), .B1(new_n1205), .B2(KEYINPUT125), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1208), .A2(new_n1211), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1206), .A2(new_n1210), .A3(KEYINPUT125), .A4(new_n1207), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT60), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1190), .A2(new_n1216), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1159), .A2(new_n1189), .A3(KEYINPUT60), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1217), .A2(new_n681), .A3(new_n1079), .A4(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1187), .A2(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(KEYINPUT124), .ZN(new_n1221));
  XNOR2_X1  g1021(.A(G384), .B(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1220), .A2(new_n1222), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n1187), .B(new_n1219), .C1(new_n1221), .C2(G384), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1201), .A2(G2897), .ZN(new_n1226));
  XNOR2_X1  g1026(.A(new_n1225), .B(new_n1226), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1155), .B1(new_n1162), .B2(new_n942), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(new_n1166), .A2(G378), .B1(new_n1198), .B2(new_n1228), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1227), .B1(new_n1229), .B2(new_n1201), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1231), .A2(new_n681), .A3(new_n1165), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1232), .A2(G378), .A3(new_n1155), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1198), .A2(new_n1228), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT62), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1201), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1225), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1235), .A2(new_n1236), .A3(new_n1237), .A4(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT61), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1230), .A2(new_n1239), .A3(new_n1240), .ZN(new_n1241));
  XNOR2_X1  g1041(.A(KEYINPUT126), .B(KEYINPUT62), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1201), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1242), .B1(new_n1243), .B2(new_n1238), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1215), .B1(new_n1241), .B2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT63), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1235), .A2(new_n1237), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1246), .B1(new_n1247), .B2(new_n1225), .ZN(new_n1248));
  AOI21_X1  g1048(.A(KEYINPUT61), .B1(new_n1247), .B2(new_n1227), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1243), .A2(KEYINPUT63), .A3(new_n1238), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1248), .A2(new_n1249), .A3(new_n1214), .A4(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1245), .A2(new_n1251), .ZN(G405));
  NAND2_X1  g1052(.A1(new_n1214), .A2(new_n1238), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1212), .A2(new_n1213), .A3(new_n1225), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(G375), .A2(new_n1198), .ZN(new_n1256));
  AND2_X1   g1056(.A1(new_n1256), .A2(new_n1233), .ZN(new_n1257));
  XNOR2_X1  g1057(.A(new_n1255), .B(new_n1257), .ZN(G402));
endmodule


