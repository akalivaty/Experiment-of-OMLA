

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581;

  AND2_X1 U320 ( .A1(n563), .A2(n387), .ZN(n359) );
  XOR2_X1 U321 ( .A(n421), .B(n428), .Z(n288) );
  XOR2_X1 U322 ( .A(G197GAT), .B(KEYINPUT21), .Z(n289) );
  XOR2_X1 U323 ( .A(G43GAT), .B(G50GAT), .Z(n290) );
  INV_X1 U324 ( .A(KEYINPUT99), .ZN(n358) );
  NOR2_X1 U325 ( .A1(n570), .A2(n507), .ZN(n508) );
  XNOR2_X1 U326 ( .A(n341), .B(n383), .ZN(n342) );
  XNOR2_X1 U327 ( .A(n343), .B(n342), .ZN(n344) );
  NOR2_X1 U328 ( .A1(n543), .A2(n542), .ZN(n564) );
  OR2_X1 U329 ( .A1(n544), .A2(n547), .ZN(n346) );
  XNOR2_X1 U330 ( .A(KEYINPUT37), .B(n411), .ZN(n487) );
  XNOR2_X1 U331 ( .A(n409), .B(n408), .ZN(n523) );
  XOR2_X1 U332 ( .A(KEYINPUT96), .B(n386), .Z(n543) );
  XNOR2_X1 U333 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n448) );
  XNOR2_X1 U334 ( .A(n449), .B(n448), .ZN(G1330GAT) );
  XOR2_X1 U335 ( .A(KEYINPUT17), .B(KEYINPUT19), .Z(n292) );
  XNOR2_X1 U336 ( .A(G183GAT), .B(KEYINPUT18), .ZN(n291) );
  XNOR2_X1 U337 ( .A(n292), .B(n291), .ZN(n355) );
  XOR2_X1 U338 ( .A(n355), .B(G71GAT), .Z(n294) );
  NAND2_X1 U339 ( .A1(G227GAT), .A2(G233GAT), .ZN(n293) );
  XNOR2_X1 U340 ( .A(n294), .B(n293), .ZN(n309) );
  XOR2_X1 U341 ( .A(G190GAT), .B(G43GAT), .Z(n296) );
  XNOR2_X1 U342 ( .A(G134GAT), .B(G99GAT), .ZN(n295) );
  XNOR2_X1 U343 ( .A(n296), .B(n295), .ZN(n300) );
  XOR2_X1 U344 ( .A(G169GAT), .B(G176GAT), .Z(n298) );
  XNOR2_X1 U345 ( .A(G127GAT), .B(KEYINPUT86), .ZN(n297) );
  XNOR2_X1 U346 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U347 ( .A(n300), .B(n299), .Z(n307) );
  XOR2_X1 U348 ( .A(G113GAT), .B(KEYINPUT85), .Z(n302) );
  XNOR2_X1 U349 ( .A(KEYINPUT0), .B(KEYINPUT84), .ZN(n301) );
  XNOR2_X1 U350 ( .A(n302), .B(n301), .ZN(n366) );
  XOR2_X1 U351 ( .A(KEYINPUT20), .B(KEYINPUT87), .Z(n304) );
  XNOR2_X1 U352 ( .A(G120GAT), .B(G15GAT), .ZN(n303) );
  XNOR2_X1 U353 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U354 ( .A(n366), .B(n305), .ZN(n306) );
  XNOR2_X1 U355 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U356 ( .A(n309), .B(n308), .Z(n515) );
  INV_X1 U357 ( .A(n515), .ZN(n547) );
  XOR2_X1 U358 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n446) );
  XOR2_X1 U359 ( .A(G64GAT), .B(G78GAT), .Z(n311) );
  XNOR2_X1 U360 ( .A(G57GAT), .B(G211GAT), .ZN(n310) );
  XNOR2_X1 U361 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U362 ( .A(n312), .B(G183GAT), .Z(n314) );
  XOR2_X1 U363 ( .A(G15GAT), .B(G22GAT), .Z(n412) );
  XNOR2_X1 U364 ( .A(G155GAT), .B(n412), .ZN(n313) );
  XNOR2_X1 U365 ( .A(n314), .B(n313), .ZN(n327) );
  XOR2_X1 U366 ( .A(G71GAT), .B(KEYINPUT13), .Z(n429) );
  XOR2_X1 U367 ( .A(KEYINPUT14), .B(n429), .Z(n316) );
  NAND2_X1 U368 ( .A1(G231GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U369 ( .A(n316), .B(n315), .ZN(n320) );
  XOR2_X1 U370 ( .A(KEYINPUT15), .B(KEYINPUT77), .Z(n318) );
  XNOR2_X1 U371 ( .A(KEYINPUT81), .B(KEYINPUT12), .ZN(n317) );
  XNOR2_X1 U372 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U373 ( .A(n320), .B(n319), .Z(n325) );
  XOR2_X1 U374 ( .A(G127GAT), .B(G1GAT), .Z(n375) );
  XOR2_X1 U375 ( .A(KEYINPUT78), .B(KEYINPUT79), .Z(n322) );
  XNOR2_X1 U376 ( .A(G8GAT), .B(KEYINPUT80), .ZN(n321) );
  XNOR2_X1 U377 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U378 ( .A(n375), .B(n323), .ZN(n324) );
  XNOR2_X1 U379 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U380 ( .A(n327), .B(n326), .ZN(n556) );
  XOR2_X1 U381 ( .A(KEYINPUT89), .B(KEYINPUT23), .Z(n329) );
  XNOR2_X1 U382 ( .A(G22GAT), .B(KEYINPUT24), .ZN(n328) );
  XNOR2_X1 U383 ( .A(n329), .B(n328), .ZN(n345) );
  XNOR2_X1 U384 ( .A(G218GAT), .B(G211GAT), .ZN(n330) );
  XNOR2_X1 U385 ( .A(n289), .B(n330), .ZN(n354) );
  XOR2_X1 U386 ( .A(n354), .B(KEYINPUT88), .Z(n332) );
  NAND2_X1 U387 ( .A1(G228GAT), .A2(G233GAT), .ZN(n331) );
  XNOR2_X1 U388 ( .A(n332), .B(n331), .ZN(n343) );
  XOR2_X1 U389 ( .A(KEYINPUT22), .B(KEYINPUT90), .Z(n334) );
  XNOR2_X1 U390 ( .A(G50GAT), .B(G204GAT), .ZN(n333) );
  XNOR2_X1 U391 ( .A(n334), .B(n333), .ZN(n337) );
  XOR2_X1 U392 ( .A(KEYINPUT70), .B(G78GAT), .Z(n336) );
  XNOR2_X1 U393 ( .A(G148GAT), .B(G106GAT), .ZN(n335) );
  XNOR2_X1 U394 ( .A(n336), .B(n335), .ZN(n426) );
  XOR2_X1 U395 ( .A(n337), .B(n426), .Z(n341) );
  XOR2_X1 U396 ( .A(KEYINPUT3), .B(G162GAT), .Z(n339) );
  XNOR2_X1 U397 ( .A(G155GAT), .B(G141GAT), .ZN(n338) );
  XNOR2_X1 U398 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U399 ( .A(KEYINPUT2), .B(n340), .Z(n383) );
  XNOR2_X1 U400 ( .A(n345), .B(n344), .ZN(n544) );
  XOR2_X1 U401 ( .A(n346), .B(KEYINPUT26), .Z(n563) );
  XOR2_X1 U402 ( .A(G204GAT), .B(G176GAT), .Z(n348) );
  XNOR2_X1 U403 ( .A(G92GAT), .B(G64GAT), .ZN(n347) );
  XNOR2_X1 U404 ( .A(n348), .B(n347), .ZN(n427) );
  XOR2_X1 U405 ( .A(G190GAT), .B(G36GAT), .Z(n394) );
  XOR2_X1 U406 ( .A(n427), .B(n394), .Z(n350) );
  NAND2_X1 U407 ( .A1(G226GAT), .A2(G233GAT), .ZN(n349) );
  XNOR2_X1 U408 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U409 ( .A(G8GAT), .B(G169GAT), .Z(n417) );
  XOR2_X1 U410 ( .A(n351), .B(n417), .Z(n353) );
  XNOR2_X1 U411 ( .A(KEYINPUT98), .B(KEYINPUT97), .ZN(n352) );
  XNOR2_X1 U412 ( .A(n353), .B(n352), .ZN(n357) );
  XOR2_X1 U413 ( .A(n355), .B(n354), .Z(n356) );
  XNOR2_X1 U414 ( .A(n357), .B(n356), .ZN(n539) );
  INV_X1 U415 ( .A(n539), .ZN(n490) );
  XNOR2_X1 U416 ( .A(KEYINPUT27), .B(n490), .ZN(n387) );
  XNOR2_X1 U417 ( .A(n359), .B(n358), .ZN(n364) );
  NAND2_X1 U418 ( .A1(n547), .A2(n490), .ZN(n360) );
  NAND2_X1 U419 ( .A1(n360), .A2(n544), .ZN(n361) );
  XNOR2_X1 U420 ( .A(n361), .B(KEYINPUT100), .ZN(n362) );
  XNOR2_X1 U421 ( .A(KEYINPUT25), .B(n362), .ZN(n363) );
  NOR2_X1 U422 ( .A1(n364), .A2(n363), .ZN(n365) );
  XNOR2_X1 U423 ( .A(n365), .B(KEYINPUT101), .ZN(n385) );
  XOR2_X1 U424 ( .A(n366), .B(KEYINPUT92), .Z(n368) );
  NAND2_X1 U425 ( .A1(G225GAT), .A2(G233GAT), .ZN(n367) );
  XNOR2_X1 U426 ( .A(n368), .B(n367), .ZN(n382) );
  XOR2_X1 U427 ( .A(KEYINPUT91), .B(KEYINPUT93), .Z(n370) );
  XNOR2_X1 U428 ( .A(KEYINPUT95), .B(KEYINPUT4), .ZN(n369) );
  XNOR2_X1 U429 ( .A(n370), .B(n369), .ZN(n374) );
  XOR2_X1 U430 ( .A(KEYINPUT94), .B(KEYINPUT1), .Z(n372) );
  XNOR2_X1 U431 ( .A(KEYINPUT6), .B(KEYINPUT5), .ZN(n371) );
  XNOR2_X1 U432 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U433 ( .A(n374), .B(n373), .Z(n380) );
  XOR2_X1 U434 ( .A(G29GAT), .B(G134GAT), .Z(n399) );
  XOR2_X1 U435 ( .A(G148GAT), .B(G85GAT), .Z(n377) );
  XOR2_X1 U436 ( .A(G120GAT), .B(G57GAT), .Z(n439) );
  XNOR2_X1 U437 ( .A(n375), .B(n439), .ZN(n376) );
  XNOR2_X1 U438 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U439 ( .A(n399), .B(n378), .ZN(n379) );
  XNOR2_X1 U440 ( .A(n380), .B(n379), .ZN(n381) );
  XNOR2_X1 U441 ( .A(n382), .B(n381), .ZN(n384) );
  XNOR2_X1 U442 ( .A(n384), .B(n383), .ZN(n386) );
  NAND2_X1 U443 ( .A1(n385), .A2(n386), .ZN(n390) );
  XNOR2_X1 U444 ( .A(KEYINPUT28), .B(n544), .ZN(n513) );
  NAND2_X1 U445 ( .A1(n543), .A2(n387), .ZN(n512) );
  NOR2_X1 U446 ( .A1(n547), .A2(n512), .ZN(n388) );
  NAND2_X1 U447 ( .A1(n513), .A2(n388), .ZN(n389) );
  NAND2_X1 U448 ( .A1(n390), .A2(n389), .ZN(n454) );
  NAND2_X1 U449 ( .A1(n556), .A2(n454), .ZN(n391) );
  XNOR2_X1 U450 ( .A(KEYINPUT107), .B(n391), .ZN(n410) );
  XOR2_X1 U451 ( .A(KEYINPUT11), .B(KEYINPUT75), .Z(n393) );
  XNOR2_X1 U452 ( .A(G218GAT), .B(KEYINPUT67), .ZN(n392) );
  XNOR2_X1 U453 ( .A(n393), .B(n392), .ZN(n395) );
  XOR2_X1 U454 ( .A(n395), .B(n394), .Z(n401) );
  XNOR2_X1 U455 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n396) );
  XNOR2_X1 U456 ( .A(n290), .B(n396), .ZN(n421) );
  XOR2_X1 U457 ( .A(G85GAT), .B(G99GAT), .Z(n428) );
  NAND2_X1 U458 ( .A1(G232GAT), .A2(G233GAT), .ZN(n397) );
  XNOR2_X1 U459 ( .A(n288), .B(n397), .ZN(n398) );
  XNOR2_X1 U460 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U461 ( .A(n401), .B(n400), .ZN(n409) );
  XOR2_X1 U462 ( .A(KEYINPUT9), .B(KEYINPUT10), .Z(n403) );
  XNOR2_X1 U463 ( .A(KEYINPUT66), .B(KEYINPUT64), .ZN(n402) );
  XNOR2_X1 U464 ( .A(n403), .B(n402), .ZN(n407) );
  XOR2_X1 U465 ( .A(G106GAT), .B(G92GAT), .Z(n405) );
  XNOR2_X1 U466 ( .A(G162GAT), .B(KEYINPUT76), .ZN(n404) );
  XNOR2_X1 U467 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U468 ( .A(n407), .B(n406), .Z(n408) );
  XNOR2_X1 U469 ( .A(KEYINPUT36), .B(n523), .ZN(n503) );
  BUF_X1 U470 ( .A(n503), .Z(n576) );
  NAND2_X1 U471 ( .A1(n410), .A2(n576), .ZN(n411) );
  XNOR2_X1 U472 ( .A(G29GAT), .B(G36GAT), .ZN(n413) );
  XNOR2_X1 U473 ( .A(n413), .B(n412), .ZN(n425) );
  XOR2_X1 U474 ( .A(G197GAT), .B(G1GAT), .Z(n415) );
  XNOR2_X1 U475 ( .A(G141GAT), .B(G113GAT), .ZN(n414) );
  XNOR2_X1 U476 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U477 ( .A(n417), .B(n416), .Z(n419) );
  NAND2_X1 U478 ( .A1(G229GAT), .A2(G233GAT), .ZN(n418) );
  XNOR2_X1 U479 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U480 ( .A(n420), .B(KEYINPUT30), .Z(n423) );
  XNOR2_X1 U481 ( .A(n421), .B(KEYINPUT29), .ZN(n422) );
  XNOR2_X1 U482 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U483 ( .A(n425), .B(n424), .ZN(n565) );
  XNOR2_X1 U484 ( .A(n427), .B(n426), .ZN(n443) );
  XOR2_X1 U485 ( .A(n429), .B(n428), .Z(n431) );
  NAND2_X1 U486 ( .A1(G230GAT), .A2(G233GAT), .ZN(n430) );
  XNOR2_X1 U487 ( .A(n431), .B(n430), .ZN(n435) );
  XOR2_X1 U488 ( .A(KEYINPUT72), .B(KEYINPUT69), .Z(n433) );
  XNOR2_X1 U489 ( .A(KEYINPUT73), .B(KEYINPUT31), .ZN(n432) );
  XNOR2_X1 U490 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U491 ( .A(n435), .B(n434), .Z(n441) );
  XOR2_X1 U492 ( .A(KEYINPUT33), .B(KEYINPUT32), .Z(n437) );
  XNOR2_X1 U493 ( .A(KEYINPUT71), .B(KEYINPUT68), .ZN(n436) );
  XNOR2_X1 U494 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U495 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U496 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U497 ( .A(n443), .B(n442), .ZN(n570) );
  NOR2_X1 U498 ( .A1(n565), .A2(n570), .ZN(n444) );
  XNOR2_X1 U499 ( .A(n444), .B(KEYINPUT74), .ZN(n455) );
  NAND2_X1 U500 ( .A1(n487), .A2(n455), .ZN(n445) );
  XNOR2_X1 U501 ( .A(n446), .B(n445), .ZN(n447) );
  XOR2_X1 U502 ( .A(KEYINPUT38), .B(n447), .Z(n472) );
  NAND2_X1 U503 ( .A1(n547), .A2(n472), .ZN(n449) );
  XOR2_X1 U504 ( .A(KEYINPUT16), .B(KEYINPUT83), .Z(n451) );
  INV_X1 U505 ( .A(n556), .ZN(n574) );
  INV_X1 U506 ( .A(n523), .ZN(n559) );
  NAND2_X1 U507 ( .A1(n574), .A2(n559), .ZN(n450) );
  XNOR2_X1 U508 ( .A(n451), .B(n450), .ZN(n452) );
  XOR2_X1 U509 ( .A(KEYINPUT82), .B(n452), .Z(n453) );
  AND2_X1 U510 ( .A1(n454), .A2(n453), .ZN(n475) );
  NAND2_X1 U511 ( .A1(n455), .A2(n475), .ZN(n456) );
  XOR2_X1 U512 ( .A(KEYINPUT102), .B(n456), .Z(n466) );
  NAND2_X1 U513 ( .A1(n466), .A2(n543), .ZN(n459) );
  XOR2_X1 U514 ( .A(G1GAT), .B(KEYINPUT103), .Z(n457) );
  XNOR2_X1 U515 ( .A(KEYINPUT34), .B(n457), .ZN(n458) );
  XNOR2_X1 U516 ( .A(n459), .B(n458), .ZN(G1324GAT) );
  NAND2_X1 U517 ( .A1(n466), .A2(n490), .ZN(n460) );
  XNOR2_X1 U518 ( .A(n460), .B(KEYINPUT104), .ZN(n461) );
  XNOR2_X1 U519 ( .A(G8GAT), .B(n461), .ZN(G1325GAT) );
  XOR2_X1 U520 ( .A(KEYINPUT35), .B(KEYINPUT106), .Z(n463) );
  NAND2_X1 U521 ( .A1(n466), .A2(n547), .ZN(n462) );
  XNOR2_X1 U522 ( .A(n463), .B(n462), .ZN(n465) );
  XOR2_X1 U523 ( .A(G15GAT), .B(KEYINPUT105), .Z(n464) );
  XNOR2_X1 U524 ( .A(n465), .B(n464), .ZN(G1326GAT) );
  INV_X1 U525 ( .A(n513), .ZN(n495) );
  NAND2_X1 U526 ( .A1(n466), .A2(n495), .ZN(n467) );
  XNOR2_X1 U527 ( .A(n467), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U528 ( .A(G29GAT), .B(KEYINPUT39), .Z(n469) );
  NAND2_X1 U529 ( .A1(n472), .A2(n543), .ZN(n468) );
  XNOR2_X1 U530 ( .A(n469), .B(n468), .ZN(G1328GAT) );
  NAND2_X1 U531 ( .A1(n472), .A2(n490), .ZN(n470) );
  XNOR2_X1 U532 ( .A(n470), .B(KEYINPUT110), .ZN(n471) );
  XNOR2_X1 U533 ( .A(G36GAT), .B(n471), .ZN(G1329GAT) );
  XOR2_X1 U534 ( .A(G50GAT), .B(KEYINPUT111), .Z(n474) );
  NAND2_X1 U535 ( .A1(n472), .A2(n495), .ZN(n473) );
  XNOR2_X1 U536 ( .A(n474), .B(n473), .ZN(G1331GAT) );
  INV_X1 U537 ( .A(n565), .ZN(n516) );
  XNOR2_X1 U538 ( .A(n570), .B(KEYINPUT41), .ZN(n552) );
  NOR2_X1 U539 ( .A1(n516), .A2(n552), .ZN(n486) );
  AND2_X1 U540 ( .A1(n486), .A2(n475), .ZN(n482) );
  NAND2_X1 U541 ( .A1(n543), .A2(n482), .ZN(n476) );
  XNOR2_X1 U542 ( .A(KEYINPUT42), .B(n476), .ZN(n477) );
  XNOR2_X1 U543 ( .A(G57GAT), .B(n477), .ZN(G1332GAT) );
  NAND2_X1 U544 ( .A1(n482), .A2(n490), .ZN(n478) );
  XNOR2_X1 U545 ( .A(n478), .B(KEYINPUT112), .ZN(n479) );
  XNOR2_X1 U546 ( .A(G64GAT), .B(n479), .ZN(G1333GAT) );
  XOR2_X1 U547 ( .A(G71GAT), .B(KEYINPUT113), .Z(n481) );
  NAND2_X1 U548 ( .A1(n482), .A2(n547), .ZN(n480) );
  XNOR2_X1 U549 ( .A(n481), .B(n480), .ZN(G1334GAT) );
  XOR2_X1 U550 ( .A(KEYINPUT114), .B(KEYINPUT43), .Z(n484) );
  NAND2_X1 U551 ( .A1(n482), .A2(n495), .ZN(n483) );
  XNOR2_X1 U552 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U553 ( .A(G78GAT), .B(n485), .ZN(G1335GAT) );
  NAND2_X1 U554 ( .A1(n487), .A2(n486), .ZN(n488) );
  XNOR2_X1 U555 ( .A(KEYINPUT115), .B(n488), .ZN(n494) );
  NAND2_X1 U556 ( .A1(n494), .A2(n543), .ZN(n489) );
  XNOR2_X1 U557 ( .A(n489), .B(G85GAT), .ZN(G1336GAT) );
  NAND2_X1 U558 ( .A1(n494), .A2(n490), .ZN(n491) );
  XNOR2_X1 U559 ( .A(n491), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U560 ( .A1(n547), .A2(n494), .ZN(n492) );
  XNOR2_X1 U561 ( .A(n492), .B(KEYINPUT116), .ZN(n493) );
  XNOR2_X1 U562 ( .A(G99GAT), .B(n493), .ZN(G1338GAT) );
  NAND2_X1 U563 ( .A1(n495), .A2(n494), .ZN(n496) );
  XNOR2_X1 U564 ( .A(n496), .B(KEYINPUT44), .ZN(n497) );
  XNOR2_X1 U565 ( .A(G106GAT), .B(n497), .ZN(G1339GAT) );
  NOR2_X1 U566 ( .A1(n565), .A2(n552), .ZN(n499) );
  XNOR2_X1 U567 ( .A(KEYINPUT117), .B(KEYINPUT46), .ZN(n498) );
  XNOR2_X1 U568 ( .A(n499), .B(n498), .ZN(n500) );
  NAND2_X1 U569 ( .A1(n500), .A2(n556), .ZN(n501) );
  NOR2_X1 U570 ( .A1(n523), .A2(n501), .ZN(n502) );
  XOR2_X1 U571 ( .A(KEYINPUT47), .B(n502), .Z(n510) );
  NAND2_X1 U572 ( .A1(n574), .A2(n503), .ZN(n504) );
  XNOR2_X1 U573 ( .A(n504), .B(KEYINPUT45), .ZN(n505) );
  XNOR2_X1 U574 ( .A(n505), .B(KEYINPUT65), .ZN(n506) );
  NAND2_X1 U575 ( .A1(n506), .A2(n565), .ZN(n507) );
  XNOR2_X1 U576 ( .A(KEYINPUT118), .B(n508), .ZN(n509) );
  NOR2_X1 U577 ( .A1(n510), .A2(n509), .ZN(n511) );
  XNOR2_X1 U578 ( .A(n511), .B(KEYINPUT48), .ZN(n540) );
  NOR2_X1 U579 ( .A1(n512), .A2(n540), .ZN(n528) );
  NAND2_X1 U580 ( .A1(n513), .A2(n528), .ZN(n514) );
  NOR2_X1 U581 ( .A1(n515), .A2(n514), .ZN(n524) );
  NAND2_X1 U582 ( .A1(n516), .A2(n524), .ZN(n517) );
  XNOR2_X1 U583 ( .A(G113GAT), .B(n517), .ZN(G1340GAT) );
  XOR2_X1 U584 ( .A(G120GAT), .B(KEYINPUT49), .Z(n520) );
  INV_X1 U585 ( .A(n552), .ZN(n518) );
  NAND2_X1 U586 ( .A1(n524), .A2(n518), .ZN(n519) );
  XNOR2_X1 U587 ( .A(n520), .B(n519), .ZN(G1341GAT) );
  NAND2_X1 U588 ( .A1(n524), .A2(n574), .ZN(n521) );
  XNOR2_X1 U589 ( .A(n521), .B(KEYINPUT50), .ZN(n522) );
  XNOR2_X1 U590 ( .A(G127GAT), .B(n522), .ZN(G1342GAT) );
  XOR2_X1 U591 ( .A(KEYINPUT119), .B(KEYINPUT51), .Z(n526) );
  NAND2_X1 U592 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U593 ( .A(n526), .B(n525), .ZN(n527) );
  XOR2_X1 U594 ( .A(G134GAT), .B(n527), .Z(G1343GAT) );
  NAND2_X1 U595 ( .A1(n528), .A2(n563), .ZN(n536) );
  NOR2_X1 U596 ( .A1(n565), .A2(n536), .ZN(n529) );
  XOR2_X1 U597 ( .A(G141GAT), .B(n529), .Z(G1344GAT) );
  XOR2_X1 U598 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n531) );
  XNOR2_X1 U599 ( .A(G148GAT), .B(KEYINPUT120), .ZN(n530) );
  XNOR2_X1 U600 ( .A(n531), .B(n530), .ZN(n533) );
  NOR2_X1 U601 ( .A1(n552), .A2(n536), .ZN(n532) );
  XOR2_X1 U602 ( .A(n533), .B(n532), .Z(G1345GAT) );
  NOR2_X1 U603 ( .A1(n556), .A2(n536), .ZN(n535) );
  XNOR2_X1 U604 ( .A(G155GAT), .B(KEYINPUT121), .ZN(n534) );
  XNOR2_X1 U605 ( .A(n535), .B(n534), .ZN(G1346GAT) );
  NOR2_X1 U606 ( .A1(n559), .A2(n536), .ZN(n537) );
  XOR2_X1 U607 ( .A(KEYINPUT122), .B(n537), .Z(n538) );
  XNOR2_X1 U608 ( .A(G162GAT), .B(n538), .ZN(G1347GAT) );
  XOR2_X1 U609 ( .A(KEYINPUT123), .B(KEYINPUT55), .Z(n546) );
  NOR2_X1 U610 ( .A1(n540), .A2(n539), .ZN(n541) );
  XOR2_X1 U611 ( .A(KEYINPUT54), .B(n541), .Z(n542) );
  NAND2_X1 U612 ( .A1(n564), .A2(n544), .ZN(n545) );
  XNOR2_X1 U613 ( .A(n546), .B(n545), .ZN(n548) );
  NAND2_X1 U614 ( .A1(n548), .A2(n547), .ZN(n558) );
  NOR2_X1 U615 ( .A1(n565), .A2(n558), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n549), .B(KEYINPUT124), .ZN(n550) );
  INV_X1 U617 ( .A(n550), .ZN(n551) );
  XNOR2_X1 U618 ( .A(G169GAT), .B(n551), .ZN(G1348GAT) );
  NOR2_X1 U619 ( .A1(n552), .A2(n558), .ZN(n554) );
  XNOR2_X1 U620 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n553) );
  XNOR2_X1 U621 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U622 ( .A(G176GAT), .B(n555), .ZN(G1349GAT) );
  NOR2_X1 U623 ( .A1(n556), .A2(n558), .ZN(n557) );
  XOR2_X1 U624 ( .A(G183GAT), .B(n557), .Z(G1350GAT) );
  NOR2_X1 U625 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U626 ( .A(G190GAT), .B(n560), .ZN(n561) );
  INV_X1 U627 ( .A(n561), .ZN(n562) );
  XNOR2_X1 U628 ( .A(KEYINPUT58), .B(n562), .ZN(G1351GAT) );
  NAND2_X1 U629 ( .A1(n564), .A2(n563), .ZN(n569) );
  NOR2_X1 U630 ( .A1(n565), .A2(n569), .ZN(n567) );
  XNOR2_X1 U631 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U633 ( .A(G197GAT), .B(n568), .ZN(G1352GAT) );
  XOR2_X1 U634 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n572) );
  INV_X1 U635 ( .A(n569), .ZN(n577) );
  NAND2_X1 U636 ( .A1(n577), .A2(n570), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(n573) );
  XOR2_X1 U638 ( .A(G204GAT), .B(n573), .Z(G1353GAT) );
  NAND2_X1 U639 ( .A1(n577), .A2(n574), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n575), .B(G211GAT), .ZN(G1354GAT) );
  XNOR2_X1 U641 ( .A(G218GAT), .B(KEYINPUT126), .ZN(n581) );
  XOR2_X1 U642 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n579) );
  NAND2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n581), .B(n580), .ZN(G1355GAT) );
endmodule

