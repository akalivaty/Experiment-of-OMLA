//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 0 0 0 1 0 0 0 0 0 1 0 1 1 0 0 1 0 0 1 0 0 1 1 0 1 1 1 0 0 1 0 1 1 1 0 0 0 1 0 1 1 0 1 1 0 1 0 0 1 1 1 0 1 1 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:29 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1146, new_n1147, new_n1148, new_n1149, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1184, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1234, new_n1235, new_n1236, new_n1237, new_n1238, new_n1239,
    new_n1240, new_n1241, new_n1242, new_n1243, new_n1244, new_n1245,
    new_n1246, new_n1247, new_n1248, new_n1249;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n203), .A2(G50), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(new_n209), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n220));
  INV_X1    g0020(.A(G238), .ZN(new_n221));
  INV_X1    g0021(.A(G87), .ZN(new_n222));
  INV_X1    g0022(.A(G250), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n220), .B1(new_n202), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n225));
  INV_X1    g0025(.A(G232), .ZN(new_n226));
  INV_X1    g0026(.A(G97), .ZN(new_n227));
  INV_X1    g0027(.A(G257), .ZN(new_n228));
  OAI221_X1 g0028(.A(new_n225), .B1(new_n201), .B2(new_n226), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n211), .B1(new_n224), .B2(new_n229), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n214), .B(new_n219), .C1(KEYINPUT1), .C2(new_n230), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n230), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(new_n226), .ZN(new_n234));
  XOR2_X1   g0034(.A(KEYINPUT2), .B(G226), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n236), .B(new_n239), .Z(G358));
  XNOR2_X1  g0040(.A(G50), .B(G68), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G58), .B(G77), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n241), .B(new_n242), .Z(new_n243));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  INV_X1    g0047(.A(KEYINPUT3), .ZN(new_n248));
  INV_X1    g0048(.A(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(KEYINPUT3), .A2(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G1698), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n252), .A2(G222), .A3(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G77), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n252), .A2(G1698), .ZN(new_n256));
  INV_X1    g0056(.A(G223), .ZN(new_n257));
  OAI221_X1 g0057(.A(new_n254), .B1(new_n255), .B2(new_n252), .C1(new_n256), .C2(new_n257), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n217), .B1(G33), .B2(G41), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n261));
  INV_X1    g0061(.A(G274), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G41), .ZN(new_n264));
  INV_X1    g0064(.A(G45), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  AND2_X1   g0066(.A1(G1), .A2(G13), .ZN(new_n267));
  NAND2_X1  g0067(.A1(G33), .A2(G41), .ZN(new_n268));
  AOI22_X1  g0068(.A1(new_n208), .A2(new_n266), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n263), .B1(new_n269), .B2(G226), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n260), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G190), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n273), .B1(G200), .B2(new_n271), .ZN(new_n274));
  OAI21_X1  g0074(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n275));
  INV_X1    g0075(.A(G150), .ZN(new_n276));
  NOR2_X1   g0076(.A1(G20), .A2(G33), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  XNOR2_X1  g0078(.A(KEYINPUT8), .B(G58), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n209), .A2(G33), .ZN(new_n280));
  OAI221_X1 g0080(.A(new_n275), .B1(new_n276), .B2(new_n278), .C1(new_n279), .C2(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(new_n217), .ZN(new_n283));
  INV_X1    g0083(.A(G50), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  AOI22_X1  g0086(.A1(new_n281), .A2(new_n283), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(new_n283), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(new_n285), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT64), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n286), .A2(new_n283), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(KEYINPUT64), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n208), .A2(G20), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n291), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n287), .B1(new_n284), .B2(new_n295), .ZN(new_n296));
  XNOR2_X1  g0096(.A(new_n296), .B(KEYINPUT9), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n274), .A2(new_n297), .ZN(new_n298));
  XNOR2_X1  g0098(.A(new_n298), .B(KEYINPUT10), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n252), .A2(G232), .A3(G1698), .ZN(new_n300));
  NAND2_X1  g0100(.A1(G33), .A2(G97), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n252), .A2(new_n253), .ZN(new_n302));
  INV_X1    g0102(.A(G226), .ZN(new_n303));
  OAI211_X1 g0103(.A(new_n300), .B(new_n301), .C1(new_n302), .C2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(new_n259), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT13), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n263), .B1(new_n269), .B2(G238), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n305), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n306), .B1(new_n305), .B2(new_n307), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(G190), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n286), .A2(new_n202), .ZN(new_n313));
  XNOR2_X1  g0113(.A(new_n313), .B(KEYINPUT12), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n292), .A2(G68), .A3(new_n294), .ZN(new_n315));
  OAI22_X1  g0115(.A1(new_n280), .A2(new_n255), .B1(new_n209), .B2(G68), .ZN(new_n316));
  OAI22_X1  g0116(.A1(new_n316), .A2(KEYINPUT71), .B1(new_n284), .B2(new_n278), .ZN(new_n317));
  AND2_X1   g0117(.A1(new_n316), .A2(KEYINPUT71), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n283), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT11), .ZN(new_n320));
  OAI211_X1 g0120(.A(new_n314), .B(new_n315), .C1(new_n319), .C2(new_n320), .ZN(new_n321));
  AND2_X1   g0121(.A1(new_n319), .A2(new_n320), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  OAI21_X1  g0123(.A(G200), .B1(new_n309), .B2(new_n310), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n312), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(G169), .ZN(new_n327));
  OAI21_X1  g0127(.A(KEYINPUT14), .B1(new_n311), .B2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT14), .ZN(new_n329));
  OAI211_X1 g0129(.A(new_n329), .B(G169), .C1(new_n309), .C2(new_n310), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n311), .A2(G179), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n328), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(new_n323), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n326), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n250), .A2(new_n209), .A3(new_n251), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(KEYINPUT7), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT7), .ZN(new_n337));
  NAND4_X1  g0137(.A1(new_n250), .A2(new_n337), .A3(new_n209), .A4(new_n251), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n336), .A2(G68), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(G58), .A2(G68), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(KEYINPUT72), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT72), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n342), .A2(G58), .A3(G68), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n341), .A2(new_n343), .A3(new_n203), .ZN(new_n344));
  AOI22_X1  g0144(.A1(new_n344), .A2(G20), .B1(G159), .B2(new_n277), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT16), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n339), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n346), .B1(new_n339), .B2(new_n345), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n283), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  XOR2_X1   g0150(.A(KEYINPUT8), .B(G58), .Z(new_n351));
  NAND4_X1  g0151(.A1(new_n291), .A2(new_n293), .A3(new_n351), .A4(new_n294), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n279), .A2(new_n286), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n257), .A2(new_n253), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n303), .A2(G1698), .ZN(new_n357));
  AND2_X1   g0157(.A1(KEYINPUT3), .A2(G33), .ZN(new_n358));
  NOR2_X1   g0158(.A1(KEYINPUT3), .A2(G33), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n356), .B(new_n357), .C1(new_n358), .C2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(G33), .A2(G87), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(new_n259), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n263), .B1(new_n269), .B2(G232), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n363), .A2(new_n272), .A3(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(G200), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n267), .A2(new_n268), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n367), .B1(new_n360), .B2(new_n361), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n367), .A2(G232), .A3(new_n261), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n266), .A2(new_n208), .A3(G274), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n366), .B1(new_n368), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n365), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n350), .A2(new_n355), .A3(new_n373), .ZN(new_n374));
  XNOR2_X1  g0174(.A(new_n374), .B(KEYINPUT17), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n339), .A2(new_n345), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(KEYINPUT16), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n288), .B1(new_n377), .B2(new_n347), .ZN(new_n378));
  AND2_X1   g0178(.A1(KEYINPUT65), .A2(G179), .ZN(new_n379));
  NOR2_X1   g0179(.A1(KEYINPUT65), .A2(G179), .ZN(new_n380));
  OR2_X1    g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n363), .A2(new_n381), .A3(new_n364), .ZN(new_n382));
  OAI21_X1  g0182(.A(G169), .B1(new_n368), .B2(new_n371), .ZN(new_n383));
  AND3_X1   g0183(.A1(new_n382), .A2(new_n383), .A3(KEYINPUT73), .ZN(new_n384));
  AOI21_X1  g0184(.A(KEYINPUT73), .B1(new_n382), .B2(new_n383), .ZN(new_n385));
  OAI22_X1  g0185(.A1(new_n378), .A2(new_n354), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(KEYINPUT18), .ZN(new_n387));
  OR2_X1    g0187(.A1(new_n386), .A2(KEYINPUT18), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n375), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n271), .A2(new_n327), .ZN(new_n391));
  OAI211_X1 g0191(.A(new_n391), .B(new_n296), .C1(new_n381), .C2(new_n271), .ZN(new_n392));
  XOR2_X1   g0192(.A(new_n392), .B(KEYINPUT66), .Z(new_n393));
  NAND4_X1  g0193(.A1(new_n299), .A2(new_n334), .A3(new_n390), .A4(new_n393), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n252), .A2(G232), .A3(new_n253), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n358), .A2(new_n359), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(G107), .ZN(new_n397));
  OAI211_X1 g0197(.A(new_n395), .B(new_n397), .C1(new_n256), .C2(new_n221), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(new_n259), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n263), .B1(new_n269), .B2(G244), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT67), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n399), .A2(KEYINPUT67), .A3(new_n400), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(new_n381), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT68), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n351), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n279), .A2(KEYINPUT68), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n278), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  XNOR2_X1  g0211(.A(KEYINPUT15), .B(G87), .ZN(new_n412));
  OAI22_X1  g0212(.A1(new_n412), .A2(new_n280), .B1(new_n209), .B2(new_n255), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n283), .B1(new_n411), .B2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT69), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  OAI211_X1 g0216(.A(KEYINPUT69), .B(new_n283), .C1(new_n411), .C2(new_n413), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n294), .A2(G77), .ZN(new_n419));
  OAI22_X1  g0219(.A1(new_n289), .A2(new_n419), .B1(G77), .B2(new_n285), .ZN(new_n420));
  INV_X1    g0220(.A(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n418), .A2(new_n421), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n407), .B(new_n422), .C1(new_n405), .C2(G169), .ZN(new_n423));
  INV_X1    g0223(.A(new_n404), .ZN(new_n424));
  AOI21_X1  g0224(.A(KEYINPUT67), .B1(new_n399), .B2(new_n400), .ZN(new_n425));
  OAI21_X1  g0225(.A(G190), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n403), .A2(G200), .A3(new_n404), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n420), .B1(new_n416), .B2(new_n417), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n426), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n423), .A2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT70), .ZN(new_n431));
  XNOR2_X1  g0231(.A(new_n430), .B(new_n431), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n394), .A2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(G116), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n286), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n208), .A2(G33), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n285), .A2(new_n436), .A3(new_n217), .A4(new_n282), .ZN(new_n437));
  AOI22_X1  g0237(.A1(new_n282), .A2(new_n217), .B1(G20), .B2(new_n434), .ZN(new_n438));
  AOI21_X1  g0238(.A(G20), .B1(G33), .B2(G283), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n439), .B1(G33), .B2(new_n227), .ZN(new_n440));
  AND3_X1   g0240(.A1(new_n438), .A2(new_n440), .A3(KEYINPUT20), .ZN(new_n441));
  AOI21_X1  g0241(.A(KEYINPUT20), .B1(new_n438), .B2(new_n440), .ZN(new_n442));
  OAI221_X1 g0242(.A(new_n435), .B1(new_n434), .B2(new_n437), .C1(new_n441), .C2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT21), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT78), .ZN(new_n445));
  XNOR2_X1  g0245(.A(KEYINPUT5), .B(G41), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n208), .A2(G45), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n367), .A2(G274), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n445), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n262), .B1(new_n267), .B2(new_n268), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n452), .A2(KEYINPUT78), .A3(new_n446), .A4(new_n448), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n259), .B1(new_n448), .B2(new_n446), .ZN(new_n454));
  AOI22_X1  g0254(.A1(new_n451), .A2(new_n453), .B1(G270), .B2(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n252), .A2(G264), .A3(G1698), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n396), .A2(G303), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n456), .B(new_n457), .C1(new_n302), .C2(new_n228), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(new_n259), .ZN(new_n459));
  AOI211_X1 g0259(.A(new_n444), .B(new_n327), .C1(new_n455), .C2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n455), .A2(new_n459), .ZN(new_n461));
  INV_X1    g0261(.A(G179), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n443), .B1(new_n460), .B2(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n443), .B1(new_n461), .B2(G200), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n465), .B1(new_n272), .B2(new_n461), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n461), .A2(G169), .A3(new_n443), .ZN(new_n467));
  AND3_X1   g0267(.A1(new_n467), .A2(KEYINPUT81), .A3(new_n444), .ZN(new_n468));
  AOI21_X1  g0268(.A(KEYINPUT81), .B1(new_n467), .B2(new_n444), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n464), .B(new_n466), .C1(new_n468), .C2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(KEYINPUT75), .B1(new_n286), .B2(new_n227), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT75), .ZN(new_n473));
  NOR3_X1   g0273(.A1(new_n285), .A2(new_n473), .A3(G97), .ZN(new_n474));
  OAI22_X1  g0274(.A1(new_n472), .A2(new_n474), .B1(new_n227), .B2(new_n437), .ZN(new_n475));
  NOR2_X1   g0275(.A1(KEYINPUT74), .A2(KEYINPUT6), .ZN(new_n476));
  AND2_X1   g0276(.A1(G97), .A2(G107), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n476), .B1(new_n477), .B2(new_n205), .ZN(new_n478));
  OR2_X1    g0278(.A1(KEYINPUT74), .A2(KEYINPUT6), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n227), .A2(KEYINPUT6), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  XNOR2_X1  g0281(.A(G97), .B(G107), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n478), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(G20), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n336), .A2(G107), .A3(new_n338), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n277), .A2(G77), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n484), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n475), .B1(new_n487), .B2(new_n283), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(KEYINPUT76), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT76), .ZN(new_n490));
  AOI22_X1  g0290(.A1(new_n483), .A2(G20), .B1(G77), .B2(new_n277), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n288), .B1(new_n491), .B2(new_n485), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n490), .B1(new_n492), .B2(new_n475), .ZN(new_n493));
  OAI211_X1 g0293(.A(G244), .B(new_n253), .C1(new_n358), .C2(new_n359), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT4), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n494), .A2(KEYINPUT77), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(KEYINPUT77), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n252), .A2(G244), .A3(new_n253), .A4(new_n497), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n252), .A2(G250), .A3(G1698), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT77), .ZN(new_n500));
  AOI22_X1  g0300(.A1(new_n500), .A2(KEYINPUT4), .B1(G33), .B2(G283), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n496), .A2(new_n498), .A3(new_n499), .A4(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(new_n259), .ZN(new_n503));
  AOI22_X1  g0303(.A1(new_n451), .A2(new_n453), .B1(G257), .B2(new_n454), .ZN(new_n504));
  AND3_X1   g0304(.A1(new_n503), .A2(new_n272), .A3(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(G200), .B1(new_n503), .B2(new_n504), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n489), .B(new_n493), .C1(new_n505), .C2(new_n506), .ZN(new_n507));
  AND3_X1   g0307(.A1(new_n503), .A2(new_n381), .A3(new_n504), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n327), .B1(new_n503), .B2(new_n504), .ZN(new_n509));
  OAI22_X1  g0309(.A1(new_n508), .A2(new_n509), .B1(new_n492), .B2(new_n475), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT79), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n447), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n208), .A2(KEYINPUT79), .A3(G45), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n367), .A2(G250), .ZN(new_n515));
  OAI22_X1  g0315(.A1(new_n514), .A2(new_n515), .B1(new_n262), .B2(new_n447), .ZN(new_n516));
  OAI211_X1 g0316(.A(G238), .B(new_n253), .C1(new_n358), .C2(new_n359), .ZN(new_n517));
  OAI211_X1 g0317(.A(G244), .B(G1698), .C1(new_n358), .C2(new_n359), .ZN(new_n518));
  NAND2_X1  g0318(.A1(G33), .A2(G116), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n516), .B1(new_n259), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(G190), .ZN(new_n522));
  AND2_X1   g0322(.A1(new_n512), .A2(new_n513), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n259), .A2(new_n223), .ZN(new_n524));
  AOI22_X1  g0324(.A1(new_n523), .A2(new_n524), .B1(G274), .B2(new_n448), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n520), .A2(new_n259), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(G200), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n252), .A2(new_n209), .A3(G68), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT19), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n209), .B1(new_n301), .B2(new_n530), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n531), .B1(G87), .B2(new_n206), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n530), .B1(new_n280), .B2(new_n227), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n529), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n534), .A2(new_n283), .B1(new_n412), .B2(new_n286), .ZN(new_n535));
  INV_X1    g0335(.A(new_n437), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(G87), .ZN(new_n537));
  XNOR2_X1  g0337(.A(new_n537), .B(KEYINPUT80), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n522), .A2(new_n528), .A3(new_n535), .A4(new_n538), .ZN(new_n539));
  AND3_X1   g0339(.A1(new_n507), .A2(new_n510), .A3(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n252), .A2(G250), .A3(new_n253), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n252), .A2(G257), .A3(G1698), .ZN(new_n542));
  NAND2_X1  g0342(.A1(G33), .A2(G294), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(new_n259), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n451), .A2(new_n453), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n449), .A2(G264), .A3(new_n367), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(G169), .ZN(new_n549));
  AOI22_X1  g0349(.A1(new_n259), .A2(new_n544), .B1(new_n451), .B2(new_n453), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n547), .A2(KEYINPUT83), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT83), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n454), .A2(new_n552), .A3(G264), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n550), .A2(new_n554), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n549), .B1(new_n462), .B2(new_n555), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n209), .B(G87), .C1(new_n358), .C2(new_n359), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(KEYINPUT22), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT22), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n252), .A2(new_n559), .A3(new_n209), .A4(G87), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT24), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n519), .A2(G20), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT23), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n564), .B1(new_n209), .B2(G107), .ZN(new_n565));
  INV_X1    g0365(.A(G107), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n566), .A2(KEYINPUT23), .A3(G20), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n563), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  AND3_X1   g0368(.A1(new_n561), .A2(new_n562), .A3(new_n568), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n562), .B1(new_n561), .B2(new_n568), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n283), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT25), .ZN(new_n572));
  AOI211_X1 g0372(.A(G107), .B(new_n285), .C1(KEYINPUT82), .C2(new_n572), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n572), .A2(KEYINPUT82), .ZN(new_n574));
  OR2_X1    g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n573), .A2(new_n574), .ZN(new_n576));
  AOI22_X1  g0376(.A1(new_n575), .A2(new_n576), .B1(new_n536), .B2(G107), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n571), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n556), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(G200), .B1(new_n550), .B2(new_n554), .ZN(new_n580));
  AND4_X1   g0380(.A1(new_n272), .A2(new_n545), .A3(new_n546), .A4(new_n547), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n571), .B(new_n577), .C1(new_n580), .C2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(new_n412), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n536), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n535), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n527), .A2(new_n327), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n525), .A2(new_n526), .A3(new_n406), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  AND3_X1   g0388(.A1(new_n579), .A2(new_n582), .A3(new_n588), .ZN(new_n589));
  AND4_X1   g0389(.A1(new_n433), .A2(new_n471), .A3(new_n540), .A4(new_n589), .ZN(G372));
  INV_X1    g0390(.A(new_n299), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n332), .A2(new_n333), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n423), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n593), .A2(new_n325), .A3(new_n375), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT18), .ZN(new_n595));
  XNOR2_X1  g0395(.A(new_n386), .B(new_n595), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n591), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT86), .ZN(new_n598));
  INV_X1    g0398(.A(new_n393), .ZN(new_n599));
  OR3_X1    g0399(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n598), .B1(new_n597), .B2(new_n599), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(new_n433), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT26), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n487), .A2(new_n283), .ZN(new_n605));
  INV_X1    g0405(.A(new_n475), .ZN(new_n606));
  AOI21_X1  g0406(.A(KEYINPUT76), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  AOI211_X1 g0407(.A(new_n490), .B(new_n475), .C1(new_n487), .C2(new_n283), .ZN(new_n608));
  OAI22_X1  g0408(.A1(new_n607), .A2(new_n608), .B1(new_n508), .B2(new_n509), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n539), .A2(new_n588), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n604), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(KEYINPUT84), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT84), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n613), .B(new_n604), .C1(new_n609), .C2(new_n610), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n503), .A2(new_n504), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(G169), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n503), .A2(new_n504), .A3(new_n381), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n488), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n618), .A2(KEYINPUT26), .A3(new_n539), .A4(new_n588), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(KEYINPUT85), .ZN(new_n620));
  INV_X1    g0420(.A(new_n610), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT85), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n621), .A2(new_n618), .A3(new_n622), .A4(KEYINPUT26), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n612), .A2(new_n614), .A3(new_n620), .A4(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n588), .ZN(new_n625));
  AND4_X1   g0425(.A1(new_n510), .A2(new_n507), .A3(new_n539), .A4(new_n582), .ZN(new_n626));
  OAI211_X1 g0426(.A(new_n579), .B(new_n464), .C1(new_n468), .C2(new_n469), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n625), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  AND2_X1   g0428(.A1(new_n624), .A2(new_n628), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n602), .B1(new_n603), .B2(new_n629), .ZN(G369));
  NAND3_X1  g0430(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n631));
  OAI21_X1  g0431(.A(G213), .B1(new_n631), .B2(KEYINPUT27), .ZN(new_n632));
  AOI21_X1  g0432(.A(KEYINPUT87), .B1(new_n631), .B2(KEYINPUT27), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n631), .A2(KEYINPUT87), .A3(KEYINPUT27), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n632), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(G343), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(new_n443), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n471), .A2(new_n639), .ZN(new_n640));
  OR2_X1    g0440(.A1(new_n468), .A2(new_n469), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(new_n464), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n640), .B1(new_n643), .B2(new_n639), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n644), .A2(G330), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n579), .A2(new_n582), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n578), .A2(new_n638), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n648), .B1(new_n579), .B2(new_n637), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n645), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n556), .A2(new_n578), .A3(new_n637), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n642), .A2(new_n646), .A3(new_n637), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n650), .A2(new_n651), .A3(new_n652), .ZN(G399));
  INV_X1    g0453(.A(new_n212), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n654), .A2(G41), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  NOR3_X1   g0456(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n656), .A2(G1), .A3(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n658), .B1(new_n215), .B2(new_n656), .ZN(new_n659));
  XNOR2_X1  g0459(.A(new_n659), .B(KEYINPUT28), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n638), .B1(new_n624), .B2(new_n628), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT29), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n626), .A2(new_n627), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(new_n588), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n610), .A2(new_n510), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(new_n604), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n609), .A2(new_n610), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n668), .B1(new_n669), .B2(new_n604), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n637), .B1(new_n666), .B2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT89), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  OAI211_X1 g0473(.A(KEYINPUT89), .B(new_n637), .C1(new_n666), .C2(new_n670), .ZN(new_n674));
  AND2_X1   g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n664), .B1(new_n675), .B2(new_n663), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT31), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n471), .A2(new_n540), .A3(new_n589), .A4(new_n637), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n521), .A2(new_n554), .A3(new_n545), .ZN(new_n679));
  NOR4_X1   g0479(.A1(new_n679), .A2(new_n615), .A3(new_n461), .A4(new_n462), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n461), .A2(new_n406), .A3(new_n527), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n555), .A2(new_n615), .ZN(new_n682));
  OAI22_X1  g0482(.A1(new_n680), .A2(KEYINPUT30), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  AND2_X1   g0483(.A1(new_n680), .A2(KEYINPUT30), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n638), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n677), .B1(new_n678), .B2(new_n685), .ZN(new_n686));
  AND2_X1   g0486(.A1(new_n685), .A2(new_n677), .ZN(new_n687));
  OAI21_X1  g0487(.A(G330), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT88), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  OAI211_X1 g0490(.A(KEYINPUT88), .B(G330), .C1(new_n686), .C2(new_n687), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n676), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT90), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n676), .A2(KEYINPUT90), .A3(new_n692), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n660), .B1(new_n697), .B2(G1), .ZN(G364));
  AND2_X1   g0498(.A1(new_n209), .A2(G13), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n208), .B1(new_n699), .B2(G45), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n655), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n644), .A2(G330), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  AOI211_X1 g0504(.A(new_n702), .B(new_n645), .C1(new_n704), .C2(KEYINPUT91), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n705), .B1(KEYINPUT91), .B2(new_n704), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n217), .B1(G20), .B2(new_n327), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n209), .A2(G190), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NOR3_X1   g0509(.A1(new_n709), .A2(G179), .A3(G200), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(G159), .ZN(new_n711));
  XOR2_X1   g0511(.A(new_n711), .B(KEYINPUT32), .Z(new_n712));
  NOR2_X1   g0512(.A1(new_n209), .A2(new_n272), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n381), .A2(new_n366), .A3(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n712), .B1(new_n201), .B2(new_n714), .ZN(new_n715));
  NOR3_X1   g0515(.A1(new_n272), .A2(G179), .A3(G200), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n716), .A2(new_n209), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(G97), .ZN(new_n719));
  NOR3_X1   g0519(.A1(new_n209), .A2(new_n272), .A3(new_n366), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n381), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n709), .A2(new_n366), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(new_n381), .ZN(new_n723));
  OAI221_X1 g0523(.A(new_n719), .B1(new_n284), .B2(new_n721), .C1(new_n202), .C2(new_n723), .ZN(new_n724));
  NOR3_X1   g0524(.A1(new_n406), .A2(G200), .A3(new_n709), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n726), .A2(new_n255), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n366), .A2(G179), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n708), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n713), .A2(new_n728), .ZN(new_n730));
  OAI221_X1 g0530(.A(new_n252), .B1(new_n729), .B2(new_n566), .C1(new_n222), .C2(new_n730), .ZN(new_n731));
  NOR4_X1   g0531(.A1(new_n715), .A2(new_n724), .A3(new_n727), .A4(new_n731), .ZN(new_n732));
  OR2_X1    g0532(.A1(new_n730), .A2(KEYINPUT93), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n730), .A2(KEYINPUT93), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n714), .ZN(new_n737));
  AOI22_X1  g0537(.A1(new_n736), .A2(G303), .B1(G322), .B2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(G311), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n738), .B1(new_n739), .B2(new_n726), .ZN(new_n740));
  INV_X1    g0540(.A(new_n729), .ZN(new_n741));
  AOI22_X1  g0541(.A1(new_n710), .A2(G329), .B1(new_n741), .B2(G283), .ZN(new_n742));
  XOR2_X1   g0542(.A(new_n742), .B(KEYINPUT94), .Z(new_n743));
  INV_X1    g0543(.A(new_n721), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n252), .B1(new_n744), .B2(G326), .ZN(new_n745));
  INV_X1    g0545(.A(G294), .ZN(new_n746));
  XOR2_X1   g0546(.A(KEYINPUT33), .B(G317), .Z(new_n747));
  OAI221_X1 g0547(.A(new_n745), .B1(new_n746), .B2(new_n717), .C1(new_n723), .C2(new_n747), .ZN(new_n748));
  NOR3_X1   g0548(.A1(new_n740), .A2(new_n743), .A3(new_n748), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n707), .B1(new_n732), .B2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(G13), .A2(G33), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(G20), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n753), .A2(new_n707), .ZN(new_n754));
  XOR2_X1   g0554(.A(new_n754), .B(KEYINPUT92), .Z(new_n755));
  NAND2_X1  g0555(.A1(new_n212), .A2(new_n252), .ZN(new_n756));
  INV_X1    g0556(.A(G355), .ZN(new_n757));
  OAI22_X1  g0557(.A1(new_n756), .A2(new_n757), .B1(G116), .B2(new_n212), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n654), .A2(new_n252), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n760), .B1(new_n265), .B2(new_n216), .ZN(new_n761));
  OR2_X1    g0561(.A1(new_n243), .A2(new_n265), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n758), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  OAI211_X1 g0563(.A(new_n750), .B(new_n702), .C1(new_n755), .C2(new_n763), .ZN(new_n764));
  XNOR2_X1  g0564(.A(new_n764), .B(KEYINPUT95), .ZN(new_n765));
  INV_X1    g0565(.A(new_n753), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n765), .B1(new_n644), .B2(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n706), .A2(new_n767), .ZN(G396));
  NAND2_X1  g0568(.A1(new_n422), .A2(new_n638), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n429), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(new_n423), .ZN(new_n771));
  INV_X1    g0571(.A(new_n405), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n428), .B1(new_n772), .B2(new_n327), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n773), .A2(new_n407), .A3(new_n637), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n771), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  XNOR2_X1  g0576(.A(new_n661), .B(new_n776), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n702), .B1(new_n692), .B2(new_n777), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n778), .B1(new_n692), .B2(new_n777), .ZN(new_n779));
  OAI22_X1  g0579(.A1(new_n735), .A2(new_n284), .B1(new_n202), .B2(new_n729), .ZN(new_n780));
  XNOR2_X1  g0580(.A(new_n780), .B(KEYINPUT96), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n396), .B1(new_n710), .B2(G132), .ZN(new_n782));
  OAI211_X1 g0582(.A(new_n781), .B(new_n782), .C1(new_n201), .C2(new_n717), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n783), .B(KEYINPUT97), .ZN(new_n784));
  INV_X1    g0584(.A(new_n723), .ZN(new_n785));
  AOI22_X1  g0585(.A1(new_n785), .A2(G150), .B1(G137), .B2(new_n744), .ZN(new_n786));
  INV_X1    g0586(.A(G143), .ZN(new_n787));
  INV_X1    g0587(.A(G159), .ZN(new_n788));
  OAI221_X1 g0588(.A(new_n786), .B1(new_n787), .B2(new_n714), .C1(new_n788), .C2(new_n726), .ZN(new_n789));
  XOR2_X1   g0589(.A(new_n789), .B(KEYINPUT34), .Z(new_n790));
  NOR2_X1   g0590(.A1(new_n784), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(G303), .ZN(new_n792));
  INV_X1    g0592(.A(G283), .ZN(new_n793));
  OAI221_X1 g0593(.A(new_n719), .B1(new_n792), .B2(new_n721), .C1(new_n793), .C2(new_n723), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n726), .A2(new_n434), .ZN(new_n795));
  OAI22_X1  g0595(.A1(new_n735), .A2(new_n566), .B1(new_n746), .B2(new_n714), .ZN(new_n796));
  INV_X1    g0596(.A(new_n710), .ZN(new_n797));
  OAI221_X1 g0597(.A(new_n396), .B1(new_n222), .B2(new_n729), .C1(new_n797), .C2(new_n739), .ZN(new_n798));
  NOR4_X1   g0598(.A1(new_n794), .A2(new_n795), .A3(new_n796), .A4(new_n798), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n707), .B1(new_n791), .B2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n702), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n707), .A2(new_n751), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n801), .B1(new_n255), .B2(new_n802), .ZN(new_n803));
  OAI211_X1 g0603(.A(new_n800), .B(new_n803), .C1(new_n776), .C2(new_n752), .ZN(new_n804));
  AND2_X1   g0604(.A1(new_n779), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(G384));
  OR2_X1    g0606(.A1(new_n483), .A2(KEYINPUT35), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n483), .A2(KEYINPUT35), .ZN(new_n808));
  NAND4_X1  g0608(.A1(new_n807), .A2(G116), .A3(new_n218), .A4(new_n808), .ZN(new_n809));
  XNOR2_X1  g0609(.A(KEYINPUT98), .B(KEYINPUT36), .ZN(new_n810));
  XNOR2_X1  g0610(.A(new_n809), .B(new_n810), .ZN(new_n811));
  NAND4_X1  g0611(.A1(new_n216), .A2(G77), .A3(new_n343), .A4(new_n341), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n284), .A2(G68), .ZN(new_n813));
  AOI211_X1 g0613(.A(new_n208), .B(G13), .C1(new_n812), .C2(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n811), .A2(new_n814), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n334), .B1(new_n323), .B2(new_n637), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n332), .A2(new_n333), .A3(new_n638), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n818), .A2(new_n776), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n686), .A2(new_n687), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n636), .B1(new_n378), .B2(new_n354), .ZN(new_n822));
  INV_X1    g0622(.A(KEYINPUT101), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  OAI211_X1 g0624(.A(KEYINPUT101), .B(new_n636), .C1(new_n378), .C2(new_n354), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n389), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n386), .A2(new_n374), .ZN(new_n828));
  OAI21_X1  g0628(.A(KEYINPUT37), .B1(new_n826), .B2(new_n828), .ZN(new_n829));
  AND2_X1   g0629(.A1(new_n386), .A2(new_n374), .ZN(new_n830));
  INV_X1    g0630(.A(KEYINPUT37), .ZN(new_n831));
  NAND4_X1  g0631(.A1(new_n830), .A2(new_n831), .A3(new_n824), .A4(new_n825), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n829), .A2(new_n832), .ZN(new_n833));
  AOI21_X1  g0633(.A(KEYINPUT38), .B1(new_n827), .B2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n386), .A2(new_n822), .A3(new_n374), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n836), .A2(KEYINPUT37), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT100), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n836), .A2(KEYINPUT100), .A3(KEYINPUT37), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n839), .A2(new_n832), .A3(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n822), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n389), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n841), .A2(new_n843), .A3(KEYINPUT38), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n835), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n821), .A2(KEYINPUT40), .A3(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT103), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND4_X1  g0648(.A1(new_n821), .A2(KEYINPUT103), .A3(KEYINPUT40), .A4(new_n845), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n841), .A2(new_n843), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT38), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(new_n844), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n821), .A2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT40), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n850), .A2(new_n857), .ZN(new_n858));
  XOR2_X1   g0658(.A(new_n858), .B(KEYINPUT104), .Z(new_n859));
  OR3_X1    g0659(.A1(new_n859), .A2(new_n603), .A3(new_n820), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n859), .B1(new_n603), .B2(new_n820), .ZN(new_n861));
  AND3_X1   g0661(.A1(new_n860), .A2(G330), .A3(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n774), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n863), .B1(new_n661), .B2(new_n776), .ZN(new_n864));
  AND2_X1   g0664(.A1(new_n816), .A2(new_n817), .ZN(new_n865));
  OAI21_X1  g0665(.A(KEYINPUT99), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT99), .ZN(new_n867));
  AOI211_X1 g0667(.A(new_n638), .B(new_n775), .C1(new_n624), .C2(new_n628), .ZN(new_n868));
  OAI211_X1 g0668(.A(new_n867), .B(new_n818), .C1(new_n868), .C2(new_n863), .ZN(new_n869));
  AND3_X1   g0669(.A1(new_n866), .A2(new_n854), .A3(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT39), .ZN(new_n871));
  AND3_X1   g0671(.A1(new_n841), .A2(new_n843), .A3(KEYINPUT38), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n871), .B1(new_n872), .B2(new_n834), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n853), .A2(KEYINPUT39), .A3(new_n844), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n592), .A2(new_n638), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  OR2_X1    g0676(.A1(new_n596), .A2(new_n636), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g0678(.A(KEYINPUT102), .B1(new_n870), .B2(new_n878), .ZN(new_n879));
  AND2_X1   g0679(.A1(new_n876), .A2(new_n877), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT102), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n866), .A2(new_n869), .A3(new_n854), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n880), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n879), .A2(new_n883), .ZN(new_n884));
  OAI211_X1 g0684(.A(new_n433), .B(new_n664), .C1(new_n675), .C2(new_n663), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(new_n602), .ZN(new_n886));
  XNOR2_X1  g0686(.A(new_n884), .B(new_n886), .ZN(new_n887));
  OAI22_X1  g0687(.A1(new_n862), .A2(new_n887), .B1(new_n208), .B2(new_n699), .ZN(new_n888));
  AND2_X1   g0688(.A1(new_n862), .A2(new_n887), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n815), .B1(new_n888), .B2(new_n889), .ZN(G367));
  NOR2_X1   g0690(.A1(new_n643), .A2(new_n638), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT106), .ZN(new_n892));
  OAI221_X1 g0692(.A(new_n652), .B1(new_n649), .B2(new_n891), .C1(new_n645), .C2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n645), .A2(new_n892), .ZN(new_n894));
  XOR2_X1   g0694(.A(new_n893), .B(new_n894), .Z(new_n895));
  OR2_X1    g0695(.A1(new_n609), .A2(new_n637), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n638), .B1(new_n607), .B2(new_n608), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n507), .A2(new_n897), .A3(new_n510), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n899), .B1(new_n652), .B2(new_n651), .ZN(new_n900));
  XNOR2_X1  g0700(.A(new_n900), .B(KEYINPUT44), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n652), .A2(new_n651), .A3(new_n899), .ZN(new_n902));
  XOR2_X1   g0702(.A(KEYINPUT105), .B(KEYINPUT45), .Z(new_n903));
  XNOR2_X1  g0703(.A(new_n902), .B(new_n903), .ZN(new_n904));
  AND3_X1   g0704(.A1(new_n901), .A2(new_n650), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n650), .B1(new_n901), .B2(new_n904), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  AOI22_X1  g0707(.A1(new_n895), .A2(new_n907), .B1(new_n695), .B2(new_n696), .ZN(new_n908));
  XOR2_X1   g0708(.A(new_n655), .B(KEYINPUT41), .Z(new_n909));
  OAI21_X1  g0709(.A(new_n700), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n652), .B1(new_n898), .B2(new_n896), .ZN(new_n911));
  XNOR2_X1  g0711(.A(new_n911), .B(KEYINPUT42), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n579), .B1(new_n896), .B2(new_n898), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n637), .B1(new_n913), .B2(new_n618), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n538), .A2(new_n535), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(new_n638), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n621), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n625), .A2(new_n916), .A3(new_n638), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(KEYINPUT43), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n915), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n920), .A2(KEYINPUT43), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(new_n924), .ZN(new_n925));
  NOR3_X1   g0725(.A1(new_n915), .A2(KEYINPUT43), .A3(new_n920), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(new_n650), .ZN(new_n928));
  AOI22_X1  g0728(.A1(new_n925), .A2(new_n927), .B1(new_n928), .B2(new_n899), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n899), .ZN(new_n930));
  NOR3_X1   g0730(.A1(new_n924), .A2(new_n930), .A3(new_n926), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n910), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n736), .A2(KEYINPUT46), .A3(G116), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n934), .B(KEYINPUT107), .ZN(new_n935));
  INV_X1    g0735(.A(new_n730), .ZN(new_n936));
  AOI21_X1  g0736(.A(KEYINPUT46), .B1(new_n936), .B2(G116), .ZN(new_n937));
  OAI22_X1  g0737(.A1(new_n721), .A2(new_n739), .B1(new_n566), .B2(new_n717), .ZN(new_n938));
  AOI211_X1 g0738(.A(new_n937), .B(new_n938), .C1(G294), .C2(new_n785), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n714), .A2(new_n792), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n741), .A2(G97), .ZN(new_n941));
  INV_X1    g0741(.A(G317), .ZN(new_n942));
  OAI211_X1 g0742(.A(new_n396), .B(new_n941), .C1(new_n797), .C2(new_n942), .ZN(new_n943));
  AOI211_X1 g0743(.A(new_n940), .B(new_n943), .C1(G283), .C2(new_n725), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n935), .A2(new_n939), .A3(new_n944), .ZN(new_n945));
  OAI22_X1  g0745(.A1(new_n721), .A2(new_n787), .B1(new_n202), .B2(new_n717), .ZN(new_n946));
  INV_X1    g0746(.A(G137), .ZN(new_n947));
  OAI22_X1  g0747(.A1(new_n797), .A2(new_n947), .B1(new_n201), .B2(new_n730), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n252), .B1(new_n729), .B2(new_n255), .ZN(new_n949));
  NOR3_X1   g0749(.A1(new_n946), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  OAI22_X1  g0750(.A1(new_n726), .A2(new_n284), .B1(new_n723), .B2(new_n788), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(KEYINPUT108), .ZN(new_n952));
  OAI211_X1 g0752(.A(new_n950), .B(new_n952), .C1(new_n276), .C2(new_n714), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n951), .A2(KEYINPUT108), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n945), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n955), .B(KEYINPUT47), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n956), .A2(new_n707), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n755), .B1(new_n654), .B2(new_n583), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n759), .A2(new_n239), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n801), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  OAI211_X1 g0760(.A(new_n957), .B(new_n960), .C1(new_n766), .C2(new_n920), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n933), .A2(new_n961), .ZN(G387));
  XNOR2_X1  g0762(.A(new_n893), .B(new_n894), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n963), .B1(new_n695), .B2(new_n696), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n695), .A2(new_n963), .A3(new_n696), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n965), .A2(new_n655), .A3(new_n966), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n649), .A2(new_n766), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n409), .A2(new_n410), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(new_n284), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n970), .B(KEYINPUT50), .Z(new_n971));
  INV_X1    g0771(.A(KEYINPUT110), .ZN(new_n972));
  AND2_X1   g0772(.A1(new_n657), .A2(KEYINPUT109), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n657), .A2(KEYINPUT109), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n265), .B1(new_n202), .B2(new_n255), .ZN(new_n975));
  NOR3_X1   g0775(.A1(new_n973), .A2(new_n974), .A3(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n971), .B1(new_n972), .B2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(new_n976), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n978), .A2(KEYINPUT110), .ZN(new_n979));
  OAI221_X1 g0779(.A(new_n759), .B1(new_n265), .B2(new_n236), .C1(new_n977), .C2(new_n979), .ZN(new_n980));
  OAI221_X1 g0780(.A(new_n980), .B1(G107), .B2(new_n212), .C1(new_n657), .C2(new_n756), .ZN(new_n981));
  INV_X1    g0781(.A(new_n755), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(new_n702), .ZN(new_n984));
  AOI22_X1  g0784(.A1(new_n785), .A2(G311), .B1(G322), .B2(new_n744), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n985), .B(KEYINPUT111), .ZN(new_n986));
  OAI221_X1 g0786(.A(new_n986), .B1(new_n792), .B2(new_n726), .C1(new_n942), .C2(new_n714), .ZN(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(new_n988));
  OR2_X1    g0788(.A1(new_n988), .A2(KEYINPUT48), .ZN(new_n989));
  OAI22_X1  g0789(.A1(new_n717), .A2(new_n793), .B1(new_n730), .B2(new_n746), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n990), .B1(new_n988), .B2(KEYINPUT48), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n989), .A2(KEYINPUT49), .A3(new_n991), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n252), .B1(new_n710), .B2(G326), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n992), .B(new_n993), .C1(new_n434), .C2(new_n729), .ZN(new_n994));
  AOI21_X1  g0794(.A(KEYINPUT49), .B1(new_n989), .B2(new_n991), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n717), .A2(new_n412), .ZN(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  OAI221_X1 g0797(.A(new_n997), .B1(new_n723), .B2(new_n279), .C1(new_n788), .C2(new_n721), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n730), .A2(new_n255), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n999), .B1(G150), .B2(new_n710), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n1000), .A2(new_n252), .A3(new_n941), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n1001), .B1(G68), .B2(new_n725), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(new_n284), .B2(new_n714), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n994), .A2(new_n995), .B1(new_n998), .B2(new_n1003), .ZN(new_n1004));
  AOI211_X1 g0804(.A(new_n968), .B(new_n984), .C1(new_n1004), .C2(new_n707), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1005), .B1(new_n895), .B2(new_n701), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n967), .A2(new_n1006), .ZN(G393));
  NAND2_X1  g0807(.A1(new_n907), .A2(new_n701), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n982), .B1(new_n227), .B2(new_n212), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n760), .A2(new_n246), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n702), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n717), .A2(new_n255), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n396), .B1(new_n741), .B2(G87), .ZN(new_n1013));
  OAI221_X1 g0813(.A(new_n1013), .B1(new_n202), .B2(new_n730), .C1(new_n797), .C2(new_n787), .ZN(new_n1014));
  AOI211_X1 g0814(.A(new_n1012), .B(new_n1014), .C1(G50), .C2(new_n785), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n714), .A2(new_n788), .B1(new_n721), .B2(new_n276), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1016), .B(KEYINPUT51), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n725), .A2(new_n969), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1015), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n710), .A2(G322), .B1(new_n936), .B2(G283), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n1020), .B(new_n396), .C1(new_n566), .C2(new_n729), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT112), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(new_n785), .A2(G303), .B1(G116), .B2(new_n718), .ZN(new_n1023));
  OAI211_X1 g0823(.A(new_n1022), .B(new_n1023), .C1(new_n746), .C2(new_n726), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n714), .A2(new_n739), .B1(new_n721), .B2(new_n942), .ZN(new_n1025));
  XOR2_X1   g0825(.A(new_n1025), .B(KEYINPUT52), .Z(new_n1026));
  OAI21_X1  g0826(.A(new_n1019), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1011), .B1(new_n1027), .B2(new_n707), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(new_n899), .B2(new_n766), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1008), .A2(new_n1029), .ZN(new_n1030));
  OR2_X1    g0830(.A1(new_n964), .A2(new_n907), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n656), .B1(new_n964), .B2(new_n907), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1030), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n1033), .ZN(G390));
  AOI21_X1  g0834(.A(new_n775), .B1(new_n816), .B2(new_n817), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n690), .A2(new_n691), .A3(new_n1035), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n673), .A2(new_n674), .A3(new_n774), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1037), .A2(new_n771), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n865), .B1(new_n688), .B2(new_n775), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1036), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n1035), .B(G330), .C1(new_n686), .C2(new_n687), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n1041), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n690), .A2(new_n691), .A3(new_n776), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1042), .B1(new_n1043), .B2(new_n865), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1040), .B1(new_n1044), .B2(new_n864), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n688), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT113), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1046), .A2(new_n1047), .A3(new_n433), .ZN(new_n1048));
  OAI21_X1  g0848(.A(KEYINPUT113), .B1(new_n603), .B2(new_n688), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  AND3_X1   g0850(.A1(new_n1050), .A2(new_n885), .A3(new_n602), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1045), .A2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1037), .A2(new_n771), .A3(new_n818), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n875), .B1(new_n835), .B2(new_n844), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n873), .A2(new_n874), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n864), .A2(new_n865), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1056), .B1(new_n1057), .B2(new_n875), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1055), .A2(new_n1036), .A3(new_n1058), .ZN(new_n1059));
  AND2_X1   g0859(.A1(new_n1055), .A2(new_n1058), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1059), .B1(new_n1060), .B2(new_n1041), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n656), .B1(new_n1052), .B2(new_n1061), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1062), .B1(new_n1052), .B2(new_n1061), .ZN(new_n1063));
  OAI211_X1 g0863(.A(new_n701), .B(new_n1059), .C1(new_n1060), .C2(new_n1041), .ZN(new_n1064));
  INV_X1    g0864(.A(KEYINPUT114), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1064), .B(new_n1065), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n802), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n702), .B1(new_n351), .B2(new_n1067), .ZN(new_n1068));
  XOR2_X1   g0868(.A(new_n1068), .B(KEYINPUT115), .Z(new_n1069));
  OAI221_X1 g0869(.A(new_n396), .B1(new_n202), .B2(new_n729), .C1(new_n797), .C2(new_n746), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(new_n725), .B2(G97), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n723), .A2(new_n566), .ZN(new_n1072));
  AOI211_X1 g0872(.A(new_n1012), .B(new_n1072), .C1(G283), .C2(new_n744), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n736), .A2(G87), .B1(G116), .B2(new_n737), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1071), .A2(new_n1073), .A3(new_n1074), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n730), .A2(new_n276), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT53), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n1076), .A2(new_n1077), .B1(new_n788), .B2(new_n717), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1078), .B1(G137), .B2(new_n785), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n729), .A2(new_n284), .ZN(new_n1080));
  AOI211_X1 g0880(.A(new_n396), .B(new_n1080), .C1(G125), .C2(new_n710), .ZN(new_n1081));
  XOR2_X1   g0881(.A(KEYINPUT54), .B(G143), .Z(new_n1082));
  AOI22_X1  g0882(.A1(new_n725), .A2(new_n1082), .B1(new_n737), .B2(G132), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n744), .A2(G128), .B1(new_n1077), .B2(new_n1076), .ZN(new_n1084));
  NAND4_X1  g0884(.A1(new_n1079), .A2(new_n1081), .A3(new_n1083), .A4(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1075), .A2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1069), .B1(new_n1086), .B2(new_n707), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1056), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1087), .B1(new_n1088), .B2(new_n752), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1063), .A2(new_n1066), .A3(new_n1089), .ZN(G378));
  NAND3_X1  g0890(.A1(new_n850), .A2(G330), .A3(new_n857), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n299), .A2(new_n392), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n296), .A2(new_n636), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1092), .B(new_n1093), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1095), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(new_n1094), .B(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(KEYINPUT119), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  AND3_X1   g0899(.A1(new_n879), .A2(new_n883), .A3(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1099), .B1(new_n879), .B2(new_n883), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1091), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1045), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1051), .B1(new_n1061), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1099), .ZN(new_n1105));
  NOR3_X1   g0905(.A1(new_n870), .A2(new_n878), .A3(KEYINPUT102), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n881), .B1(new_n880), .B2(new_n882), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1105), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  AND3_X1   g0908(.A1(new_n850), .A2(G330), .A3(new_n857), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n879), .A2(new_n883), .A3(new_n1099), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1108), .A2(new_n1109), .A3(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1102), .A2(new_n1104), .A3(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(KEYINPUT57), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND4_X1  g0914(.A1(new_n1102), .A2(new_n1111), .A3(new_n1104), .A4(KEYINPUT57), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1114), .A2(new_n655), .A3(new_n1115), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1102), .A2(new_n701), .A3(new_n1111), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1097), .A2(new_n751), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n702), .B1(G50), .B2(new_n1067), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n721), .A2(new_n434), .B1(new_n202), .B2(new_n717), .ZN(new_n1120));
  XNOR2_X1  g0920(.A(new_n1120), .B(KEYINPUT116), .ZN(new_n1121));
  NOR3_X1   g0921(.A1(new_n999), .A2(G41), .A3(new_n252), .ZN(new_n1122));
  OAI221_X1 g0922(.A(new_n1122), .B1(new_n201), .B2(new_n729), .C1(new_n793), .C2(new_n797), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n726), .A2(new_n412), .B1(new_n566), .B2(new_n714), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n723), .A2(new_n227), .ZN(new_n1125));
  NOR4_X1   g0925(.A1(new_n1121), .A2(new_n1123), .A3(new_n1124), .A4(new_n1125), .ZN(new_n1126));
  OR2_X1    g0926(.A1(new_n1126), .A2(KEYINPUT58), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(new_n725), .A2(G137), .B1(new_n737), .B2(G128), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n785), .A2(G132), .B1(G150), .B2(new_n718), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(new_n744), .A2(G125), .B1(new_n936), .B2(new_n1082), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1128), .A2(new_n1129), .A3(new_n1130), .ZN(new_n1131));
  OR2_X1    g0931(.A1(new_n1131), .A2(KEYINPUT59), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1131), .A2(KEYINPUT59), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n249), .B(new_n264), .C1(new_n729), .C2(new_n788), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(KEYINPUT117), .B(G124), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1134), .B1(new_n710), .B2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1132), .A2(new_n1133), .A3(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1126), .A2(KEYINPUT58), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n284), .B1(new_n358), .B2(G41), .ZN(new_n1139));
  NAND4_X1  g0939(.A1(new_n1127), .A2(new_n1137), .A3(new_n1138), .A4(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1119), .B1(new_n1140), .B2(new_n707), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1118), .A2(new_n1141), .ZN(new_n1142));
  XNOR2_X1  g0942(.A(new_n1142), .B(KEYINPUT118), .ZN(new_n1143));
  AND2_X1   g0943(.A1(new_n1117), .A2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1116), .A2(new_n1144), .ZN(G375));
  XOR2_X1   g0945(.A(new_n700), .B(KEYINPUT120), .Z(new_n1146));
  NAND2_X1  g0946(.A1(new_n1045), .A2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n801), .B1(new_n202), .B2(new_n802), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n710), .A2(G128), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n1149), .B(new_n252), .C1(new_n201), .C2(new_n729), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n726), .A2(new_n276), .B1(new_n947), .B2(new_n714), .ZN(new_n1151));
  AOI211_X1 g0951(.A(new_n1150), .B(new_n1151), .C1(G159), .C2(new_n736), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n785), .A2(new_n1082), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n744), .A2(G132), .B1(G50), .B2(new_n718), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1152), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1155));
  OAI221_X1 g0955(.A(new_n997), .B1(new_n723), .B2(new_n434), .C1(new_n746), .C2(new_n721), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(new_n736), .A2(G97), .B1(G283), .B2(new_n737), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n396), .B1(new_n729), .B2(new_n255), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1158), .B1(G303), .B2(new_n710), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n1157), .B(new_n1159), .C1(new_n566), .C2(new_n726), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1155), .B1(new_n1156), .B2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(KEYINPUT121), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(new_n707), .ZN(new_n1165));
  OAI221_X1 g0965(.A(new_n1148), .B1(new_n1163), .B2(new_n1165), .C1(new_n818), .C2(new_n752), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1147), .A2(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(KEYINPUT122), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1147), .A2(KEYINPUT122), .A3(new_n1166), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  OR2_X1    g0971(.A1(new_n1045), .A2(new_n1051), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n909), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1172), .A2(new_n1173), .A3(new_n1052), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1171), .A2(new_n1174), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(new_n1175), .B(KEYINPUT123), .ZN(G381));
  NAND4_X1  g0976(.A1(new_n967), .A2(new_n706), .A3(new_n767), .A4(new_n1006), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1033), .A2(new_n805), .ZN(new_n1178));
  NOR4_X1   g0978(.A1(G381), .A2(G387), .A3(new_n1177), .A4(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(G378), .ZN(new_n1180));
  OR2_X1    g0980(.A1(G375), .A2(KEYINPUT124), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(G375), .A2(KEYINPUT124), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1179), .A2(new_n1180), .A3(new_n1181), .A4(new_n1182), .ZN(G407));
  NAND3_X1  g0983(.A1(new_n1181), .A2(new_n1180), .A3(new_n1182), .ZN(new_n1184));
  OAI211_X1 g0984(.A(G407), .B(G213), .C1(G343), .C2(new_n1184), .ZN(G409));
  INV_X1    g0985(.A(G343), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1186), .A2(G213), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1052), .A2(KEYINPUT60), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1189), .A2(new_n1172), .ZN(new_n1190));
  INV_X1    g0990(.A(KEYINPUT60), .ZN(new_n1191));
  NOR3_X1   g0991(.A1(new_n1045), .A2(new_n1051), .A3(new_n1191), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n1192), .A2(new_n656), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1190), .A2(new_n1193), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1194), .A2(new_n1171), .A3(G384), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(G384), .B1(new_n1194), .B2(new_n1171), .ZN(new_n1197));
  OAI211_X1 g0997(.A(G2897), .B(new_n1188), .C1(new_n1196), .C2(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1197), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1188), .A2(G2897), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1199), .A2(new_n1195), .A3(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1198), .A2(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1116), .A2(G378), .A3(new_n1144), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1102), .A2(new_n1111), .A3(new_n1146), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n1142), .B(new_n1205), .C1(new_n1112), .C2(new_n909), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1180), .A2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1204), .A2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1208), .A2(new_n1187), .ZN(new_n1209));
  AOI21_X1  g1009(.A(KEYINPUT61), .B1(new_n1203), .B2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT63), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1199), .A2(new_n1195), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1211), .B1(new_n1209), .B2(new_n1212), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(G390), .A2(new_n933), .A3(new_n961), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(G387), .A2(new_n1033), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(G393), .A2(G396), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1216), .A2(new_n1177), .ZN(new_n1217));
  AND4_X1   g1017(.A1(KEYINPUT125), .A2(new_n1214), .A3(new_n1215), .A4(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT125), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1219), .B1(G387), .B2(new_n1033), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n1220), .A2(new_n1217), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1221));
  OR2_X1    g1021(.A1(new_n1218), .A2(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1188), .B1(new_n1204), .B2(new_n1207), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1223), .A2(KEYINPUT63), .A3(new_n1224), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n1210), .A2(new_n1213), .A3(new_n1222), .A4(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT62), .ZN(new_n1227));
  AND3_X1   g1027(.A1(new_n1223), .A2(new_n1227), .A3(new_n1224), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT61), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1229), .B1(new_n1223), .B2(new_n1202), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1227), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1231));
  NOR3_X1   g1031(.A1(new_n1228), .A2(new_n1230), .A3(new_n1231), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1226), .B1(new_n1232), .B2(new_n1222), .ZN(G405));
  AND3_X1   g1033(.A1(new_n1116), .A2(G378), .A3(new_n1144), .ZN(new_n1234));
  AOI21_X1  g1034(.A(G378), .B1(new_n1116), .B2(new_n1144), .ZN(new_n1235));
  NOR3_X1   g1035(.A1(new_n1234), .A2(new_n1235), .A3(new_n1224), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(G375), .A2(new_n1180), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1212), .B1(new_n1237), .B2(new_n1204), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1222), .B1(new_n1236), .B2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT127), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  OAI211_X1 g1041(.A(new_n1222), .B(KEYINPUT127), .C1(new_n1236), .C2(new_n1238), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n1218), .A2(new_n1221), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1224), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1237), .A2(new_n1204), .A3(new_n1212), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1243), .A2(new_n1244), .A3(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT126), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1243), .A2(new_n1244), .A3(new_n1245), .A4(KEYINPUT126), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(new_n1241), .A2(new_n1242), .B1(new_n1248), .B2(new_n1249), .ZN(G402));
endmodule


