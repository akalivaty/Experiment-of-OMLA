//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 0 0 0 1 0 1 1 1 0 1 1 1 1 0 0 1 0 1 0 1 1 0 0 1 0 1 0 0 0 0 1 1 0 0 1 1 0 0 0 1 1 0 1 0 1 0 0 1 1 0 1 0 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:51 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n558,
    new_n559, new_n560, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n571, new_n572, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n611,
    new_n613, new_n614, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1175, new_n1176, new_n1177;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g018(.A(KEYINPUT65), .B(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(G234));
  NAND2_X1  g024(.A1(new_n447), .A2(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT67), .Z(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  OAI21_X1  g039(.A(KEYINPUT68), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT68), .ZN(new_n469));
  NAND2_X1  g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n465), .A2(new_n471), .A3(G125), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  XOR2_X1   g048(.A(new_n473), .B(KEYINPUT69), .Z(new_n474));
  AOI21_X1  g049(.A(new_n462), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(new_n476));
  AOI21_X1  g051(.A(G2105), .B1(new_n468), .B2(new_n470), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n477), .A2(KEYINPUT70), .A3(G137), .ZN(new_n478));
  OAI211_X1 g053(.A(G137), .B(new_n462), .C1(new_n463), .C2(new_n464), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT70), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n467), .A2(G2105), .ZN(new_n482));
  AOI22_X1  g057(.A1(new_n478), .A2(new_n481), .B1(G101), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n476), .A2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G160));
  NAND2_X1  g060(.A1(new_n468), .A2(new_n470), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(new_n462), .ZN(new_n487));
  INV_X1    g062(.A(G136), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n462), .A2(G112), .ZN(new_n489));
  OAI21_X1  g064(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n490));
  OAI22_X1  g065(.A1(new_n487), .A2(new_n488), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n463), .A2(new_n464), .ZN(new_n492));
  OAI21_X1  g067(.A(KEYINPUT71), .B1(new_n492), .B2(new_n462), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT71), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n486), .A2(new_n494), .A3(G2105), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n491), .B1(G124), .B2(new_n496), .ZN(new_n497));
  XNOR2_X1  g072(.A(new_n497), .B(KEYINPUT72), .ZN(G162));
  OAI21_X1  g073(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n499));
  INV_X1    g074(.A(G114), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n499), .B1(new_n500), .B2(G2105), .ZN(new_n501));
  AND2_X1   g076(.A1(G126), .A2(G2105), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n502), .B1(new_n463), .B2(new_n464), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT73), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n486), .A2(KEYINPUT73), .A3(new_n502), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n501), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(G138), .ZN(new_n508));
  NOR3_X1   g083(.A1(new_n508), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n465), .A2(new_n471), .A3(new_n509), .ZN(new_n510));
  OAI211_X1 g085(.A(G138), .B(new_n462), .C1(new_n463), .C2(new_n464), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(KEYINPUT4), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n507), .A2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(new_n514), .ZN(G164));
  INV_X1    g090(.A(G50), .ZN(new_n516));
  AND2_X1   g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  NOR2_X1   g092(.A1(KEYINPUT6), .A2(G651), .ZN(new_n518));
  OR2_X1    g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G543), .ZN(new_n520));
  XNOR2_X1  g095(.A(KEYINPUT5), .B(G543), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(G88), .ZN(new_n523));
  OAI22_X1  g098(.A1(new_n516), .A2(new_n520), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n521), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n525));
  INV_X1    g100(.A(G651), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n524), .A2(new_n527), .ZN(G166));
  AND2_X1   g103(.A1(new_n519), .A2(G89), .ZN(new_n529));
  AND2_X1   g104(.A1(G63), .A2(G651), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n521), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n517), .A2(new_n518), .ZN(new_n532));
  INV_X1    g107(.A(G543), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(KEYINPUT7), .ZN(new_n536));
  OR2_X1    g111(.A1(new_n535), .A2(KEYINPUT7), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n534), .A2(G51), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n531), .A2(KEYINPUT74), .A3(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(new_n539), .ZN(new_n540));
  AOI21_X1  g115(.A(KEYINPUT74), .B1(new_n531), .B2(new_n538), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n540), .A2(new_n541), .ZN(G286));
  INV_X1    g117(.A(G286), .ZN(G168));
  INV_X1    g118(.A(G52), .ZN(new_n544));
  INV_X1    g119(.A(G90), .ZN(new_n545));
  OAI22_X1  g120(.A1(new_n544), .A2(new_n520), .B1(new_n522), .B2(new_n545), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n521), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n547), .A2(new_n526), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n546), .A2(new_n548), .ZN(G171));
  INV_X1    g124(.A(G43), .ZN(new_n550));
  INV_X1    g125(.A(G81), .ZN(new_n551));
  OAI22_X1  g126(.A1(new_n550), .A2(new_n520), .B1(new_n522), .B2(new_n551), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n521), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n553), .A2(new_n526), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  NAND4_X1  g131(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT75), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND4_X1  g135(.A1(G319), .A2(G483), .A3(G661), .A4(new_n560), .ZN(G188));
  NAND2_X1  g136(.A1(new_n534), .A2(G53), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT9), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n562), .B(new_n563), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n521), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n565));
  INV_X1    g140(.A(G91), .ZN(new_n566));
  OAI22_X1  g141(.A1(new_n526), .A2(new_n565), .B1(new_n522), .B2(new_n566), .ZN(new_n567));
  NOR2_X1   g142(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(new_n568), .ZN(G299));
  INV_X1    g144(.A(G171), .ZN(G301));
  OR2_X1    g145(.A1(G166), .A2(KEYINPUT76), .ZN(new_n571));
  NAND2_X1  g146(.A1(G166), .A2(KEYINPUT76), .ZN(new_n572));
  AND2_X1   g147(.A1(new_n571), .A2(new_n572), .ZN(G303));
  INV_X1    g148(.A(G49), .ZN(new_n574));
  OR3_X1    g149(.A1(new_n520), .A2(KEYINPUT77), .A3(new_n574), .ZN(new_n575));
  OAI21_X1  g150(.A(KEYINPUT77), .B1(new_n520), .B2(new_n574), .ZN(new_n576));
  INV_X1    g151(.A(new_n522), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n577), .A2(G87), .ZN(new_n578));
  OAI21_X1  g153(.A(G651), .B1(new_n521), .B2(G74), .ZN(new_n579));
  NAND4_X1  g154(.A1(new_n575), .A2(new_n576), .A3(new_n578), .A4(new_n579), .ZN(G288));
  AOI22_X1  g155(.A1(new_n521), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n581), .A2(new_n526), .ZN(new_n582));
  INV_X1    g157(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n577), .A2(G86), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n534), .A2(G48), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(G305));
  INV_X1    g161(.A(G85), .ZN(new_n587));
  XOR2_X1   g162(.A(KEYINPUT78), .B(G47), .Z(new_n588));
  OAI22_X1  g163(.A1(new_n587), .A2(new_n522), .B1(new_n520), .B2(new_n588), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n521), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n590), .A2(new_n526), .ZN(new_n591));
  OR3_X1    g166(.A1(new_n589), .A2(KEYINPUT79), .A3(new_n591), .ZN(new_n592));
  OAI21_X1  g167(.A(KEYINPUT79), .B1(new_n589), .B2(new_n591), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(G290));
  NAND2_X1  g169(.A1(G301), .A2(G868), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n521), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n596));
  INV_X1    g171(.A(G54), .ZN(new_n597));
  OAI22_X1  g172(.A1(new_n526), .A2(new_n596), .B1(new_n520), .B2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT80), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  OAI221_X1 g175(.A(KEYINPUT80), .B1(new_n520), .B2(new_n597), .C1(new_n526), .C2(new_n596), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT10), .ZN(new_n602));
  INV_X1    g177(.A(G92), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n522), .B2(new_n603), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n577), .A2(KEYINPUT10), .A3(G92), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n600), .A2(new_n601), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n595), .B1(new_n606), .B2(G868), .ZN(G284));
  OAI21_X1  g182(.A(new_n595), .B1(new_n606), .B2(G868), .ZN(G321));
  MUX2_X1   g183(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g184(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g185(.A(G559), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n606), .B1(new_n611), .B2(G860), .ZN(G148));
  NAND2_X1  g187(.A1(new_n606), .A2(new_n611), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n613), .A2(G868), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n614), .B1(G868), .B2(new_n555), .ZN(G323));
  XNOR2_X1  g190(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g191(.A1(new_n465), .A2(new_n471), .A3(new_n482), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT12), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT13), .ZN(new_n619));
  INV_X1    g194(.A(G2100), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(KEYINPUT81), .Z(new_n622));
  INV_X1    g197(.A(G135), .ZN(new_n623));
  NOR2_X1   g198(.A1(new_n462), .A2(G111), .ZN(new_n624));
  OAI21_X1  g199(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n625));
  OAI22_X1  g200(.A1(new_n487), .A2(new_n623), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  AOI21_X1  g201(.A(new_n626), .B1(G123), .B2(new_n496), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(KEYINPUT82), .Z(new_n628));
  INV_X1    g203(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n629), .A2(G2096), .ZN(new_n630));
  OR2_X1    g205(.A1(new_n629), .A2(G2096), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n619), .A2(new_n620), .ZN(new_n632));
  NAND4_X1  g207(.A1(new_n622), .A2(new_n630), .A3(new_n631), .A4(new_n632), .ZN(G156));
  XOR2_X1   g208(.A(G2451), .B(G2454), .Z(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT16), .ZN(new_n635));
  XNOR2_X1  g210(.A(G1341), .B(G1348), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  INV_X1    g212(.A(KEYINPUT14), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2427), .B(G2438), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2430), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT15), .B(G2435), .ZN(new_n641));
  AOI21_X1  g216(.A(new_n638), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  OAI21_X1  g217(.A(new_n642), .B1(new_n641), .B2(new_n640), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n637), .B(new_n643), .Z(new_n644));
  XNOR2_X1  g219(.A(G2443), .B(G2446), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n644), .A2(new_n645), .ZN(new_n647));
  AND3_X1   g222(.A1(new_n646), .A2(G14), .A3(new_n647), .ZN(G401));
  XNOR2_X1  g223(.A(G2072), .B(G2078), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT17), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2067), .B(G2678), .ZN(new_n651));
  XOR2_X1   g226(.A(G2084), .B(G2090), .Z(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  NOR3_X1   g228(.A1(new_n650), .A2(new_n651), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT83), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n650), .A2(new_n651), .ZN(new_n656));
  OAI211_X1 g231(.A(new_n656), .B(new_n653), .C1(new_n649), .C2(new_n651), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n652), .A2(new_n649), .A3(new_n651), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(KEYINPUT18), .Z(new_n659));
  NAND3_X1  g234(.A1(new_n655), .A2(new_n657), .A3(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(G2096), .B(G2100), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(G227));
  XOR2_X1   g237(.A(KEYINPUT84), .B(KEYINPUT19), .Z(new_n663));
  XNOR2_X1  g238(.A(G1971), .B(G1976), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1956), .B(G2474), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1961), .B(G1966), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT20), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n666), .A2(new_n667), .ZN(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n665), .A2(new_n672), .ZN(new_n673));
  OR2_X1    g248(.A1(new_n672), .A2(new_n668), .ZN(new_n674));
  OAI211_X1 g249(.A(new_n670), .B(new_n673), .C1(new_n665), .C2(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n675), .B(KEYINPUT85), .Z(new_n676));
  XNOR2_X1  g251(.A(G1991), .B(G1996), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1981), .B(G1986), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  OR2_X1    g256(.A1(new_n676), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n676), .A2(new_n681), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n682), .A2(new_n683), .ZN(G229));
  INV_X1    g259(.A(G29), .ZN(new_n685));
  AND2_X1   g260(.A1(new_n685), .A2(G32), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n496), .A2(G129), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT92), .ZN(new_n688));
  NAND3_X1  g263(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT93), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT26), .ZN(new_n691));
  AOI22_X1  g266(.A1(new_n477), .A2(G141), .B1(G105), .B2(new_n482), .ZN(new_n692));
  AND2_X1   g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n688), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT94), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n686), .B1(new_n695), .B2(G29), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT27), .B(G1996), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT95), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n696), .B(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(KEYINPUT24), .ZN(new_n700));
  INV_X1    g275(.A(G34), .ZN(new_n701));
  AOI21_X1  g276(.A(G29), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(new_n700), .B2(new_n701), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n704), .B1(new_n484), .B2(G29), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(G2084), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n707), .B(KEYINPUT90), .Z(new_n708));
  NOR2_X1   g283(.A1(G29), .A2(G33), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT89), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(KEYINPUT25), .Z(new_n712));
  INV_X1    g287(.A(G139), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n712), .B1(new_n713), .B2(new_n487), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n465), .A2(new_n471), .A3(G127), .ZN(new_n715));
  NAND2_X1  g290(.A1(G115), .A2(G2104), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n462), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n714), .A2(new_n717), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n710), .B1(new_n718), .B2(G29), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G2072), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(KEYINPUT91), .Z(new_n721));
  XOR2_X1   g296(.A(KEYINPUT31), .B(G11), .Z(new_n722));
  INV_X1    g297(.A(KEYINPUT30), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n685), .B1(new_n723), .B2(G28), .ZN(new_n724));
  INV_X1    g299(.A(new_n724), .ZN(new_n725));
  OR2_X1    g300(.A1(new_n725), .A2(KEYINPUT96), .ZN(new_n726));
  AOI22_X1  g301(.A1(new_n725), .A2(KEYINPUT96), .B1(new_n723), .B2(G28), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n722), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(new_n629), .B2(new_n685), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT97), .ZN(new_n730));
  AND4_X1   g305(.A1(new_n699), .A2(new_n708), .A3(new_n721), .A4(new_n730), .ZN(new_n731));
  NOR2_X1   g306(.A1(G16), .A2(G19), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(new_n555), .B2(G16), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT88), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(G1341), .Z(new_n735));
  INV_X1    g310(.A(G16), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n736), .A2(G21), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(G168), .B2(new_n736), .ZN(new_n738));
  OR2_X1    g313(.A1(new_n738), .A2(G1966), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n739), .A2(KEYINPUT98), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n736), .A2(G4), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(new_n606), .B2(new_n736), .ZN(new_n742));
  OR2_X1    g317(.A1(new_n742), .A2(G1348), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n742), .A2(G1348), .ZN(new_n744));
  NAND4_X1  g319(.A1(new_n735), .A2(new_n740), .A3(new_n743), .A4(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n738), .A2(G1966), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n685), .A2(G26), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(KEYINPUT28), .Z(new_n748));
  AND2_X1   g323(.A1(new_n496), .A2(G128), .ZN(new_n749));
  OAI21_X1  g324(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n750));
  INV_X1    g325(.A(G116), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n750), .B1(new_n751), .B2(G2105), .ZN(new_n752));
  INV_X1    g327(.A(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(G140), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n753), .B1(new_n487), .B2(new_n754), .ZN(new_n755));
  OR2_X1    g330(.A1(new_n749), .A2(new_n755), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n748), .B1(new_n756), .B2(G29), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(G2067), .ZN(new_n758));
  OAI211_X1 g333(.A(new_n746), .B(new_n758), .C1(G2072), .C2(new_n719), .ZN(new_n759));
  NOR2_X1   g334(.A1(G164), .A2(new_n685), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(G27), .B2(new_n685), .ZN(new_n761));
  INV_X1    g336(.A(G2078), .ZN(new_n762));
  OR2_X1    g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g338(.A1(G5), .A2(G16), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(G171), .B2(G16), .ZN(new_n765));
  OR2_X1    g340(.A1(new_n765), .A2(G1961), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n761), .A2(new_n762), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n765), .A2(G1961), .ZN(new_n768));
  NAND4_X1  g343(.A1(new_n763), .A2(new_n766), .A3(new_n767), .A4(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n736), .A2(G20), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT99), .Z(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT23), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(G299), .B2(G16), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(G1956), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(G2084), .B2(new_n706), .ZN(new_n775));
  NOR4_X1   g350(.A1(new_n745), .A2(new_n759), .A3(new_n769), .A4(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(G162), .A2(G29), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G29), .B2(G35), .ZN(new_n778));
  XOR2_X1   g353(.A(KEYINPUT29), .B(G2090), .Z(new_n779));
  OAI22_X1  g354(.A1(new_n739), .A2(KEYINPUT98), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(new_n778), .B2(new_n779), .ZN(new_n781));
  AND3_X1   g356(.A1(new_n731), .A2(new_n776), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n736), .A2(G23), .ZN(new_n783));
  INV_X1    g358(.A(G288), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n783), .B1(new_n784), .B2(new_n736), .ZN(new_n785));
  XNOR2_X1  g360(.A(KEYINPUT33), .B(G1976), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n736), .A2(G22), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G166), .B2(new_n736), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(G1971), .Z(new_n790));
  MUX2_X1   g365(.A(G6), .B(G305), .S(G16), .Z(new_n791));
  XOR2_X1   g366(.A(KEYINPUT32), .B(G1981), .Z(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n787), .A2(new_n790), .A3(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(KEYINPUT34), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  AND2_X1   g371(.A1(new_n736), .A2(G24), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(G290), .B2(G16), .ZN(new_n798));
  INV_X1    g373(.A(G1986), .ZN(new_n799));
  AND2_X1   g374(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NOR2_X1   g375(.A1(G25), .A2(G29), .ZN(new_n801));
  AND2_X1   g376(.A1(new_n496), .A2(G119), .ZN(new_n802));
  INV_X1    g377(.A(G131), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n462), .A2(G107), .ZN(new_n804));
  OAI21_X1  g379(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n805));
  OAI22_X1  g380(.A1(new_n487), .A2(new_n803), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n802), .A2(new_n806), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n801), .B1(new_n807), .B2(G29), .ZN(new_n808));
  XNOR2_X1  g383(.A(KEYINPUT35), .B(G1991), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT86), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n808), .B(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n798), .A2(new_n799), .ZN(new_n812));
  NOR4_X1   g387(.A1(new_n800), .A2(new_n811), .A3(new_n812), .A4(KEYINPUT87), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n796), .A2(new_n813), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT36), .ZN(new_n815));
  INV_X1    g390(.A(KEYINPUT100), .ZN(new_n816));
  AND3_X1   g391(.A1(new_n782), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n816), .B1(new_n782), .B2(new_n815), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n817), .A2(new_n818), .ZN(G311));
  NAND2_X1  g394(.A1(new_n782), .A2(new_n815), .ZN(G150));
  AOI22_X1  g395(.A1(new_n521), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n821));
  OR2_X1    g396(.A1(new_n821), .A2(new_n526), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n577), .A2(G93), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n534), .A2(G55), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n822), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT101), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND4_X1  g402(.A1(new_n822), .A2(new_n823), .A3(KEYINPUT101), .A4(new_n824), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n827), .A2(new_n555), .A3(new_n828), .ZN(new_n829));
  OAI211_X1 g404(.A(new_n825), .B(new_n826), .C1(new_n554), .C2(new_n552), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT38), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n606), .A2(G559), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n832), .B(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(KEYINPUT39), .ZN(new_n835));
  AOI21_X1  g410(.A(G860), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n836), .B1(new_n835), .B2(new_n834), .ZN(new_n837));
  XOR2_X1   g412(.A(new_n837), .B(KEYINPUT102), .Z(new_n838));
  NAND2_X1  g413(.A1(new_n825), .A2(G860), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n839), .B(KEYINPUT37), .Z(new_n840));
  NAND2_X1  g415(.A1(new_n838), .A2(new_n840), .ZN(G145));
  XNOR2_X1  g416(.A(new_n628), .B(new_n484), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(G162), .ZN(new_n843));
  INV_X1    g418(.A(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT103), .ZN(new_n845));
  AND3_X1   g420(.A1(new_n510), .A2(new_n512), .A3(new_n845), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n845), .B1(new_n510), .B2(new_n512), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n507), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT104), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  OAI211_X1 g425(.A(KEYINPUT104), .B(new_n507), .C1(new_n846), .C2(new_n847), .ZN(new_n851));
  AND3_X1   g426(.A1(new_n850), .A2(new_n756), .A3(new_n851), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n756), .B1(new_n850), .B2(new_n851), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n694), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n850), .A2(new_n851), .ZN(new_n855));
  INV_X1    g430(.A(new_n756), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(new_n694), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n850), .A2(new_n756), .A3(new_n851), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n857), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n854), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n861), .A2(KEYINPUT94), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT94), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n854), .A2(new_n860), .A3(new_n863), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n862), .A2(new_n718), .A3(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(new_n718), .ZN(new_n866));
  AOI21_X1  g441(.A(KEYINPUT105), .B1(new_n861), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n807), .B(KEYINPUT106), .ZN(new_n869));
  XOR2_X1   g444(.A(new_n869), .B(new_n618), .Z(new_n870));
  NAND2_X1  g445(.A1(new_n496), .A2(G130), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n477), .A2(G142), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n462), .A2(G118), .ZN(new_n873));
  OAI21_X1  g448(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n874));
  OAI211_X1 g449(.A(new_n871), .B(new_n872), .C1(new_n873), .C2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n870), .B(new_n875), .ZN(new_n876));
  NAND4_X1  g451(.A1(new_n862), .A2(KEYINPUT105), .A3(new_n718), .A4(new_n864), .ZN(new_n877));
  AND3_X1   g452(.A1(new_n868), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n876), .B1(new_n868), .B2(new_n877), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n844), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n868), .A2(new_n877), .ZN(new_n881));
  INV_X1    g456(.A(new_n876), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n868), .A2(new_n876), .A3(new_n877), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n883), .A2(new_n843), .A3(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(G37), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n880), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g463(.A(G166), .ZN(new_n889));
  XNOR2_X1  g464(.A(G290), .B(new_n889), .ZN(new_n890));
  XOR2_X1   g465(.A(G288), .B(G305), .Z(new_n891));
  XNOR2_X1  g466(.A(new_n890), .B(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(KEYINPUT42), .ZN(new_n893));
  AND2_X1   g468(.A1(new_n829), .A2(new_n830), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(new_n613), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n600), .A2(new_n601), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n605), .A2(new_n604), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(G299), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n606), .A2(new_n568), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(KEYINPUT41), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT41), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n899), .A2(new_n903), .A3(new_n900), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n895), .A2(new_n905), .ZN(new_n906));
  OR2_X1    g481(.A1(new_n906), .A2(KEYINPUT107), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(KEYINPUT107), .ZN(new_n908));
  OAI211_X1 g483(.A(new_n907), .B(new_n908), .C1(new_n895), .C2(new_n901), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT108), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n893), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n909), .A2(new_n910), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NOR3_X1   g488(.A1(new_n909), .A2(new_n910), .A3(new_n893), .ZN(new_n914));
  OAI21_X1  g489(.A(G868), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(G868), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n825), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n915), .A2(new_n917), .ZN(G295));
  NAND2_X1  g493(.A1(new_n915), .A2(new_n917), .ZN(G331));
  INV_X1    g494(.A(KEYINPUT109), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n920), .B1(new_n540), .B2(new_n541), .ZN(new_n921));
  INV_X1    g496(.A(new_n541), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n922), .A2(KEYINPUT109), .A3(new_n539), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n921), .A2(new_n923), .A3(G171), .ZN(new_n924));
  NAND3_X1  g499(.A1(G286), .A2(KEYINPUT109), .A3(G301), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n894), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n894), .B1(new_n924), .B2(new_n925), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n905), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n924), .A2(new_n925), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n930), .A2(new_n831), .ZN(new_n931));
  NAND4_X1  g506(.A1(new_n931), .A2(new_n899), .A3(new_n900), .A4(new_n926), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n929), .A2(new_n932), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n933), .A2(new_n892), .ZN(new_n934));
  AOI21_X1  g509(.A(G37), .B1(new_n933), .B2(new_n892), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n934), .B1(new_n935), .B2(KEYINPUT110), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT110), .ZN(new_n937));
  INV_X1    g512(.A(new_n892), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n938), .B1(new_n929), .B2(new_n932), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n937), .B1(new_n939), .B2(G37), .ZN(new_n940));
  AOI21_X1  g515(.A(KEYINPUT43), .B1(new_n936), .B2(new_n940), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n886), .B1(new_n933), .B2(new_n892), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT111), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n904), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(new_n902), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n904), .A2(new_n943), .ZN(new_n946));
  OAI22_X1  g521(.A1(new_n945), .A2(new_n946), .B1(new_n927), .B2(new_n928), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n938), .B1(new_n947), .B2(new_n932), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT43), .ZN(new_n949));
  NOR3_X1   g524(.A1(new_n942), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  OAI21_X1  g525(.A(KEYINPUT44), .B1(new_n941), .B2(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n949), .B1(new_n936), .B2(new_n940), .ZN(new_n952));
  NOR3_X1   g527(.A1(new_n942), .A2(new_n948), .A3(KEYINPUT43), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n951), .B1(new_n954), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g530(.A(G1384), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n850), .A2(new_n956), .A3(new_n851), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT45), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n478), .A2(new_n481), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n482), .A2(G101), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(G40), .ZN(new_n962));
  NOR3_X1   g537(.A1(new_n961), .A2(new_n475), .A3(new_n962), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n957), .A2(new_n958), .A3(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT112), .ZN(new_n966));
  INV_X1    g541(.A(G1996), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n965), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  OAI21_X1  g543(.A(KEYINPUT112), .B1(new_n964), .B2(G1996), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(new_n695), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  XOR2_X1   g547(.A(new_n756), .B(G2067), .Z(new_n973));
  OAI21_X1  g548(.A(new_n973), .B1(new_n858), .B2(new_n967), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(new_n965), .ZN(new_n975));
  AND2_X1   g550(.A1(new_n972), .A2(new_n975), .ZN(new_n976));
  XOR2_X1   g551(.A(new_n807), .B(new_n810), .Z(new_n977));
  NAND2_X1  g552(.A1(new_n965), .A2(new_n977), .ZN(new_n978));
  NOR2_X1   g553(.A1(G290), .A2(G1986), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n799), .B1(new_n592), .B2(new_n593), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n965), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n976), .A2(new_n978), .A3(new_n981), .ZN(new_n982));
  XOR2_X1   g557(.A(new_n982), .B(KEYINPUT113), .Z(new_n983));
  NAND3_X1  g558(.A1(new_n571), .A2(G8), .A3(new_n572), .ZN(new_n984));
  XNOR2_X1  g559(.A(new_n984), .B(KEYINPUT55), .ZN(new_n985));
  INV_X1    g560(.A(new_n985), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n958), .A2(G1384), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n850), .A2(new_n851), .A3(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n476), .A2(G40), .A3(new_n483), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n514), .A2(new_n956), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n989), .B1(new_n958), .B2(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(G1971), .B1(new_n988), .B2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT114), .ZN(new_n993));
  AND2_X1   g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  AOI21_X1  g569(.A(KEYINPUT50), .B1(new_n848), .B2(new_n956), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n514), .A2(KEYINPUT50), .A3(new_n956), .ZN(new_n996));
  INV_X1    g571(.A(new_n996), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n963), .B1(new_n995), .B2(new_n997), .ZN(new_n998));
  OAI22_X1  g573(.A1(new_n992), .A2(new_n993), .B1(G2090), .B2(new_n998), .ZN(new_n999));
  OAI211_X1 g574(.A(new_n986), .B(G8), .C1(new_n994), .C2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n963), .A2(new_n956), .A3(new_n848), .ZN(new_n1002));
  AND2_X1   g577(.A1(new_n1002), .A2(G8), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n784), .A2(G1976), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(KEYINPUT52), .ZN(new_n1006));
  INV_X1    g581(.A(G1976), .ZN(new_n1007));
  AOI21_X1  g582(.A(KEYINPUT52), .B1(G288), .B2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1003), .A2(new_n1004), .A3(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(G86), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n585), .B1(new_n522), .B2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g586(.A(G1981), .B1(new_n1011), .B2(new_n582), .ZN(new_n1012));
  INV_X1    g587(.A(G1981), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n583), .A2(new_n584), .A3(new_n1013), .A4(new_n585), .ZN(new_n1014));
  AND3_X1   g589(.A1(new_n1012), .A2(new_n1014), .A3(KEYINPUT49), .ZN(new_n1015));
  AOI21_X1  g590(.A(KEYINPUT49), .B1(new_n1012), .B2(new_n1014), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  AND3_X1   g592(.A1(new_n1003), .A2(new_n1017), .A3(KEYINPUT115), .ZN(new_n1018));
  AOI21_X1  g593(.A(KEYINPUT115), .B1(new_n1003), .B2(new_n1017), .ZN(new_n1019));
  OAI211_X1 g594(.A(new_n1006), .B(new_n1009), .C1(new_n1018), .C2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1020), .ZN(new_n1021));
  OAI211_X1 g596(.A(new_n1007), .B(new_n784), .C1(new_n1018), .C2(new_n1019), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(new_n1014), .ZN(new_n1023));
  AOI22_X1  g598(.A1(new_n1001), .A2(new_n1021), .B1(new_n1023), .B2(new_n1003), .ZN(new_n1024));
  INV_X1    g599(.A(G1966), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT116), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1026), .B1(new_n514), .B2(new_n987), .ZN(new_n1027));
  INV_X1    g602(.A(new_n987), .ZN(new_n1028));
  AOI211_X1 g603(.A(KEYINPUT116), .B(new_n1028), .C1(new_n507), .C2(new_n513), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n963), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(KEYINPUT45), .B1(new_n848), .B2(new_n956), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1025), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n989), .A2(G2084), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1033), .B1(new_n995), .B2(new_n997), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1032), .A2(G168), .A3(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(G8), .ZN(new_n1036));
  AOI21_X1  g611(.A(G168), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1037));
  OAI21_X1  g612(.A(KEYINPUT51), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT122), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT51), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1035), .A2(new_n1040), .A3(G8), .ZN(new_n1041));
  AND3_X1   g616(.A1(new_n1038), .A2(new_n1039), .A3(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1039), .B1(new_n1038), .B2(new_n1041), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT54), .ZN(new_n1045));
  XNOR2_X1  g620(.A(KEYINPUT123), .B(G1961), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n998), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT53), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1049), .A2(G2078), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1050), .ZN(new_n1051));
  NOR3_X1   g626(.A1(new_n1030), .A2(new_n1051), .A3(new_n1031), .ZN(new_n1052));
  OAI21_X1  g627(.A(KEYINPUT124), .B1(new_n1048), .B2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1052), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT124), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1054), .A2(new_n1055), .A3(new_n1047), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1053), .A2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n988), .A2(new_n991), .A3(new_n762), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(new_n1049), .ZN(new_n1059));
  AOI21_X1  g634(.A(G301), .B1(new_n1057), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1047), .A2(KEYINPUT125), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n957), .A2(new_n958), .ZN(new_n1062));
  NOR3_X1   g637(.A1(new_n475), .A2(new_n962), .A3(new_n1051), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1063), .B1(KEYINPUT126), .B2(new_n483), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1064), .B1(KEYINPUT126), .B2(new_n483), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1062), .A2(new_n988), .A3(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT125), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n998), .A2(new_n1067), .A3(new_n1046), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1061), .A2(new_n1059), .A3(new_n1066), .A4(new_n1068), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1069), .A2(G171), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1045), .B1(new_n1060), .B2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1057), .A2(G301), .A3(new_n1059), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1069), .A2(G171), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(KEYINPUT127), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT127), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1069), .A2(new_n1075), .A3(G171), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1072), .A2(new_n1074), .A3(KEYINPUT54), .A4(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT50), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1078), .B1(new_n848), .B2(new_n956), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n514), .A2(new_n1078), .A3(new_n956), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n963), .A2(new_n1080), .ZN(new_n1081));
  NOR3_X1   g656(.A1(new_n1079), .A2(new_n1081), .A3(G2090), .ZN(new_n1082));
  OAI21_X1  g657(.A(G8), .B1(new_n992), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(new_n985), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1021), .A2(new_n1000), .A3(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1085), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1044), .A2(new_n1071), .A3(new_n1077), .A4(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(G1348), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n998), .A2(new_n1088), .ZN(new_n1089));
  OR2_X1    g664(.A1(new_n1002), .A2(G2067), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n898), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  XNOR2_X1  g666(.A(KEYINPUT56), .B(G2072), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n988), .A2(new_n991), .A3(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT120), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n988), .A2(new_n991), .A3(KEYINPUT120), .A4(new_n1092), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  XNOR2_X1  g672(.A(KEYINPUT118), .B(G1956), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1098), .B1(new_n1079), .B2(new_n1081), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(KEYINPUT119), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT119), .ZN(new_n1101));
  OAI211_X1 g676(.A(new_n1101), .B(new_n1098), .C1(new_n1079), .C2(new_n1081), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1097), .A2(new_n1103), .ZN(new_n1104));
  XNOR2_X1  g679(.A(new_n568), .B(KEYINPUT57), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1091), .B1(new_n1104), .B2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1097), .A2(new_n1105), .A3(new_n1103), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1108), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1111));
  AOI21_X1  g686(.A(KEYINPUT61), .B1(new_n1111), .B2(new_n1108), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n988), .A2(new_n991), .A3(new_n967), .ZN(new_n1113));
  XOR2_X1   g688(.A(KEYINPUT58), .B(G1341), .Z(new_n1114));
  NAND2_X1  g689(.A1(new_n1002), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(new_n555), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(KEYINPUT59), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT59), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1116), .A2(new_n1119), .A3(new_n555), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n848), .A2(new_n956), .ZN(new_n1122));
  NOR3_X1   g697(.A1(new_n1122), .A2(G2067), .A3(new_n989), .ZN(new_n1123));
  AOI211_X1 g698(.A(new_n606), .B(new_n1123), .C1(new_n1088), .C2(new_n998), .ZN(new_n1124));
  OAI21_X1  g699(.A(KEYINPUT60), .B1(new_n1124), .B2(new_n1091), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n898), .A2(KEYINPUT60), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1089), .A2(new_n1090), .A3(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1121), .A2(new_n1125), .A3(new_n1127), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1112), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1108), .A2(KEYINPUT121), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT121), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1097), .A2(new_n1131), .A3(new_n1103), .A4(new_n1105), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1130), .A2(new_n1111), .A3(KEYINPUT61), .A4(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1110), .B1(new_n1129), .B2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1024), .B1(new_n1087), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT62), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1136), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1038), .A2(new_n1041), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1138), .A2(KEYINPUT122), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1038), .A2(new_n1039), .A3(new_n1041), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1139), .A2(KEYINPUT62), .A3(new_n1140), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1137), .A2(new_n1141), .A3(new_n1086), .A4(new_n1060), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT63), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1144), .A2(G8), .A3(G168), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1143), .B1(new_n1085), .B2(new_n1145), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1145), .A2(new_n1143), .ZN(new_n1147));
  OAI21_X1  g722(.A(G8), .B1(new_n999), .B2(new_n994), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1020), .B1(new_n1148), .B2(new_n985), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT117), .ZN(new_n1150));
  OAI211_X1 g725(.A(new_n1000), .B(new_n1147), .C1(new_n1149), .C2(new_n1150), .ZN(new_n1151));
  AND2_X1   g726(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1146), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1142), .A2(new_n1153), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n983), .B1(new_n1135), .B2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n964), .B1(new_n973), .B2(new_n858), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT46), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n970), .A2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n968), .A2(KEYINPUT46), .A3(new_n969), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1156), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT47), .ZN(new_n1161));
  AND2_X1   g736(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n976), .A2(new_n978), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n965), .A2(new_n979), .ZN(new_n1165));
  XOR2_X1   g740(.A(new_n1165), .B(KEYINPUT48), .Z(new_n1166));
  OAI22_X1  g741(.A1(new_n1162), .A2(new_n1163), .B1(new_n1164), .B2(new_n1166), .ZN(new_n1167));
  NOR3_X1   g742(.A1(new_n802), .A2(new_n810), .A3(new_n806), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n976), .A2(new_n1168), .ZN(new_n1169));
  OR2_X1    g744(.A1(new_n756), .A2(G2067), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n964), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n1167), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1155), .A2(new_n1172), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g748(.A1(G401), .A2(new_n460), .A3(G227), .ZN(new_n1175));
  NAND3_X1  g749(.A1(new_n1175), .A2(new_n683), .A3(new_n682), .ZN(new_n1176));
  INV_X1    g750(.A(new_n1176), .ZN(new_n1177));
  OAI211_X1 g751(.A(new_n887), .B(new_n1177), .C1(new_n952), .C2(new_n953), .ZN(G225));
  INV_X1    g752(.A(G225), .ZN(G308));
endmodule


