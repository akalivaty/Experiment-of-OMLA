

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740;

  INV_X2 U366 ( .A(G953), .ZN(n734) );
  XNOR2_X2 U367 ( .A(n485), .B(KEYINPUT101), .ZN(n516) );
  NAND2_X2 U368 ( .A1(n599), .A2(n598), .ZN(n601) );
  XNOR2_X1 U369 ( .A(n646), .B(G146), .ZN(n426) );
  OR2_X1 U370 ( .A1(n538), .A2(n698), .ZN(n694) );
  XNOR2_X2 U371 ( .A(n419), .B(KEYINPUT105), .ZN(n506) );
  XNOR2_X1 U372 ( .A(n514), .B(n513), .ZN(n523) );
  OR2_X2 U373 ( .A1(n546), .A2(n545), .ZN(n547) );
  AND2_X2 U374 ( .A1(n583), .A2(n582), .ZN(n584) );
  NAND2_X2 U375 ( .A1(n585), .A2(n584), .ZN(n586) );
  AND2_X2 U376 ( .A1(n523), .A2(n522), .ZN(n672) );
  XOR2_X2 U377 ( .A(G110), .B(G101), .Z(n411) );
  XNOR2_X2 U378 ( .A(n414), .B(n345), .ZN(n615) );
  XNOR2_X2 U379 ( .A(n393), .B(KEYINPUT76), .ZN(n482) );
  INV_X1 U380 ( .A(n567), .ZN(n550) );
  NOR2_X2 U381 ( .A1(n482), .A2(n575), .ZN(n407) );
  INV_X2 U382 ( .A(n700), .ZN(n575) );
  INV_X1 U383 ( .A(n469), .ZN(n700) );
  NAND2_X1 U384 ( .A1(n355), .A2(n697), .ZN(n634) );
  XNOR2_X1 U385 ( .A(n353), .B(n397), .ZN(n422) );
  NOR2_X2 U386 ( .A1(n694), .A2(n468), .ZN(n576) );
  XNOR2_X1 U387 ( .A(n426), .B(n368), .ZN(n442) );
  INV_X1 U388 ( .A(KEYINPUT10), .ZN(n368) );
  XNOR2_X1 U389 ( .A(n398), .B(KEYINPUT3), .ZN(n353) );
  XNOR2_X1 U390 ( .A(n440), .B(n366), .ZN(n441) );
  XNOR2_X1 U391 ( .A(n423), .B(n424), .ZN(n352) );
  XNOR2_X1 U392 ( .A(n459), .B(n458), .ZN(n465) );
  OR2_X1 U393 ( .A1(n611), .A2(G902), .ZN(n458) );
  AND2_X1 U394 ( .A1(n481), .A2(n480), .ZN(n492) );
  OR2_X1 U395 ( .A1(n695), .A2(n360), .ZN(n362) );
  INV_X1 U396 ( .A(n694), .ZN(n359) );
  OR2_X2 U397 ( .A1(n364), .A2(n562), .ZN(n583) );
  INV_X1 U398 ( .A(KEYINPUT88), .ZN(n363) );
  XNOR2_X1 U399 ( .A(n486), .B(n436), .ZN(n531) );
  XNOR2_X1 U400 ( .A(G107), .B(G104), .ZN(n410) );
  NAND2_X1 U401 ( .A1(n484), .A2(n550), .ZN(n485) );
  AND2_X1 U402 ( .A1(n518), .A2(n683), .ZN(n486) );
  XNOR2_X1 U403 ( .A(n537), .B(n536), .ZN(n539) );
  AND2_X1 U404 ( .A1(n506), .A2(n531), .ZN(n622) );
  XNOR2_X1 U405 ( .A(n450), .B(G475), .ZN(n451) );
  AND2_X1 U406 ( .A1(n539), .A2(n695), .ZN(n568) );
  XNOR2_X1 U407 ( .A(G119), .B(G110), .ZN(n374) );
  XNOR2_X1 U408 ( .A(n358), .B(n357), .ZN(n611) );
  XNOR2_X1 U409 ( .A(n457), .B(n344), .ZN(n357) );
  XNOR2_X1 U410 ( .A(n640), .B(n350), .ZN(n605) );
  XNOR2_X1 U411 ( .A(n351), .B(n428), .ZN(n350) );
  BUF_X1 U412 ( .A(n622), .Z(n629) );
  XNOR2_X1 U413 ( .A(n356), .B(KEYINPUT67), .ZN(n355) );
  NAND2_X1 U414 ( .A1(n568), .A2(n575), .ZN(n356) );
  AND2_X1 U415 ( .A1(n501), .A2(n465), .ZN(n666) );
  AND2_X1 U416 ( .A1(n523), .A2(n346), .ZN(n343) );
  XOR2_X1 U417 ( .A(G107), .B(KEYINPUT9), .Z(n344) );
  XOR2_X1 U418 ( .A(n422), .B(n402), .Z(n345) );
  AND2_X1 U419 ( .A1(n522), .A2(n593), .ZN(n346) );
  XOR2_X1 U420 ( .A(KEYINPUT69), .B(KEYINPUT1), .Z(n347) );
  XOR2_X1 U421 ( .A(n558), .B(KEYINPUT35), .Z(n348) );
  AND2_X1 U422 ( .A1(n562), .A2(KEYINPUT88), .ZN(n349) );
  XNOR2_X1 U423 ( .A(n425), .B(n352), .ZN(n351) );
  XNOR2_X2 U424 ( .A(n354), .B(n422), .ZN(n640) );
  XNOR2_X2 U425 ( .A(n421), .B(n420), .ZN(n354) );
  XNOR2_X2 U426 ( .A(n411), .B(n410), .ZN(n421) );
  NAND2_X1 U427 ( .A1(n672), .A2(KEYINPUT2), .ZN(n524) );
  XNOR2_X1 U428 ( .A(n456), .B(n455), .ZN(n358) );
  NAND2_X1 U429 ( .A1(n359), .A2(n549), .ZN(n360) );
  NAND2_X1 U430 ( .A1(n572), .A2(KEYINPUT99), .ZN(n361) );
  OR2_X2 U431 ( .A1(n695), .A2(n694), .ZN(n572) );
  NAND2_X1 U432 ( .A1(n362), .A2(n361), .ZN(n551) );
  NAND2_X1 U433 ( .A1(n364), .A2(n363), .ZN(n560) );
  NAND2_X1 U434 ( .A1(n364), .A2(n349), .ZN(n564) );
  XNOR2_X1 U435 ( .A(n364), .B(n657), .ZN(G24) );
  XNOR2_X2 U436 ( .A(n559), .B(n348), .ZN(n364) );
  BUF_X1 U437 ( .A(n718), .Z(n725) );
  BUF_X1 U438 ( .A(n490), .Z(n468) );
  XNOR2_X2 U439 ( .A(n547), .B(KEYINPUT32), .ZN(n645) );
  AND2_X1 U440 ( .A1(G221), .A2(n453), .ZN(n365) );
  AND2_X1 U441 ( .A1(n439), .A2(G214), .ZN(n366) );
  XOR2_X1 U442 ( .A(n373), .B(KEYINPUT91), .Z(n367) );
  INV_X1 U443 ( .A(KEYINPUT46), .ZN(n508) );
  INV_X1 U444 ( .A(KEYINPUT66), .ZN(n600) );
  XNOR2_X1 U445 ( .A(n553), .B(n552), .ZN(n678) );
  NAND2_X1 U446 ( .A1(n678), .A2(n578), .ZN(n555) );
  XNOR2_X1 U447 ( .A(n452), .B(n451), .ZN(n501) );
  INV_X1 U448 ( .A(KEYINPUT63), .ZN(n620) );
  INV_X2 U449 ( .A(G125), .ZN(n646) );
  XNOR2_X1 U450 ( .A(G140), .B(G137), .ZN(n409) );
  XNOR2_X1 U451 ( .A(n442), .B(n409), .ZN(n731) );
  NAND2_X1 U452 ( .A1(n734), .A2(G234), .ZN(n370) );
  XNOR2_X1 U453 ( .A(KEYINPUT71), .B(KEYINPUT8), .ZN(n369) );
  XNOR2_X1 U454 ( .A(n370), .B(n369), .ZN(n453) );
  XNOR2_X1 U455 ( .A(n731), .B(n365), .ZN(n376) );
  XOR2_X1 U456 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n372) );
  XNOR2_X1 U457 ( .A(G128), .B(KEYINPUT92), .ZN(n371) );
  XNOR2_X1 U458 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U459 ( .A(n367), .B(n374), .ZN(n375) );
  XNOR2_X1 U460 ( .A(n376), .B(n375), .ZN(n726) );
  NOR2_X1 U461 ( .A1(n726), .A2(G902), .ZN(n382) );
  XOR2_X1 U462 ( .A(KEYINPUT25), .B(KEYINPUT80), .Z(n380) );
  XOR2_X1 U463 ( .A(KEYINPUT20), .B(KEYINPUT93), .Z(n378) );
  XNOR2_X1 U464 ( .A(KEYINPUT15), .B(G902), .ZN(n429) );
  NAND2_X1 U465 ( .A1(G234), .A2(n429), .ZN(n377) );
  XNOR2_X1 U466 ( .A(n378), .B(n377), .ZN(n383) );
  NAND2_X1 U467 ( .A1(n383), .A2(G217), .ZN(n379) );
  XNOR2_X1 U468 ( .A(n380), .B(n379), .ZN(n381) );
  XNOR2_X1 U469 ( .A(n382), .B(n381), .ZN(n538) );
  AND2_X1 U470 ( .A1(n383), .A2(G221), .ZN(n385) );
  INV_X1 U471 ( .A(KEYINPUT21), .ZN(n384) );
  XNOR2_X1 U472 ( .A(n385), .B(n384), .ZN(n698) );
  NOR2_X1 U473 ( .A1(G900), .A2(n734), .ZN(n386) );
  NAND2_X1 U474 ( .A1(G902), .A2(n386), .ZN(n387) );
  NAND2_X1 U475 ( .A1(n734), .A2(G952), .ZN(n526) );
  AND2_X1 U476 ( .A1(n387), .A2(n526), .ZN(n390) );
  NAND2_X1 U477 ( .A1(G237), .A2(G234), .ZN(n389) );
  INV_X1 U478 ( .A(KEYINPUT14), .ZN(n388) );
  XNOR2_X1 U479 ( .A(n389), .B(n388), .ZN(n714) );
  NOR2_X1 U480 ( .A1(n390), .A2(n714), .ZN(n472) );
  INV_X1 U481 ( .A(n472), .ZN(n391) );
  NOR2_X1 U482 ( .A1(n698), .A2(n391), .ZN(n392) );
  NAND2_X1 U483 ( .A1(n538), .A2(n392), .ZN(n393) );
  XNOR2_X2 U484 ( .A(G143), .B(KEYINPUT65), .ZN(n394) );
  XNOR2_X2 U485 ( .A(n394), .B(G128), .ZN(n425) );
  XNOR2_X2 U486 ( .A(n425), .B(G134), .ZN(n456) );
  XNOR2_X2 U487 ( .A(KEYINPUT64), .B(KEYINPUT4), .ZN(n427) );
  XNOR2_X1 U488 ( .A(n427), .B(KEYINPUT73), .ZN(n395) );
  XNOR2_X1 U489 ( .A(KEYINPUT72), .B(G131), .ZN(n445) );
  XNOR2_X1 U490 ( .A(n395), .B(n445), .ZN(n396) );
  XNOR2_X2 U491 ( .A(n456), .B(n396), .ZN(n733) );
  XNOR2_X2 U492 ( .A(n733), .B(G146), .ZN(n414) );
  XNOR2_X1 U493 ( .A(G119), .B(G113), .ZN(n397) );
  XNOR2_X1 U494 ( .A(G116), .B(KEYINPUT77), .ZN(n398) );
  NOR2_X1 U495 ( .A1(G953), .A2(G237), .ZN(n439) );
  NAND2_X1 U496 ( .A1(n439), .A2(G210), .ZN(n399) );
  XNOR2_X1 U497 ( .A(n399), .B(G101), .ZN(n401) );
  XNOR2_X1 U498 ( .A(KEYINPUT5), .B(G137), .ZN(n400) );
  XNOR2_X1 U499 ( .A(n401), .B(n400), .ZN(n402) );
  INV_X1 U500 ( .A(n615), .ZN(n404) );
  INV_X1 U501 ( .A(G902), .ZN(n403) );
  NAND2_X1 U502 ( .A1(n404), .A2(n403), .ZN(n406) );
  INV_X1 U503 ( .A(G472), .ZN(n405) );
  XNOR2_X1 U504 ( .A(n406), .B(n405), .ZN(n469) );
  XNOR2_X1 U505 ( .A(n407), .B(KEYINPUT28), .ZN(n418) );
  NAND2_X1 U506 ( .A1(n734), .A2(G227), .ZN(n408) );
  XNOR2_X1 U507 ( .A(n409), .B(n408), .ZN(n412) );
  XNOR2_X1 U508 ( .A(n412), .B(n421), .ZN(n413) );
  XNOR2_X1 U509 ( .A(n414), .B(n413), .ZN(n719) );
  OR2_X2 U510 ( .A1(n719), .A2(G902), .ZN(n416) );
  INV_X1 U511 ( .A(G469), .ZN(n415) );
  XNOR2_X2 U512 ( .A(n416), .B(n415), .ZN(n490) );
  XOR2_X1 U513 ( .A(n468), .B(KEYINPUT104), .Z(n417) );
  NAND2_X1 U514 ( .A1(n418), .A2(n417), .ZN(n419) );
  XNOR2_X1 U515 ( .A(KEYINPUT16), .B(G122), .ZN(n420) );
  XNOR2_X1 U516 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n424) );
  NAND2_X1 U517 ( .A1(n734), .A2(G224), .ZN(n423) );
  XNOR2_X1 U518 ( .A(n427), .B(n426), .ZN(n428) );
  INV_X1 U519 ( .A(n429), .ZN(n591) );
  OR2_X2 U520 ( .A1(n605), .A2(n591), .ZN(n434) );
  INV_X1 U521 ( .A(G237), .ZN(n430) );
  NAND2_X1 U522 ( .A1(n403), .A2(n430), .ZN(n435) );
  NAND2_X1 U523 ( .A1(n435), .A2(G210), .ZN(n432) );
  INV_X1 U524 ( .A(KEYINPUT84), .ZN(n431) );
  XNOR2_X1 U525 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X2 U526 ( .A(n434), .B(n433), .ZN(n518) );
  AND2_X1 U527 ( .A1(n435), .A2(G214), .ZN(n502) );
  INV_X1 U528 ( .A(n502), .ZN(n683) );
  XNOR2_X1 U529 ( .A(KEYINPUT79), .B(KEYINPUT19), .ZN(n436) );
  XOR2_X1 U530 ( .A(KEYINPUT12), .B(KEYINPUT95), .Z(n438) );
  XNOR2_X1 U531 ( .A(G140), .B(KEYINPUT94), .ZN(n437) );
  XNOR2_X1 U532 ( .A(n438), .B(n437), .ZN(n440) );
  XNOR2_X1 U533 ( .A(n442), .B(n441), .ZN(n449) );
  XNOR2_X1 U534 ( .A(G143), .B(G122), .ZN(n443) );
  XOR2_X1 U535 ( .A(n443), .B(KEYINPUT11), .Z(n444) );
  XNOR2_X1 U536 ( .A(n445), .B(n444), .ZN(n447) );
  XOR2_X1 U537 ( .A(G104), .B(G113), .Z(n446) );
  XNOR2_X1 U538 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U539 ( .A(n449), .B(n448), .ZN(n651) );
  NOR2_X1 U540 ( .A1(G902), .A2(n651), .ZN(n452) );
  XNOR2_X1 U541 ( .A(KEYINPUT96), .B(KEYINPUT13), .ZN(n450) );
  XNOR2_X1 U542 ( .A(G478), .B(KEYINPUT97), .ZN(n459) );
  NAND2_X1 U543 ( .A1(n453), .A2(G217), .ZN(n457) );
  XOR2_X1 U544 ( .A(KEYINPUT7), .B(G122), .Z(n454) );
  XOR2_X1 U545 ( .A(n454), .B(G116), .Z(n455) );
  INV_X1 U546 ( .A(n666), .ZN(n460) );
  OR2_X1 U547 ( .A1(n501), .A2(n465), .ZN(n628) );
  AND2_X1 U548 ( .A1(n460), .A2(n628), .ZN(n688) );
  INV_X1 U549 ( .A(n688), .ZN(n478) );
  NOR2_X1 U550 ( .A1(KEYINPUT47), .A2(KEYINPUT85), .ZN(n461) );
  NAND2_X1 U551 ( .A1(n478), .A2(n461), .ZN(n463) );
  NAND2_X1 U552 ( .A1(n688), .A2(KEYINPUT85), .ZN(n462) );
  NAND2_X1 U553 ( .A1(n463), .A2(n462), .ZN(n464) );
  NAND2_X1 U554 ( .A1(n622), .A2(n464), .ZN(n477) );
  INV_X1 U555 ( .A(n465), .ZN(n500) );
  NAND2_X1 U556 ( .A1(n501), .A2(n500), .ZN(n467) );
  INV_X1 U557 ( .A(KEYINPUT100), .ZN(n466) );
  XNOR2_X1 U558 ( .A(n467), .B(n466), .ZN(n556) );
  AND2_X1 U559 ( .A1(n556), .A2(n518), .ZN(n476) );
  XNOR2_X1 U560 ( .A(n576), .B(KEYINPUT102), .ZN(n475) );
  OR2_X1 U561 ( .A1(n469), .A2(n502), .ZN(n471) );
  XNOR2_X1 U562 ( .A(KEYINPUT103), .B(KEYINPUT30), .ZN(n470) );
  XNOR2_X1 U563 ( .A(n471), .B(n470), .ZN(n473) );
  AND2_X1 U564 ( .A1(n473), .A2(n472), .ZN(n474) );
  AND2_X1 U565 ( .A1(n475), .A2(n474), .ZN(n494) );
  NAND2_X1 U566 ( .A1(n476), .A2(n494), .ZN(n665) );
  AND2_X1 U567 ( .A1(n477), .A2(n665), .ZN(n481) );
  NAND2_X1 U568 ( .A1(n622), .A2(n478), .ZN(n479) );
  NAND2_X1 U569 ( .A1(n479), .A2(KEYINPUT47), .ZN(n480) );
  INV_X1 U570 ( .A(n482), .ZN(n483) );
  AND2_X1 U571 ( .A1(n483), .A2(n666), .ZN(n484) );
  XNOR2_X2 U572 ( .A(n700), .B(KEYINPUT6), .ZN(n567) );
  XNOR2_X1 U573 ( .A(n516), .B(KEYINPUT108), .ZN(n487) );
  NAND2_X1 U574 ( .A1(n487), .A2(n486), .ZN(n489) );
  INV_X1 U575 ( .A(KEYINPUT36), .ZN(n488) );
  XNOR2_X1 U576 ( .A(n489), .B(n488), .ZN(n491) );
  XNOR2_X2 U577 ( .A(n490), .B(n347), .ZN(n695) );
  INV_X1 U578 ( .A(n695), .ZN(n540) );
  NAND2_X1 U579 ( .A1(n491), .A2(n540), .ZN(n649) );
  NAND2_X1 U580 ( .A1(n492), .A2(n649), .ZN(n493) );
  XNOR2_X1 U581 ( .A(n493), .B(KEYINPUT75), .ZN(n511) );
  XNOR2_X1 U582 ( .A(n518), .B(KEYINPUT38), .ZN(n503) );
  INV_X1 U583 ( .A(n503), .ZN(n684) );
  NAND2_X1 U584 ( .A1(n494), .A2(n684), .ZN(n496) );
  INV_X1 U585 ( .A(KEYINPUT39), .ZN(n495) );
  XNOR2_X1 U586 ( .A(n496), .B(n495), .ZN(n521) );
  INV_X1 U587 ( .A(n521), .ZN(n497) );
  NAND2_X1 U588 ( .A1(n497), .A2(n666), .ZN(n499) );
  XNOR2_X1 U589 ( .A(KEYINPUT106), .B(KEYINPUT40), .ZN(n498) );
  XNOR2_X1 U590 ( .A(n499), .B(n498), .ZN(n650) );
  OR2_X1 U591 ( .A1(n501), .A2(n500), .ZN(n686) );
  OR2_X1 U592 ( .A1(n503), .A2(n502), .ZN(n687) );
  NOR2_X1 U593 ( .A1(n686), .A2(n687), .ZN(n505) );
  XNOR2_X1 U594 ( .A(KEYINPUT107), .B(KEYINPUT41), .ZN(n504) );
  XNOR2_X1 U595 ( .A(n505), .B(n504), .ZN(n707) );
  NAND2_X1 U596 ( .A1(n506), .A2(n707), .ZN(n507) );
  XNOR2_X1 U597 ( .A(n507), .B(KEYINPUT42), .ZN(n632) );
  NAND2_X1 U598 ( .A1(n650), .A2(n632), .ZN(n509) );
  XNOR2_X1 U599 ( .A(n509), .B(n508), .ZN(n510) );
  NAND2_X1 U600 ( .A1(n511), .A2(n510), .ZN(n514) );
  INV_X1 U601 ( .A(KEYINPUT74), .ZN(n512) );
  XNOR2_X1 U602 ( .A(n512), .B(KEYINPUT48), .ZN(n513) );
  AND2_X1 U603 ( .A1(n695), .A2(n683), .ZN(n515) );
  NAND2_X1 U604 ( .A1(n516), .A2(n515), .ZN(n517) );
  XNOR2_X1 U605 ( .A(n517), .B(KEYINPUT43), .ZN(n520) );
  INV_X1 U606 ( .A(n518), .ZN(n519) );
  NAND2_X1 U607 ( .A1(n520), .A2(n519), .ZN(n627) );
  OR2_X1 U608 ( .A1(n521), .A2(n628), .ZN(n625) );
  AND2_X1 U609 ( .A1(n627), .A2(n625), .ZN(n522) );
  XNOR2_X1 U610 ( .A(n524), .B(KEYINPUT86), .ZN(n588) );
  NOR2_X1 U611 ( .A1(n686), .A2(n698), .ZN(n534) );
  NOR2_X1 U612 ( .A1(G898), .A2(n734), .ZN(n525) );
  XOR2_X1 U613 ( .A(KEYINPUT89), .B(n525), .Z(n639) );
  NAND2_X1 U614 ( .A1(n639), .A2(G902), .ZN(n527) );
  NAND2_X1 U615 ( .A1(n527), .A2(n526), .ZN(n529) );
  INV_X1 U616 ( .A(n714), .ZN(n528) );
  AND2_X1 U617 ( .A1(n529), .A2(n528), .ZN(n530) );
  NAND2_X1 U618 ( .A1(n531), .A2(n530), .ZN(n533) );
  INV_X1 U619 ( .A(KEYINPUT0), .ZN(n532) );
  XNOR2_X2 U620 ( .A(n533), .B(n532), .ZN(n573) );
  NAND2_X1 U621 ( .A1(n534), .A2(n573), .ZN(n537) );
  INV_X1 U622 ( .A(KEYINPUT68), .ZN(n535) );
  XNOR2_X1 U623 ( .A(n535), .B(KEYINPUT22), .ZN(n536) );
  BUF_X1 U624 ( .A(n538), .Z(n697) );
  INV_X1 U625 ( .A(n539), .ZN(n546) );
  NAND2_X1 U626 ( .A1(n540), .A2(n697), .ZN(n541) );
  XNOR2_X1 U627 ( .A(n541), .B(KEYINPUT98), .ZN(n543) );
  XNOR2_X1 U628 ( .A(n567), .B(KEYINPUT83), .ZN(n542) );
  OR2_X1 U629 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U630 ( .A(n544), .B(KEYINPUT82), .ZN(n545) );
  NAND2_X1 U631 ( .A1(n634), .A2(n645), .ZN(n548) );
  INV_X1 U632 ( .A(KEYINPUT44), .ZN(n562) );
  AND2_X1 U633 ( .A1(n548), .A2(n562), .ZN(n561) );
  INV_X1 U634 ( .A(KEYINPUT99), .ZN(n549) );
  NAND2_X1 U635 ( .A1(n551), .A2(n550), .ZN(n553) );
  XNOR2_X1 U636 ( .A(KEYINPUT78), .B(KEYINPUT33), .ZN(n552) );
  XNOR2_X1 U637 ( .A(n573), .B(KEYINPUT90), .ZN(n578) );
  INV_X1 U638 ( .A(KEYINPUT34), .ZN(n554) );
  XNOR2_X1 U639 ( .A(n555), .B(n554), .ZN(n557) );
  NAND2_X1 U640 ( .A1(n557), .A2(n556), .ZN(n559) );
  INV_X1 U641 ( .A(KEYINPUT81), .ZN(n558) );
  NAND2_X1 U642 ( .A1(n561), .A2(n560), .ZN(n566) );
  AND2_X1 U643 ( .A1(n634), .A2(n645), .ZN(n563) );
  NAND2_X1 U644 ( .A1(n564), .A2(n563), .ZN(n565) );
  NAND2_X1 U645 ( .A1(n566), .A2(n565), .ZN(n585) );
  NAND2_X1 U646 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U647 ( .A(n569), .B(KEYINPUT87), .ZN(n571) );
  INV_X1 U648 ( .A(n697), .ZN(n570) );
  AND2_X1 U649 ( .A1(n571), .A2(n570), .ZN(n658) );
  NOR2_X1 U650 ( .A1(n572), .A2(n575), .ZN(n704) );
  NAND2_X1 U651 ( .A1(n704), .A2(n573), .ZN(n574) );
  XNOR2_X1 U652 ( .A(n574), .B(KEYINPUT31), .ZN(n669) );
  AND2_X1 U653 ( .A1(n576), .A2(n575), .ZN(n577) );
  AND2_X1 U654 ( .A1(n578), .A2(n577), .ZN(n661) );
  OR2_X1 U655 ( .A1(n669), .A2(n661), .ZN(n580) );
  XNOR2_X1 U656 ( .A(n688), .B(KEYINPUT85), .ZN(n579) );
  AND2_X1 U657 ( .A1(n580), .A2(n579), .ZN(n581) );
  NOR2_X1 U658 ( .A1(n658), .A2(n581), .ZN(n582) );
  XNOR2_X2 U659 ( .A(n586), .B(KEYINPUT45), .ZN(n673) );
  INV_X1 U660 ( .A(n673), .ZN(n587) );
  NOR2_X2 U661 ( .A1(n588), .A2(n587), .ZN(n676) );
  NAND2_X1 U662 ( .A1(n591), .A2(KEYINPUT2), .ZN(n590) );
  INV_X1 U663 ( .A(KEYINPUT70), .ZN(n589) );
  NAND2_X1 U664 ( .A1(n590), .A2(n589), .ZN(n594) );
  INV_X1 U665 ( .A(n594), .ZN(n592) );
  OR2_X1 U666 ( .A1(n592), .A2(n591), .ZN(n593) );
  NAND2_X1 U667 ( .A1(n343), .A2(n673), .ZN(n599) );
  INV_X1 U668 ( .A(n593), .ZN(n597) );
  NAND2_X1 U669 ( .A1(KEYINPUT2), .A2(KEYINPUT70), .ZN(n595) );
  AND2_X1 U670 ( .A1(n595), .A2(n594), .ZN(n596) );
  OR2_X1 U671 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X2 U672 ( .A(n601), .B(n600), .ZN(n602) );
  NOR2_X4 U673 ( .A1(n676), .A2(n602), .ZN(n718) );
  NAND2_X1 U674 ( .A1(n718), .A2(G210), .ZN(n607) );
  XOR2_X1 U675 ( .A(KEYINPUT117), .B(KEYINPUT54), .Z(n603) );
  XOR2_X1 U676 ( .A(n603), .B(KEYINPUT55), .Z(n604) );
  XNOR2_X1 U677 ( .A(n605), .B(n604), .ZN(n606) );
  XNOR2_X1 U678 ( .A(n607), .B(n606), .ZN(n609) );
  INV_X1 U679 ( .A(G952), .ZN(n608) );
  AND2_X1 U680 ( .A1(n608), .A2(G953), .ZN(n730) );
  NOR2_X2 U681 ( .A1(n609), .A2(n730), .ZN(n610) );
  XNOR2_X1 U682 ( .A(n610), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U683 ( .A1(n718), .A2(G478), .ZN(n612) );
  XNOR2_X1 U684 ( .A(n612), .B(n611), .ZN(n613) );
  NOR2_X2 U685 ( .A1(n613), .A2(n730), .ZN(n614) );
  XNOR2_X1 U686 ( .A(n614), .B(KEYINPUT120), .ZN(G63) );
  NAND2_X1 U687 ( .A1(n718), .A2(G472), .ZN(n618) );
  XOR2_X1 U688 ( .A(KEYINPUT109), .B(KEYINPUT62), .Z(n616) );
  XNOR2_X1 U689 ( .A(n615), .B(n616), .ZN(n617) );
  XNOR2_X1 U690 ( .A(n618), .B(n617), .ZN(n619) );
  NOR2_X2 U691 ( .A1(n619), .A2(n730), .ZN(n621) );
  XNOR2_X1 U692 ( .A(n621), .B(n620), .ZN(G57) );
  NAND2_X1 U693 ( .A1(n629), .A2(n666), .ZN(n624) );
  XOR2_X1 U694 ( .A(G146), .B(KEYINPUT111), .Z(n623) );
  XNOR2_X1 U695 ( .A(n624), .B(n623), .ZN(G48) );
  XNOR2_X1 U696 ( .A(n625), .B(G134), .ZN(G36) );
  XNOR2_X1 U697 ( .A(G140), .B(KEYINPUT114), .ZN(n626) );
  XNOR2_X1 U698 ( .A(n627), .B(n626), .ZN(G42) );
  XNOR2_X1 U699 ( .A(G128), .B(KEYINPUT29), .ZN(n631) );
  INV_X1 U700 ( .A(n628), .ZN(n670) );
  NAND2_X1 U701 ( .A1(n629), .A2(n670), .ZN(n630) );
  XOR2_X1 U702 ( .A(n631), .B(n630), .Z(G30) );
  XOR2_X1 U703 ( .A(G137), .B(KEYINPUT126), .Z(n633) );
  XOR2_X1 U704 ( .A(n633), .B(n632), .Z(G39) );
  XNOR2_X1 U705 ( .A(n634), .B(G110), .ZN(G12) );
  NAND2_X1 U706 ( .A1(n673), .A2(n734), .ZN(n638) );
  NAND2_X1 U707 ( .A1(G953), .A2(G224), .ZN(n635) );
  XNOR2_X1 U708 ( .A(KEYINPUT61), .B(n635), .ZN(n636) );
  NAND2_X1 U709 ( .A1(n636), .A2(G898), .ZN(n637) );
  NAND2_X1 U710 ( .A1(n638), .A2(n637), .ZN(n643) );
  NOR2_X1 U711 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U712 ( .A(n641), .B(KEYINPUT122), .ZN(n642) );
  XNOR2_X1 U713 ( .A(n643), .B(n642), .ZN(G69) );
  XNOR2_X1 U714 ( .A(G119), .B(KEYINPUT125), .ZN(n644) );
  XOR2_X1 U715 ( .A(n645), .B(n644), .Z(G21) );
  XOR2_X1 U716 ( .A(KEYINPUT37), .B(KEYINPUT113), .Z(n647) );
  XNOR2_X1 U717 ( .A(n647), .B(n646), .ZN(n648) );
  XNOR2_X1 U718 ( .A(n649), .B(n648), .ZN(G27) );
  XNOR2_X1 U719 ( .A(n650), .B(G131), .ZN(G33) );
  NAND2_X1 U720 ( .A1(n718), .A2(G475), .ZN(n653) );
  XOR2_X1 U721 ( .A(KEYINPUT59), .B(n651), .Z(n652) );
  XNOR2_X1 U722 ( .A(n653), .B(n652), .ZN(n654) );
  NOR2_X2 U723 ( .A1(n654), .A2(n730), .ZN(n656) );
  XOR2_X1 U724 ( .A(KEYINPUT119), .B(KEYINPUT60), .Z(n655) );
  XNOR2_X1 U725 ( .A(n656), .B(n655), .ZN(G60) );
  XNOR2_X1 U726 ( .A(G122), .B(KEYINPUT124), .ZN(n657) );
  XOR2_X1 U727 ( .A(G101), .B(n658), .Z(G3) );
  NAND2_X1 U728 ( .A1(n661), .A2(n666), .ZN(n659) );
  XNOR2_X1 U729 ( .A(n659), .B(KEYINPUT110), .ZN(n660) );
  XNOR2_X1 U730 ( .A(G104), .B(n660), .ZN(G6) );
  XOR2_X1 U731 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n663) );
  NAND2_X1 U732 ( .A1(n661), .A2(n670), .ZN(n662) );
  XNOR2_X1 U733 ( .A(n663), .B(n662), .ZN(n664) );
  XNOR2_X1 U734 ( .A(G107), .B(n664), .ZN(G9) );
  XNOR2_X1 U735 ( .A(G143), .B(n665), .ZN(G45) );
  NAND2_X1 U736 ( .A1(n666), .A2(n669), .ZN(n667) );
  XNOR2_X1 U737 ( .A(n667), .B(KEYINPUT112), .ZN(n668) );
  XNOR2_X1 U738 ( .A(G113), .B(n668), .ZN(G15) );
  NAND2_X1 U739 ( .A1(n670), .A2(n669), .ZN(n671) );
  XNOR2_X1 U740 ( .A(n671), .B(G116), .ZN(G18) );
  AND2_X1 U741 ( .A1(n672), .A2(n673), .ZN(n674) );
  NOR2_X1 U742 ( .A1(n674), .A2(KEYINPUT2), .ZN(n675) );
  NOR2_X1 U743 ( .A1(n676), .A2(n675), .ZN(n677) );
  NOR2_X1 U744 ( .A1(n677), .A2(G953), .ZN(n682) );
  BUF_X1 U745 ( .A(n678), .Z(n679) );
  NAND2_X1 U746 ( .A1(n679), .A2(n707), .ZN(n680) );
  XNOR2_X1 U747 ( .A(n680), .B(KEYINPUT116), .ZN(n681) );
  NAND2_X1 U748 ( .A1(n682), .A2(n681), .ZN(n716) );
  INV_X1 U749 ( .A(n679), .ZN(n692) );
  NOR2_X1 U750 ( .A1(n684), .A2(n683), .ZN(n685) );
  NOR2_X1 U751 ( .A1(n686), .A2(n685), .ZN(n690) );
  NOR2_X1 U752 ( .A1(n688), .A2(n687), .ZN(n689) );
  NOR2_X1 U753 ( .A1(n690), .A2(n689), .ZN(n691) );
  NOR2_X1 U754 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U755 ( .A(n693), .B(KEYINPUT115), .ZN(n710) );
  NAND2_X1 U756 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U757 ( .A(n696), .B(KEYINPUT50), .ZN(n703) );
  NAND2_X1 U758 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U759 ( .A(KEYINPUT49), .B(n699), .ZN(n701) );
  NOR2_X1 U760 ( .A1(n701), .A2(n700), .ZN(n702) );
  AND2_X1 U761 ( .A1(n703), .A2(n702), .ZN(n705) );
  NOR2_X1 U762 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U763 ( .A(KEYINPUT51), .B(n706), .ZN(n708) );
  NAND2_X1 U764 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U765 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U766 ( .A(KEYINPUT52), .B(n711), .ZN(n712) );
  NAND2_X1 U767 ( .A1(n712), .A2(G952), .ZN(n713) );
  NOR2_X1 U768 ( .A1(n714), .A2(n713), .ZN(n715) );
  NOR2_X1 U769 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U770 ( .A(KEYINPUT53), .B(n717), .ZN(G75) );
  NAND2_X1 U771 ( .A1(n725), .A2(G469), .ZN(n723) );
  XOR2_X1 U772 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n720) );
  XNOR2_X1 U773 ( .A(n720), .B(KEYINPUT118), .ZN(n721) );
  XNOR2_X1 U774 ( .A(n719), .B(n721), .ZN(n722) );
  XNOR2_X1 U775 ( .A(n723), .B(n722), .ZN(n724) );
  NOR2_X1 U776 ( .A1(n730), .A2(n724), .ZN(G54) );
  NAND2_X1 U777 ( .A1(n725), .A2(G217), .ZN(n728) );
  XOR2_X1 U778 ( .A(n726), .B(KEYINPUT121), .Z(n727) );
  XNOR2_X1 U779 ( .A(n728), .B(n727), .ZN(n729) );
  NOR2_X1 U780 ( .A1(n730), .A2(n729), .ZN(G66) );
  XNOR2_X1 U781 ( .A(n731), .B(KEYINPUT123), .ZN(n732) );
  XNOR2_X1 U782 ( .A(n733), .B(n732), .ZN(n736) );
  XOR2_X1 U783 ( .A(n736), .B(n672), .Z(n735) );
  NAND2_X1 U784 ( .A1(n735), .A2(n734), .ZN(n740) );
  XNOR2_X1 U785 ( .A(G227), .B(n736), .ZN(n737) );
  NAND2_X1 U786 ( .A1(n737), .A2(G900), .ZN(n738) );
  NAND2_X1 U787 ( .A1(n738), .A2(G953), .ZN(n739) );
  NAND2_X1 U788 ( .A1(n740), .A2(n739), .ZN(G72) );
endmodule

