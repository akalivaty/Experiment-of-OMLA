//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 1 1 1 0 1 1 0 0 0 1 1 1 1 0 0 1 1 0 0 0 1 1 1 1 0 1 0 1 0 1 1 1 0 0 1 1 0 0 0 0 0 0 1 1 0 0 0 1 0 0 0 0 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:35 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1225,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  INV_X1    g0003(.A(G77), .ZN(new_n204));
  NAND4_X1  g0004(.A1(new_n201), .A2(new_n202), .A3(new_n203), .A4(new_n204), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT64), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XOR2_X1   g0010(.A(KEYINPUT65), .B(KEYINPUT0), .Z(new_n211));
  XNOR2_X1  g0011(.A(new_n210), .B(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT67), .ZN(new_n214));
  INV_X1    g0014(.A(G232), .ZN(new_n215));
  INV_X1    g0015(.A(G238), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n214), .B1(new_n202), .B2(new_n215), .C1(new_n203), .C2(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  XOR2_X1   g0018(.A(KEYINPUT68), .B(G244), .Z(new_n219));
  AOI22_X1  g0019(.A1(new_n219), .A2(G77), .B1(G107), .B2(G264), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(KEYINPUT69), .ZN(new_n222));
  NAND3_X1  g0022(.A1(new_n218), .A2(new_n220), .A3(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n223), .A2(new_n208), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT1), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  INV_X1    g0026(.A(G20), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT66), .ZN(new_n229));
  OAI21_X1  g0029(.A(G50), .B1(G58), .B2(G68), .ZN(new_n230));
  INV_X1    g0030(.A(new_n230), .ZN(new_n231));
  AOI211_X1 g0031(.A(new_n212), .B(new_n225), .C1(new_n229), .C2(new_n231), .ZN(G361));
  XNOR2_X1  g0032(.A(KEYINPUT2), .B(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  INV_X1    g0037(.A(G264), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n236), .B(new_n240), .ZN(G358));
  XOR2_X1   g0041(.A(G68), .B(G77), .Z(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G58), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G107), .B(G116), .Z(new_n245));
  XNOR2_X1  g0045(.A(G87), .B(G97), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  NAND3_X1  g0048(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(KEYINPUT72), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT72), .ZN(new_n251));
  NAND4_X1  g0051(.A1(new_n251), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n250), .A2(new_n226), .A3(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G116), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(G20), .ZN(new_n255));
  NAND2_X1  g0055(.A1(G33), .A2(G283), .ZN(new_n256));
  INV_X1    g0056(.A(G97), .ZN(new_n257));
  OAI211_X1 g0057(.A(new_n256), .B(new_n227), .C1(G33), .C2(new_n257), .ZN(new_n258));
  NAND4_X1  g0058(.A1(new_n253), .A2(KEYINPUT20), .A3(new_n255), .A4(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT85), .ZN(new_n260));
  OR2_X1    g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n253), .A2(new_n255), .A3(new_n258), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT20), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n259), .A2(new_n260), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n261), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G33), .ZN(new_n267));
  INV_X1    g0067(.A(G1), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(KEYINPUT71), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT71), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(G1), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n267), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n227), .B1(new_n269), .B2(new_n271), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n272), .B1(G13), .B2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(new_n253), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G116), .ZN(new_n278));
  INV_X1    g0078(.A(G13), .ZN(new_n279));
  AOI211_X1 g0079(.A(new_n279), .B(new_n227), .C1(new_n269), .C2(new_n271), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(new_n254), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n266), .A2(new_n278), .A3(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G169), .ZN(new_n283));
  INV_X1    g0083(.A(G45), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n284), .B1(new_n269), .B2(new_n271), .ZN(new_n285));
  INV_X1    g0085(.A(G41), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(KEYINPUT5), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(KEYINPUT70), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT70), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G41), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT5), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n288), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n285), .A2(new_n287), .A3(new_n292), .ZN(new_n293));
  OAI211_X1 g0093(.A(G1), .B(G13), .C1(new_n267), .C2(new_n286), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(G274), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT78), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n297), .A2(KEYINPUT3), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT3), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n299), .A2(KEYINPUT78), .ZN(new_n300));
  OAI21_X1  g0100(.A(G33), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G257), .ZN(new_n302));
  INV_X1    g0102(.A(G1698), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n238), .A2(G1698), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT77), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n306), .B1(new_n299), .B2(G33), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n267), .A2(KEYINPUT77), .A3(KEYINPUT3), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n301), .A2(new_n304), .A3(new_n305), .A4(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n267), .A2(KEYINPUT3), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n299), .A2(G33), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(G303), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n310), .A2(new_n314), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n226), .B1(G33), .B2(G41), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n296), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  AND3_X1   g0117(.A1(new_n293), .A2(G270), .A3(new_n294), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n283), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n282), .A2(KEYINPUT21), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n282), .A2(new_n320), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT21), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n294), .B1(new_n310), .B2(new_n314), .ZN(new_n325));
  NOR3_X1   g0125(.A1(new_n325), .A2(new_n318), .A3(new_n296), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n282), .A2(G179), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n317), .A2(new_n319), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(G200), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n326), .A2(G190), .ZN(new_n330));
  XNOR2_X1  g0130(.A(new_n259), .B(KEYINPUT85), .ZN(new_n331));
  AOI22_X1  g0131(.A1(new_n331), .A2(new_n264), .B1(new_n254), .B2(new_n280), .ZN(new_n332));
  NAND4_X1  g0132(.A1(new_n329), .A2(new_n330), .A3(new_n332), .A4(new_n278), .ZN(new_n333));
  AND4_X1   g0133(.A1(new_n321), .A2(new_n324), .A3(new_n327), .A4(new_n333), .ZN(new_n334));
  AND2_X1   g0134(.A1(new_n311), .A2(new_n312), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n303), .A2(G222), .ZN(new_n336));
  INV_X1    g0136(.A(G223), .ZN(new_n337));
  OAI211_X1 g0137(.A(new_n335), .B(new_n336), .C1(new_n337), .C2(new_n303), .ZN(new_n338));
  OAI211_X1 g0138(.A(new_n338), .B(new_n316), .C1(G77), .C2(new_n335), .ZN(new_n339));
  AND2_X1   g0139(.A1(new_n288), .A2(new_n290), .ZN(new_n340));
  OAI211_X1 g0140(.A(new_n268), .B(G274), .C1(new_n340), .C2(G45), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n286), .B1(new_n269), .B2(new_n271), .ZN(new_n343));
  NOR3_X1   g0143(.A1(new_n285), .A2(new_n343), .A3(new_n316), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n342), .B1(G226), .B2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(G200), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT75), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT10), .ZN(new_n348));
  OAI22_X1  g0148(.A1(new_n345), .A2(new_n346), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n349), .B1(G190), .B2(new_n345), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n253), .A2(new_n273), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(G50), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n269), .A2(new_n271), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n353), .A2(G13), .A3(G20), .ZN(new_n354));
  INV_X1    g0154(.A(G150), .ZN(new_n355));
  NOR2_X1   g0155(.A1(G20), .A2(G33), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  NOR3_X1   g0157(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n358));
  OAI22_X1  g0158(.A1(new_n355), .A2(new_n357), .B1(new_n358), .B2(new_n227), .ZN(new_n359));
  XNOR2_X1  g0159(.A(KEYINPUT8), .B(G58), .ZN(new_n360));
  XOR2_X1   g0160(.A(new_n360), .B(KEYINPUT73), .Z(new_n361));
  NOR2_X1   g0161(.A1(new_n267), .A2(G20), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n359), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  OAI221_X1 g0163(.A(new_n352), .B1(G50), .B2(new_n354), .C1(new_n363), .C2(new_n275), .ZN(new_n364));
  XNOR2_X1  g0164(.A(new_n364), .B(KEYINPUT9), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n350), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n366), .A2(new_n347), .A3(new_n348), .ZN(new_n367));
  OAI211_X1 g0167(.A(new_n350), .B(new_n365), .C1(KEYINPUT75), .C2(KEYINPUT10), .ZN(new_n368));
  OR2_X1    g0168(.A1(new_n345), .A2(G169), .ZN(new_n369));
  INV_X1    g0169(.A(G179), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n345), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n369), .A2(new_n364), .A3(new_n371), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n367), .A2(new_n368), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n351), .A2(G77), .ZN(new_n374));
  XOR2_X1   g0174(.A(KEYINPUT15), .B(G87), .Z(new_n375));
  INV_X1    g0175(.A(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n362), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  OAI22_X1  g0178(.A1(new_n360), .A2(new_n357), .B1(new_n227), .B2(new_n204), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n253), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  OAI211_X1 g0180(.A(new_n374), .B(new_n380), .C1(G77), .C2(new_n354), .ZN(new_n381));
  AOI21_X1  g0181(.A(G45), .B1(new_n288), .B2(new_n290), .ZN(new_n382));
  INV_X1    g0182(.A(G274), .ZN(new_n383));
  NOR3_X1   g0183(.A1(new_n382), .A2(G1), .A3(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n384), .B1(new_n344), .B2(new_n219), .ZN(new_n385));
  NAND2_X1  g0185(.A1(G238), .A2(G1698), .ZN(new_n386));
  OAI211_X1 g0186(.A(new_n335), .B(new_n386), .C1(new_n215), .C2(G1698), .ZN(new_n387));
  OAI211_X1 g0187(.A(new_n387), .B(new_n316), .C1(G107), .C2(new_n335), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n385), .A2(new_n388), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n381), .B1(new_n389), .B2(G200), .ZN(new_n390));
  XNOR2_X1  g0190(.A(new_n390), .B(KEYINPUT74), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n385), .A2(new_n388), .A3(G190), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n373), .A2(new_n394), .ZN(new_n395));
  XNOR2_X1  g0195(.A(G58), .B(G68), .ZN(new_n396));
  AOI22_X1  g0196(.A1(new_n396), .A2(G20), .B1(G159), .B2(new_n356), .ZN(new_n397));
  AOI21_X1  g0197(.A(KEYINPUT7), .B1(new_n313), .B2(new_n227), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n299), .A2(KEYINPUT78), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n297), .A2(KEYINPUT3), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n399), .A2(new_n400), .A3(new_n267), .ZN(new_n401));
  AOI21_X1  g0201(.A(G20), .B1(new_n401), .B2(new_n312), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n398), .B1(new_n402), .B2(KEYINPUT7), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n397), .B1(new_n403), .B2(new_n203), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT16), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  XOR2_X1   g0206(.A(KEYINPUT79), .B(KEYINPUT7), .Z(new_n407));
  AND2_X1   g0207(.A1(new_n307), .A2(new_n308), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n267), .B1(new_n399), .B2(new_n400), .ZN(new_n409));
  OAI211_X1 g0209(.A(new_n227), .B(new_n407), .C1(new_n408), .C2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(KEYINPUT79), .A2(KEYINPUT7), .ZN(new_n411));
  AOI21_X1  g0211(.A(G20), .B1(new_n301), .B2(new_n309), .ZN(new_n412));
  OAI211_X1 g0212(.A(new_n410), .B(G68), .C1(new_n411), .C2(new_n412), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n413), .A2(KEYINPUT16), .A3(new_n397), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n406), .A2(new_n414), .A3(new_n253), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n337), .A2(new_n303), .ZN(new_n416));
  OR2_X1    g0216(.A1(new_n303), .A2(G226), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n301), .A2(new_n309), .A3(new_n416), .A4(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(G33), .A2(G87), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(new_n316), .ZN(new_n421));
  INV_X1    g0221(.A(G190), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n384), .B1(new_n344), .B2(G232), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n421), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n294), .B1(new_n418), .B2(new_n419), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n353), .A2(G45), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n353), .A2(G41), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n426), .A2(new_n427), .A3(G232), .A4(new_n294), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(new_n341), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n346), .B1(new_n425), .B2(new_n429), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n424), .A2(new_n430), .A3(KEYINPUT80), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n361), .A2(new_n354), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n432), .B1(new_n351), .B2(new_n361), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n425), .A2(new_n429), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT80), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n434), .A2(new_n435), .A3(new_n422), .ZN(new_n436));
  AND4_X1   g0236(.A1(new_n415), .A2(new_n431), .A3(new_n433), .A4(new_n436), .ZN(new_n437));
  XNOR2_X1  g0237(.A(KEYINPUT81), .B(KEYINPUT17), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n415), .A2(new_n431), .A3(new_n433), .A4(new_n436), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT81), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n441), .A2(KEYINPUT17), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n415), .A2(new_n433), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n434), .A2(G179), .ZN(new_n445));
  OAI21_X1  g0245(.A(G169), .B1(new_n425), .B2(new_n429), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  AND3_X1   g0247(.A1(new_n444), .A2(KEYINPUT18), .A3(new_n447), .ZN(new_n448));
  AOI21_X1  g0248(.A(KEYINPUT18), .B1(new_n444), .B2(new_n447), .ZN(new_n449));
  OAI211_X1 g0249(.A(new_n439), .B(new_n443), .C1(new_n448), .C2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(KEYINPUT82), .ZN(new_n452));
  NOR2_X1   g0252(.A1(G226), .A2(G1698), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n453), .B1(new_n215), .B2(G1698), .ZN(new_n454));
  AOI22_X1  g0254(.A1(new_n335), .A2(new_n454), .B1(G33), .B2(G97), .ZN(new_n455));
  OR2_X1    g0255(.A1(new_n455), .A2(new_n294), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT13), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n344), .A2(G238), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n456), .A2(new_n457), .A3(new_n458), .A4(new_n341), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n341), .B1(new_n455), .B2(new_n294), .ZN(new_n460));
  NOR4_X1   g0260(.A1(new_n285), .A2(new_n343), .A3(new_n216), .A4(new_n316), .ZN(new_n461));
  OAI21_X1  g0261(.A(KEYINPUT13), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n459), .A2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT14), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n465), .A2(KEYINPUT76), .ZN(new_n466));
  NOR3_X1   g0266(.A1(new_n464), .A2(new_n283), .A3(new_n466), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n463), .A2(new_n370), .ZN(new_n468));
  INV_X1    g0268(.A(new_n466), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n469), .B1(new_n463), .B2(G169), .ZN(new_n470));
  NOR3_X1   g0270(.A1(new_n467), .A2(new_n468), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n280), .A2(new_n203), .ZN(new_n472));
  XNOR2_X1  g0272(.A(new_n472), .B(KEYINPUT12), .ZN(new_n473));
  OAI22_X1  g0273(.A1(new_n377), .A2(new_n204), .B1(new_n227), .B2(G68), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n357), .A2(new_n201), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n253), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT11), .ZN(new_n477));
  OR2_X1    g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n476), .A2(new_n477), .B1(G68), .B2(new_n351), .ZN(new_n479));
  AND3_X1   g0279(.A1(new_n473), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  OR2_X1    g0280(.A1(new_n471), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n464), .A2(G190), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n482), .B(new_n480), .C1(new_n346), .C2(new_n464), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n389), .A2(new_n283), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n385), .A2(new_n388), .A3(new_n370), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n484), .A2(new_n381), .A3(new_n485), .ZN(new_n486));
  AND3_X1   g0286(.A1(new_n481), .A2(new_n483), .A3(new_n486), .ZN(new_n487));
  OR2_X1    g0287(.A1(new_n451), .A2(KEYINPUT82), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n395), .A2(new_n452), .A3(new_n487), .A4(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(G87), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n491), .A2(G20), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n301), .A2(KEYINPUT22), .A3(new_n309), .A4(new_n492), .ZN(new_n493));
  OR3_X1    g0293(.A1(new_n227), .A2(KEYINPUT23), .A3(G107), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n362), .A2(G116), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT22), .ZN(new_n496));
  INV_X1    g0296(.A(new_n492), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n496), .B1(new_n313), .B2(new_n497), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n493), .A2(new_n494), .A3(new_n495), .A4(new_n498), .ZN(new_n499));
  OAI22_X1  g0299(.A1(new_n227), .A2(G107), .B1(KEYINPUT86), .B2(KEYINPUT23), .ZN(new_n500));
  AND2_X1   g0300(.A1(KEYINPUT86), .A2(KEYINPUT23), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT87), .ZN(new_n502));
  OR3_X1    g0302(.A1(new_n500), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n502), .B1(new_n500), .B2(new_n501), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(new_n505), .ZN(new_n506));
  OAI21_X1  g0306(.A(KEYINPUT24), .B1(new_n499), .B2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(new_n507), .ZN(new_n508));
  NOR3_X1   g0308(.A1(new_n499), .A2(new_n506), .A3(KEYINPUT24), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n253), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT25), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n511), .B1(new_n354), .B2(G107), .ZN(new_n512));
  INV_X1    g0312(.A(G107), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n280), .A2(KEYINPUT25), .A3(new_n513), .ZN(new_n514));
  AOI22_X1  g0314(.A1(new_n277), .A2(G107), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  OR2_X1    g0315(.A1(G250), .A2(G1698), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n302), .A2(G1698), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n301), .A2(new_n309), .A3(new_n516), .A4(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(G33), .A2(G294), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n316), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n293), .A2(G264), .A3(new_n294), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n521), .A2(KEYINPUT88), .A3(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT88), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n294), .B1(new_n518), .B2(new_n519), .ZN(new_n525));
  AND3_X1   g0325(.A1(new_n293), .A2(G264), .A3(new_n294), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n316), .A2(new_n383), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n528), .A2(new_n285), .A3(new_n287), .A4(new_n292), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n523), .A2(new_n527), .A3(G179), .A4(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n521), .A2(new_n529), .A3(new_n522), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(G169), .ZN(new_n532));
  AOI22_X1  g0332(.A1(new_n510), .A2(new_n515), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(new_n515), .ZN(new_n534));
  INV_X1    g0334(.A(new_n509), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n507), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n534), .B1(new_n536), .B2(new_n253), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n523), .A2(new_n529), .A3(new_n527), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n346), .ZN(new_n539));
  NOR4_X1   g0339(.A1(new_n525), .A2(new_n526), .A3(G190), .A4(new_n296), .ZN(new_n540));
  INV_X1    g0340(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n533), .B1(new_n537), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n513), .A2(KEYINPUT6), .A3(G97), .ZN(new_n544));
  XOR2_X1   g0344(.A(G97), .B(G107), .Z(new_n545));
  OAI21_X1  g0345(.A(new_n544), .B1(new_n545), .B2(KEYINPUT6), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(G20), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n356), .A2(G77), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n547), .B(new_n548), .C1(new_n403), .C2(new_n513), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n253), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n354), .A2(G97), .ZN(new_n551));
  INV_X1    g0351(.A(new_n551), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n552), .B1(new_n276), .B2(new_n257), .ZN(new_n553));
  INV_X1    g0353(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n550), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n293), .A2(G257), .A3(new_n294), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(new_n529), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n301), .A2(G244), .A3(new_n309), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT4), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(G250), .ZN(new_n561));
  OAI21_X1  g0361(.A(KEYINPUT4), .B1(new_n313), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(G1698), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n559), .A2(G1698), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n564), .A2(new_n311), .A3(new_n312), .A4(G244), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n256), .ZN(new_n566));
  INV_X1    g0366(.A(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n560), .A2(new_n563), .A3(new_n567), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n557), .B1(new_n568), .B2(new_n316), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n370), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n566), .B1(new_n558), .B2(new_n559), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n294), .B1(new_n571), .B2(new_n563), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n283), .B1(new_n572), .B2(new_n557), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n555), .A2(new_n570), .A3(new_n573), .ZN(new_n574));
  OAI21_X1  g0374(.A(G200), .B1(new_n572), .B2(new_n557), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n553), .B1(new_n549), .B2(new_n253), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n568), .A2(new_n316), .ZN(new_n577));
  INV_X1    g0377(.A(new_n557), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n575), .B(new_n576), .C1(new_n579), .C2(new_n422), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n574), .A2(new_n580), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n301), .A2(new_n227), .A3(G68), .A4(new_n309), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT19), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n362), .A2(new_n583), .A3(G97), .ZN(new_n584));
  AOI21_X1  g0384(.A(G20), .B1(G33), .B2(G97), .ZN(new_n585));
  NOR2_X1   g0385(.A1(G97), .A2(G107), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n585), .B1(new_n491), .B2(new_n586), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n584), .B1(new_n587), .B2(new_n583), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n582), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(new_n253), .ZN(new_n590));
  INV_X1    g0390(.A(new_n272), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n275), .A2(new_n354), .A3(new_n591), .A4(new_n375), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT84), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n354), .A2(new_n375), .ZN(new_n595));
  INV_X1    g0395(.A(new_n595), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n274), .A2(KEYINPUT84), .A3(new_n275), .A4(new_n375), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n590), .A2(new_n594), .A3(new_n596), .A4(new_n597), .ZN(new_n598));
  XNOR2_X1  g0398(.A(KEYINPUT71), .B(G1), .ZN(new_n599));
  OAI211_X1 g0399(.A(G250), .B(new_n294), .C1(new_n599), .C2(new_n284), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(KEYINPUT83), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n528), .A2(new_n285), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT83), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n426), .A2(new_n603), .A3(G250), .A4(new_n294), .ZN(new_n604));
  AND3_X1   g0404(.A1(new_n601), .A2(new_n602), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n216), .A2(new_n303), .ZN(new_n606));
  OR2_X1    g0406(.A1(new_n303), .A2(G244), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n301), .A2(new_n309), .A3(new_n606), .A4(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(G33), .A2(G116), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n316), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n605), .A2(new_n611), .A3(new_n370), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n601), .A2(new_n604), .A3(new_n602), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n294), .B1(new_n608), .B2(new_n609), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n283), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n598), .A2(new_n612), .A3(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n605), .A2(new_n611), .A3(G190), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n275), .B1(new_n582), .B2(new_n588), .ZN(new_n618));
  NOR4_X1   g0418(.A1(new_n280), .A2(new_n253), .A3(new_n272), .A4(new_n491), .ZN(new_n619));
  NOR3_X1   g0419(.A1(new_n618), .A2(new_n619), .A3(new_n595), .ZN(new_n620));
  OAI21_X1  g0420(.A(G200), .B1(new_n613), .B2(new_n614), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n617), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n616), .A2(new_n622), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n581), .A2(new_n623), .ZN(new_n624));
  AND4_X1   g0424(.A1(new_n334), .A2(new_n490), .A3(new_n543), .A4(new_n624), .ZN(G372));
  INV_X1    g0425(.A(new_n372), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n448), .A2(new_n449), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n471), .A2(new_n480), .ZN(new_n629));
  INV_X1    g0429(.A(new_n486), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n629), .B1(new_n483), .B2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(new_n438), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n443), .B1(new_n440), .B2(new_n632), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n628), .B1(new_n631), .B2(new_n633), .ZN(new_n634));
  AND2_X1   g0434(.A1(new_n367), .A2(new_n368), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n626), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n613), .A2(KEYINPUT89), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT89), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n601), .A2(new_n604), .A3(new_n638), .A4(new_n602), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n637), .A2(new_n611), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(G200), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n641), .A2(new_n617), .A3(new_n620), .ZN(new_n642));
  AND2_X1   g0442(.A1(new_n598), .A2(new_n612), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n640), .A2(new_n283), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n510), .A2(new_n515), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n540), .B1(new_n538), .B2(new_n346), .ZN(new_n647));
  OAI211_X1 g0447(.A(new_n642), .B(new_n645), .C1(new_n646), .C2(new_n647), .ZN(new_n648));
  OAI21_X1  g0448(.A(KEYINPUT90), .B1(new_n648), .B2(new_n581), .ZN(new_n649));
  INV_X1    g0449(.A(new_n581), .ZN(new_n650));
  AND2_X1   g0450(.A1(new_n642), .A2(new_n645), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n542), .A2(new_n537), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT90), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n650), .A2(new_n651), .A3(new_n652), .A4(new_n653), .ZN(new_n654));
  AND2_X1   g0454(.A1(new_n324), .A2(new_n327), .ZN(new_n655));
  INV_X1    g0455(.A(new_n533), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n655), .A2(new_n656), .A3(new_n321), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n649), .A2(new_n654), .A3(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT26), .ZN(new_n659));
  INV_X1    g0459(.A(new_n574), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n651), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(KEYINPUT26), .B1(new_n574), .B2(new_n623), .ZN(new_n662));
  AND3_X1   g0462(.A1(new_n661), .A2(new_n645), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n658), .A2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n636), .B1(new_n489), .B2(new_n665), .ZN(G369));
  INV_X1    g0466(.A(G330), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n655), .A2(new_n321), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n279), .A2(G20), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  OR3_X1    g0470(.A1(new_n599), .A2(new_n670), .A3(KEYINPUT27), .ZN(new_n671));
  OAI21_X1  g0471(.A(KEYINPUT27), .B1(new_n599), .B2(new_n670), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n671), .A2(new_n672), .A3(G213), .ZN(new_n673));
  INV_X1    g0473(.A(G343), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n282), .A2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n668), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n334), .A2(new_n676), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(KEYINPUT91), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT91), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n678), .A2(new_n682), .A3(new_n679), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n667), .B1(new_n681), .B2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n675), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n543), .B1(new_n537), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n533), .A2(new_n675), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n684), .A2(KEYINPUT92), .A3(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  AOI21_X1  g0490(.A(KEYINPUT92), .B1(new_n684), .B2(new_n688), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n668), .A2(new_n685), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n693), .A2(KEYINPUT93), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT93), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n695), .B1(new_n668), .B2(new_n685), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n688), .B1(new_n694), .B2(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n656), .A2(new_n675), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n692), .A2(new_n701), .ZN(G399));
  INV_X1    g0502(.A(new_n209), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n340), .A2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(G1), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n586), .A2(new_n491), .A3(new_n254), .ZN(new_n707));
  OAI22_X1  g0507(.A1(new_n706), .A2(new_n707), .B1(new_n230), .B2(new_n705), .ZN(new_n708));
  XNOR2_X1  g0508(.A(new_n708), .B(KEYINPUT28), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n659), .B1(new_n574), .B2(new_n623), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(KEYINPUT95), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n660), .A2(new_n642), .A3(KEYINPUT26), .A4(new_n645), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT95), .ZN(new_n713));
  OAI211_X1 g0513(.A(new_n713), .B(new_n659), .C1(new_n574), .C2(new_n623), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n711), .A2(new_n712), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(new_n645), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(KEYINPUT96), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n657), .A2(new_n652), .A3(new_n650), .A4(new_n651), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT96), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n715), .A2(new_n719), .A3(new_n645), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n717), .A2(new_n718), .A3(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n721), .A2(KEYINPUT29), .A3(new_n685), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n664), .A2(new_n685), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT29), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n723), .A2(KEYINPUT94), .A3(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT94), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n675), .B1(new_n658), .B2(new_n663), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n726), .B1(new_n727), .B2(KEYINPUT29), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n722), .A2(new_n725), .A3(new_n728), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n543), .A2(new_n334), .A3(new_n624), .A4(new_n685), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n317), .A2(G179), .A3(new_n319), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n579), .A2(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n613), .A2(new_n614), .ZN(new_n733));
  AND3_X1   g0533(.A1(new_n523), .A2(new_n527), .A3(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n732), .A2(new_n734), .A3(KEYINPUT30), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT30), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n569), .A2(G179), .A3(new_n326), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n523), .A2(new_n527), .A3(new_n733), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n736), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n735), .A2(new_n739), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n538), .A2(new_n370), .A3(new_n328), .A4(new_n640), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n741), .A2(new_n569), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n675), .B1(new_n740), .B2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT31), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  OAI211_X1 g0545(.A(KEYINPUT31), .B(new_n675), .C1(new_n740), .C2(new_n742), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n730), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(G330), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n729), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n709), .B1(new_n750), .B2(G1), .ZN(G364));
  NOR2_X1   g0551(.A1(G13), .A2(G33), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n753), .A2(G20), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n681), .A2(new_n683), .A3(new_n754), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n226), .B1(G20), .B2(new_n283), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n408), .A2(new_n409), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(new_n703), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n244), .A2(new_n284), .ZN(new_n761));
  AOI211_X1 g0561(.A(new_n760), .B(new_n761), .C1(new_n284), .C2(new_n231), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n335), .A2(G355), .A3(new_n209), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n763), .B1(G116), .B2(new_n209), .ZN(new_n764));
  XOR2_X1   g0564(.A(new_n764), .B(KEYINPUT97), .Z(new_n765));
  OAI21_X1  g0565(.A(new_n757), .B1(new_n762), .B2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n422), .A2(G200), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(new_n370), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(G20), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(G294), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n422), .A2(new_n346), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n227), .A2(G179), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(G303), .ZN(new_n777));
  NAND2_X1  g0577(.A1(G20), .A2(G179), .ZN(new_n778));
  XOR2_X1   g0578(.A(new_n778), .B(KEYINPUT98), .Z(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(new_n422), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(new_n346), .ZN(new_n781));
  XNOR2_X1  g0581(.A(KEYINPUT33), .B(G317), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n774), .A2(new_n422), .A3(G200), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(G283), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n779), .A2(new_n773), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(G326), .ZN(new_n789));
  AND4_X1   g0589(.A1(new_n777), .A2(new_n783), .A3(new_n786), .A4(new_n789), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n774), .A2(new_n422), .A3(new_n346), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n335), .B1(new_n792), .B2(G329), .ZN(new_n793));
  INV_X1    g0593(.A(G311), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n780), .A2(G200), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  OAI211_X1 g0596(.A(new_n790), .B(new_n793), .C1(new_n794), .C2(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n779), .A2(new_n767), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  AOI211_X1 g0599(.A(new_n772), .B(new_n797), .C1(G322), .C2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n781), .ZN(new_n801));
  OAI22_X1  g0601(.A1(new_n801), .A2(new_n203), .B1(new_n798), .B2(new_n202), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  OAI221_X1 g0603(.A(new_n803), .B1(new_n201), .B2(new_n787), .C1(new_n204), .C2(new_n796), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n770), .A2(new_n257), .ZN(new_n805));
  OAI221_X1 g0605(.A(new_n335), .B1(new_n775), .B2(new_n491), .C1(new_n513), .C2(new_n784), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n792), .A2(G159), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n807), .B(KEYINPUT32), .ZN(new_n808));
  NOR4_X1   g0608(.A1(new_n804), .A2(new_n805), .A3(new_n806), .A4(new_n808), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n756), .B1(new_n800), .B2(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n669), .A2(G45), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n705), .A2(G1), .A3(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  NAND4_X1  g0613(.A1(new_n755), .A2(new_n766), .A3(new_n810), .A4(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n681), .A2(new_n683), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n815), .A2(G330), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(new_n812), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n815), .A2(G330), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n814), .B1(new_n817), .B2(new_n818), .ZN(G396));
  NAND2_X1  g0619(.A1(new_n785), .A2(G87), .ZN(new_n820));
  INV_X1    g0620(.A(G303), .ZN(new_n821));
  OAI221_X1 g0621(.A(new_n820), .B1(new_n821), .B2(new_n787), .C1(new_n796), .C2(new_n254), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(G283), .ZN(new_n824));
  OAI221_X1 g0624(.A(new_n313), .B1(new_n794), .B2(new_n791), .C1(new_n801), .C2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n799), .A2(G294), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n805), .B1(G107), .B2(new_n776), .ZN(new_n828));
  NAND4_X1  g0628(.A1(new_n823), .A2(new_n826), .A3(new_n827), .A4(new_n828), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n775), .A2(new_n201), .ZN(new_n830));
  INV_X1    g0630(.A(G143), .ZN(new_n831));
  OAI22_X1  g0631(.A1(new_n801), .A2(new_n355), .B1(new_n798), .B2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(G137), .ZN(new_n834));
  INV_X1    g0634(.A(G159), .ZN(new_n835));
  OAI221_X1 g0635(.A(new_n833), .B1(new_n834), .B2(new_n787), .C1(new_n835), .C2(new_n796), .ZN(new_n836));
  XOR2_X1   g0636(.A(new_n836), .B(KEYINPUT34), .Z(new_n837));
  AOI211_X1 g0637(.A(new_n830), .B(new_n837), .C1(G132), .C2(new_n792), .ZN(new_n838));
  OAI221_X1 g0638(.A(new_n838), .B1(new_n202), .B2(new_n770), .C1(new_n203), .C2(new_n784), .ZN(new_n839));
  INV_X1    g0639(.A(new_n758), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n829), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  XNOR2_X1  g0641(.A(new_n486), .B(KEYINPUT100), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n393), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n381), .A2(new_n675), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  OAI22_X1  g0645(.A1(new_n843), .A2(new_n845), .B1(new_n486), .B2(new_n685), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  AOI22_X1  g0647(.A1(new_n841), .A2(new_n756), .B1(new_n752), .B2(new_n847), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n756), .A2(new_n752), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n812), .B1(new_n204), .B2(new_n849), .ZN(new_n850));
  XNOR2_X1  g0650(.A(new_n850), .B(KEYINPUT99), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n848), .A2(new_n851), .ZN(new_n852));
  AOI211_X1 g0652(.A(new_n675), .B(new_n843), .C1(new_n658), .C2(new_n663), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n853), .B1(new_n723), .B2(new_n847), .ZN(new_n854));
  XNOR2_X1  g0654(.A(new_n854), .B(new_n748), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(new_n812), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n852), .A2(new_n856), .ZN(G384));
  NAND4_X1  g0657(.A1(new_n490), .A2(new_n722), .A3(new_n728), .A4(new_n725), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(new_n636), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n413), .A2(new_n397), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(new_n405), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n861), .A2(new_n253), .A3(new_n414), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n673), .B1(new_n862), .B2(new_n433), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n863), .B1(new_n627), .B2(new_n633), .ZN(new_n864));
  INV_X1    g0664(.A(new_n447), .ZN(new_n865));
  AOI22_X1  g0665(.A1(new_n865), .A2(new_n673), .B1(new_n862), .B2(new_n433), .ZN(new_n866));
  OAI21_X1  g0666(.A(KEYINPUT37), .B1(new_n866), .B2(new_n437), .ZN(new_n867));
  XNOR2_X1  g0667(.A(new_n673), .B(KEYINPUT102), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n444), .B1(new_n447), .B2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT37), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n869), .A2(new_n870), .A3(new_n440), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n867), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(KEYINPUT38), .B1(new_n864), .B2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(new_n873), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n864), .A2(KEYINPUT38), .A3(new_n872), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n629), .A2(new_n675), .ZN(new_n877));
  OR2_X1    g0677(.A1(new_n480), .A2(new_n685), .ZN(new_n878));
  OAI211_X1 g0678(.A(new_n483), .B(new_n878), .C1(new_n471), .C2(new_n480), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n842), .A2(new_n675), .ZN(new_n881));
  OAI211_X1 g0681(.A(new_n876), .B(new_n880), .C1(new_n853), .C2(new_n881), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n874), .A2(KEYINPUT39), .A3(new_n875), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT39), .ZN(new_n884));
  AND3_X1   g0684(.A1(new_n864), .A2(KEYINPUT38), .A3(new_n872), .ZN(new_n885));
  XOR2_X1   g0685(.A(KEYINPUT103), .B(KEYINPUT38), .Z(new_n886));
  INV_X1    g0686(.A(new_n886), .ZN(new_n887));
  AND2_X1   g0687(.A1(new_n444), .A2(new_n868), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n450), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n869), .A2(new_n440), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(KEYINPUT37), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(new_n871), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n887), .B1(new_n889), .B2(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n884), .B1(new_n885), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n629), .A2(new_n685), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n883), .A2(new_n894), .A3(new_n896), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n628), .A2(new_n868), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  AND3_X1   g0699(.A1(new_n882), .A2(new_n897), .A3(new_n899), .ZN(new_n900));
  XNOR2_X1  g0700(.A(new_n859), .B(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT104), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n902), .B1(new_n885), .B2(new_n893), .ZN(new_n903));
  AND3_X1   g0703(.A1(new_n747), .A2(new_n880), .A3(new_n846), .ZN(new_n904));
  AOI22_X1  g0704(.A1(new_n450), .A2(new_n888), .B1(new_n891), .B2(new_n871), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n875), .B(KEYINPUT104), .C1(new_n905), .C2(new_n887), .ZN(new_n906));
  NAND4_X1  g0706(.A1(new_n903), .A2(KEYINPUT40), .A3(new_n904), .A4(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT40), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n885), .A2(new_n873), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n747), .A2(new_n880), .A3(new_n846), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n908), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n907), .A2(G330), .A3(new_n911), .ZN(new_n912));
  OR2_X1    g0712(.A1(new_n489), .A2(new_n748), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n907), .A2(new_n747), .A3(new_n911), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n914), .B1(new_n489), .B2(new_n915), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n901), .B(new_n916), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n917), .B1(new_n353), .B2(new_n669), .ZN(new_n918));
  XOR2_X1   g0718(.A(new_n546), .B(KEYINPUT101), .Z(new_n919));
  AOI21_X1  g0719(.A(new_n254), .B1(new_n919), .B2(KEYINPUT35), .ZN(new_n920));
  OAI211_X1 g0720(.A(new_n920), .B(new_n229), .C1(KEYINPUT35), .C2(new_n919), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n921), .B(KEYINPUT36), .ZN(new_n922));
  OAI21_X1  g0722(.A(G77), .B1(new_n202), .B2(new_n203), .ZN(new_n923));
  OAI22_X1  g0723(.A1(new_n923), .A2(new_n230), .B1(G50), .B2(new_n203), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n924), .A2(new_n279), .A3(new_n599), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n918), .A2(new_n922), .A3(new_n925), .ZN(G367));
  OAI221_X1 g0726(.A(new_n757), .B1(new_n209), .B2(new_n376), .C1(new_n240), .C2(new_n760), .ZN(new_n927));
  OAI221_X1 g0727(.A(new_n335), .B1(new_n834), .B2(new_n791), .C1(new_n787), .C2(new_n831), .ZN(new_n928));
  AOI22_X1  g0728(.A1(new_n795), .A2(G50), .B1(G77), .B2(new_n785), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n769), .A2(G68), .ZN(new_n930));
  OAI211_X1 g0730(.A(new_n929), .B(new_n930), .C1(new_n835), .C2(new_n801), .ZN(new_n931));
  AOI211_X1 g0731(.A(new_n928), .B(new_n931), .C1(G58), .C2(new_n776), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(new_n355), .B2(new_n798), .ZN(new_n933));
  XOR2_X1   g0733(.A(new_n933), .B(KEYINPUT108), .Z(new_n934));
  AOI22_X1  g0734(.A1(new_n795), .A2(G283), .B1(G107), .B2(new_n769), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(KEYINPUT107), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n785), .A2(G97), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n936), .A2(new_n840), .A3(new_n937), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n775), .A2(new_n254), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n939), .B(KEYINPUT46), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n792), .A2(G317), .ZN(new_n941));
  OAI221_X1 g0741(.A(new_n941), .B1(new_n821), .B2(new_n798), .C1(new_n801), .C2(new_n771), .ZN(new_n942));
  NOR3_X1   g0742(.A1(new_n938), .A2(new_n940), .A3(new_n942), .ZN(new_n943));
  OAI221_X1 g0743(.A(new_n943), .B1(KEYINPUT107), .B2(new_n935), .C1(new_n794), .C2(new_n787), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n934), .A2(new_n944), .ZN(new_n945));
  XOR2_X1   g0745(.A(new_n945), .B(KEYINPUT47), .Z(new_n946));
  INV_X1    g0746(.A(new_n756), .ZN(new_n947));
  OAI211_X1 g0747(.A(new_n813), .B(new_n927), .C1(new_n946), .C2(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n651), .B1(new_n620), .B2(new_n685), .ZN(new_n949));
  OR3_X1    g0749(.A1(new_n645), .A2(new_n620), .A3(new_n685), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NOR3_X1   g0751(.A1(new_n951), .A2(G20), .A3(new_n753), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n948), .A2(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n650), .B1(new_n576), .B2(new_n685), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n660), .A2(new_n675), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n697), .A2(new_n957), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n958), .B(KEYINPUT42), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n574), .B1(new_n954), .B2(new_n656), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(new_n685), .ZN(new_n961));
  AOI22_X1  g0761(.A1(new_n959), .A2(new_n961), .B1(KEYINPUT43), .B2(new_n951), .ZN(new_n962));
  OR2_X1    g0762(.A1(new_n951), .A2(KEYINPUT43), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n962), .B(new_n963), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n692), .A2(new_n957), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n964), .B(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT44), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(KEYINPUT105), .ZN(new_n968));
  AND3_X1   g0768(.A1(new_n700), .A2(new_n957), .A3(new_n968), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n967), .A2(KEYINPUT105), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n697), .A2(new_n699), .A3(new_n956), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT45), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND4_X1  g0774(.A1(new_n697), .A2(KEYINPUT45), .A3(new_n699), .A4(new_n956), .ZN(new_n975));
  AOI22_X1  g0775(.A1(new_n969), .A2(new_n971), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(KEYINPUT106), .B1(new_n690), .B2(new_n691), .ZN(new_n977));
  INV_X1    g0777(.A(new_n691), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT106), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n978), .A2(new_n979), .A3(new_n689), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n970), .B1(new_n701), .B2(new_n956), .ZN(new_n981));
  NAND4_X1  g0781(.A1(new_n976), .A2(new_n977), .A3(new_n980), .A4(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n974), .A2(new_n975), .ZN(new_n983));
  NAND4_X1  g0783(.A1(new_n700), .A2(new_n971), .A3(new_n957), .A4(new_n968), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n983), .A2(new_n981), .A3(new_n984), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n985), .A2(new_n979), .A3(new_n692), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n982), .A2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n688), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n816), .A2(new_n988), .ZN(new_n989));
  OR2_X1    g0789(.A1(new_n694), .A2(new_n696), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n815), .A2(G330), .A3(new_n688), .ZN(new_n991));
  AND3_X1   g0791(.A1(new_n989), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n990), .B1(new_n989), .B2(new_n991), .ZN(new_n993));
  NOR3_X1   g0793(.A1(new_n992), .A2(new_n749), .A3(new_n993), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n749), .B1(new_n987), .B2(new_n994), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n704), .B(KEYINPUT41), .ZN(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  OAI211_X1 g0797(.A(G1), .B(new_n811), .C1(new_n995), .C2(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n953), .B1(new_n966), .B2(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(new_n999), .ZN(G387));
  NOR2_X1   g0800(.A1(new_n992), .A2(new_n993), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n811), .A2(G1), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  XOR2_X1   g0803(.A(new_n1003), .B(KEYINPUT109), .Z(new_n1004));
  NOR2_X1   g0804(.A1(new_n775), .A2(new_n204), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n937), .B1(new_n787), .B2(new_n835), .ZN(new_n1006));
  AOI211_X1 g0806(.A(new_n1005), .B(new_n1006), .C1(new_n361), .C2(new_n781), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n792), .A2(G150), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n769), .A2(new_n375), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1009), .B1(new_n798), .B2(new_n201), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT110), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n840), .B1(new_n795), .B2(G68), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n1007), .A2(new_n1008), .A3(new_n1011), .A4(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(G317), .ZN(new_n1014));
  OAI22_X1  g0814(.A1(new_n801), .A2(new_n794), .B1(new_n798), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(G322), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n1016), .B1(new_n821), .B2(new_n796), .C1(new_n1017), .C2(new_n787), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT48), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n1019), .B1(new_n824), .B2(new_n770), .C1(new_n771), .C2(new_n775), .ZN(new_n1020));
  XOR2_X1   g0820(.A(new_n1020), .B(KEYINPUT49), .Z(new_n1021));
  AOI21_X1  g0821(.A(new_n758), .B1(G326), .B2(new_n792), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1022), .B1(new_n254), .B2(new_n784), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1013), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1024), .A2(new_n756), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n360), .A2(G50), .ZN(new_n1026));
  XOR2_X1   g0826(.A(new_n1026), .B(KEYINPUT50), .Z(new_n1027));
  NOR2_X1   g0827(.A1(new_n203), .A2(new_n204), .ZN(new_n1028));
  NOR4_X1   g0828(.A1(new_n1027), .A2(G45), .A3(new_n1028), .A4(new_n707), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n759), .B1(new_n236), .B2(new_n284), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n335), .A2(new_n707), .A3(new_n209), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1029), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n209), .A2(G107), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n757), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n812), .B1(new_n988), .B2(new_n754), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1025), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n1001), .A2(new_n750), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1001), .A2(new_n750), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1038), .A2(new_n704), .ZN(new_n1039));
  OAI211_X1 g0839(.A(new_n1004), .B(new_n1036), .C1(new_n1037), .C2(new_n1039), .ZN(G393));
  INV_X1    g0840(.A(KEYINPUT111), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n987), .A2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n982), .A2(new_n986), .A3(KEYINPUT111), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1042), .A2(new_n1002), .A3(new_n1043), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n770), .A2(new_n254), .B1(new_n775), .B2(new_n824), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n794), .A2(new_n798), .B1(new_n787), .B2(new_n1014), .ZN(new_n1046));
  XOR2_X1   g0846(.A(new_n1046), .B(KEYINPUT52), .Z(new_n1047));
  AOI211_X1 g0847(.A(new_n1045), .B(new_n1047), .C1(G322), .C2(new_n792), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n1048), .B(new_n313), .C1(new_n513), .C2(new_n784), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1049), .B1(G294), .B2(new_n795), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1050), .B1(new_n821), .B2(new_n801), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT114), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n201), .A2(new_n801), .B1(new_n796), .B2(new_n360), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT113), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n820), .B1(new_n203), .B2(new_n775), .C1(new_n831), .C2(new_n791), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1055), .B1(G77), .B2(new_n769), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n355), .A2(new_n787), .B1(new_n798), .B2(new_n835), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1057), .B(KEYINPUT51), .ZN(new_n1058));
  AND4_X1   g0858(.A1(new_n758), .A2(new_n1054), .A3(new_n1056), .A4(new_n1058), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n756), .B1(new_n1052), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n957), .A2(new_n754), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n757), .B1(new_n257), .B2(new_n209), .C1(new_n760), .C2(new_n247), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1062), .A2(new_n813), .ZN(new_n1063));
  XOR2_X1   g0863(.A(new_n1063), .B(KEYINPUT112), .Z(new_n1064));
  NAND3_X1  g0864(.A1(new_n1060), .A2(new_n1061), .A3(new_n1064), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1038), .A2(new_n982), .A3(new_n986), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1066), .A2(KEYINPUT115), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n987), .A2(new_n994), .ZN(new_n1068));
  INV_X1    g0868(.A(KEYINPUT115), .ZN(new_n1069));
  NAND4_X1  g0869(.A1(new_n1038), .A2(new_n982), .A3(new_n986), .A4(new_n1069), .ZN(new_n1070));
  NAND4_X1  g0870(.A1(new_n1067), .A2(new_n704), .A3(new_n1068), .A4(new_n1070), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n1071), .A2(KEYINPUT116), .ZN(new_n1072));
  INV_X1    g0872(.A(KEYINPUT116), .ZN(new_n1073));
  AND2_X1   g0873(.A1(new_n1068), .A2(new_n1070), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n705), .B1(new_n1066), .B2(KEYINPUT115), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1073), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n1044), .B(new_n1065), .C1(new_n1072), .C2(new_n1076), .ZN(G390));
  NAND4_X1  g0877(.A1(new_n747), .A2(new_n880), .A3(new_n846), .A4(G330), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1078), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n903), .A2(new_n906), .A3(new_n895), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n843), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n721), .A2(new_n685), .A3(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n881), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1080), .B1(new_n1084), .B2(new_n880), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n880), .B1(new_n853), .B2(new_n881), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n1086), .A2(new_n895), .B1(new_n894), .B2(new_n883), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1079), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n883), .A2(new_n894), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n880), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n727), .A2(new_n1081), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1090), .B1(new_n1091), .B2(new_n1083), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1089), .B1(new_n1092), .B2(new_n896), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1090), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n1093), .B(new_n1078), .C1(new_n1094), .C2(new_n1080), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1088), .A2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n747), .A2(new_n846), .A3(G330), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1097), .A2(new_n1090), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(new_n1078), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1091), .A2(new_n1083), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(KEYINPUT117), .ZN(new_n1102));
  NAND4_X1  g0902(.A1(new_n1082), .A2(new_n1083), .A3(new_n1078), .A4(new_n1098), .ZN(new_n1103));
  INV_X1    g0903(.A(KEYINPUT117), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1099), .A2(new_n1104), .A3(new_n1100), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1102), .A2(new_n1103), .A3(new_n1105), .ZN(new_n1106));
  AND3_X1   g0906(.A1(new_n858), .A2(new_n636), .A3(new_n913), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1096), .A2(new_n1108), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n1088), .A2(new_n1095), .A3(new_n1107), .A4(new_n1106), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1109), .A2(new_n704), .A3(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1088), .A2(new_n1002), .A3(new_n1095), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1089), .A2(new_n752), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n849), .ZN(new_n1114));
  OR2_X1    g0914(.A1(new_n361), .A2(new_n1114), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n784), .A2(new_n201), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n775), .A2(new_n355), .ZN(new_n1117));
  XOR2_X1   g0917(.A(new_n1117), .B(KEYINPUT53), .Z(new_n1118));
  AOI211_X1 g0918(.A(new_n1116), .B(new_n1118), .C1(G128), .C2(new_n788), .ZN(new_n1119));
  OAI221_X1 g0919(.A(new_n1119), .B1(new_n834), .B2(new_n801), .C1(new_n835), .C2(new_n770), .ZN(new_n1120));
  AND2_X1   g0920(.A1(new_n792), .A2(G125), .ZN(new_n1121));
  XNOR2_X1  g0921(.A(KEYINPUT54), .B(G143), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n796), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(G132), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n335), .B1(new_n798), .B2(new_n1124), .ZN(new_n1125));
  NOR4_X1   g0925(.A1(new_n1120), .A2(new_n1121), .A3(new_n1123), .A4(new_n1125), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n792), .A2(G294), .B1(new_n776), .B2(G87), .ZN(new_n1127));
  OAI211_X1 g0927(.A(new_n1127), .B(new_n313), .C1(new_n254), .C2(new_n798), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n795), .A2(G97), .B1(G77), .B2(new_n769), .ZN(new_n1129));
  OAI221_X1 g0929(.A(new_n1129), .B1(new_n203), .B2(new_n784), .C1(new_n824), .C2(new_n787), .ZN(new_n1130));
  AOI211_X1 g0930(.A(new_n1128), .B(new_n1130), .C1(G107), .C2(new_n781), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n756), .B1(new_n1126), .B2(new_n1131), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n1113), .A2(new_n813), .A3(new_n1115), .A4(new_n1132), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1111), .A2(new_n1112), .A3(new_n1133), .ZN(G378));
  NAND2_X1  g0934(.A1(new_n1110), .A2(new_n1107), .ZN(new_n1135));
  INV_X1    g0935(.A(KEYINPUT120), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1110), .A2(KEYINPUT120), .A3(new_n1107), .ZN(new_n1138));
  INV_X1    g0938(.A(KEYINPUT119), .ZN(new_n1139));
  XOR2_X1   g0939(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1140));
  INV_X1    g0940(.A(new_n1140), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n635), .A2(new_n372), .A3(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n673), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n364), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n373), .A2(new_n1140), .ZN(new_n1146));
  AND3_X1   g0946(.A1(new_n1142), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1145), .B1(new_n1142), .B2(new_n1146), .ZN(new_n1148));
  OR2_X1    g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n912), .A2(new_n1149), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1151));
  NAND4_X1  g0951(.A1(new_n1151), .A2(new_n907), .A3(G330), .A4(new_n911), .ZN(new_n1152));
  AND3_X1   g0952(.A1(new_n1150), .A2(new_n1152), .A3(new_n900), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n900), .B1(new_n1150), .B2(new_n1152), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1139), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1150), .A2(new_n1152), .A3(new_n900), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1156), .A2(KEYINPUT119), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(new_n1137), .A2(new_n1138), .B1(new_n1155), .B2(new_n1157), .ZN(new_n1158));
  OAI21_X1  g0958(.A(KEYINPUT121), .B1(new_n1158), .B2(KEYINPUT57), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1160), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n705), .B1(new_n1161), .B2(KEYINPUT57), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1163));
  AND3_X1   g0963(.A1(new_n1110), .A2(KEYINPUT120), .A3(new_n1107), .ZN(new_n1164));
  AOI21_X1  g0964(.A(KEYINPUT120), .B1(new_n1110), .B2(new_n1107), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1163), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT121), .ZN(new_n1167));
  INV_X1    g0967(.A(KEYINPUT57), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1166), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1159), .A2(new_n1162), .A3(new_n1169), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1151), .A2(new_n753), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n799), .A2(G107), .ZN(new_n1172));
  OR2_X1    g0972(.A1(new_n1172), .A2(KEYINPUT118), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n758), .A2(new_n340), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n795), .A2(new_n375), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n1173), .A2(new_n930), .A3(new_n1174), .A4(new_n1175), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n1172), .A2(KEYINPUT118), .B1(G283), .B2(new_n792), .ZN(new_n1177));
  OAI221_X1 g0977(.A(new_n1177), .B1(new_n202), .B2(new_n784), .C1(new_n204), .C2(new_n775), .ZN(new_n1178));
  AOI211_X1 g0978(.A(new_n1176), .B(new_n1178), .C1(G116), .C2(new_n788), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1179), .B1(new_n257), .B2(new_n801), .ZN(new_n1180));
  XNOR2_X1  g0980(.A(new_n1180), .B(KEYINPUT58), .ZN(new_n1181));
  AOI211_X1 g0981(.A(G50), .B(new_n1174), .C1(new_n267), .C2(new_n286), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(G132), .A2(new_n781), .B1(new_n795), .B2(G137), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n775), .A2(new_n1122), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1184), .B1(new_n788), .B2(G125), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n1183), .B(new_n1185), .C1(new_n355), .C2(new_n770), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1186), .B1(G128), .B2(new_n799), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(new_n1187), .B(KEYINPUT59), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(new_n785), .A2(G159), .B1(new_n792), .B2(G124), .ZN(new_n1189));
  AND3_X1   g0989(.A1(new_n1189), .A2(new_n267), .A3(new_n286), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1182), .B1(new_n1188), .B2(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n947), .B1(new_n1181), .B2(new_n1191), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n1114), .A2(G50), .ZN(new_n1193));
  NOR4_X1   g0993(.A1(new_n1171), .A2(new_n812), .A3(new_n1192), .A4(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(new_n1163), .B2(new_n1002), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1170), .A2(new_n1195), .ZN(G375));
  OR2_X1    g0996(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1197), .A2(new_n996), .A3(new_n1108), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n335), .B1(new_n799), .B2(G283), .ZN(new_n1199));
  OAI211_X1 g0999(.A(new_n1199), .B(new_n1009), .C1(new_n801), .C2(new_n254), .ZN(new_n1200));
  OAI22_X1  g1000(.A1(new_n796), .A2(new_n513), .B1(new_n787), .B2(new_n771), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  OAI221_X1 g1002(.A(new_n1202), .B1(new_n204), .B2(new_n784), .C1(new_n257), .C2(new_n775), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n1200), .B(new_n1203), .C1(G303), .C2(new_n792), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n788), .A2(G132), .B1(G58), .B2(new_n785), .ZN(new_n1205));
  OAI221_X1 g1005(.A(new_n1205), .B1(new_n835), .B2(new_n775), .C1(new_n801), .C2(new_n1122), .ZN(new_n1206));
  AND2_X1   g1006(.A1(new_n792), .A2(G128), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n796), .A2(new_n355), .ZN(new_n1208));
  OAI221_X1 g1008(.A(new_n758), .B1(new_n770), .B2(new_n201), .C1(new_n798), .C2(new_n834), .ZN(new_n1209));
  NOR4_X1   g1009(.A1(new_n1206), .A2(new_n1207), .A3(new_n1208), .A4(new_n1209), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n756), .B1(new_n1204), .B2(new_n1210), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n813), .B(new_n1211), .C1(new_n880), .C2(new_n753), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1212), .B1(new_n203), .B2(new_n849), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(new_n1106), .B2(new_n1002), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1198), .A2(new_n1214), .ZN(G381));
  NOR2_X1   g1015(.A1(G375), .A2(G378), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1065), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1071), .A2(KEYINPUT116), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1074), .A2(new_n1073), .A3(new_n1075), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1217), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1220), .A2(new_n999), .A3(new_n1044), .ZN(new_n1221));
  OR3_X1    g1021(.A1(G393), .A2(G396), .A3(G381), .ZN(new_n1222));
  NOR3_X1   g1022(.A1(new_n1221), .A2(new_n1222), .A3(G384), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1216), .A2(new_n1223), .ZN(G407));
  OAI21_X1  g1024(.A(new_n1216), .B1(new_n1223), .B2(new_n674), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1225), .A2(G213), .ZN(G409));
  AND3_X1   g1026(.A1(new_n1166), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1167), .B1(new_n1166), .B2(new_n1168), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1160), .ZN(new_n1229));
  OAI211_X1 g1029(.A(KEYINPUT57), .B(new_n1229), .C1(new_n1164), .C2(new_n1165), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1230), .A2(new_n704), .ZN(new_n1231));
  NOR3_X1   g1031(.A1(new_n1227), .A2(new_n1228), .A3(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1195), .ZN(new_n1233));
  OAI21_X1  g1033(.A(G378), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(G213), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n1235), .A2(G343), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1158), .A2(new_n996), .ZN(new_n1238));
  INV_X1    g1038(.A(G378), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1194), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1229), .A2(new_n1002), .ZN(new_n1241));
  NAND4_X1  g1041(.A1(new_n1238), .A2(new_n1239), .A3(new_n1240), .A4(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT60), .ZN(new_n1243));
  OR3_X1    g1043(.A1(new_n1106), .A2(new_n1107), .A3(new_n1243), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1243), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1245));
  NAND4_X1  g1045(.A1(new_n1244), .A2(new_n704), .A3(new_n1108), .A4(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(new_n1214), .ZN(new_n1247));
  INV_X1    g1047(.A(G384), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1246), .A2(G384), .A3(new_n1214), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1251), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1234), .A2(new_n1237), .A3(new_n1242), .A4(new_n1252), .ZN(new_n1253));
  AND2_X1   g1053(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1234), .A2(new_n1237), .A3(new_n1242), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT122), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1251), .A2(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1249), .A2(KEYINPUT122), .A3(new_n1250), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1258), .A2(G2897), .A3(new_n1236), .A4(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1236), .A2(G2897), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1251), .A2(new_n1257), .A3(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1260), .A2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1256), .A2(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT61), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1236), .B1(G375), .B2(G378), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n1254), .A2(new_n1267), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1266), .A2(new_n1242), .A3(new_n1252), .A4(new_n1268), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1255), .A2(new_n1264), .A3(new_n1265), .A4(new_n1269), .ZN(new_n1270));
  XNOR2_X1  g1070(.A(G393), .B(G396), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1271), .ZN(new_n1272));
  OAI21_X1  g1072(.A(KEYINPUT124), .B1(G390), .B2(G387), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n999), .B1(new_n1220), .B2(new_n1044), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1272), .B1(new_n1273), .B2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT126), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(G390), .A2(G387), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1277), .A2(new_n1221), .A3(new_n1271), .A4(KEYINPUT124), .ZN(new_n1278));
  AND3_X1   g1078(.A1(new_n1275), .A2(new_n1276), .A3(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1276), .B1(new_n1275), .B2(new_n1278), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1270), .A2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1275), .A2(new_n1278), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1239), .B1(new_n1170), .B2(new_n1195), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1242), .ZN(new_n1285));
  NOR4_X1   g1085(.A1(new_n1284), .A2(new_n1236), .A3(new_n1285), .A4(new_n1251), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1283), .B1(new_n1286), .B2(KEYINPUT63), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT123), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1263), .A2(new_n1288), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1260), .A2(KEYINPUT123), .A3(new_n1262), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1289), .A2(new_n1256), .A3(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT63), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1253), .A2(new_n1292), .ZN(new_n1293));
  NAND4_X1  g1093(.A1(new_n1287), .A2(new_n1265), .A3(new_n1291), .A4(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1282), .A2(new_n1294), .ZN(G405));
  XNOR2_X1  g1095(.A(new_n1251), .B(KEYINPUT127), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1296), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1297), .B1(new_n1275), .B2(new_n1278), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1298), .ZN(new_n1299));
  NOR2_X1   g1099(.A1(new_n1216), .A2(new_n1284), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1275), .A2(new_n1278), .A3(new_n1297), .ZN(new_n1301));
  AND3_X1   g1101(.A1(new_n1299), .A2(new_n1300), .A3(new_n1301), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1300), .B1(new_n1299), .B2(new_n1301), .ZN(new_n1303));
  NOR2_X1   g1103(.A1(new_n1302), .A2(new_n1303), .ZN(G402));
endmodule


