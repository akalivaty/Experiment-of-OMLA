//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 0 0 0 0 1 1 0 1 1 0 0 0 0 1 1 1 0 0 0 1 1 1 0 1 1 0 0 1 0 0 0 1 0 0 1 0 0 0 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:17 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n698, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n714, new_n715, new_n716, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n734, new_n735, new_n736,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n922, new_n923, new_n924, new_n925, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017;
  INV_X1    g000(.A(G140), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G125), .ZN(new_n188));
  INV_X1    g002(.A(G125), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G140), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n188), .A2(new_n190), .A3(KEYINPUT16), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT16), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n192), .A2(new_n187), .A3(G125), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT76), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  NAND4_X1  g009(.A1(new_n192), .A2(new_n187), .A3(KEYINPUT76), .A4(G125), .ZN(new_n196));
  NAND4_X1  g010(.A1(new_n191), .A2(new_n195), .A3(G146), .A4(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(KEYINPUT77), .ZN(new_n198));
  AND2_X1   g012(.A1(new_n195), .A2(new_n196), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT77), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n199), .A2(new_n200), .A3(G146), .A4(new_n191), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n191), .A2(new_n195), .A3(new_n196), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT78), .ZN(new_n203));
  INV_X1    g017(.A(G146), .ZN(new_n204));
  AND3_X1   g018(.A1(new_n202), .A2(new_n203), .A3(new_n204), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n203), .B1(new_n202), .B2(new_n204), .ZN(new_n206));
  OAI211_X1 g020(.A(new_n198), .B(new_n201), .C1(new_n205), .C2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT92), .ZN(new_n208));
  INV_X1    g022(.A(G237), .ZN(new_n209));
  INV_X1    g023(.A(G953), .ZN(new_n210));
  NAND4_X1  g024(.A1(new_n209), .A2(new_n210), .A3(G143), .A4(G214), .ZN(new_n211));
  XNOR2_X1  g025(.A(KEYINPUT66), .B(G143), .ZN(new_n212));
  AND3_X1   g026(.A1(new_n209), .A2(new_n210), .A3(G214), .ZN(new_n213));
  OAI211_X1 g027(.A(new_n208), .B(new_n211), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n213), .A2(KEYINPUT92), .A3(G143), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT17), .ZN(new_n217));
  XNOR2_X1  g031(.A(KEYINPUT68), .B(G131), .ZN(new_n218));
  INV_X1    g032(.A(new_n218), .ZN(new_n219));
  NOR3_X1   g033(.A1(new_n216), .A2(new_n217), .A3(new_n219), .ZN(new_n220));
  OAI21_X1  g034(.A(KEYINPUT96), .B1(new_n207), .B2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT93), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n222), .B1(new_n216), .B2(new_n219), .ZN(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  AND2_X1   g038(.A1(new_n214), .A2(new_n215), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(new_n218), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n216), .A2(new_n222), .A3(new_n219), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n224), .A2(new_n217), .A3(new_n226), .A4(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(new_n206), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n202), .A2(new_n203), .A3(new_n204), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n225), .A2(KEYINPUT17), .A3(new_n218), .ZN(new_n232));
  XNOR2_X1  g046(.A(new_n197), .B(new_n200), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT96), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n231), .A2(new_n232), .A3(new_n233), .A4(new_n234), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n221), .A2(new_n228), .A3(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(KEYINPUT18), .A2(G131), .ZN(new_n237));
  XNOR2_X1  g051(.A(new_n216), .B(new_n237), .ZN(new_n238));
  AND2_X1   g052(.A1(new_n188), .A2(new_n190), .ZN(new_n239));
  XNOR2_X1  g053(.A(new_n239), .B(G146), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  XOR2_X1   g056(.A(G113), .B(G122), .Z(new_n243));
  XNOR2_X1  g057(.A(new_n243), .B(KEYINPUT95), .ZN(new_n244));
  INV_X1    g058(.A(G104), .ZN(new_n245));
  XNOR2_X1  g059(.A(new_n244), .B(new_n245), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n236), .A2(new_n242), .A3(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n246), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT19), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n239), .B1(KEYINPUT94), .B2(new_n249), .ZN(new_n250));
  XNOR2_X1  g064(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n250), .B1(new_n239), .B2(new_n251), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n197), .B1(new_n252), .B2(G146), .ZN(new_n253));
  AOI211_X1 g067(.A(KEYINPUT93), .B(new_n218), .C1(new_n214), .C2(new_n215), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n223), .A2(new_n254), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n253), .B1(new_n255), .B2(new_n226), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n248), .B1(new_n256), .B2(new_n241), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n247), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT20), .ZN(new_n259));
  NOR2_X1   g073(.A1(G475), .A2(G902), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n258), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n259), .B1(new_n258), .B2(new_n260), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT97), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n261), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NAND4_X1  g078(.A1(new_n258), .A2(KEYINPUT97), .A3(new_n259), .A4(new_n260), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(G475), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n236), .A2(new_n242), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(new_n248), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(new_n247), .ZN(new_n270));
  INV_X1    g084(.A(G902), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n267), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n266), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(KEYINPUT98), .ZN(new_n275));
  INV_X1    g089(.A(G128), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(G143), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n277), .B1(new_n212), .B2(new_n276), .ZN(new_n278));
  XNOR2_X1  g092(.A(new_n278), .B(G134), .ZN(new_n279));
  XOR2_X1   g093(.A(G116), .B(G122), .Z(new_n280));
  OAI21_X1  g094(.A(new_n279), .B1(G107), .B2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(G116), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n282), .A2(KEYINPUT14), .A3(G122), .ZN(new_n283));
  OAI211_X1 g097(.A(G107), .B(new_n283), .C1(new_n280), .C2(KEYINPUT14), .ZN(new_n284));
  XNOR2_X1  g098(.A(new_n284), .B(KEYINPUT99), .ZN(new_n285));
  INV_X1    g099(.A(G143), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(KEYINPUT66), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT66), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(G143), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT13), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n290), .A2(new_n291), .A3(G128), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n292), .B1(new_n278), .B2(new_n291), .ZN(new_n293));
  INV_X1    g107(.A(G134), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  XNOR2_X1  g109(.A(new_n280), .B(G107), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n296), .B1(G134), .B2(new_n278), .ZN(new_n297));
  OAI22_X1  g111(.A1(new_n281), .A2(new_n285), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  XOR2_X1   g112(.A(KEYINPUT9), .B(G234), .Z(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(G217), .ZN(new_n301));
  NOR3_X1   g115(.A1(new_n300), .A2(new_n301), .A3(G953), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  OR2_X1    g117(.A1(new_n298), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n298), .A2(new_n303), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(new_n271), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT15), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n307), .A2(new_n308), .A3(G478), .ZN(new_n309));
  INV_X1    g123(.A(G478), .ZN(new_n310));
  OAI211_X1 g124(.A(new_n306), .B(new_n271), .C1(KEYINPUT15), .C2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n210), .A2(G952), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n314), .B1(G234), .B2(G237), .ZN(new_n315));
  XOR2_X1   g129(.A(KEYINPUT21), .B(G898), .Z(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(G234), .A2(G237), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n318), .A2(G902), .A3(G953), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n315), .B1(new_n317), .B2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT98), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n266), .A2(new_n323), .A3(new_n273), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n275), .A2(new_n313), .A3(new_n322), .A4(new_n324), .ZN(new_n325));
  OAI21_X1  g139(.A(G214), .B1(G237), .B2(G902), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT87), .ZN(new_n328));
  OAI21_X1  g142(.A(KEYINPUT3), .B1(new_n245), .B2(G107), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT80), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n245), .A2(G107), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT3), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n245), .A2(G107), .ZN(new_n335));
  OAI211_X1 g149(.A(KEYINPUT80), .B(KEYINPUT3), .C1(new_n245), .C2(G107), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n331), .A2(new_n334), .A3(new_n335), .A4(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(G101), .ZN(new_n338));
  INV_X1    g152(.A(G107), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n339), .A2(G104), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n340), .B1(new_n333), .B2(new_n332), .ZN(new_n341));
  INV_X1    g155(.A(G101), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n341), .A2(new_n342), .A3(new_n331), .A4(new_n336), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n338), .A2(KEYINPUT4), .A3(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT4), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n337), .A2(new_n345), .A3(G101), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  XOR2_X1   g161(.A(KEYINPUT2), .B(G113), .Z(new_n348));
  NAND2_X1  g162(.A1(new_n282), .A2(G119), .ZN(new_n349));
  INV_X1    g163(.A(G119), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n350), .A2(KEYINPUT71), .A3(G116), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT71), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n352), .B1(new_n282), .B2(G119), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n348), .A2(new_n349), .A3(new_n351), .A4(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT72), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n353), .A2(new_n349), .A3(new_n351), .ZN(new_n356));
  XNOR2_X1  g170(.A(KEYINPUT2), .B(G113), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n354), .A2(new_n355), .A3(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n356), .A2(KEYINPUT72), .A3(new_n357), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n328), .B1(new_n347), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n339), .A2(G104), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n342), .B1(new_n363), .B2(new_n335), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(KEYINPUT81), .ZN(new_n365));
  OAI21_X1  g179(.A(G101), .B1(new_n332), .B2(new_n340), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT81), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n343), .A2(new_n365), .A3(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT82), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  XNOR2_X1  g185(.A(new_n364), .B(new_n367), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n372), .A2(KEYINPUT82), .A3(new_n343), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n353), .A2(new_n351), .A3(KEYINPUT5), .A4(new_n349), .ZN(new_n374));
  OR3_X1    g188(.A1(new_n282), .A2(KEYINPUT5), .A3(G119), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n374), .A2(G113), .A3(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT88), .ZN(new_n377));
  OR2_X1    g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n356), .A2(new_n357), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n379), .B1(new_n376), .B2(new_n377), .ZN(new_n380));
  NAND4_X1  g194(.A1(new_n371), .A2(new_n373), .A3(new_n378), .A4(new_n380), .ZN(new_n381));
  AND2_X1   g195(.A1(new_n359), .A2(new_n360), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n382), .A2(KEYINPUT87), .A3(new_n346), .A4(new_n344), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n362), .A2(new_n381), .A3(new_n383), .ZN(new_n384));
  XOR2_X1   g198(.A(G110), .B(G122), .Z(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT89), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(KEYINPUT6), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(new_n385), .ZN(new_n390));
  NAND4_X1  g204(.A1(new_n362), .A2(new_n383), .A3(new_n390), .A4(new_n381), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n384), .A2(new_n387), .A3(KEYINPUT6), .A4(new_n385), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n389), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n286), .A2(G146), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n394), .B1(new_n290), .B2(G146), .ZN(new_n395));
  OR2_X1    g209(.A1(KEYINPUT0), .A2(G128), .ZN(new_n396));
  NAND2_X1  g210(.A1(KEYINPUT0), .A2(G128), .ZN(new_n397));
  XNOR2_X1  g211(.A(new_n397), .B(KEYINPUT65), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n395), .A2(new_n396), .A3(new_n398), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n286), .A2(G146), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n400), .B1(new_n290), .B2(G146), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n401), .A2(KEYINPUT0), .A3(G128), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n189), .B1(new_n399), .B2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT70), .ZN(new_n405));
  INV_X1    g219(.A(new_n400), .ZN(new_n406));
  OAI211_X1 g220(.A(G128), .B(new_n406), .C1(new_n212), .C2(new_n204), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n405), .B1(new_n407), .B2(KEYINPUT1), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT1), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n401), .A2(KEYINPUT70), .A3(new_n409), .A4(G128), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  OAI21_X1  g225(.A(G128), .B1(new_n400), .B2(new_n409), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n395), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n404), .B1(new_n414), .B2(G125), .ZN(new_n415));
  INV_X1    g229(.A(G224), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n416), .A2(G953), .ZN(new_n417));
  XNOR2_X1  g231(.A(new_n415), .B(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n393), .A2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT91), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n371), .A2(new_n373), .A3(new_n354), .A4(new_n376), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n378), .A2(new_n380), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(new_n369), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  XOR2_X1   g238(.A(new_n385), .B(KEYINPUT8), .Z(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n391), .A2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT90), .ZN(new_n428));
  AOI22_X1  g242(.A1(new_n408), .A2(new_n410), .B1(new_n395), .B2(new_n412), .ZN(new_n429));
  AOI211_X1 g243(.A(new_n428), .B(new_n403), .C1(new_n429), .C2(new_n189), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n429), .A2(new_n428), .A3(new_n189), .ZN(new_n431));
  OAI21_X1  g245(.A(KEYINPUT7), .B1(new_n416), .B2(G953), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  OAI22_X1  g247(.A1(new_n430), .A2(new_n433), .B1(new_n415), .B2(new_n432), .ZN(new_n434));
  OAI211_X1 g248(.A(new_n420), .B(new_n271), .C1(new_n427), .C2(new_n434), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n271), .B1(new_n427), .B2(new_n434), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(KEYINPUT91), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n419), .A2(new_n435), .A3(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(G210), .B1(G237), .B2(G902), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  AOI22_X1  g255(.A1(new_n393), .A2(new_n418), .B1(new_n436), .B2(KEYINPUT91), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n442), .A2(new_n439), .A3(new_n435), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n327), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  OAI21_X1  g258(.A(G221), .B1(new_n300), .B2(G902), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n369), .A2(new_n370), .ZN(new_n447));
  AOI21_X1  g261(.A(KEYINPUT82), .B1(new_n372), .B2(new_n343), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n429), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  OAI21_X1  g263(.A(KEYINPUT1), .B1(new_n290), .B2(G146), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(G128), .ZN(new_n451));
  INV_X1    g265(.A(new_n401), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n411), .A2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n369), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n449), .A2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT84), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT11), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n459), .B1(new_n294), .B2(G137), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT67), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n294), .A2(G137), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(KEYINPUT11), .ZN(new_n464));
  INV_X1    g278(.A(G137), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n465), .A2(G134), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  OAI211_X1 g281(.A(KEYINPUT67), .B(new_n459), .C1(new_n294), .C2(G137), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n462), .A2(new_n464), .A3(new_n467), .A4(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT69), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n466), .B1(KEYINPUT11), .B2(new_n463), .ZN(new_n472));
  NAND4_X1  g286(.A1(new_n472), .A2(KEYINPUT69), .A3(new_n462), .A4(new_n468), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n471), .A2(G131), .A3(new_n473), .ZN(new_n474));
  OR2_X1    g288(.A1(new_n469), .A2(new_n218), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n457), .A2(new_n458), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(KEYINPUT12), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n469), .A2(new_n218), .ZN(new_n479));
  AND2_X1   g293(.A1(new_n473), .A2(G131), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n479), .B1(new_n480), .B2(new_n471), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT83), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n476), .A2(KEYINPUT83), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT10), .ZN(new_n486));
  AOI22_X1  g300(.A1(new_n408), .A2(new_n410), .B1(new_n452), .B2(new_n451), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n486), .B1(new_n487), .B2(new_n369), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n344), .A2(new_n402), .A3(new_n399), .A4(new_n346), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n414), .A2(KEYINPUT10), .A3(new_n371), .A4(new_n373), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n485), .A2(new_n488), .A3(new_n489), .A4(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT12), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n457), .A2(new_n458), .A3(new_n492), .A4(new_n476), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n478), .A2(new_n491), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(KEYINPUT85), .ZN(new_n495));
  XNOR2_X1  g309(.A(G110), .B(G140), .ZN(new_n496));
  AND2_X1   g310(.A1(new_n210), .A2(G227), .ZN(new_n497));
  XOR2_X1   g311(.A(new_n496), .B(new_n497), .Z(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT85), .ZN(new_n500));
  NAND4_X1  g314(.A1(new_n478), .A2(new_n500), .A3(new_n491), .A4(new_n493), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n495), .A2(new_n499), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n491), .A2(new_n498), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT86), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n490), .A2(new_n488), .A3(new_n489), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(new_n476), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n491), .A2(KEYINPUT86), .A3(new_n498), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n505), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n502), .A2(G469), .A3(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(G469), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n511), .A2(new_n271), .ZN(new_n512));
  NAND4_X1  g326(.A1(new_n478), .A2(new_n491), .A3(new_n498), .A4(new_n493), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n507), .A2(new_n491), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(new_n499), .ZN(new_n515));
  AOI21_X1  g329(.A(G902), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n512), .B1(new_n516), .B2(new_n511), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n446), .B1(new_n510), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n444), .A2(new_n518), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n325), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n210), .A2(G221), .A3(G234), .ZN(new_n521));
  XNOR2_X1  g335(.A(new_n521), .B(KEYINPUT79), .ZN(new_n522));
  XOR2_X1   g336(.A(new_n522), .B(KEYINPUT22), .Z(new_n523));
  XNOR2_X1  g337(.A(new_n523), .B(new_n465), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n276), .A2(G119), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n350), .A2(G128), .ZN(new_n527));
  AND2_X1   g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  XOR2_X1   g342(.A(KEYINPUT24), .B(G110), .Z(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT74), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n526), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(KEYINPUT23), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT23), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n526), .A2(new_n531), .A3(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n533), .A2(new_n527), .A3(new_n535), .ZN(new_n536));
  XOR2_X1   g350(.A(new_n536), .B(KEYINPUT75), .Z(new_n537));
  INV_X1    g351(.A(G110), .ZN(new_n538));
  OAI211_X1 g352(.A(new_n530), .B(new_n207), .C1(new_n537), .C2(new_n538), .ZN(new_n539));
  OAI22_X1  g353(.A1(new_n536), .A2(G110), .B1(new_n528), .B2(new_n529), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n239), .A2(new_n204), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n540), .A2(new_n197), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n539), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n525), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n524), .A2(new_n539), .A3(new_n542), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n544), .A2(new_n545), .A3(new_n271), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n301), .B1(G234), .B2(new_n271), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT25), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n546), .B(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n548), .B1(new_n550), .B2(new_n547), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  XNOR2_X1  g366(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n553), .B(G101), .ZN(new_n554));
  INV_X1    g368(.A(G210), .ZN(new_n555));
  NOR3_X1   g369(.A1(new_n555), .A2(G237), .A3(G953), .ZN(new_n556));
  XOR2_X1   g370(.A(new_n554), .B(new_n556), .Z(new_n557));
  OAI21_X1  g371(.A(G131), .B1(new_n463), .B2(new_n466), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n475), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n399), .A2(new_n402), .ZN(new_n560));
  OAI221_X1 g374(.A(new_n361), .B1(new_n429), .B2(new_n559), .C1(new_n481), .C2(new_n560), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n561), .B(KEYINPUT28), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n429), .A2(new_n559), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n560), .B1(new_n474), .B2(new_n475), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n382), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n557), .B1(new_n562), .B2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT64), .ZN(new_n567));
  OAI211_X1 g381(.A(new_n567), .B(KEYINPUT30), .C1(new_n563), .C2(new_n564), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  OAI22_X1  g383(.A1(new_n481), .A2(new_n560), .B1(new_n429), .B2(new_n559), .ZN(new_n570));
  AOI21_X1  g384(.A(KEYINPUT30), .B1(new_n570), .B2(new_n567), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n382), .B1(new_n569), .B2(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n572), .A2(new_n557), .A3(new_n561), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT31), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n561), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n567), .B1(new_n563), .B2(new_n564), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT30), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(new_n568), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n576), .B1(new_n580), .B2(new_n382), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n581), .A2(KEYINPUT31), .A3(new_n557), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n566), .B1(new_n575), .B2(new_n582), .ZN(new_n583));
  NOR2_X1   g397(.A1(G472), .A2(G902), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  OAI21_X1  g399(.A(KEYINPUT32), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n566), .ZN(new_n587));
  AOI21_X1  g401(.A(KEYINPUT31), .B1(new_n581), .B2(new_n557), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n361), .B1(new_n579), .B2(new_n568), .ZN(new_n589));
  INV_X1    g403(.A(new_n557), .ZN(new_n590));
  NOR4_X1   g404(.A1(new_n589), .A2(new_n574), .A3(new_n590), .A4(new_n576), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n587), .B1(new_n588), .B2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT32), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n592), .A2(new_n593), .A3(new_n584), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n586), .A2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(G472), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n561), .A2(new_n565), .A3(KEYINPUT73), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT73), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n570), .A2(new_n598), .A3(new_n382), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n597), .A2(KEYINPUT28), .A3(new_n599), .ZN(new_n600));
  OR2_X1    g414(.A1(new_n576), .A2(KEYINPUT28), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n600), .A2(KEYINPUT29), .A3(new_n557), .A4(new_n601), .ZN(new_n602));
  AND2_X1   g416(.A1(new_n602), .A2(new_n271), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT29), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n590), .B1(new_n562), .B2(new_n565), .ZN(new_n605));
  NOR3_X1   g419(.A1(new_n589), .A2(new_n557), .A3(new_n576), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n604), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n596), .B1(new_n603), .B2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n552), .B1(new_n595), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n520), .A2(new_n610), .ZN(new_n611));
  XOR2_X1   g425(.A(KEYINPUT100), .B(G101), .Z(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(G3));
  NAND2_X1  g427(.A1(new_n444), .A2(new_n322), .ZN(new_n614));
  OAI21_X1  g428(.A(G472), .B1(new_n583), .B2(G902), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n592), .A2(new_n584), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n510), .A2(new_n517), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(new_n445), .ZN(new_n619));
  NOR4_X1   g433(.A1(new_n614), .A2(new_n617), .A3(new_n619), .A4(new_n552), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n306), .A2(KEYINPUT33), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT33), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n304), .A2(new_n622), .A3(new_n305), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n621), .A2(new_n623), .A3(G478), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n306), .A2(new_n310), .A3(new_n271), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n310), .A2(new_n271), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n624), .A2(new_n625), .A3(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(KEYINPUT101), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n323), .B1(new_n266), .B2(new_n273), .ZN(new_n630));
  AOI211_X1 g444(.A(KEYINPUT98), .B(new_n272), .C1(new_n264), .C2(new_n265), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n629), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(KEYINPUT102), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT102), .ZN(new_n634));
  OAI211_X1 g448(.A(new_n634), .B(new_n629), .C1(new_n630), .C2(new_n631), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n620), .A2(new_n633), .A3(new_n635), .ZN(new_n636));
  XOR2_X1   g450(.A(KEYINPUT34), .B(G104), .Z(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G6));
  NAND2_X1  g452(.A1(new_n273), .A2(new_n312), .ZN(new_n639));
  INV_X1    g453(.A(new_n261), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n640), .A2(new_n262), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n620), .A2(new_n642), .ZN(new_n643));
  XOR2_X1   g457(.A(KEYINPUT35), .B(G107), .Z(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G9));
  NOR3_X1   g459(.A1(new_n630), .A2(new_n631), .A3(new_n321), .ZN(new_n646));
  AND2_X1   g460(.A1(new_n444), .A2(new_n518), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n543), .B(KEYINPUT103), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n525), .A2(KEYINPUT36), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n547), .A2(G902), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n550), .A2(new_n547), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  AND3_X1   g468(.A1(new_n615), .A2(new_n616), .A3(new_n654), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n646), .A2(new_n647), .A3(new_n655), .A4(new_n313), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(KEYINPUT37), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(new_n538), .ZN(G12));
  NAND3_X1  g472(.A1(new_n444), .A2(new_n518), .A3(new_n654), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n608), .B1(new_n586), .B2(new_n594), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(G900), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n315), .B1(new_n320), .B2(new_n662), .ZN(new_n663));
  NOR3_X1   g477(.A1(new_n639), .A2(new_n641), .A3(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(G128), .ZN(G30));
  OAI21_X1  g480(.A(new_n557), .B1(new_n589), .B2(new_n576), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n597), .A2(new_n599), .ZN(new_n668));
  AOI21_X1  g482(.A(G902), .B1(new_n668), .B2(new_n590), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n596), .B1(new_n667), .B2(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  NOR3_X1   g485(.A1(new_n583), .A2(KEYINPUT32), .A3(new_n585), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n593), .B1(new_n592), .B2(new_n584), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n671), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT105), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n670), .B1(new_n586), .B2(new_n594), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(KEYINPUT105), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n654), .B1(new_n676), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n275), .A2(new_n324), .ZN(new_n680));
  XOR2_X1   g494(.A(new_n663), .B(KEYINPUT39), .Z(new_n681));
  AND2_X1   g495(.A1(new_n518), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n679), .A2(new_n312), .A3(new_n680), .A4(new_n685), .ZN(new_n686));
  OR2_X1    g500(.A1(new_n682), .A2(new_n684), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n441), .A2(new_n443), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT104), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n688), .B(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(KEYINPUT38), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n688), .B(KEYINPUT104), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT38), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n687), .A2(new_n691), .A3(new_n694), .A4(new_n326), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n686), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(new_n290), .ZN(G45));
  INV_X1    g511(.A(new_n663), .ZN(new_n698));
  OAI211_X1 g512(.A(new_n629), .B(new_n698), .C1(new_n630), .C2(new_n631), .ZN(new_n699));
  INV_X1    g513(.A(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n661), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G146), .ZN(G48));
  NOR3_X1   g516(.A1(new_n660), .A2(new_n552), .A3(new_n321), .ZN(new_n703));
  AND2_X1   g517(.A1(new_n513), .A2(new_n515), .ZN(new_n704));
  OAI21_X1  g518(.A(G469), .B1(new_n704), .B2(G902), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n516), .A2(new_n511), .ZN(new_n706));
  AND3_X1   g520(.A1(new_n705), .A2(new_n445), .A3(new_n706), .ZN(new_n707));
  AND2_X1   g521(.A1(new_n707), .A2(new_n444), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n703), .A2(new_n633), .A3(new_n635), .A4(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(KEYINPUT41), .B(G113), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n709), .B(new_n710), .ZN(G15));
  NAND4_X1  g525(.A1(new_n610), .A2(new_n322), .A3(new_n642), .A4(new_n708), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G116), .ZN(G18));
  AND3_X1   g527(.A1(new_n707), .A2(new_n444), .A3(new_n654), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n609), .B1(new_n672), .B2(new_n673), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n714), .A2(new_n646), .A3(new_n715), .A4(new_n313), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G119), .ZN(G21));
  OAI211_X1 g531(.A(new_n707), .B(new_n312), .C1(new_n630), .C2(new_n631), .ZN(new_n718));
  INV_X1    g532(.A(new_n718), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n557), .B1(new_n600), .B2(new_n601), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n720), .B1(new_n575), .B2(new_n582), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT108), .ZN(new_n722));
  XOR2_X1   g536(.A(new_n584), .B(KEYINPUT107), .Z(new_n723));
  NOR3_X1   g537(.A1(new_n721), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(new_n720), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n725), .B1(new_n588), .B2(new_n591), .ZN(new_n726));
  INV_X1    g540(.A(new_n723), .ZN(new_n727));
  AOI21_X1  g541(.A(KEYINPUT108), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  OAI211_X1 g542(.A(new_n551), .B(new_n615), .C1(new_n724), .C2(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(new_n729), .ZN(new_n730));
  INV_X1    g544(.A(new_n614), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n719), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G122), .ZN(G24));
  OAI211_X1 g547(.A(new_n615), .B(new_n654), .C1(new_n724), .C2(new_n728), .ZN(new_n734));
  INV_X1    g548(.A(new_n734), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n700), .A2(new_n735), .A3(new_n708), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G125), .ZN(G27));
  INV_X1    g551(.A(KEYINPUT42), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n446), .A2(new_n327), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n441), .A2(new_n443), .A3(new_n739), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n498), .B1(new_n494), .B2(KEYINPUT85), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n741), .A2(KEYINPUT109), .A3(new_n501), .ZN(new_n742));
  INV_X1    g556(.A(new_n742), .ZN(new_n743));
  AOI21_X1  g557(.A(KEYINPUT109), .B1(new_n741), .B2(new_n501), .ZN(new_n744));
  OAI211_X1 g558(.A(G469), .B(new_n509), .C1(new_n743), .C2(new_n744), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n740), .B1(new_n745), .B2(new_n517), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n746), .A2(new_n715), .A3(new_n551), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n738), .B1(new_n747), .B2(new_n699), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n700), .A2(KEYINPUT42), .A3(new_n610), .A4(new_n746), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G131), .ZN(G33));
  NAND3_X1  g565(.A1(new_n610), .A2(new_n664), .A3(new_n746), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(KEYINPUT110), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT110), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n610), .A2(new_n754), .A3(new_n664), .A4(new_n746), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G134), .ZN(G36));
  INV_X1    g571(.A(new_n509), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT109), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n502), .A2(new_n759), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n758), .B1(new_n760), .B2(new_n742), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(KEYINPUT45), .ZN(new_n762));
  AOI21_X1  g576(.A(KEYINPUT45), .B1(new_n502), .B2(new_n509), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n763), .A2(new_n511), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n512), .B1(new_n762), .B2(new_n764), .ZN(new_n765));
  AND2_X1   g579(.A1(new_n765), .A2(KEYINPUT46), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n706), .B1(new_n765), .B2(KEYINPUT46), .ZN(new_n767));
  OAI211_X1 g581(.A(new_n445), .B(new_n681), .C1(new_n766), .C2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(new_n617), .ZN(new_n769));
  INV_X1    g583(.A(new_n654), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT43), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT111), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n771), .B1(new_n680), .B2(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(new_n629), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n680), .A2(new_n774), .ZN(new_n775));
  OR2_X1    g589(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n773), .A2(new_n775), .ZN(new_n777));
  AOI211_X1 g591(.A(new_n769), .B(new_n770), .C1(new_n776), .C2(new_n777), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n768), .B1(new_n778), .B2(KEYINPUT44), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n441), .A2(new_n326), .A3(new_n443), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n776), .A2(new_n777), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n781), .A2(new_n617), .A3(new_n654), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT44), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n780), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n779), .A2(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(G137), .ZN(G39));
  OAI21_X1  g600(.A(new_n445), .B1(new_n766), .B2(new_n767), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT47), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  OAI211_X1 g603(.A(KEYINPUT47), .B(new_n445), .C1(new_n766), .C2(new_n767), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(new_n780), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n700), .A2(new_n660), .A3(new_n552), .A4(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(KEYINPUT112), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n791), .A2(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(G140), .ZN(G42));
  NAND2_X1  g610(.A1(new_n705), .A2(new_n706), .ZN(new_n797));
  INV_X1    g611(.A(new_n315), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n740), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n781), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n800), .A2(new_n610), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT48), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n801), .B(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n730), .A2(new_n315), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n804), .B1(new_n776), .B2(new_n777), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n805), .A2(new_n708), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n803), .A2(new_n314), .A3(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT54), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT53), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n748), .A2(new_n749), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n709), .A2(new_n712), .A3(new_n716), .A4(new_n732), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n661), .B1(new_n700), .B2(new_n664), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n813), .A2(new_n736), .ZN(new_n814));
  OAI211_X1 g628(.A(new_n312), .B(new_n444), .C1(new_n630), .C2(new_n631), .ZN(new_n815));
  INV_X1    g629(.A(new_n517), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n816), .B1(new_n761), .B2(G469), .ZN(new_n817));
  NOR4_X1   g631(.A1(new_n815), .A2(new_n817), .A3(new_n446), .A4(new_n663), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(new_n679), .ZN(new_n819));
  AOI21_X1  g633(.A(KEYINPUT52), .B1(new_n814), .B2(new_n819), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n677), .A2(KEYINPUT105), .ZN(new_n821));
  AOI211_X1 g635(.A(new_n675), .B(new_n670), .C1(new_n586), .C2(new_n594), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n770), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  AND4_X1   g637(.A1(new_n439), .A2(new_n419), .A3(new_n435), .A4(new_n437), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n439), .B1(new_n442), .B2(new_n435), .ZN(new_n825));
  OAI211_X1 g639(.A(new_n312), .B(new_n326), .C1(new_n824), .C2(new_n825), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n826), .B1(new_n324), .B2(new_n275), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n745), .A2(new_n517), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n827), .A2(new_n445), .A3(new_n698), .A4(new_n828), .ZN(new_n829));
  OAI211_X1 g643(.A(new_n813), .B(new_n736), .C1(new_n823), .C2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT52), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n812), .B1(new_n820), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n632), .A2(KEYINPUT113), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT113), .ZN(new_n835));
  OAI211_X1 g649(.A(new_n835), .B(new_n629), .C1(new_n630), .C2(new_n631), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n837), .A2(new_n620), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n838), .A2(new_n611), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n617), .A2(new_n619), .ZN(new_n840));
  INV_X1    g654(.A(new_n826), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n840), .A2(new_n646), .A3(new_n841), .A4(new_n551), .ZN(new_n842));
  AOI21_X1  g656(.A(KEYINPUT114), .B1(new_n842), .B2(new_n656), .ZN(new_n843));
  INV_X1    g657(.A(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n842), .A2(new_n656), .A3(KEYINPUT114), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n839), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NOR4_X1   g660(.A1(new_n770), .A2(new_n780), .A3(new_n312), .A4(new_n272), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n619), .A2(new_n641), .A3(new_n663), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n847), .A2(new_n715), .A3(new_n848), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n700), .A2(new_n735), .A3(new_n746), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n756), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n846), .A2(new_n851), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n809), .B1(new_n833), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n830), .A2(new_n831), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n819), .A2(KEYINPUT52), .A3(new_n736), .A4(new_n813), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n809), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  AOI22_X1  g670(.A1(new_n837), .A2(new_n620), .B1(new_n520), .B2(new_n610), .ZN(new_n857));
  AND3_X1   g671(.A1(new_n842), .A2(new_n656), .A3(KEYINPUT114), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n857), .B1(new_n858), .B2(new_n843), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n756), .A2(new_n849), .A3(new_n850), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n856), .A2(new_n861), .A3(new_n812), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n808), .B1(new_n853), .B2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(new_n863), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n821), .A2(new_n822), .A3(new_n552), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n865), .A2(new_n633), .A3(new_n635), .A4(new_n799), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n732), .A2(new_n712), .A3(new_n716), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n867), .A2(new_n750), .A3(new_n709), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT115), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n867), .A2(new_n750), .A3(KEYINPUT115), .A4(new_n709), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n856), .A2(new_n861), .A3(new_n870), .A4(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n853), .A2(new_n808), .A3(new_n872), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n807), .A2(new_n864), .A3(new_n866), .A4(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n800), .A2(new_n735), .ZN(new_n875));
  INV_X1    g689(.A(new_n680), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n865), .A2(new_n876), .A3(new_n774), .A4(new_n799), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n691), .A2(new_n694), .ZN(new_n878));
  AND3_X1   g692(.A1(new_n878), .A2(new_n327), .A3(new_n707), .ZN(new_n879));
  AOI21_X1  g693(.A(KEYINPUT116), .B1(new_n805), .B2(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT50), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  AOI211_X1 g696(.A(KEYINPUT116), .B(KEYINPUT50), .C1(new_n805), .C2(new_n879), .ZN(new_n883));
  OAI211_X1 g697(.A(new_n875), .B(new_n877), .C1(new_n882), .C2(new_n883), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n797), .A2(new_n445), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n805), .B1(new_n791), .B2(new_n885), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n886), .A2(new_n780), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT51), .ZN(new_n888));
  OR3_X1    g702(.A1(new_n884), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n888), .B1(new_n884), .B2(new_n887), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  OAI22_X1  g705(.A1(new_n874), .A2(new_n891), .B1(G952), .B2(G953), .ZN(new_n892));
  INV_X1    g706(.A(new_n739), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n775), .B1(KEYINPUT49), .B2(new_n797), .ZN(new_n894));
  AOI211_X1 g708(.A(new_n893), .B(new_n894), .C1(KEYINPUT49), .C2(new_n797), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n895), .A2(new_n878), .A3(new_n865), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n892), .A2(new_n896), .ZN(G75));
  NOR2_X1   g711(.A1(new_n210), .A2(G952), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n898), .B(KEYINPUT117), .ZN(new_n899));
  AND2_X1   g713(.A1(new_n856), .A2(new_n861), .ZN(new_n900));
  AND2_X1   g714(.A1(new_n870), .A2(new_n871), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n854), .A2(new_n855), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n861), .A2(new_n902), .A3(new_n812), .ZN(new_n903));
  AOI22_X1  g717(.A1(new_n900), .A2(new_n901), .B1(new_n903), .B2(new_n809), .ZN(new_n904));
  NOR3_X1   g718(.A1(new_n904), .A2(new_n555), .A3(new_n271), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n393), .B(new_n418), .Z(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(KEYINPUT55), .ZN(new_n907));
  OR3_X1    g721(.A1(new_n905), .A2(KEYINPUT56), .A3(new_n907), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n907), .B1(new_n905), .B2(KEYINPUT56), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n899), .B1(new_n908), .B2(new_n909), .ZN(G51));
  INV_X1    g724(.A(new_n704), .ZN(new_n911));
  INV_X1    g725(.A(new_n512), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(KEYINPUT57), .ZN(new_n913));
  AND3_X1   g727(.A1(new_n853), .A2(new_n808), .A3(new_n872), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n808), .B1(new_n853), .B2(new_n872), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n913), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n912), .A2(KEYINPUT57), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n911), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n853), .A2(new_n872), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n919), .A2(G902), .A3(new_n762), .A4(new_n764), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n898), .B1(new_n918), .B2(new_n920), .ZN(G54));
  NAND4_X1  g735(.A1(new_n919), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n922));
  INV_X1    g736(.A(new_n258), .ZN(new_n923));
  AND2_X1   g737(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n922), .A2(new_n923), .ZN(new_n925));
  NOR3_X1   g739(.A1(new_n924), .A2(new_n925), .A3(new_n898), .ZN(G60));
  INV_X1    g740(.A(KEYINPUT119), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n621), .A2(new_n623), .ZN(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  XNOR2_X1  g743(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n627), .B(new_n930), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(new_n932), .ZN(new_n933));
  AND4_X1   g747(.A1(new_n861), .A2(new_n856), .A3(new_n870), .A4(new_n871), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n868), .B1(new_n854), .B2(new_n855), .ZN(new_n935));
  AOI21_X1  g749(.A(KEYINPUT53), .B1(new_n935), .B2(new_n861), .ZN(new_n936));
  OAI21_X1  g750(.A(KEYINPUT54), .B1(new_n934), .B2(new_n936), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n933), .B1(new_n937), .B2(new_n873), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n927), .B1(new_n938), .B2(new_n899), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n932), .B1(new_n914), .B2(new_n915), .ZN(new_n940));
  INV_X1    g754(.A(new_n899), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n940), .A2(KEYINPUT119), .A3(new_n941), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n914), .A2(new_n863), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n929), .B1(new_n943), .B2(new_n931), .ZN(new_n944));
  AND3_X1   g758(.A1(new_n939), .A2(new_n942), .A3(new_n944), .ZN(G63));
  NAND2_X1  g759(.A1(G217), .A2(G902), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n946), .B(KEYINPUT60), .ZN(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  OAI211_X1 g762(.A(new_n650), .B(new_n948), .C1(new_n934), .C2(new_n936), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(KEYINPUT120), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n947), .B1(new_n853), .B2(new_n872), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT120), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n951), .A2(new_n952), .A3(new_n650), .ZN(new_n953));
  AND2_X1   g767(.A1(new_n544), .A2(new_n545), .ZN(new_n954));
  INV_X1    g768(.A(new_n954), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n955), .B1(new_n904), .B2(new_n947), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n950), .A2(new_n953), .A3(new_n956), .A4(new_n941), .ZN(new_n957));
  INV_X1    g771(.A(KEYINPUT61), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n954), .B1(new_n919), .B2(new_n948), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n958), .B1(new_n960), .B2(KEYINPUT121), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT121), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n962), .B1(new_n951), .B2(new_n954), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n961), .A2(new_n941), .A3(new_n949), .A4(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n959), .A2(new_n964), .ZN(G66));
  OAI21_X1  g779(.A(G953), .B1(new_n317), .B2(new_n416), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n859), .A2(new_n811), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n966), .B1(new_n967), .B2(G953), .ZN(new_n968));
  INV_X1    g782(.A(new_n393), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n969), .B1(G898), .B2(new_n210), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n970), .B(KEYINPUT122), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n968), .B(new_n971), .ZN(G69));
  NAND3_X1  g786(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n580), .B(KEYINPUT123), .Z(new_n974));
  XNOR2_X1  g788(.A(new_n974), .B(new_n252), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n837), .B1(new_n312), .B2(new_n876), .ZN(new_n976));
  INV_X1    g790(.A(new_n610), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n682), .A2(new_n792), .ZN(new_n978));
  NOR3_X1   g792(.A1(new_n976), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n979), .B1(new_n791), .B2(new_n794), .ZN(new_n980));
  AND2_X1   g794(.A1(new_n785), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n814), .B1(new_n686), .B2(new_n695), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n982), .A2(KEYINPUT62), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT124), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n983), .B(new_n984), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n982), .A2(KEYINPUT62), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n986), .B(KEYINPUT125), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n981), .A2(new_n985), .A3(new_n987), .ZN(new_n988));
  OAI211_X1 g802(.A(new_n973), .B(new_n975), .C1(new_n988), .C2(G953), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n814), .A2(new_n750), .ZN(new_n990));
  INV_X1    g804(.A(new_n990), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n792), .B1(new_n778), .B2(KEYINPUT44), .ZN(new_n992));
  NAND4_X1  g806(.A1(new_n781), .A2(KEYINPUT44), .A3(new_n617), .A4(new_n654), .ZN(new_n993));
  INV_X1    g807(.A(new_n768), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  OAI211_X1 g809(.A(new_n795), .B(new_n991), .C1(new_n992), .C2(new_n995), .ZN(new_n996));
  NOR2_X1   g810(.A1(new_n977), .A2(new_n815), .ZN(new_n997));
  AOI22_X1  g811(.A1(new_n994), .A2(new_n997), .B1(new_n755), .B2(new_n753), .ZN(new_n998));
  INV_X1    g812(.A(new_n998), .ZN(new_n999));
  OAI21_X1  g813(.A(KEYINPUT126), .B1(new_n996), .B2(new_n999), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n990), .B1(new_n779), .B2(new_n784), .ZN(new_n1001));
  INV_X1    g815(.A(KEYINPUT126), .ZN(new_n1002));
  NAND4_X1  g816(.A1(new_n1001), .A2(new_n1002), .A3(new_n795), .A4(new_n998), .ZN(new_n1003));
  AOI21_X1  g817(.A(G953), .B1(new_n1000), .B2(new_n1003), .ZN(new_n1004));
  OR2_X1    g818(.A1(new_n1004), .A2(new_n975), .ZN(new_n1005));
  NOR3_X1   g819(.A1(new_n662), .A2(new_n210), .A3(G227), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n989), .B1(new_n1005), .B2(new_n1006), .ZN(G72));
  INV_X1    g821(.A(new_n606), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n1000), .A2(new_n1003), .A3(new_n967), .ZN(new_n1009));
  XNOR2_X1  g823(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n1010));
  NAND2_X1  g824(.A1(G472), .A2(G902), .ZN(new_n1011));
  XNOR2_X1  g825(.A(new_n1010), .B(new_n1011), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n1008), .B1(new_n1009), .B2(new_n1012), .ZN(new_n1013));
  NAND4_X1  g827(.A1(new_n981), .A2(new_n985), .A3(new_n967), .A4(new_n987), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n667), .B1(new_n1014), .B2(new_n1012), .ZN(new_n1015));
  NAND3_X1  g829(.A1(new_n1008), .A2(new_n667), .A3(new_n1012), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n1016), .B1(new_n853), .B2(new_n862), .ZN(new_n1017));
  NOR4_X1   g831(.A1(new_n1013), .A2(new_n1015), .A3(new_n898), .A4(new_n1017), .ZN(G57));
endmodule


