//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 1 1 0 0 1 1 0 1 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 1 1 0 0 1 0 1 1 0 1 1 1 1 0 0 0 0 0 0 1 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:30 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n774, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n862,
    new_n863, new_n865, new_n866, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n922, new_n923, new_n924,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n957, new_n958, new_n959, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n984, new_n985, new_n986, new_n987,
    new_n989, new_n990;
  XNOR2_X1  g000(.A(G57gat), .B(G64gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT90), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT9), .ZN(new_n205));
  INV_X1    g004(.A(G71gat), .ZN(new_n206));
  INV_X1    g005(.A(G78gat), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n205), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(G71gat), .B(G78gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n204), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT88), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  OR2_X1    g011(.A1(new_n209), .A2(new_n211), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT89), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n202), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(new_n208), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n202), .A2(new_n214), .ZN(new_n217));
  OAI211_X1 g016(.A(new_n212), .B(new_n213), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  AND2_X1   g017(.A1(new_n210), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(G85gat), .A2(G92gat), .ZN(new_n220));
  XNOR2_X1  g019(.A(new_n220), .B(KEYINPUT7), .ZN(new_n221));
  NAND2_X1  g020(.A1(G99gat), .A2(G106gat), .ZN(new_n222));
  INV_X1    g021(.A(G85gat), .ZN(new_n223));
  INV_X1    g022(.A(G92gat), .ZN(new_n224));
  AOI22_X1  g023(.A1(KEYINPUT8), .A2(new_n222), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n221), .A2(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(G99gat), .B(G106gat), .ZN(new_n227));
  XNOR2_X1  g026(.A(new_n226), .B(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n219), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(new_n228), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n210), .A2(new_n218), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT10), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n229), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(new_n229), .ZN(new_n235));
  AOI22_X1  g034(.A1(new_n234), .A2(KEYINPUT94), .B1(new_n235), .B2(KEYINPUT10), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT94), .ZN(new_n237));
  NAND4_X1  g036(.A1(new_n229), .A2(new_n232), .A3(new_n237), .A4(new_n233), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(G230gat), .A2(G233gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n240), .B1(new_n229), .B2(new_n232), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n242), .B(KEYINPUT95), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  XNOR2_X1  g043(.A(G120gat), .B(G148gat), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n245), .B(G176gat), .ZN(new_n246));
  INV_X1    g045(.A(G204gat), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n246), .B(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n244), .A2(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n241), .A2(new_n248), .A3(new_n243), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(G229gat), .A2(G233gat), .ZN(new_n254));
  XOR2_X1   g053(.A(new_n254), .B(KEYINPUT87), .Z(new_n255));
  XNOR2_X1  g054(.A(G15gat), .B(G22gat), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT16), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n256), .B1(new_n257), .B2(G1gat), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n258), .B1(G1gat), .B2(new_n256), .ZN(new_n259));
  XOR2_X1   g058(.A(new_n259), .B(G8gat), .Z(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  XNOR2_X1  g060(.A(G43gat), .B(G50gat), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n262), .A2(KEYINPUT15), .ZN(new_n263));
  INV_X1    g062(.A(G29gat), .ZN(new_n264));
  INV_X1    g063(.A(G36gat), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n264), .A2(new_n265), .A3(KEYINPUT14), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT14), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n267), .B1(G29gat), .B2(G36gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(G29gat), .A2(G36gat), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n266), .A2(new_n268), .A3(KEYINPUT85), .A4(new_n269), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n263), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n262), .A2(KEYINPUT15), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n270), .A2(KEYINPUT15), .A3(new_n262), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n261), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT17), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n278), .B(KEYINPUT86), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n273), .A2(KEYINPUT17), .A3(new_n274), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n260), .A2(new_n280), .ZN(new_n281));
  OAI211_X1 g080(.A(new_n255), .B(new_n276), .C1(new_n279), .C2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT18), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT86), .ZN(new_n285));
  XNOR2_X1  g084(.A(new_n278), .B(new_n285), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n286), .A2(new_n260), .A3(new_n280), .ZN(new_n287));
  NAND4_X1  g086(.A1(new_n287), .A2(KEYINPUT18), .A3(new_n255), .A4(new_n276), .ZN(new_n288));
  XOR2_X1   g087(.A(new_n260), .B(new_n275), .Z(new_n289));
  XOR2_X1   g088(.A(new_n255), .B(KEYINPUT13), .Z(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n284), .A2(new_n288), .A3(new_n291), .ZN(new_n292));
  XNOR2_X1  g091(.A(G113gat), .B(G141gat), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n293), .B(KEYINPUT11), .ZN(new_n294));
  INV_X1    g093(.A(G169gat), .ZN(new_n295));
  XNOR2_X1  g094(.A(new_n294), .B(new_n295), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n296), .B(G197gat), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n297), .B(KEYINPUT12), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n292), .A2(new_n299), .ZN(new_n300));
  NAND4_X1  g099(.A1(new_n284), .A2(new_n288), .A3(new_n298), .A4(new_n291), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n253), .A2(new_n302), .ZN(new_n303));
  XNOR2_X1  g102(.A(KEYINPUT92), .B(G183gat), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n219), .A2(KEYINPUT21), .ZN(new_n306));
  XNOR2_X1  g105(.A(G127gat), .B(G155gat), .ZN(new_n307));
  XNOR2_X1  g106(.A(new_n306), .B(new_n307), .ZN(new_n308));
  XNOR2_X1  g107(.A(new_n308), .B(G211gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(G231gat), .A2(G233gat), .ZN(new_n310));
  XNOR2_X1  g109(.A(new_n310), .B(KEYINPUT91), .ZN(new_n311));
  XNOR2_X1  g110(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n312));
  XOR2_X1   g111(.A(new_n311), .B(new_n312), .Z(new_n313));
  NAND2_X1  g112(.A1(new_n309), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(G211gat), .ZN(new_n315));
  XNOR2_X1  g114(.A(new_n308), .B(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(new_n313), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n261), .B1(new_n219), .B2(KEYINPUT21), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  AND3_X1   g119(.A1(new_n314), .A2(new_n318), .A3(new_n320), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n320), .B1(new_n314), .B2(new_n318), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n305), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n314), .A2(new_n318), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(new_n319), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n314), .A2(new_n318), .A3(new_n320), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n325), .A2(new_n304), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n323), .A2(new_n327), .ZN(new_n328));
  XOR2_X1   g127(.A(G190gat), .B(G218gat), .Z(new_n329));
  INV_X1    g128(.A(KEYINPUT93), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT41), .ZN(new_n331));
  NAND2_X1  g130(.A1(G232gat), .A2(G233gat), .ZN(new_n332));
  OAI22_X1  g131(.A1(new_n329), .A2(new_n330), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n333), .B1(new_n228), .B2(new_n275), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n230), .A2(new_n280), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n334), .B1(new_n279), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n329), .A2(new_n330), .ZN(new_n337));
  XNOR2_X1  g136(.A(new_n336), .B(new_n337), .ZN(new_n338));
  XOR2_X1   g137(.A(G134gat), .B(G162gat), .Z(new_n339));
  NAND2_X1  g138(.A1(new_n332), .A2(new_n331), .ZN(new_n340));
  XNOR2_X1  g139(.A(new_n339), .B(new_n340), .ZN(new_n341));
  XOR2_X1   g140(.A(new_n338), .B(new_n341), .Z(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n328), .A2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT35), .ZN(new_n345));
  NAND2_X1  g144(.A1(G228gat), .A2(G233gat), .ZN(new_n346));
  INV_X1    g145(.A(G197gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(new_n247), .ZN(new_n348));
  NAND2_X1  g147(.A1(G197gat), .A2(G204gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(G211gat), .A2(G218gat), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT22), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n350), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT72), .ZN(new_n355));
  INV_X1    g154(.A(G218gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n315), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(new_n351), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n354), .A2(new_n355), .A3(new_n359), .ZN(new_n360));
  AOI22_X1  g159(.A1(new_n348), .A2(new_n349), .B1(new_n352), .B2(new_n351), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n357), .A2(new_n355), .A3(new_n351), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n360), .A2(new_n363), .ZN(new_n364));
  XNOR2_X1  g163(.A(G141gat), .B(G148gat), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(KEYINPUT74), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT74), .ZN(new_n367));
  INV_X1    g166(.A(G141gat), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n368), .A2(G148gat), .ZN(new_n369));
  INV_X1    g168(.A(G148gat), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n370), .A2(G141gat), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n367), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(G155gat), .A2(G162gat), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(KEYINPUT2), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n366), .A2(new_n372), .A3(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(G155gat), .ZN(new_n376));
  INV_X1    g175(.A(G162gat), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  AND2_X1   g177(.A1(new_n378), .A2(new_n373), .ZN(new_n379));
  INV_X1    g178(.A(new_n369), .ZN(new_n380));
  XNOR2_X1  g179(.A(KEYINPUT75), .B(G141gat), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n380), .B1(new_n381), .B2(new_n370), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n373), .B1(new_n378), .B2(KEYINPUT2), .ZN(new_n383));
  AOI22_X1  g182(.A1(new_n375), .A2(new_n379), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  XOR2_X1   g183(.A(KEYINPUT77), .B(KEYINPUT3), .Z(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT29), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n364), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT80), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n354), .A2(new_n389), .A3(new_n358), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n354), .A2(new_n389), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n359), .B1(new_n361), .B2(KEYINPUT80), .ZN(new_n392));
  OAI211_X1 g191(.A(new_n387), .B(new_n390), .C1(new_n391), .C2(new_n392), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n384), .B1(new_n393), .B2(new_n385), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n346), .B1(new_n388), .B2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(G22gat), .ZN(new_n396));
  INV_X1    g195(.A(new_n364), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n374), .B1(new_n365), .B2(KEYINPUT74), .ZN(new_n398));
  NOR3_X1   g197(.A1(new_n369), .A2(new_n371), .A3(new_n367), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n379), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n382), .A2(new_n383), .ZN(new_n401));
  AND3_X1   g200(.A1(new_n400), .A2(new_n401), .A3(new_n385), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n397), .B1(new_n402), .B2(KEYINPUT29), .ZN(new_n403));
  INV_X1    g202(.A(new_n346), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n400), .A2(new_n401), .ZN(new_n405));
  AOI21_X1  g204(.A(KEYINPUT29), .B1(new_n360), .B2(new_n363), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n405), .B1(new_n406), .B2(KEYINPUT3), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n403), .A2(new_n404), .A3(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n395), .A2(new_n396), .A3(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT81), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  XNOR2_X1  g210(.A(G78gat), .B(G106gat), .ZN(new_n412));
  INV_X1    g211(.A(G50gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n412), .B(new_n413), .ZN(new_n414));
  XOR2_X1   g213(.A(KEYINPUT79), .B(KEYINPUT31), .Z(new_n415));
  XNOR2_X1  g214(.A(new_n414), .B(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n394), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n404), .B1(new_n417), .B2(new_n403), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n407), .A2(new_n404), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n388), .A2(new_n419), .ZN(new_n420));
  OAI21_X1  g219(.A(G22gat), .B1(new_n418), .B2(new_n420), .ZN(new_n421));
  AOI22_X1  g220(.A1(new_n411), .A2(new_n416), .B1(new_n421), .B2(new_n409), .ZN(new_n422));
  AND4_X1   g221(.A1(KEYINPUT81), .A2(new_n421), .A3(new_n409), .A4(new_n416), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT70), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT1), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n426), .B1(G113gat), .B2(G120gat), .ZN(new_n427));
  AND2_X1   g226(.A1(G113gat), .A2(G120gat), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n425), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  XNOR2_X1  g228(.A(G127gat), .B(G134gat), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(G113gat), .ZN(new_n433));
  INV_X1    g232(.A(G120gat), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(G113gat), .A2(G120gat), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n435), .A2(KEYINPUT70), .A3(new_n426), .A4(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n430), .B1(new_n429), .B2(new_n437), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n432), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT28), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT68), .ZN(new_n441));
  INV_X1    g240(.A(G183gat), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(KEYINPUT27), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT27), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(G183gat), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n441), .B1(new_n443), .B2(new_n445), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n441), .B1(new_n444), .B2(G183gat), .ZN(new_n447));
  INV_X1    g246(.A(G190gat), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n440), .B1(new_n446), .B2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT69), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n444), .A2(G183gat), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n442), .A2(KEYINPUT27), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n454), .A2(KEYINPUT28), .A3(new_n448), .ZN(new_n455));
  AND3_X1   g254(.A1(new_n450), .A2(new_n451), .A3(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n451), .B1(new_n450), .B2(new_n455), .ZN(new_n457));
  NAND2_X1  g256(.A1(G183gat), .A2(G190gat), .ZN(new_n458));
  NAND2_X1  g257(.A1(G169gat), .A2(G176gat), .ZN(new_n459));
  NOR2_X1   g258(.A1(G169gat), .A2(G176gat), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT26), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n459), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NOR3_X1   g261(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n458), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NOR3_X1   g263(.A1(new_n456), .A2(new_n457), .A3(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT24), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n458), .A2(KEYINPUT66), .A3(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n466), .B1(new_n458), .B2(KEYINPUT66), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n442), .A2(new_n448), .ZN(new_n470));
  INV_X1    g269(.A(new_n470), .ZN(new_n471));
  NOR3_X1   g270(.A1(new_n468), .A2(new_n469), .A3(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT25), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n473), .B1(new_n460), .B2(KEYINPUT23), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT23), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n475), .B1(G169gat), .B2(G176gat), .ZN(new_n476));
  AOI21_X1  g275(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n477));
  NAND3_X1  g276(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  OAI211_X1 g278(.A(new_n474), .B(new_n476), .C1(new_n477), .C2(new_n479), .ZN(new_n480));
  OAI21_X1  g279(.A(KEYINPUT67), .B1(new_n472), .B2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(G176gat), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n295), .A2(new_n482), .A3(KEYINPUT23), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n483), .A2(new_n476), .A3(KEYINPUT25), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n479), .A2(new_n477), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT67), .ZN(new_n487));
  INV_X1    g286(.A(new_n469), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n488), .A2(new_n467), .A3(new_n470), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n486), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n458), .A2(new_n466), .ZN(new_n491));
  NAND3_X1  g290(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n491), .A2(new_n470), .A3(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT64), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n491), .A2(new_n470), .A3(KEYINPUT64), .A4(new_n492), .ZN(new_n496));
  AND3_X1   g295(.A1(new_n483), .A2(new_n476), .A3(new_n459), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n495), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  AOI22_X1  g297(.A1(new_n481), .A2(new_n490), .B1(new_n473), .B2(new_n498), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n439), .B1(new_n465), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(G227gat), .A2(G233gat), .ZN(new_n501));
  INV_X1    g300(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n498), .A2(new_n473), .ZN(new_n503));
  NOR3_X1   g302(.A1(new_n472), .A2(new_n480), .A3(KEYINPUT67), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n487), .B1(new_n486), .B2(new_n489), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n503), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  OAI21_X1  g305(.A(KEYINPUT68), .B1(new_n452), .B2(new_n453), .ZN(new_n507));
  AOI21_X1  g306(.A(G190gat), .B1(new_n443), .B2(new_n441), .ZN(new_n508));
  AOI21_X1  g307(.A(KEYINPUT28), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NOR4_X1   g308(.A1(new_n452), .A2(new_n453), .A3(new_n440), .A4(G190gat), .ZN(new_n510));
  OAI21_X1  g309(.A(KEYINPUT69), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n450), .A2(new_n451), .A3(new_n455), .ZN(new_n512));
  INV_X1    g311(.A(new_n464), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n511), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n429), .A2(new_n437), .ZN(new_n515));
  INV_X1    g314(.A(new_n430), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(new_n431), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n506), .A2(new_n514), .A3(new_n518), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n500), .A2(new_n502), .A3(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT33), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  XOR2_X1   g321(.A(G15gat), .B(G43gat), .Z(new_n523));
  XNOR2_X1  g322(.A(G71gat), .B(G99gat), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n523), .B(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n522), .A2(new_n525), .ZN(new_n526));
  AND3_X1   g325(.A1(new_n506), .A2(new_n514), .A3(new_n518), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n518), .B1(new_n506), .B2(new_n514), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n501), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n529), .A2(KEYINPUT34), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n500), .A2(new_n519), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT34), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n531), .A2(new_n532), .A3(new_n501), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n520), .A2(KEYINPUT32), .ZN(new_n534));
  AND3_X1   g333(.A1(new_n530), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n534), .B1(new_n530), .B2(new_n533), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n526), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  AND2_X1   g336(.A1(new_n520), .A2(KEYINPUT32), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n532), .B1(new_n531), .B2(new_n501), .ZN(new_n539));
  AOI211_X1 g338(.A(KEYINPUT34), .B(new_n502), .C1(new_n500), .C2(new_n519), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n526), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n530), .A2(new_n533), .A3(new_n534), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  NAND4_X1  g343(.A1(new_n424), .A2(new_n537), .A3(KEYINPUT84), .A4(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT76), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n517), .A2(new_n547), .A3(new_n431), .ZN(new_n548));
  OAI21_X1  g347(.A(KEYINPUT76), .B1(new_n432), .B2(new_n438), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n405), .A2(KEYINPUT3), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n550), .A2(new_n551), .A3(new_n386), .ZN(new_n552));
  NAND2_X1  g351(.A1(G225gat), .A2(G233gat), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n554), .A2(KEYINPUT5), .ZN(new_n555));
  NAND4_X1  g354(.A1(new_n400), .A2(new_n517), .A3(new_n401), .A4(new_n431), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(KEYINPUT4), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT78), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT4), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n384), .A2(new_n439), .A3(new_n559), .ZN(new_n560));
  AND3_X1   g359(.A1(new_n557), .A2(new_n558), .A3(new_n560), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n558), .B1(new_n557), .B2(new_n560), .ZN(new_n562));
  OAI211_X1 g361(.A(new_n552), .B(new_n555), .C1(new_n561), .C2(new_n562), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n384), .B1(new_n549), .B2(new_n548), .ZN(new_n564));
  INV_X1    g363(.A(new_n556), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n554), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n556), .A2(KEYINPUT4), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n559), .B1(new_n384), .B2(new_n439), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n553), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  AND3_X1   g368(.A1(new_n550), .A2(new_n551), .A3(new_n386), .ZN(new_n570));
  OAI211_X1 g369(.A(KEYINPUT5), .B(new_n566), .C1(new_n569), .C2(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(G1gat), .B(G29gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n572), .B(KEYINPUT0), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n573), .B(G57gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n574), .B(new_n223), .ZN(new_n575));
  AND3_X1   g374(.A1(new_n563), .A2(new_n571), .A3(new_n575), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n575), .B1(new_n563), .B2(new_n571), .ZN(new_n577));
  NOR3_X1   g376(.A1(new_n576), .A2(new_n577), .A3(KEYINPUT6), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT6), .ZN(new_n579));
  AOI211_X1 g378(.A(new_n579), .B(new_n575), .C1(new_n563), .C2(new_n571), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(G226gat), .A2(G233gat), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n506), .A2(new_n514), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n583), .B1(new_n584), .B2(new_n387), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n450), .A2(new_n455), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n464), .B1(new_n586), .B2(KEYINPUT69), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n481), .A2(new_n490), .ZN(new_n588));
  AOI22_X1  g387(.A1(new_n512), .A2(new_n587), .B1(new_n588), .B2(new_n503), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n589), .A2(new_n582), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n397), .B1(new_n585), .B2(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(G8gat), .B(G36gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n592), .B(G64gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(new_n224), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n364), .B1(new_n589), .B2(new_n582), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT73), .ZN(new_n596));
  NOR3_X1   g395(.A1(new_n595), .A2(new_n585), .A3(new_n596), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n582), .B1(new_n589), .B2(KEYINPUT29), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n397), .B1(new_n584), .B2(new_n583), .ZN(new_n599));
  AOI21_X1  g398(.A(KEYINPUT73), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  OAI211_X1 g399(.A(new_n591), .B(new_n594), .C1(new_n597), .C2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT30), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n596), .B1(new_n595), .B2(new_n585), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n598), .A2(KEYINPUT73), .A3(new_n599), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n584), .A2(new_n583), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n598), .A2(new_n606), .ZN(new_n607));
  AOI22_X1  g406(.A1(new_n604), .A2(new_n605), .B1(new_n607), .B2(new_n397), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n608), .A2(KEYINPUT30), .A3(new_n594), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n591), .B1(new_n597), .B2(new_n600), .ZN(new_n610));
  INV_X1    g409(.A(new_n594), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n603), .A2(new_n609), .A3(new_n612), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n581), .A2(new_n613), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n345), .B1(new_n546), .B2(new_n614), .ZN(new_n615));
  NOR4_X1   g414(.A1(new_n545), .A2(new_n581), .A3(new_n613), .A4(KEYINPUT35), .ZN(new_n616));
  OR2_X1    g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT39), .ZN(new_n618));
  OAI21_X1  g417(.A(KEYINPUT78), .B1(new_n567), .B2(new_n568), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n557), .A2(new_n558), .A3(new_n560), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n570), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT82), .ZN(new_n622));
  NOR3_X1   g421(.A1(new_n621), .A2(new_n622), .A3(new_n553), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n552), .B1(new_n561), .B2(new_n562), .ZN(new_n624));
  AOI21_X1  g423(.A(KEYINPUT82), .B1(new_n624), .B2(new_n554), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n618), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n622), .B1(new_n621), .B2(new_n553), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n624), .A2(KEYINPUT82), .A3(new_n554), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n564), .A2(new_n565), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n618), .B1(new_n629), .B2(new_n553), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n627), .A2(new_n628), .A3(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n626), .A2(new_n575), .A3(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT40), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n577), .ZN(new_n635));
  NAND4_X1  g434(.A1(new_n626), .A2(KEYINPUT40), .A3(new_n575), .A4(new_n631), .ZN(new_n636));
  NAND4_X1  g435(.A1(new_n634), .A2(new_n635), .A3(new_n613), .A4(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n604), .A2(new_n605), .ZN(new_n638));
  AOI21_X1  g437(.A(KEYINPUT37), .B1(new_n607), .B2(new_n397), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n594), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n598), .A2(new_n599), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n591), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g441(.A(KEYINPUT38), .B1(new_n642), .B2(KEYINPUT37), .ZN(new_n643));
  AOI22_X1  g442(.A1(new_n640), .A2(new_n643), .B1(new_n608), .B2(new_n594), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT38), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n610), .A2(KEYINPUT37), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n645), .B1(new_n646), .B2(new_n640), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT83), .ZN(new_n648));
  OAI211_X1 g447(.A(new_n581), .B(new_n644), .C1(new_n647), .C2(new_n648), .ZN(new_n649));
  AOI211_X1 g448(.A(KEYINPUT83), .B(new_n645), .C1(new_n646), .C2(new_n640), .ZN(new_n650));
  OAI211_X1 g449(.A(new_n637), .B(new_n424), .C1(new_n649), .C2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n424), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n652), .B1(new_n581), .B2(new_n613), .ZN(new_n653));
  NOR3_X1   g452(.A1(new_n535), .A2(new_n536), .A3(new_n526), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n542), .B1(new_n541), .B2(new_n543), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT71), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT36), .ZN(new_n657));
  OAI22_X1  g456(.A1(new_n654), .A2(new_n655), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  XOR2_X1   g457(.A(KEYINPUT71), .B(KEYINPUT36), .Z(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n537), .A2(new_n544), .A3(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n651), .A2(new_n653), .A3(new_n662), .ZN(new_n663));
  AOI211_X1 g462(.A(new_n303), .B(new_n344), .C1(new_n617), .C2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(new_n581), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(G1gat), .ZN(G1324gat));
  OR2_X1    g465(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n667));
  NAND2_X1  g466(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n668));
  NAND4_X1  g467(.A1(new_n664), .A2(new_n613), .A3(new_n667), .A4(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT42), .ZN(new_n670));
  OR2_X1    g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n664), .ZN(new_n672));
  INV_X1    g471(.A(new_n613), .ZN(new_n673));
  OAI21_X1  g472(.A(G8gat), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n669), .A2(new_n670), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n671), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(KEYINPUT96), .ZN(G1325gat));
  INV_X1    g476(.A(G15gat), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n654), .A2(new_n655), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n664), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  AND3_X1   g479(.A1(new_n537), .A2(new_n544), .A3(new_n660), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n656), .A2(new_n657), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n682), .B1(new_n537), .B2(new_n544), .ZN(new_n683));
  OAI21_X1  g482(.A(KEYINPUT97), .B1(new_n681), .B2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT97), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n658), .A2(new_n685), .A3(new_n661), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT98), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n687), .B(new_n688), .ZN(new_n689));
  AND2_X1   g488(.A1(new_n664), .A2(new_n689), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n680), .B1(new_n690), .B2(new_n678), .ZN(G1326gat));
  NAND2_X1  g490(.A1(new_n664), .A2(new_n652), .ZN(new_n692));
  XOR2_X1   g491(.A(KEYINPUT43), .B(G22gat), .Z(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(KEYINPUT99), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n692), .B(new_n694), .ZN(G1327gat));
  INV_X1    g494(.A(KEYINPUT44), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n342), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n615), .A2(new_n616), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n651), .A2(new_n687), .A3(new_n653), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n698), .B1(new_n699), .B2(KEYINPUT100), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT100), .ZN(new_n701));
  NAND4_X1  g500(.A1(new_n651), .A2(new_n687), .A3(new_n701), .A4(new_n653), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n697), .B1(new_n700), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n617), .A2(new_n663), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n696), .B1(new_n704), .B2(new_n342), .ZN(new_n705));
  OR2_X1    g504(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n328), .A2(new_n303), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(new_n581), .ZN(new_n709));
  OAI21_X1  g508(.A(G29gat), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  AND3_X1   g509(.A1(new_n704), .A2(new_n342), .A3(new_n707), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n711), .A2(new_n264), .A3(new_n581), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n712), .B(KEYINPUT45), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n710), .A2(new_n713), .ZN(G1328gat));
  NAND3_X1  g513(.A1(new_n711), .A2(new_n265), .A3(new_n613), .ZN(new_n715));
  XOR2_X1   g514(.A(KEYINPUT101), .B(KEYINPUT46), .Z(new_n716));
  XNOR2_X1  g515(.A(new_n715), .B(new_n716), .ZN(new_n717));
  AND2_X1   g516(.A1(new_n706), .A2(new_n707), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(new_n613), .ZN(new_n719));
  INV_X1    g518(.A(new_n719), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n717), .B1(new_n720), .B2(new_n265), .ZN(G1329gat));
  INV_X1    g520(.A(G43gat), .ZN(new_n722));
  AND3_X1   g521(.A1(new_n711), .A2(new_n722), .A3(new_n679), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT47), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(new_n687), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n718), .A2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(new_n727), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n725), .B1(new_n728), .B2(new_n722), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n718), .A2(new_n689), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n723), .B1(new_n730), .B2(G43gat), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n729), .B1(KEYINPUT47), .B2(new_n731), .ZN(G1330gat));
  NAND3_X1  g531(.A1(new_n711), .A2(new_n413), .A3(new_n652), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n718), .A2(new_n652), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT102), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n735), .B1(new_n708), .B2(new_n424), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(G50gat), .ZN(new_n738));
  OAI211_X1 g537(.A(KEYINPUT48), .B(new_n733), .C1(new_n736), .C2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n734), .A2(G50gat), .ZN(new_n740));
  AND2_X1   g539(.A1(new_n740), .A2(new_n733), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n739), .B1(KEYINPUT48), .B2(new_n741), .ZN(G1331gat));
  NAND2_X1  g541(.A1(new_n700), .A2(new_n702), .ZN(new_n743));
  NOR3_X1   g542(.A1(new_n344), .A2(new_n253), .A3(new_n302), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT103), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n743), .A2(KEYINPUT103), .A3(new_n744), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  XOR2_X1   g548(.A(new_n581), .B(KEYINPUT104), .Z(new_n750));
  INV_X1    g549(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  XOR2_X1   g551(.A(KEYINPUT105), .B(G57gat), .Z(new_n753));
  XNOR2_X1  g552(.A(new_n752), .B(new_n753), .ZN(G1332gat));
  OR2_X1    g553(.A1(new_n673), .A2(KEYINPUT106), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n673), .A2(KEYINPUT106), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n749), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g558(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n760));
  AND2_X1   g559(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n759), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n762), .B1(new_n759), .B2(new_n760), .ZN(G1333gat));
  INV_X1    g562(.A(new_n689), .ZN(new_n764));
  NOR3_X1   g563(.A1(new_n749), .A2(new_n206), .A3(new_n764), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n747), .A2(new_n679), .A3(new_n748), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT107), .ZN(new_n767));
  OR2_X1    g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  AOI21_X1  g567(.A(G71gat), .B1(new_n766), .B2(new_n767), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n765), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  XNOR2_X1  g569(.A(KEYINPUT108), .B(KEYINPUT50), .ZN(new_n771));
  INV_X1    g570(.A(new_n771), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n770), .B(new_n772), .ZN(G1334gat));
  NOR2_X1   g572(.A1(new_n749), .A2(new_n424), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(new_n207), .ZN(G1335gat));
  NOR3_X1   g574(.A1(new_n253), .A2(new_n709), .A3(G85gat), .ZN(new_n776));
  INV_X1    g575(.A(new_n328), .ZN(new_n777));
  INV_X1    g576(.A(new_n302), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n779), .A2(new_n343), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n743), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n781), .B(KEYINPUT51), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(KEYINPUT110), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT51), .ZN(new_n784));
  OR3_X1    g583(.A1(new_n781), .A2(KEYINPUT110), .A3(new_n784), .ZN(new_n785));
  AND3_X1   g584(.A1(new_n783), .A2(KEYINPUT111), .A3(new_n785), .ZN(new_n786));
  AOI21_X1  g585(.A(KEYINPUT111), .B1(new_n783), .B2(new_n785), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n776), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n779), .A2(new_n253), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n789), .B1(new_n703), .B2(new_n705), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT109), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  OAI211_X1 g591(.A(KEYINPUT109), .B(new_n789), .C1(new_n703), .C2(new_n705), .ZN(new_n793));
  AND3_X1   g592(.A1(new_n792), .A2(new_n581), .A3(new_n793), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n788), .B1(new_n223), .B2(new_n794), .ZN(G1336gat));
  NAND3_X1  g594(.A1(new_n706), .A2(new_n757), .A3(new_n789), .ZN(new_n796));
  AOI21_X1  g595(.A(KEYINPUT52), .B1(new_n796), .B2(G92gat), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n783), .A2(new_n785), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n757), .A2(new_n224), .A3(new_n252), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n797), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n792), .A2(new_n613), .A3(new_n793), .ZN(new_n801));
  AND3_X1   g600(.A1(new_n801), .A2(KEYINPUT112), .A3(G92gat), .ZN(new_n802));
  AOI21_X1  g601(.A(KEYINPUT112), .B1(new_n801), .B2(G92gat), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n782), .A2(new_n799), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n802), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT52), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n800), .B1(new_n805), .B2(new_n806), .ZN(G1337gat));
  INV_X1    g606(.A(new_n679), .ZN(new_n808));
  NOR3_X1   g607(.A1(new_n808), .A2(new_n253), .A3(G99gat), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n809), .B1(new_n786), .B2(new_n787), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n792), .A2(new_n689), .A3(new_n793), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(G99gat), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n810), .A2(new_n812), .ZN(G1338gat));
  XOR2_X1   g612(.A(KEYINPUT113), .B(G106gat), .Z(new_n814));
  NAND3_X1  g613(.A1(new_n706), .A2(new_n652), .A3(new_n789), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n814), .B1(new_n815), .B2(KEYINPUT114), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n816), .B1(KEYINPUT114), .B2(new_n815), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT53), .ZN(new_n818));
  NOR3_X1   g617(.A1(new_n253), .A2(G106gat), .A3(new_n424), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n783), .A2(new_n785), .A3(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n817), .A2(new_n818), .A3(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(new_n782), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n792), .A2(new_n652), .A3(new_n793), .ZN(new_n823));
  INV_X1    g622(.A(new_n814), .ZN(new_n824));
  AOI22_X1  g623(.A1(new_n822), .A2(new_n819), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n821), .B1(new_n818), .B2(new_n825), .ZN(G1339gat));
  INV_X1    g625(.A(new_n240), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n236), .A2(new_n827), .A3(new_n238), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n241), .A2(KEYINPUT54), .A3(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n827), .B1(new_n236), .B2(new_n238), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT54), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n248), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n829), .A2(KEYINPUT55), .A3(new_n832), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n833), .A2(new_n251), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n255), .B1(new_n287), .B2(new_n276), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n289), .A2(new_n290), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n297), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  AND2_X1   g636(.A1(new_n301), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n829), .A2(new_n832), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT55), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n834), .A2(new_n342), .A3(new_n838), .A4(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n841), .A2(new_n251), .A3(new_n302), .A4(new_n833), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n252), .A2(new_n838), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n342), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n777), .B1(new_n843), .B2(new_n846), .ZN(new_n847));
  NAND4_X1  g646(.A1(new_n328), .A2(new_n343), .A3(new_n253), .A4(new_n778), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(new_n750), .ZN(new_n850));
  NOR3_X1   g649(.A1(new_n850), .A2(new_n652), .A3(new_n808), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(new_n758), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n433), .B1(new_n852), .B2(new_n778), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n652), .B1(new_n847), .B2(new_n848), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n757), .A2(new_n709), .ZN(new_n855));
  INV_X1    g654(.A(new_n855), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n856), .A2(new_n808), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n854), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n302), .A2(G113gat), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n853), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  XNOR2_X1  g659(.A(new_n860), .B(KEYINPUT115), .ZN(G1340gat));
  NOR3_X1   g660(.A1(new_n858), .A2(new_n434), .A3(new_n253), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n851), .A2(new_n252), .A3(new_n758), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n862), .B1(new_n863), .B2(new_n434), .ZN(G1341gat));
  OAI21_X1  g663(.A(G127gat), .B1(new_n858), .B2(new_n777), .ZN(new_n865));
  OR2_X1    g664(.A1(new_n777), .A2(G127gat), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n865), .B1(new_n852), .B2(new_n866), .ZN(G1342gat));
  NOR3_X1   g666(.A1(new_n343), .A2(G134gat), .A3(new_n613), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n851), .A2(new_n868), .ZN(new_n869));
  OR2_X1    g668(.A1(new_n869), .A2(KEYINPUT56), .ZN(new_n870));
  OAI21_X1  g669(.A(G134gat), .B1(new_n858), .B2(new_n343), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n869), .A2(KEYINPUT56), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n870), .A2(new_n871), .A3(new_n872), .ZN(G1343gat));
  INV_X1    g672(.A(KEYINPUT118), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n850), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n689), .A2(new_n424), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n849), .A2(KEYINPUT118), .A3(new_n750), .ZN(new_n877));
  NAND4_X1  g676(.A1(new_n875), .A2(new_n758), .A3(new_n876), .A4(new_n877), .ZN(new_n878));
  NOR3_X1   g677(.A1(new_n878), .A2(G141gat), .A3(new_n778), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n424), .A2(KEYINPUT57), .ZN(new_n880));
  AOI211_X1 g679(.A(new_n726), .B(new_n856), .C1(new_n849), .C2(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(KEYINPUT116), .B1(new_n839), .B2(new_n840), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT116), .ZN(new_n883));
  AOI211_X1 g682(.A(new_n883), .B(KEYINPUT55), .C1(new_n829), .C2(new_n832), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n834), .B1(new_n882), .B2(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT117), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  OAI211_X1 g686(.A(new_n834), .B(KEYINPUT117), .C1(new_n882), .C2(new_n884), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n887), .A2(new_n302), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n342), .B1(new_n889), .B2(new_n845), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n777), .B1(new_n890), .B2(new_n843), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n424), .B1(new_n891), .B2(new_n848), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT57), .ZN(new_n893));
  OAI211_X1 g692(.A(new_n302), .B(new_n881), .C1(new_n892), .C2(new_n893), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n879), .B1(new_n894), .B2(new_n381), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT119), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n896), .B1(new_n894), .B2(new_n381), .ZN(new_n897));
  NOR3_X1   g696(.A1(new_n895), .A2(new_n897), .A3(KEYINPUT58), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT58), .ZN(new_n899));
  AOI221_X4 g698(.A(new_n879), .B1(new_n896), .B2(new_n899), .C1(new_n381), .C2(new_n894), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n898), .A2(new_n900), .ZN(G1344gat));
  INV_X1    g700(.A(KEYINPUT59), .ZN(new_n902));
  XNOR2_X1  g701(.A(new_n848), .B(KEYINPUT121), .ZN(new_n903));
  AND2_X1   g702(.A1(new_n888), .A2(new_n302), .ZN(new_n904));
  AOI22_X1  g703(.A1(new_n904), .A2(new_n887), .B1(new_n252), .B2(new_n838), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n842), .B1(new_n905), .B2(new_n342), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n903), .B1(new_n906), .B2(new_n777), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n893), .B1(new_n907), .B2(new_n424), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n849), .A2(KEYINPUT57), .A3(new_n652), .ZN(new_n909));
  XNOR2_X1  g708(.A(new_n909), .B(KEYINPUT120), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  NAND4_X1  g710(.A1(new_n911), .A2(new_n252), .A3(new_n687), .A4(new_n855), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n902), .B1(new_n912), .B2(G148gat), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n881), .B1(new_n892), .B2(new_n893), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n914), .A2(new_n253), .ZN(new_n915));
  NOR3_X1   g714(.A1(new_n915), .A2(KEYINPUT59), .A3(new_n370), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n252), .A2(new_n370), .ZN(new_n917));
  OAI22_X1  g716(.A1(new_n913), .A2(new_n916), .B1(new_n878), .B2(new_n917), .ZN(G1345gat));
  OAI21_X1  g717(.A(G155gat), .B1(new_n914), .B2(new_n777), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n328), .A2(new_n376), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n919), .B1(new_n878), .B2(new_n920), .ZN(G1346gat));
  OAI21_X1  g720(.A(G162gat), .B1(new_n914), .B2(new_n343), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n342), .A2(new_n377), .A3(new_n673), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n922), .B1(new_n923), .B2(new_n924), .ZN(G1347gat));
  AOI21_X1  g724(.A(new_n581), .B1(new_n847), .B2(new_n848), .ZN(new_n926));
  NOR3_X1   g725(.A1(new_n758), .A2(new_n652), .A3(new_n808), .ZN(new_n927));
  AND2_X1   g726(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g727(.A(G169gat), .B1(new_n928), .B2(new_n302), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n751), .A2(new_n613), .A3(new_n679), .ZN(new_n930));
  INV_X1    g729(.A(new_n930), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n854), .A2(new_n931), .ZN(new_n932));
  NOR3_X1   g731(.A1(new_n932), .A2(new_n295), .A3(new_n778), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n929), .A2(new_n933), .ZN(G1348gat));
  NAND3_X1  g733(.A1(new_n928), .A2(new_n482), .A3(new_n252), .ZN(new_n935));
  OAI21_X1  g734(.A(G176gat), .B1(new_n932), .B2(new_n253), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(G1349gat));
  AND2_X1   g736(.A1(new_n328), .A2(new_n454), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n928), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n939), .A2(KEYINPUT122), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT122), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n928), .A2(new_n941), .A3(new_n938), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT124), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n854), .A2(new_n328), .A3(new_n931), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n442), .B1(new_n945), .B2(KEYINPUT123), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n946), .B1(KEYINPUT123), .B2(new_n945), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n943), .A2(new_n944), .A3(new_n947), .ZN(new_n948));
  INV_X1    g747(.A(new_n948), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n944), .B1(new_n943), .B2(new_n947), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT60), .ZN(new_n951));
  NOR3_X1   g750(.A1(new_n949), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n943), .A2(new_n947), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(KEYINPUT124), .ZN(new_n954));
  AOI21_X1  g753(.A(KEYINPUT60), .B1(new_n954), .B2(new_n948), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n952), .A2(new_n955), .ZN(G1350gat));
  OAI21_X1  g755(.A(G190gat), .B1(new_n932), .B2(new_n343), .ZN(new_n957));
  XNOR2_X1  g756(.A(new_n957), .B(KEYINPUT61), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n928), .A2(new_n448), .A3(new_n342), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n958), .A2(new_n959), .ZN(G1351gat));
  NOR3_X1   g759(.A1(new_n689), .A2(new_n673), .A3(new_n750), .ZN(new_n961));
  XNOR2_X1  g760(.A(new_n961), .B(KEYINPUT126), .ZN(new_n962));
  AND2_X1   g761(.A1(new_n911), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n963), .A2(new_n302), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n964), .A2(G197gat), .ZN(new_n965));
  AND3_X1   g764(.A1(new_n876), .A2(new_n757), .A3(new_n926), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n966), .A2(new_n347), .A3(new_n302), .ZN(new_n967));
  XOR2_X1   g766(.A(new_n967), .B(KEYINPUT125), .Z(new_n968));
  NAND2_X1  g767(.A1(new_n965), .A2(new_n968), .ZN(G1352gat));
  NAND3_X1  g768(.A1(new_n966), .A2(new_n247), .A3(new_n252), .ZN(new_n970));
  XOR2_X1   g769(.A(new_n970), .B(KEYINPUT62), .Z(new_n971));
  XOR2_X1   g770(.A(new_n848), .B(KEYINPUT121), .Z(new_n972));
  NAND2_X1  g771(.A1(new_n891), .A2(new_n972), .ZN(new_n973));
  AOI21_X1  g772(.A(KEYINPUT57), .B1(new_n973), .B2(new_n652), .ZN(new_n974));
  INV_X1    g773(.A(KEYINPUT120), .ZN(new_n975));
  XNOR2_X1  g774(.A(new_n909), .B(new_n975), .ZN(new_n976));
  OAI211_X1 g775(.A(new_n252), .B(new_n962), .C1(new_n974), .C2(new_n976), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n977), .A2(G204gat), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n971), .A2(new_n978), .ZN(new_n979));
  INV_X1    g778(.A(KEYINPUT127), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n971), .A2(new_n978), .A3(KEYINPUT127), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n981), .A2(new_n982), .ZN(G1353gat));
  NAND3_X1  g782(.A1(new_n966), .A2(new_n315), .A3(new_n328), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n911), .A2(new_n328), .A3(new_n962), .ZN(new_n985));
  AND3_X1   g784(.A1(new_n985), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n986));
  AOI21_X1  g785(.A(KEYINPUT63), .B1(new_n985), .B2(G211gat), .ZN(new_n987));
  OAI21_X1  g786(.A(new_n984), .B1(new_n986), .B2(new_n987), .ZN(G1354gat));
  AOI21_X1  g787(.A(G218gat), .B1(new_n966), .B2(new_n342), .ZN(new_n989));
  NOR2_X1   g788(.A1(new_n343), .A2(new_n356), .ZN(new_n990));
  AOI21_X1  g789(.A(new_n989), .B1(new_n963), .B2(new_n990), .ZN(G1355gat));
endmodule


