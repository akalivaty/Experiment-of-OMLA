//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 1 1 1 1 0 0 0 1 1 0 0 1 1 1 0 0 0 0 1 0 0 1 0 1 0 0 0 1 0 1 0 1 0 0 0 1 0 1 1 0 0 0 1 0 1 0 1 1 1 0 0 0 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:31 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n449, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n558, new_n560, new_n561, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n615, new_n616,
    new_n619, new_n621, new_n622, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n855, new_n856, new_n857,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT64), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT65), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT66), .Z(G217));
  NOR4_X1   g025(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT67), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n453), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n453), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  NAND2_X1  g035(.A1(G113), .A2(G2104), .ZN(new_n461));
  XOR2_X1   g036(.A(new_n461), .B(KEYINPUT68), .Z(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  AND3_X1   g041(.A1(new_n464), .A2(new_n466), .A3(G125), .ZN(new_n467));
  OAI21_X1  g042(.A(G2105), .B1(new_n462), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n464), .A2(new_n466), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n463), .A2(G2105), .ZN(new_n471));
  AOI22_X1  g046(.A1(new_n470), .A2(G137), .B1(G101), .B2(new_n471), .ZN(new_n472));
  AND2_X1   g047(.A1(new_n468), .A2(new_n472), .ZN(G160));
  NAND2_X1  g048(.A1(new_n470), .A2(G136), .ZN(new_n474));
  INV_X1    g049(.A(G2105), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n469), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  NOR2_X1   g052(.A1(G100), .A2(G2105), .ZN(new_n478));
  OAI21_X1  g053(.A(G2104), .B1(new_n475), .B2(G112), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n474), .B(new_n477), .C1(new_n478), .C2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G162));
  INV_X1    g056(.A(KEYINPUT69), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n471), .A2(G102), .ZN(new_n483));
  NAND2_X1  g058(.A1(G114), .A2(G2104), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  XNOR2_X1  g060(.A(KEYINPUT3), .B(G2104), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n485), .B1(new_n486), .B2(G126), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n483), .B1(new_n487), .B2(new_n475), .ZN(new_n488));
  NAND4_X1  g063(.A1(new_n464), .A2(new_n466), .A3(G138), .A4(new_n475), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n486), .A2(KEYINPUT4), .A3(G138), .A4(new_n475), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n482), .B1(new_n488), .B2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(new_n483), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n464), .A2(new_n466), .A3(G126), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(new_n484), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n495), .B1(new_n497), .B2(G2105), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n498), .A2(KEYINPUT69), .A3(new_n491), .A4(new_n492), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n494), .A2(new_n499), .ZN(G164));
  INV_X1    g075(.A(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT5), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G543), .ZN(new_n504));
  AND2_X1   g079(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  XNOR2_X1  g080(.A(KEYINPUT6), .B(G651), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(G88), .ZN(new_n508));
  INV_X1    g083(.A(G50), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n506), .A2(G543), .ZN(new_n510));
  OAI22_X1  g085(.A1(new_n507), .A2(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G651), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n505), .A2(G62), .ZN(new_n513));
  NAND2_X1  g088(.A1(G75), .A2(G543), .ZN(new_n514));
  XNOR2_X1  g089(.A(new_n514), .B(KEYINPUT70), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n512), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n511), .A2(new_n516), .ZN(G166));
  NAND2_X1  g092(.A1(new_n505), .A2(KEYINPUT71), .ZN(new_n518));
  AOI21_X1  g093(.A(KEYINPUT71), .B1(new_n502), .B2(new_n504), .ZN(new_n519));
  INV_X1    g094(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n521), .A2(G63), .A3(G651), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n510), .A2(KEYINPUT72), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT72), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n506), .A2(new_n524), .A3(G543), .ZN(new_n525));
  XOR2_X1   g100(.A(KEYINPUT73), .B(G51), .Z(new_n526));
  NAND3_X1  g101(.A1(new_n523), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n505), .A2(G89), .A3(new_n506), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT74), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n530), .B(KEYINPUT7), .ZN(new_n531));
  AND3_X1   g106(.A1(new_n528), .A2(new_n529), .A3(new_n531), .ZN(new_n532));
  AOI21_X1  g107(.A(new_n529), .B1(new_n528), .B2(new_n531), .ZN(new_n533));
  OAI211_X1 g108(.A(new_n522), .B(new_n527), .C1(new_n532), .C2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(KEYINPUT75), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n528), .A2(new_n531), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(KEYINPUT74), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n528), .A2(new_n529), .A3(new_n531), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT75), .ZN(new_n540));
  NAND4_X1  g115(.A1(new_n539), .A2(new_n540), .A3(new_n527), .A4(new_n522), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n535), .A2(new_n541), .ZN(G168));
  AOI22_X1  g117(.A1(new_n521), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n543), .A2(new_n512), .ZN(new_n544));
  AND2_X1   g119(.A1(new_n505), .A2(new_n506), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G90), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n523), .A2(new_n525), .ZN(new_n547));
  INV_X1    g122(.A(G52), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n544), .A2(new_n549), .ZN(G171));
  NAND2_X1  g125(.A1(new_n545), .A2(G81), .ZN(new_n551));
  INV_X1    g126(.A(G43), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n551), .B1(new_n547), .B2(new_n552), .ZN(new_n553));
  AOI22_X1  g128(.A1(new_n521), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  AOI21_X1  g130(.A(new_n553), .B1(new_n555), .B2(G651), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  AND3_X1   g132(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G36), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n558), .A2(new_n561), .ZN(G188));
  NAND2_X1  g137(.A1(new_n545), .A2(G91), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT76), .ZN(new_n564));
  INV_X1    g139(.A(new_n510), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G53), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT9), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n505), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT77), .ZN(new_n569));
  OAI211_X1 g144(.A(new_n564), .B(new_n567), .C1(new_n512), .C2(new_n569), .ZN(G299));
  OR2_X1    g145(.A1(new_n544), .A2(new_n549), .ZN(G301));
  INV_X1    g146(.A(G168), .ZN(G286));
  INV_X1    g147(.A(G166), .ZN(G303));
  INV_X1    g148(.A(G74), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n518), .A2(new_n574), .A3(new_n520), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT78), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n575), .A2(new_n576), .A3(G651), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n565), .A2(G49), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n576), .B1(new_n575), .B2(G651), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(G87), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n507), .A2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n581), .A2(new_n584), .ZN(G288));
  INV_X1    g160(.A(KEYINPUT79), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n505), .A2(new_n586), .A3(G61), .ZN(new_n587));
  NAND2_X1  g162(.A1(G73), .A2(G543), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n502), .A2(new_n504), .ZN(new_n589));
  INV_X1    g164(.A(G61), .ZN(new_n590));
  OAI21_X1  g165(.A(KEYINPUT79), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n587), .A2(new_n588), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n592), .A2(G651), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n545), .A2(G86), .ZN(new_n594));
  AND3_X1   g169(.A1(new_n506), .A2(G48), .A3(G543), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n593), .A2(new_n594), .A3(new_n596), .ZN(G305));
  AOI22_X1  g172(.A1(new_n521), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n598), .A2(new_n512), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n545), .A2(G85), .ZN(new_n600));
  INV_X1    g175(.A(G47), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n547), .B2(new_n601), .ZN(new_n602));
  OR2_X1    g177(.A1(new_n599), .A2(new_n602), .ZN(G290));
  NAND2_X1  g178(.A1(G301), .A2(G868), .ZN(new_n604));
  INV_X1    g179(.A(G92), .ZN(new_n605));
  NOR2_X1   g180(.A1(new_n507), .A2(new_n605), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(KEYINPUT10), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n523), .A2(G54), .A3(new_n525), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n505), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n609));
  OR2_X1    g184(.A1(new_n609), .A2(new_n512), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n607), .A2(new_n608), .A3(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n604), .B1(G868), .B2(new_n612), .ZN(G284));
  OAI21_X1  g188(.A(new_n604), .B1(G868), .B2(new_n612), .ZN(G321));
  NAND2_X1  g189(.A1(G286), .A2(G868), .ZN(new_n615));
  XOR2_X1   g190(.A(G299), .B(KEYINPUT80), .Z(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n616), .B2(G868), .ZN(G297));
  XNOR2_X1  g192(.A(G297), .B(KEYINPUT81), .ZN(G280));
  INV_X1    g193(.A(G559), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n612), .B1(new_n619), .B2(G860), .ZN(G148));
  NAND2_X1  g195(.A1(new_n612), .A2(new_n619), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n621), .A2(G868), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(G868), .B2(new_n556), .ZN(G323));
  XNOR2_X1  g198(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g199(.A1(new_n486), .A2(new_n471), .ZN(new_n625));
  XOR2_X1   g200(.A(new_n625), .B(KEYINPUT12), .Z(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(KEYINPUT13), .Z(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2100), .ZN(new_n628));
  OR2_X1    g203(.A1(new_n475), .A2(G111), .ZN(new_n629));
  INV_X1    g204(.A(KEYINPUT82), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n463), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  OAI221_X1 g206(.A(new_n631), .B1(new_n630), .B2(new_n629), .C1(G99), .C2(G2105), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n470), .A2(G135), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n476), .A2(G123), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n632), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n635), .B(G2096), .Z(new_n636));
  NAND2_X1  g211(.A1(new_n628), .A2(new_n636), .ZN(G156));
  XOR2_X1   g212(.A(G2451), .B(G2454), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT16), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2443), .ZN(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(G2427), .B(G2430), .Z(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(KEYINPUT15), .B(G2435), .Z(new_n644));
  INV_X1    g219(.A(KEYINPUT83), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT15), .B(G2435), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n647), .A2(KEYINPUT83), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n646), .A2(G2438), .A3(new_n648), .ZN(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  AOI21_X1  g225(.A(G2438), .B1(new_n646), .B2(new_n648), .ZN(new_n651));
  OAI21_X1  g226(.A(new_n643), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n646), .A2(new_n648), .ZN(new_n653));
  INV_X1    g228(.A(G2438), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n655), .A2(new_n642), .A3(new_n649), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n652), .A2(new_n656), .A3(KEYINPUT14), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n657), .A2(G1348), .ZN(new_n658));
  INV_X1    g233(.A(G2446), .ZN(new_n659));
  INV_X1    g234(.A(G1348), .ZN(new_n660));
  NAND4_X1  g235(.A1(new_n652), .A2(new_n656), .A3(KEYINPUT14), .A4(new_n660), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n658), .A2(new_n659), .A3(new_n661), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(KEYINPUT84), .B(G1341), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n659), .B1(new_n658), .B2(new_n661), .ZN(new_n666));
  NOR3_X1   g241(.A1(new_n663), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n658), .A2(new_n661), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n668), .A2(G2446), .ZN(new_n669));
  AOI21_X1  g244(.A(new_n664), .B1(new_n669), .B2(new_n662), .ZN(new_n670));
  OAI21_X1  g245(.A(new_n641), .B1(new_n667), .B2(new_n670), .ZN(new_n671));
  OAI21_X1  g246(.A(new_n665), .B1(new_n663), .B2(new_n666), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n669), .A2(new_n664), .A3(new_n662), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n672), .A2(new_n640), .A3(new_n673), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n671), .A2(G14), .A3(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(KEYINPUT85), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND4_X1  g252(.A1(new_n671), .A2(KEYINPUT85), .A3(G14), .A4(new_n674), .ZN(new_n678));
  AND2_X1   g253(.A1(new_n677), .A2(new_n678), .ZN(G401));
  XOR2_X1   g254(.A(G2084), .B(G2090), .Z(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(G2067), .B(G2678), .Z(new_n682));
  OR2_X1    g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n681), .A2(new_n682), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n683), .A2(new_n684), .A3(KEYINPUT17), .ZN(new_n685));
  INV_X1    g260(.A(KEYINPUT18), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(G2072), .B(G2078), .Z(new_n688));
  AOI21_X1  g263(.A(new_n688), .B1(new_n683), .B2(KEYINPUT18), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n687), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(G2096), .B(G2100), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(G227));
  XNOR2_X1  g267(.A(G1971), .B(G1976), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT19), .ZN(new_n694));
  XOR2_X1   g269(.A(G1956), .B(G2474), .Z(new_n695));
  XOR2_X1   g270(.A(G1961), .B(G1966), .Z(new_n696));
  OR2_X1    g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n694), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n695), .A2(new_n696), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n694), .A2(new_n699), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n698), .B1(KEYINPUT20), .B2(new_n700), .ZN(new_n701));
  NAND3_X1  g276(.A1(new_n694), .A2(new_n697), .A3(new_n699), .ZN(new_n702));
  OAI211_X1 g277(.A(new_n701), .B(new_n702), .C1(KEYINPUT20), .C2(new_n700), .ZN(new_n703));
  XOR2_X1   g278(.A(G1991), .B(G1996), .Z(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT86), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n703), .B(new_n705), .ZN(new_n706));
  XOR2_X1   g281(.A(G1981), .B(G1986), .Z(new_n707));
  AND2_X1   g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n706), .A2(new_n707), .ZN(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n710));
  INV_X1    g285(.A(new_n710), .ZN(new_n711));
  OR3_X1    g286(.A1(new_n708), .A2(new_n709), .A3(new_n711), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n711), .B1(new_n708), .B2(new_n709), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n712), .A2(new_n713), .ZN(G229));
  INV_X1    g289(.A(G29), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n715), .A2(G25), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n470), .A2(G131), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n476), .A2(G119), .ZN(new_n718));
  NOR2_X1   g293(.A1(G95), .A2(G2105), .ZN(new_n719));
  OAI21_X1  g294(.A(G2104), .B1(new_n475), .B2(G107), .ZN(new_n720));
  OAI211_X1 g295(.A(new_n717), .B(new_n718), .C1(new_n719), .C2(new_n720), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT87), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n716), .B1(new_n723), .B2(new_n715), .ZN(new_n724));
  XNOR2_X1  g299(.A(KEYINPUT35), .B(G1991), .ZN(new_n725));
  INV_X1    g300(.A(new_n725), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n724), .B(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(G1986), .ZN(new_n728));
  INV_X1    g303(.A(G16), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n729), .A2(G24), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n599), .A2(new_n602), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n730), .B1(new_n731), .B2(new_n729), .ZN(new_n732));
  INV_X1    g307(.A(new_n732), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n727), .B1(new_n728), .B2(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n729), .A2(G23), .ZN(new_n735));
  INV_X1    g310(.A(new_n735), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(G288), .B2(G16), .ZN(new_n737));
  INV_X1    g312(.A(KEYINPUT33), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(new_n739), .ZN(new_n740));
  AOI211_X1 g315(.A(KEYINPUT33), .B(new_n736), .C1(G288), .C2(G16), .ZN(new_n741));
  INV_X1    g316(.A(new_n741), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n740), .A2(G1976), .A3(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(G1976), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(new_n739), .B2(new_n741), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n729), .A2(G22), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(G166), .B2(new_n729), .ZN(new_n747));
  OR2_X1    g322(.A1(new_n747), .A2(G1971), .ZN(new_n748));
  AND2_X1   g323(.A1(new_n729), .A2(G6), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(G305), .B2(G16), .ZN(new_n750));
  XOR2_X1   g325(.A(KEYINPUT32), .B(G1981), .Z(new_n751));
  OR2_X1    g326(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n750), .A2(new_n751), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n747), .A2(G1971), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n752), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(new_n755), .ZN(new_n756));
  NAND4_X1  g331(.A1(new_n743), .A2(new_n745), .A3(new_n748), .A4(new_n756), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n734), .B1(new_n757), .B2(KEYINPUT34), .ZN(new_n758));
  OR2_X1    g333(.A1(new_n732), .A2(G1986), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n739), .A2(new_n741), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n755), .B1(new_n760), .B2(G1976), .ZN(new_n761));
  INV_X1    g336(.A(KEYINPUT34), .ZN(new_n762));
  NAND4_X1  g337(.A1(new_n761), .A2(new_n762), .A3(new_n748), .A4(new_n745), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n758), .A2(new_n759), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n764), .A2(KEYINPUT36), .ZN(new_n765));
  INV_X1    g340(.A(KEYINPUT36), .ZN(new_n766));
  NAND4_X1  g341(.A1(new_n758), .A2(new_n766), .A3(new_n759), .A4(new_n763), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(G299), .A2(G16), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n729), .A2(G20), .ZN(new_n770));
  NAND3_X1  g345(.A1(new_n769), .A2(KEYINPUT23), .A3(new_n770), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(KEYINPUT23), .B2(new_n770), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(G1956), .ZN(new_n773));
  OAI21_X1  g348(.A(KEYINPUT93), .B1(G5), .B2(G16), .ZN(new_n774));
  OR3_X1    g349(.A1(KEYINPUT93), .A2(G5), .A3(G16), .ZN(new_n775));
  OAI211_X1 g350(.A(new_n774), .B(new_n775), .C1(G301), .C2(new_n729), .ZN(new_n776));
  INV_X1    g351(.A(G1961), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n715), .A2(G35), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G162), .B2(new_n715), .ZN(new_n780));
  XOR2_X1   g355(.A(new_n780), .B(KEYINPUT95), .Z(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT29), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n778), .B1(new_n782), .B2(G2090), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n715), .A2(G33), .ZN(new_n784));
  AOI22_X1  g359(.A1(new_n486), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT89), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n786), .A2(G2105), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n470), .A2(G139), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n471), .A2(G103), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(KEYINPUT25), .Z(new_n790));
  AND3_X1   g365(.A1(new_n787), .A2(new_n788), .A3(new_n790), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n784), .B1(new_n791), .B2(new_n715), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(G2072), .Z(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(new_n777), .B2(new_n776), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n715), .A2(G26), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n470), .A2(G140), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n476), .A2(G128), .ZN(new_n797));
  OR2_X1    g372(.A1(G104), .A2(G2105), .ZN(new_n798));
  OAI211_X1 g373(.A(new_n798), .B(G2104), .C1(G116), .C2(new_n475), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n796), .A2(new_n797), .A3(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(new_n800), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n795), .B1(new_n801), .B2(new_n715), .ZN(new_n802));
  MUX2_X1   g377(.A(new_n795), .B(new_n802), .S(KEYINPUT28), .Z(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(G2067), .ZN(new_n804));
  NOR3_X1   g379(.A1(new_n783), .A2(new_n794), .A3(new_n804), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n612), .A2(new_n729), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(G4), .B2(new_n729), .ZN(new_n807));
  INV_X1    g382(.A(G27), .ZN(new_n808));
  OAI21_X1  g383(.A(KEYINPUT94), .B1(new_n808), .B2(G29), .ZN(new_n809));
  OR3_X1    g384(.A1(new_n808), .A2(KEYINPUT94), .A3(G29), .ZN(new_n810));
  OAI211_X1 g385(.A(new_n809), .B(new_n810), .C1(G164), .C2(new_n715), .ZN(new_n811));
  OAI22_X1  g386(.A1(new_n807), .A2(new_n660), .B1(G2078), .B2(new_n811), .ZN(new_n812));
  AND2_X1   g387(.A1(KEYINPUT24), .A2(G34), .ZN(new_n813));
  NOR2_X1   g388(.A1(KEYINPUT24), .A2(G34), .ZN(new_n814));
  NOR3_X1   g389(.A1(new_n813), .A2(new_n814), .A3(G29), .ZN(new_n815));
  INV_X1    g390(.A(new_n815), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(G160), .B2(new_n715), .ZN(new_n817));
  OR2_X1    g392(.A1(new_n817), .A2(G2084), .ZN(new_n818));
  XNOR2_X1  g393(.A(KEYINPUT31), .B(G11), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n817), .A2(G2084), .ZN(new_n820));
  INV_X1    g395(.A(new_n635), .ZN(new_n821));
  INV_X1    g396(.A(G28), .ZN(new_n822));
  OR2_X1    g397(.A1(new_n822), .A2(KEYINPUT30), .ZN(new_n823));
  AOI21_X1  g398(.A(G29), .B1(new_n822), .B2(KEYINPUT30), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT92), .ZN(new_n825));
  AOI22_X1  g400(.A1(new_n821), .A2(G29), .B1(new_n823), .B2(new_n825), .ZN(new_n826));
  NAND4_X1  g401(.A1(new_n818), .A2(new_n819), .A3(new_n820), .A4(new_n826), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n827), .B1(new_n811), .B2(G2078), .ZN(new_n828));
  NOR2_X1   g403(.A1(G29), .A2(G32), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n476), .A2(G129), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT90), .ZN(new_n831));
  NAND3_X1  g406(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n832));
  XOR2_X1   g407(.A(new_n832), .B(KEYINPUT26), .Z(new_n833));
  AOI22_X1  g408(.A1(new_n470), .A2(G141), .B1(G105), .B2(new_n471), .ZN(new_n834));
  AND3_X1   g409(.A1(new_n831), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n829), .B1(new_n835), .B2(G29), .ZN(new_n836));
  XNOR2_X1  g411(.A(KEYINPUT27), .B(G1996), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n836), .B(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n828), .A2(new_n838), .ZN(new_n839));
  AOI211_X1 g414(.A(new_n812), .B(new_n839), .C1(new_n660), .C2(new_n807), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n782), .A2(G2090), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n729), .A2(G19), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n842), .B1(new_n556), .B2(new_n729), .ZN(new_n843));
  XNOR2_X1  g418(.A(KEYINPUT88), .B(G1341), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n843), .B(new_n844), .ZN(new_n845));
  NAND4_X1  g420(.A1(new_n805), .A2(new_n840), .A3(new_n841), .A4(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n729), .A2(G21), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n847), .B1(G168), .B2(new_n729), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(G1966), .ZN(new_n849));
  XOR2_X1   g424(.A(new_n849), .B(KEYINPUT91), .Z(new_n850));
  OAI21_X1  g425(.A(new_n850), .B1(G1966), .B2(new_n848), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n846), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n768), .A2(new_n773), .A3(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(new_n853), .ZN(G311));
  NAND2_X1  g429(.A1(new_n853), .A2(KEYINPUT96), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT96), .ZN(new_n856));
  NAND4_X1  g431(.A1(new_n768), .A2(new_n856), .A3(new_n852), .A4(new_n773), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n855), .A2(new_n857), .ZN(G150));
  NAND2_X1  g433(.A1(new_n545), .A2(G93), .ZN(new_n859));
  INV_X1    g434(.A(G55), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n859), .B1(new_n547), .B2(new_n860), .ZN(new_n861));
  AND3_X1   g436(.A1(new_n502), .A2(new_n504), .A3(KEYINPUT71), .ZN(new_n862));
  OAI21_X1  g437(.A(G67), .B1(new_n862), .B2(new_n519), .ZN(new_n863));
  NAND2_X1  g438(.A1(G80), .A2(G543), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n512), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  OAI21_X1  g440(.A(KEYINPUT97), .B1(new_n861), .B2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  NOR3_X1   g442(.A1(new_n861), .A2(new_n865), .A3(KEYINPUT97), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(G860), .ZN(new_n870));
  XOR2_X1   g445(.A(new_n870), .B(KEYINPUT37), .Z(new_n871));
  NOR2_X1   g446(.A1(new_n611), .A2(new_n619), .ZN(new_n872));
  XOR2_X1   g447(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n873));
  XNOR2_X1  g448(.A(new_n872), .B(new_n873), .ZN(new_n874));
  OAI221_X1 g449(.A(new_n551), .B1(new_n547), .B2(new_n552), .C1(new_n554), .C2(new_n512), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n875), .B1(new_n867), .B2(new_n868), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n556), .B1(new_n865), .B2(new_n861), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n874), .B(new_n878), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n871), .B1(new_n879), .B2(G860), .ZN(G145));
  XNOR2_X1  g455(.A(G160), .B(KEYINPUT98), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT99), .ZN(new_n883));
  AND3_X1   g458(.A1(new_n491), .A2(new_n492), .A3(new_n883), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n883), .B1(new_n491), .B2(new_n492), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n498), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n886), .A2(new_n801), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n493), .A2(KEYINPUT99), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n491), .A2(new_n492), .A3(new_n883), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n890), .A2(new_n498), .A3(new_n800), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n887), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n831), .A2(new_n833), .A3(new_n834), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n835), .A2(new_n887), .A3(new_n891), .ZN(new_n895));
  INV_X1    g470(.A(new_n626), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(G162), .B(new_n635), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n896), .B1(new_n894), .B2(new_n895), .ZN(new_n901));
  NOR3_X1   g476(.A1(new_n898), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n894), .A2(new_n895), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n903), .A2(new_n626), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n899), .B1(new_n904), .B2(new_n897), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n470), .A2(G142), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n476), .A2(G130), .ZN(new_n907));
  OR2_X1    g482(.A1(G106), .A2(G2105), .ZN(new_n908));
  OAI211_X1 g483(.A(new_n908), .B(G2104), .C1(G118), .C2(new_n475), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n906), .A2(new_n907), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n791), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n787), .A2(new_n788), .A3(new_n790), .ZN(new_n912));
  INV_X1    g487(.A(new_n910), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n911), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(new_n723), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n911), .A2(new_n914), .A3(new_n722), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NOR3_X1   g493(.A1(new_n902), .A2(new_n905), .A3(new_n918), .ZN(new_n919));
  AND2_X1   g494(.A1(new_n916), .A2(new_n917), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n900), .B1(new_n898), .B2(new_n901), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n904), .A2(new_n899), .A3(new_n897), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n920), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n882), .B1(new_n919), .B2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(G37), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n918), .B1(new_n902), .B2(new_n905), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n921), .A2(new_n920), .A3(new_n922), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n926), .A2(new_n881), .A3(new_n927), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n924), .A2(new_n925), .A3(new_n928), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n929), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g505(.A1(new_n869), .A2(G868), .ZN(new_n931));
  NAND3_X1  g506(.A1(G290), .A2(new_n584), .A3(new_n581), .ZN(new_n932));
  NAND2_X1  g507(.A1(G288), .A2(new_n731), .ZN(new_n933));
  AOI21_X1  g508(.A(KEYINPUT101), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  XNOR2_X1  g509(.A(G305), .B(G166), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n932), .A2(new_n933), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT101), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n932), .A2(new_n933), .A3(KEYINPUT101), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n936), .B1(new_n941), .B2(new_n935), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n942), .B(KEYINPUT42), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n612), .B(G299), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT41), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  XNOR2_X1  g521(.A(G299), .B(new_n611), .ZN(new_n947));
  XNOR2_X1  g522(.A(KEYINPUT100), .B(KEYINPUT41), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n946), .A2(new_n949), .ZN(new_n950));
  XNOR2_X1  g525(.A(new_n878), .B(new_n621), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n952), .B1(new_n947), .B2(new_n951), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT102), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n943), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n953), .A2(new_n954), .ZN(new_n956));
  XOR2_X1   g531(.A(new_n955), .B(new_n956), .Z(new_n957));
  AOI21_X1  g532(.A(new_n931), .B1(new_n957), .B2(G868), .ZN(G295));
  AOI21_X1  g533(.A(new_n931), .B1(new_n957), .B2(G868), .ZN(G331));
  NAND3_X1  g534(.A1(G171), .A2(new_n535), .A3(new_n541), .ZN(new_n960));
  INV_X1    g535(.A(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(G171), .B1(new_n541), .B2(new_n535), .ZN(new_n962));
  INV_X1    g537(.A(new_n868), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n556), .B1(new_n963), .B2(new_n866), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n861), .A2(new_n865), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n875), .A2(new_n965), .ZN(new_n966));
  OAI22_X1  g541(.A1(new_n961), .A2(new_n962), .B1(new_n964), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(G168), .A2(G301), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n968), .A2(new_n876), .A3(new_n877), .A4(new_n960), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT103), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n967), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  OAI211_X1 g546(.A(new_n878), .B(KEYINPUT103), .C1(new_n961), .C2(new_n962), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n947), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  AOI22_X1  g548(.A1(new_n946), .A2(new_n949), .B1(new_n967), .B2(new_n969), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n941), .A2(new_n935), .ZN(new_n976));
  INV_X1    g551(.A(new_n936), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  AOI21_X1  g553(.A(G37), .B1(new_n975), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n947), .A2(new_n945), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n944), .A2(new_n948), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n971), .A2(new_n972), .A3(new_n980), .A4(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n967), .A2(new_n969), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n982), .B1(new_n947), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(new_n942), .ZN(new_n985));
  AND3_X1   g560(.A1(new_n979), .A2(KEYINPUT43), .A3(new_n985), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n942), .B1(new_n973), .B2(new_n974), .ZN(new_n987));
  AOI21_X1  g562(.A(KEYINPUT43), .B1(new_n979), .B2(new_n987), .ZN(new_n988));
  OAI21_X1  g563(.A(KEYINPUT44), .B1(new_n986), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n971), .A2(new_n972), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(new_n944), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n950), .A2(new_n983), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n991), .A2(new_n978), .A3(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n993), .A2(new_n925), .A3(new_n987), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(KEYINPUT43), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT43), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n979), .A2(new_n996), .A3(new_n985), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n989), .B1(new_n999), .B2(KEYINPUT44), .ZN(G397));
  NOR2_X1   g575(.A1(new_n800), .A2(G2067), .ZN(new_n1001));
  INV_X1    g576(.A(G1384), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n886), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT45), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g580(.A(KEYINPUT104), .B(G40), .ZN(new_n1006));
  AND3_X1   g581(.A1(new_n468), .A2(new_n472), .A3(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n1005), .A2(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g584(.A(new_n800), .B(G2067), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  XNOR2_X1  g586(.A(new_n1011), .B(KEYINPUT105), .ZN(new_n1012));
  XNOR2_X1  g587(.A(new_n893), .B(G1996), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1012), .B1(new_n1009), .B2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n722), .A2(new_n725), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1001), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1005), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(new_n1007), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1018), .A2(G1996), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT126), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(KEYINPUT46), .ZN(new_n1022));
  XNOR2_X1  g597(.A(new_n1020), .B(new_n1022), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1009), .B1(new_n893), .B2(new_n1010), .ZN(new_n1024));
  OAI211_X1 g599(.A(new_n1023), .B(new_n1024), .C1(new_n1021), .C2(KEYINPUT46), .ZN(new_n1025));
  XOR2_X1   g600(.A(new_n1025), .B(KEYINPUT47), .Z(new_n1026));
  NOR2_X1   g601(.A1(new_n723), .A2(new_n726), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1009), .B1(new_n1027), .B2(new_n1015), .ZN(new_n1028));
  AND2_X1   g603(.A1(new_n1014), .A2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1009), .A2(new_n728), .A3(new_n731), .ZN(new_n1030));
  XNOR2_X1  g605(.A(new_n1030), .B(KEYINPUT48), .ZN(new_n1031));
  AOI211_X1 g606(.A(new_n1019), .B(new_n1026), .C1(new_n1029), .C2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT63), .ZN(new_n1033));
  INV_X1    g608(.A(G1981), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n593), .A2(new_n1034), .A3(new_n594), .A4(new_n596), .ZN(new_n1035));
  XNOR2_X1  g610(.A(KEYINPUT108), .B(G86), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n507), .A2(new_n1036), .ZN(new_n1037));
  AOI211_X1 g612(.A(new_n595), .B(new_n1037), .C1(G651), .C2(new_n592), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1035), .B1(new_n1038), .B2(new_n1034), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT49), .ZN(new_n1040));
  OR2_X1    g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n886), .A2(new_n1007), .A3(new_n1002), .ZN(new_n1042));
  XNOR2_X1  g617(.A(KEYINPUT106), .B(G8), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1044), .ZN(new_n1045));
  AND3_X1   g620(.A1(new_n1039), .A2(KEYINPUT109), .A3(new_n1040), .ZN(new_n1046));
  AOI21_X1  g621(.A(KEYINPUT109), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1047));
  OAI211_X1 g622(.A(new_n1041), .B(new_n1045), .C1(new_n1046), .C2(new_n1047), .ZN(new_n1048));
  NOR4_X1   g623(.A1(new_n579), .A2(new_n580), .A3(new_n744), .A4(new_n583), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT107), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT52), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1045), .A2(new_n1050), .A3(new_n1053), .ZN(new_n1054));
  OAI22_X1  g629(.A1(new_n1044), .A2(new_n1049), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1055));
  NAND3_X1  g630(.A1(G288), .A2(new_n1052), .A3(new_n744), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1054), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  AND2_X1   g632(.A1(new_n1048), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(G303), .A2(G8), .ZN(new_n1059));
  XOR2_X1   g634(.A(new_n1059), .B(KEYINPUT55), .Z(new_n1060));
  AOI21_X1  g635(.A(G1384), .B1(new_n890), .B2(new_n498), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(KEYINPUT45), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n494), .A2(new_n499), .A3(new_n1002), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(new_n1004), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1062), .A2(new_n1007), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(G1971), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT50), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1061), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1063), .A2(KEYINPUT50), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1070), .A2(new_n1007), .A3(new_n1071), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n1072), .A2(G2090), .ZN(new_n1073));
  OAI211_X1 g648(.A(G8), .B(new_n1060), .C1(new_n1068), .C2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1043), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT112), .ZN(new_n1076));
  OAI211_X1 g651(.A(new_n1076), .B(new_n1007), .C1(new_n1061), .C2(new_n1069), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1007), .A2(new_n1069), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1042), .A2(KEYINPUT112), .A3(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(G2090), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n494), .A2(new_n499), .A3(new_n1069), .A4(new_n1002), .ZN(new_n1082));
  XNOR2_X1  g657(.A(new_n1082), .B(KEYINPUT113), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1080), .A2(new_n1081), .A3(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1075), .B1(new_n1084), .B2(new_n1067), .ZN(new_n1085));
  OAI211_X1 g660(.A(new_n1058), .B(new_n1074), .C1(new_n1060), .C2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(G1966), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1007), .B1(new_n1063), .B2(new_n1004), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1087), .B1(new_n1017), .B2(new_n1088), .ZN(new_n1089));
  XNOR2_X1  g664(.A(KEYINPUT114), .B(G2084), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1070), .A2(new_n1007), .A3(new_n1071), .A4(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1075), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(G168), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1033), .B1(new_n1086), .B2(new_n1093), .ZN(new_n1094));
  AND2_X1   g669(.A1(new_n1058), .A2(new_n1074), .ZN(new_n1095));
  OAI21_X1  g670(.A(G8), .B1(new_n1068), .B2(new_n1073), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1060), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1033), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1095), .A2(new_n1098), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1094), .B1(new_n1093), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1074), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(new_n1058), .ZN(new_n1102));
  NOR2_X1   g677(.A1(G288), .A2(G1976), .ZN(new_n1103));
  XNOR2_X1  g678(.A(new_n1103), .B(KEYINPUT111), .ZN(new_n1104));
  AND2_X1   g679(.A1(new_n1104), .A2(new_n1048), .ZN(new_n1105));
  XNOR2_X1  g680(.A(new_n1035), .B(KEYINPUT110), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1045), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1017), .A2(new_n1088), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT53), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1109), .A2(G2078), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1111));
  XNOR2_X1  g686(.A(KEYINPUT123), .B(KEYINPUT53), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1112), .B1(new_n1065), .B2(G2078), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1072), .A2(new_n777), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1111), .A2(new_n1113), .A3(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(G171), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT122), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1117), .B1(G168), .B2(new_n1075), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n535), .A2(new_n541), .A3(KEYINPUT122), .A4(new_n1043), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1118), .A2(G8), .A3(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1089), .A2(new_n1118), .A3(new_n1091), .A4(new_n1119), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1122), .A2(KEYINPUT51), .A3(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT51), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1118), .A2(new_n1125), .A3(new_n1119), .ZN(new_n1126));
  OR2_X1    g701(.A1(new_n1092), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1124), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT62), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1116), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  OR2_X1    g705(.A1(new_n1085), .A2(new_n1060), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1124), .A2(new_n1127), .A3(KEYINPUT62), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1130), .A2(new_n1131), .A3(new_n1095), .A4(new_n1132), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1100), .A2(new_n1102), .A3(new_n1107), .A4(new_n1133), .ZN(new_n1134));
  XOR2_X1   g709(.A(KEYINPUT56), .B(G2072), .Z(new_n1135));
  OR2_X1    g710(.A1(new_n1065), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT115), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1080), .A2(new_n1083), .ZN(new_n1138));
  INV_X1    g713(.A(G1956), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1137), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  AOI211_X1 g715(.A(KEYINPUT115), .B(G1956), .C1(new_n1080), .C2(new_n1083), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1136), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT57), .ZN(new_n1143));
  OAI21_X1  g718(.A(G299), .B1(KEYINPUT116), .B2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(KEYINPUT116), .ZN(new_n1145));
  XOR2_X1   g720(.A(new_n1145), .B(KEYINPUT117), .Z(new_n1146));
  XOR2_X1   g721(.A(new_n1144), .B(new_n1146), .Z(new_n1147));
  INV_X1    g722(.A(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1142), .A2(new_n1148), .ZN(new_n1149));
  OAI211_X1 g724(.A(new_n1147), .B(new_n1136), .C1(new_n1140), .C2(new_n1141), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1149), .A2(KEYINPUT61), .A3(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1151), .A2(KEYINPUT120), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT61), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1042), .A2(G2067), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1156), .B1(new_n1072), .B2(new_n660), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n1157), .A2(KEYINPUT60), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT60), .ZN(new_n1159));
  AOI211_X1 g734(.A(new_n1159), .B(new_n1156), .C1(new_n1072), .C2(new_n660), .ZN(new_n1160));
  INV_X1    g735(.A(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT121), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n611), .B1(new_n1160), .B2(KEYINPUT121), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1158), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1161), .A2(new_n1162), .A3(new_n611), .ZN(new_n1166));
  XOR2_X1   g741(.A(KEYINPUT58), .B(G1341), .Z(new_n1167));
  NAND2_X1  g742(.A1(new_n1042), .A2(new_n1167), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1168), .B1(new_n1065), .B2(G1996), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1169), .A2(KEYINPUT119), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT119), .ZN(new_n1171));
  OAI211_X1 g746(.A(new_n1171), .B(new_n1168), .C1(new_n1065), .C2(G1996), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1170), .A2(new_n556), .A3(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1173), .A2(KEYINPUT59), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT59), .ZN(new_n1175));
  NAND4_X1  g750(.A1(new_n1170), .A2(new_n1175), .A3(new_n556), .A4(new_n1172), .ZN(new_n1176));
  AOI22_X1  g751(.A1(new_n1165), .A2(new_n1166), .B1(new_n1174), .B2(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT120), .ZN(new_n1178));
  NAND4_X1  g753(.A1(new_n1149), .A2(new_n1178), .A3(KEYINPUT61), .A4(new_n1150), .ZN(new_n1179));
  NAND4_X1  g754(.A1(new_n1152), .A2(new_n1155), .A3(new_n1177), .A4(new_n1179), .ZN(new_n1180));
  OAI21_X1  g755(.A(KEYINPUT118), .B1(new_n1157), .B2(new_n611), .ZN(new_n1181));
  OR3_X1    g756(.A1(new_n1157), .A2(KEYINPUT118), .A3(new_n611), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1149), .A2(new_n1181), .A3(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1183), .A2(new_n1150), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1180), .A2(new_n1184), .ZN(new_n1185));
  NOR2_X1   g760(.A1(new_n1115), .A2(G171), .ZN(new_n1186));
  INV_X1    g761(.A(KEYINPUT54), .ZN(new_n1187));
  NOR2_X1   g762(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  AND2_X1   g763(.A1(new_n1005), .A2(G40), .ZN(new_n1189));
  NAND4_X1  g764(.A1(new_n1189), .A2(G160), .A3(new_n1062), .A4(new_n1110), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1190), .A2(new_n1113), .A3(new_n1114), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1191), .A2(KEYINPUT124), .ZN(new_n1192));
  INV_X1    g767(.A(KEYINPUT124), .ZN(new_n1193));
  NAND4_X1  g768(.A1(new_n1190), .A2(new_n1113), .A3(new_n1193), .A4(new_n1114), .ZN(new_n1194));
  NAND3_X1  g769(.A1(new_n1192), .A2(G171), .A3(new_n1194), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1128), .B1(new_n1188), .B2(new_n1195), .ZN(new_n1196));
  NAND4_X1  g771(.A1(new_n1190), .A2(new_n1113), .A3(G301), .A4(new_n1114), .ZN(new_n1197));
  AOI21_X1  g772(.A(KEYINPUT54), .B1(new_n1116), .B2(new_n1197), .ZN(new_n1198));
  NOR2_X1   g773(.A1(new_n1086), .A2(new_n1198), .ZN(new_n1199));
  INV_X1    g774(.A(KEYINPUT125), .ZN(new_n1200));
  AND3_X1   g775(.A1(new_n1196), .A2(new_n1199), .A3(new_n1200), .ZN(new_n1201));
  AOI21_X1  g776(.A(new_n1200), .B1(new_n1196), .B2(new_n1199), .ZN(new_n1202));
  NOR2_X1   g777(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  AOI21_X1  g778(.A(new_n1134), .B1(new_n1185), .B2(new_n1203), .ZN(new_n1204));
  XNOR2_X1  g779(.A(new_n731), .B(G1986), .ZN(new_n1205));
  OAI21_X1  g780(.A(new_n1029), .B1(new_n1018), .B2(new_n1205), .ZN(new_n1206));
  OAI21_X1  g781(.A(new_n1032), .B1(new_n1204), .B2(new_n1206), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g782(.A1(G227), .A2(new_n459), .ZN(new_n1209));
  AOI21_X1  g783(.A(G229), .B1(new_n677), .B2(new_n678), .ZN(new_n1210));
  AND2_X1   g784(.A1(new_n1210), .A2(new_n929), .ZN(new_n1211));
  AND4_X1   g785(.A1(KEYINPUT127), .A2(new_n998), .A3(new_n1209), .A4(new_n1211), .ZN(new_n1212));
  INV_X1    g786(.A(new_n1209), .ZN(new_n1213));
  AOI21_X1  g787(.A(new_n1213), .B1(new_n995), .B2(new_n997), .ZN(new_n1214));
  AOI21_X1  g788(.A(KEYINPUT127), .B1(new_n1214), .B2(new_n1211), .ZN(new_n1215));
  NOR2_X1   g789(.A1(new_n1212), .A2(new_n1215), .ZN(G308));
  INV_X1    g790(.A(KEYINPUT127), .ZN(new_n1217));
  AND3_X1   g791(.A1(new_n979), .A2(new_n996), .A3(new_n985), .ZN(new_n1218));
  AOI21_X1  g792(.A(new_n996), .B1(new_n979), .B2(new_n987), .ZN(new_n1219));
  OAI21_X1  g793(.A(new_n1209), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  INV_X1    g794(.A(new_n1211), .ZN(new_n1221));
  OAI21_X1  g795(.A(new_n1217), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1222));
  NAND3_X1  g796(.A1(new_n1214), .A2(KEYINPUT127), .A3(new_n1211), .ZN(new_n1223));
  NAND2_X1  g797(.A1(new_n1222), .A2(new_n1223), .ZN(G225));
endmodule


