//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 0 0 1 1 0 0 1 1 0 0 1 1 0 0 1 0 0 0 1 0 1 0 1 1 1 1 1 1 0 1 1 0 0 0 1 1 0 0 0 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n744, new_n745, new_n746, new_n748, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n778, new_n779, new_n780, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n839, new_n841, new_n842,
    new_n844, new_n845, new_n846, new_n847, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n931, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n946, new_n948,
    new_n949, new_n950, new_n951, new_n953, new_n954, new_n955, new_n956,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n986, new_n987;
  INV_X1    g000(.A(KEYINPUT22), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT72), .B(G218gat), .ZN(new_n203));
  INV_X1    g002(.A(G211gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n202), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  XOR2_X1   g004(.A(G197gat), .B(G204gat), .Z(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  XOR2_X1   g007(.A(G211gat), .B(G218gat), .Z(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(new_n209), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n205), .A2(new_n211), .A3(new_n207), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(G183gat), .A2(G190gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT24), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND3_X1  g015(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n217));
  OAI211_X1 g016(.A(new_n216), .B(new_n217), .C1(G183gat), .C2(G190gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(G169gat), .A2(G176gat), .ZN(new_n219));
  XNOR2_X1  g018(.A(new_n219), .B(KEYINPUT64), .ZN(new_n220));
  NOR2_X1   g019(.A1(G169gat), .A2(G176gat), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT23), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g022(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n218), .A2(new_n220), .A3(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT25), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  XNOR2_X1  g027(.A(KEYINPUT65), .B(G190gat), .ZN(new_n229));
  OAI211_X1 g028(.A(new_n216), .B(new_n217), .C1(new_n229), .C2(G183gat), .ZN(new_n230));
  OR2_X1    g029(.A1(new_n219), .A2(KEYINPUT64), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n219), .A2(KEYINPUT64), .ZN(new_n232));
  AOI22_X1  g031(.A1(new_n231), .A2(new_n232), .B1(new_n223), .B2(new_n224), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n230), .A2(new_n233), .A3(KEYINPUT25), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n228), .A2(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(KEYINPUT27), .B(G183gat), .ZN(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  OAI21_X1  g036(.A(KEYINPUT28), .B1(new_n237), .B2(new_n229), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n221), .B(KEYINPUT26), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(new_n220), .ZN(new_n240));
  XOR2_X1   g039(.A(KEYINPUT65), .B(G190gat), .Z(new_n241));
  INV_X1    g040(.A(KEYINPUT28), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n241), .A2(new_n242), .A3(new_n236), .ZN(new_n243));
  NAND4_X1  g042(.A1(new_n238), .A2(new_n240), .A3(new_n214), .A4(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(G226gat), .ZN(new_n245));
  INV_X1    g044(.A(G233gat), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n235), .A2(new_n244), .A3(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT29), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n250), .B1(new_n245), .B2(new_n246), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n251), .B1(new_n235), .B2(new_n244), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n213), .B1(new_n249), .B2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n252), .ZN(new_n254));
  INV_X1    g053(.A(new_n213), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n254), .A2(new_n255), .A3(new_n248), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n253), .A2(new_n256), .A3(KEYINPUT73), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT73), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n254), .A2(new_n258), .A3(new_n255), .A4(new_n248), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n257), .A2(KEYINPUT37), .A3(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(G8gat), .B(G36gat), .ZN(new_n261));
  XNOR2_X1  g060(.A(G64gat), .B(G92gat), .ZN(new_n262));
  XNOR2_X1  g061(.A(new_n261), .B(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n260), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT87), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n260), .A2(KEYINPUT87), .A3(new_n263), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n257), .A2(new_n259), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT37), .ZN(new_n269));
  AOI21_X1  g068(.A(KEYINPUT86), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT86), .ZN(new_n271));
  AOI211_X1 g070(.A(new_n271), .B(KEYINPUT37), .C1(new_n257), .C2(new_n259), .ZN(new_n272));
  OAI211_X1 g071(.A(new_n266), .B(new_n267), .C1(new_n270), .C2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(KEYINPUT38), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT88), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(G1gat), .B(G29gat), .ZN(new_n277));
  INV_X1    g076(.A(G85gat), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n277), .B(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(KEYINPUT0), .B(G57gat), .ZN(new_n280));
  XOR2_X1   g079(.A(new_n279), .B(new_n280), .Z(new_n281));
  XNOR2_X1  g080(.A(G127gat), .B(G134gat), .ZN(new_n282));
  INV_X1    g081(.A(G120gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(G113gat), .ZN(new_n284));
  INV_X1    g083(.A(G113gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(G120gat), .ZN(new_n286));
  AOI21_X1  g085(.A(KEYINPUT1), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT66), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  AOI211_X1 g088(.A(KEYINPUT66), .B(KEYINPUT1), .C1(new_n284), .C2(new_n286), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n282), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(G141gat), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n292), .A2(G148gat), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(KEYINPUT75), .B(G141gat), .ZN(new_n295));
  INV_X1    g094(.A(G148gat), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n294), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(G155gat), .A2(G162gat), .ZN(new_n298));
  INV_X1    g097(.A(G155gat), .ZN(new_n299));
  INV_X1    g098(.A(G162gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n298), .B1(new_n301), .B2(KEYINPUT2), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT2), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n296), .A2(G141gat), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n303), .B1(new_n293), .B2(new_n304), .ZN(new_n305));
  AND2_X1   g104(.A1(new_n301), .A2(new_n298), .ZN(new_n306));
  AOI22_X1  g105(.A1(new_n297), .A2(new_n302), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n287), .A2(new_n288), .ZN(new_n308));
  INV_X1    g107(.A(new_n282), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n291), .A2(new_n307), .A3(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n297), .A2(new_n302), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n305), .A2(new_n306), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(KEYINPUT3), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n291), .A2(new_n310), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT3), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n307), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n316), .A2(new_n317), .A3(new_n319), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n312), .B1(new_n320), .B2(KEYINPUT4), .ZN(new_n321));
  XNOR2_X1  g120(.A(G113gat), .B(G120gat), .ZN(new_n322));
  OAI21_X1  g121(.A(KEYINPUT66), .B1(new_n322), .B2(KEYINPUT1), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n309), .B1(new_n308), .B2(new_n323), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n290), .A2(new_n282), .ZN(new_n325));
  OAI21_X1  g124(.A(KEYINPUT67), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT67), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n291), .A2(new_n327), .A3(new_n310), .ZN(new_n328));
  NAND4_X1  g127(.A1(new_n326), .A2(new_n328), .A3(KEYINPUT4), .A4(new_n307), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(G225gat), .A2(G233gat), .ZN(new_n331));
  XOR2_X1   g130(.A(new_n331), .B(KEYINPUT76), .Z(new_n332));
  NOR3_X1   g131(.A1(new_n321), .A2(new_n330), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n315), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(new_n311), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(new_n332), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(KEYINPUT5), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n333), .A2(new_n337), .ZN(new_n338));
  AND2_X1   g137(.A1(new_n316), .A2(new_n317), .ZN(new_n339));
  AOI22_X1  g138(.A1(new_n339), .A2(new_n319), .B1(new_n312), .B2(KEYINPUT4), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT5), .ZN(new_n341));
  INV_X1    g140(.A(new_n332), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n326), .A2(new_n328), .A3(new_n307), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT4), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n340), .A2(new_n341), .A3(new_n342), .A4(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n281), .B1(new_n338), .B2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT6), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n253), .A2(new_n256), .A3(KEYINPUT85), .ZN(new_n352));
  OAI211_X1 g151(.A(new_n352), .B(KEYINPUT37), .C1(KEYINPUT85), .C2(new_n253), .ZN(new_n353));
  XOR2_X1   g152(.A(new_n263), .B(KEYINPUT74), .Z(new_n354));
  NOR2_X1   g153(.A1(new_n354), .A2(KEYINPUT38), .ZN(new_n355));
  OAI211_X1 g154(.A(new_n353), .B(new_n355), .C1(new_n270), .C2(new_n272), .ZN(new_n356));
  AND2_X1   g155(.A1(new_n320), .A2(KEYINPUT4), .ZN(new_n357));
  OAI211_X1 g156(.A(new_n329), .B(new_n342), .C1(new_n357), .C2(new_n312), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n358), .A2(KEYINPUT5), .A3(new_n336), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT77), .ZN(new_n360));
  INV_X1    g159(.A(new_n281), .ZN(new_n361));
  NAND4_X1  g160(.A1(new_n359), .A2(new_n360), .A3(new_n346), .A4(new_n361), .ZN(new_n362));
  OAI211_X1 g161(.A(new_n346), .B(new_n361), .C1(new_n333), .C2(new_n337), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(KEYINPUT77), .ZN(new_n364));
  NAND4_X1  g163(.A1(new_n362), .A2(new_n364), .A3(new_n348), .A4(new_n349), .ZN(new_n365));
  INV_X1    g164(.A(new_n263), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n268), .A2(new_n366), .ZN(new_n367));
  AND4_X1   g166(.A1(new_n351), .A2(new_n356), .A3(new_n365), .A4(new_n367), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n273), .A2(KEYINPUT88), .A3(KEYINPUT38), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n276), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  AOI21_X1  g169(.A(KEYINPUT29), .B1(new_n210), .B2(new_n212), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n315), .B1(new_n371), .B2(KEYINPUT3), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(KEYINPUT83), .ZN(new_n373));
  INV_X1    g172(.A(G228gat), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n374), .A2(new_n246), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n213), .B1(new_n250), .B2(new_n319), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT83), .ZN(new_n378));
  OAI211_X1 g177(.A(new_n378), .B(new_n315), .C1(new_n371), .C2(KEYINPUT3), .ZN(new_n379));
  NAND4_X1  g178(.A1(new_n373), .A2(new_n375), .A3(new_n377), .A4(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT82), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n210), .A2(new_n381), .A3(new_n212), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n211), .B1(new_n205), .B2(new_n207), .ZN(new_n383));
  AOI21_X1  g182(.A(KEYINPUT29), .B1(new_n383), .B2(KEYINPUT82), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n307), .B1(new_n385), .B2(new_n318), .ZN(new_n386));
  OAI22_X1  g185(.A1(new_n386), .A2(new_n376), .B1(new_n374), .B2(new_n246), .ZN(new_n387));
  INV_X1    g186(.A(G22gat), .ZN(new_n388));
  AND3_X1   g187(.A1(new_n380), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n388), .B1(new_n380), .B2(new_n387), .ZN(new_n390));
  OAI21_X1  g189(.A(KEYINPUT81), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  XNOR2_X1  g190(.A(KEYINPUT79), .B(KEYINPUT31), .ZN(new_n392));
  XNOR2_X1  g191(.A(G50gat), .B(G78gat), .ZN(new_n393));
  XOR2_X1   g192(.A(new_n392), .B(new_n393), .Z(new_n394));
  NAND2_X1  g193(.A1(new_n391), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n394), .ZN(new_n396));
  OAI211_X1 g195(.A(KEYINPUT81), .B(new_n396), .C1(new_n389), .C2(new_n390), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  XNOR2_X1  g197(.A(KEYINPUT80), .B(G106gat), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n395), .A2(new_n397), .A3(new_n399), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT39), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n335), .A2(new_n332), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n403), .B1(new_n404), .B2(KEYINPUT84), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n342), .B1(new_n340), .B2(new_n345), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT84), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n405), .B1(new_n408), .B2(new_n404), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n281), .B1(new_n406), .B2(new_n403), .ZN(new_n410));
  AND3_X1   g209(.A1(new_n409), .A2(KEYINPUT40), .A3(new_n410), .ZN(new_n411));
  AOI21_X1  g210(.A(KEYINPUT40), .B1(new_n409), .B2(new_n410), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  OR2_X1    g212(.A1(new_n367), .A2(KEYINPUT30), .ZN(new_n414));
  OAI211_X1 g213(.A(new_n367), .B(KEYINPUT30), .C1(new_n268), .C2(new_n354), .ZN(new_n415));
  AND3_X1   g214(.A1(new_n414), .A2(new_n415), .A3(new_n348), .ZN(new_n416));
  AOI22_X1  g215(.A1(new_n401), .A2(new_n402), .B1(new_n413), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n370), .A2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT71), .ZN(new_n419));
  XNOR2_X1  g218(.A(KEYINPUT68), .B(G15gat), .ZN(new_n420));
  INV_X1    g219(.A(G43gat), .ZN(new_n421));
  XNOR2_X1  g220(.A(new_n420), .B(new_n421), .ZN(new_n422));
  XOR2_X1   g221(.A(G71gat), .B(G99gat), .Z(new_n423));
  XNOR2_X1  g222(.A(new_n422), .B(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(G227gat), .A2(G233gat), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n326), .A2(new_n328), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n235), .A2(new_n244), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n326), .A2(new_n328), .A3(new_n235), .A4(new_n244), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n425), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n424), .B1(new_n430), .B2(KEYINPUT33), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT32), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n428), .A2(new_n429), .ZN(new_n435));
  INV_X1    g234(.A(new_n425), .ZN(new_n436));
  AOI221_X4 g235(.A(new_n432), .B1(KEYINPUT33), .B2(new_n424), .C1(new_n435), .C2(new_n436), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n419), .B1(new_n434), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n435), .A2(new_n436), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(KEYINPUT32), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT33), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n440), .A2(new_n442), .A3(new_n424), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n431), .A2(new_n433), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n443), .A2(new_n444), .A3(KEYINPUT71), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n436), .B1(new_n435), .B2(KEYINPUT70), .ZN(new_n446));
  AND2_X1   g245(.A1(KEYINPUT70), .A2(KEYINPUT34), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n446), .B1(new_n435), .B2(new_n447), .ZN(new_n448));
  AND2_X1   g247(.A1(KEYINPUT69), .A2(KEYINPUT34), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n428), .A2(new_n425), .A3(new_n429), .ZN(new_n450));
  NOR2_X1   g249(.A1(KEYINPUT69), .A2(KEYINPUT34), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n449), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n448), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n438), .A2(new_n445), .A3(new_n453), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n434), .A2(new_n437), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n455), .A2(KEYINPUT71), .A3(new_n448), .A4(new_n452), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n454), .A2(new_n456), .A3(KEYINPUT36), .ZN(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(KEYINPUT36), .B1(new_n454), .B2(new_n456), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  AND3_X1   g259(.A1(new_n395), .A2(new_n397), .A3(new_n399), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n399), .B1(new_n395), .B2(new_n397), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n348), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n364), .A2(new_n362), .A3(new_n349), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n464), .B1(new_n465), .B2(KEYINPUT78), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT78), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n364), .A2(new_n362), .A3(new_n467), .A4(new_n349), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n350), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  AND2_X1   g268(.A1(new_n414), .A2(new_n415), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n463), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  AND3_X1   g270(.A1(new_n418), .A2(new_n460), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n466), .A2(new_n468), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(new_n351), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n454), .A2(new_n456), .ZN(new_n475));
  INV_X1    g274(.A(new_n470), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n401), .A2(new_n402), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n474), .A2(new_n475), .A3(new_n476), .A4(new_n477), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n475), .B1(new_n461), .B2(new_n462), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n479), .A2(new_n470), .ZN(new_n480));
  AOI21_X1  g279(.A(KEYINPUT35), .B1(new_n351), .B2(new_n365), .ZN(new_n481));
  AOI22_X1  g280(.A1(new_n478), .A2(KEYINPUT35), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n472), .A2(new_n482), .ZN(new_n483));
  XNOR2_X1  g282(.A(G169gat), .B(G197gat), .ZN(new_n484));
  XNOR2_X1  g283(.A(G113gat), .B(G141gat), .ZN(new_n485));
  XNOR2_X1  g284(.A(new_n484), .B(new_n485), .ZN(new_n486));
  XNOR2_X1  g285(.A(KEYINPUT89), .B(KEYINPUT11), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n486), .B(new_n487), .ZN(new_n488));
  XOR2_X1   g287(.A(new_n488), .B(KEYINPUT12), .Z(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  OAI21_X1  g289(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n491));
  INV_X1    g290(.A(new_n491), .ZN(new_n492));
  NOR3_X1   g291(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n493));
  OAI21_X1  g292(.A(KEYINPUT91), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT14), .ZN(new_n495));
  INV_X1    g294(.A(G29gat), .ZN(new_n496));
  INV_X1    g295(.A(G36gat), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n495), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT91), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n498), .A2(new_n499), .A3(new_n491), .ZN(new_n500));
  NAND2_X1  g299(.A1(G29gat), .A2(G36gat), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n494), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  XNOR2_X1  g301(.A(G43gat), .B(G50gat), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(KEYINPUT15), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(new_n501), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n506), .B1(new_n503), .B2(KEYINPUT15), .ZN(new_n507));
  INV_X1    g306(.A(G50gat), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(G43gat), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n421), .A2(G50gat), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT15), .ZN(new_n512));
  AOI22_X1  g311(.A1(new_n511), .A2(new_n512), .B1(new_n491), .B2(new_n498), .ZN(new_n513));
  AOI22_X1  g312(.A1(new_n502), .A2(new_n505), .B1(new_n507), .B2(new_n513), .ZN(new_n514));
  XNOR2_X1  g313(.A(G15gat), .B(G22gat), .ZN(new_n515));
  INV_X1    g314(.A(G1gat), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(KEYINPUT16), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n518), .B1(G1gat), .B2(new_n515), .ZN(new_n519));
  OR2_X1    g318(.A1(new_n519), .A2(G8gat), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(G8gat), .ZN(new_n521));
  AND3_X1   g320(.A1(new_n514), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n514), .B1(new_n521), .B2(new_n520), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(G229gat), .A2(G233gat), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n525), .B(KEYINPUT13), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(new_n523), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT17), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT92), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n529), .B1(new_n514), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n498), .A2(new_n491), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n506), .B1(new_n532), .B2(KEYINPUT91), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n504), .B1(new_n533), .B2(new_n500), .ZN(new_n534));
  AND2_X1   g333(.A1(new_n513), .A2(new_n507), .ZN(new_n535));
  OAI211_X1 g334(.A(KEYINPUT92), .B(KEYINPUT17), .C1(new_n534), .C2(new_n535), .ZN(new_n536));
  AND2_X1   g335(.A1(new_n531), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n520), .A2(new_n521), .ZN(new_n538));
  OAI211_X1 g337(.A(new_n525), .B(new_n528), .C1(new_n537), .C2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT18), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n527), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n538), .B1(new_n531), .B2(new_n536), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n542), .A2(new_n523), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n543), .A2(KEYINPUT18), .A3(new_n525), .ZN(new_n544));
  AOI211_X1 g343(.A(KEYINPUT90), .B(new_n490), .C1(new_n541), .C2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n539), .A2(new_n540), .ZN(new_n546));
  INV_X1    g345(.A(new_n527), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n546), .A2(new_n544), .A3(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT90), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n489), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n545), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n483), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(G231gat), .A2(G233gat), .ZN(new_n554));
  XOR2_X1   g353(.A(new_n554), .B(G183gat), .Z(new_n555));
  XNOR2_X1  g354(.A(new_n555), .B(new_n204), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  XOR2_X1   g356(.A(G127gat), .B(G155gat), .Z(new_n558));
  INV_X1    g357(.A(new_n538), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT94), .ZN(new_n560));
  INV_X1    g359(.A(G57gat), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(G64gat), .ZN(new_n562));
  INV_X1    g361(.A(G64gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(G57gat), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(G71gat), .A2(G78gat), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT9), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(G71gat), .B(G78gat), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n565), .A2(new_n570), .A3(new_n568), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n572), .A2(KEYINPUT93), .A3(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  AOI21_X1  g374(.A(KEYINPUT93), .B1(new_n572), .B2(new_n573), .ZN(new_n576));
  OAI21_X1  g375(.A(KEYINPUT21), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n559), .A2(new_n560), .A3(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n560), .B1(new_n559), .B2(new_n577), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n558), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n580), .ZN(new_n582));
  INV_X1    g381(.A(new_n558), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n582), .A2(new_n578), .A3(new_n583), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n557), .B1(new_n581), .B2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n575), .A2(new_n576), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT21), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n589), .B(new_n590), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n581), .A2(new_n584), .A3(new_n557), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n586), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n591), .ZN(new_n594));
  INV_X1    g393(.A(new_n592), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n594), .B1(new_n595), .B2(new_n585), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(G190gat), .B(G218gat), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n514), .B1(KEYINPUT96), .B2(KEYINPUT17), .ZN(new_n599));
  XNOR2_X1  g398(.A(G99gat), .B(G106gat), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(G99gat), .A2(G106gat), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n602), .A2(KEYINPUT95), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT95), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n604), .A2(G99gat), .A3(G106gat), .ZN(new_n605));
  AND3_X1   g404(.A1(new_n603), .A2(new_n605), .A3(KEYINPUT8), .ZN(new_n606));
  NAND2_X1  g405(.A1(G85gat), .A2(G92gat), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT7), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  OR2_X1    g408(.A1(G85gat), .A2(G92gat), .ZN(new_n610));
  NAND3_X1  g409(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n601), .B1(new_n606), .B2(new_n612), .ZN(new_n613));
  AND2_X1   g412(.A1(new_n609), .A2(new_n610), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n603), .A2(new_n605), .A3(KEYINPUT8), .ZN(new_n615));
  NAND4_X1  g414(.A1(new_n614), .A2(new_n615), .A3(new_n600), .A4(new_n611), .ZN(new_n616));
  AND2_X1   g415(.A1(new_n613), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n599), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(G232gat), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n619), .A2(new_n246), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n620), .A2(KEYINPUT41), .ZN(new_n621));
  AND2_X1   g420(.A1(new_n618), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n613), .A2(new_n616), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n624), .A2(KEYINPUT96), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n537), .A2(new_n625), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n598), .B1(new_n623), .B2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n598), .ZN(new_n628));
  OAI211_X1 g427(.A(new_n622), .B(new_n628), .C1(new_n537), .C2(new_n625), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT97), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n620), .A2(KEYINPUT41), .ZN(new_n632));
  XNOR2_X1  g431(.A(G134gat), .B(G162gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n630), .A2(new_n631), .A3(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n634), .B(KEYINPUT97), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n627), .A2(new_n629), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(G120gat), .B(G148gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(G176gat), .B(G204gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n639), .B(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(G230gat), .A2(G233gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(KEYINPUT99), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT93), .ZN(new_n644));
  AND3_X1   g443(.A1(new_n565), .A2(new_n570), .A3(new_n568), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n570), .B1(new_n568), .B2(new_n565), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n644), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n624), .A2(new_n647), .A3(new_n574), .ZN(new_n648));
  NAND4_X1  g447(.A1(new_n613), .A2(new_n616), .A3(new_n572), .A4(new_n573), .ZN(new_n649));
  XOR2_X1   g448(.A(KEYINPUT98), .B(KEYINPUT10), .Z(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n648), .A2(new_n649), .A3(new_n651), .ZN(new_n652));
  OAI211_X1 g451(.A(new_n617), .B(KEYINPUT10), .C1(new_n575), .C2(new_n576), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n643), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n643), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n655), .B1(new_n648), .B2(new_n649), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n641), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT100), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n654), .A2(new_n656), .ZN(new_n659));
  INV_X1    g458(.A(new_n641), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n658), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NOR4_X1   g460(.A1(new_n654), .A2(KEYINPUT100), .A3(new_n656), .A4(new_n641), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n657), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n597), .A2(new_n638), .A3(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT101), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND4_X1  g466(.A1(new_n597), .A2(KEYINPUT101), .A3(new_n638), .A4(new_n664), .ZN(new_n668));
  AND2_X1   g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n553), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n670), .A2(new_n474), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(new_n516), .ZN(G1324gat));
  INV_X1    g471(.A(new_n670), .ZN(new_n673));
  XOR2_X1   g472(.A(KEYINPUT16), .B(G8gat), .Z(new_n674));
  NAND3_X1  g473(.A1(new_n673), .A2(new_n470), .A3(new_n674), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n675), .A2(KEYINPUT42), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT42), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n673), .A2(new_n470), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n677), .B1(new_n678), .B2(G8gat), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n676), .B1(new_n675), .B2(new_n679), .ZN(G1325gat));
  INV_X1    g479(.A(G15gat), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT102), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n682), .B1(new_n458), .B2(new_n459), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT36), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n475), .A2(new_n684), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n685), .A2(KEYINPUT102), .A3(new_n457), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  NOR3_X1   g486(.A1(new_n670), .A2(new_n681), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n673), .A2(new_n475), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n688), .B1(new_n681), .B2(new_n689), .ZN(G1326gat));
  NOR2_X1   g489(.A1(new_n670), .A2(new_n477), .ZN(new_n691));
  XOR2_X1   g490(.A(KEYINPUT43), .B(G22gat), .Z(new_n692));
  XNOR2_X1  g491(.A(new_n691), .B(new_n692), .ZN(G1327gat));
  INV_X1    g492(.A(new_n597), .ZN(new_n694));
  INV_X1    g493(.A(new_n638), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n694), .A2(new_n695), .A3(new_n664), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(KEYINPUT103), .ZN(new_n697));
  NAND4_X1  g496(.A1(new_n553), .A2(new_n496), .A3(new_n469), .A4(new_n697), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(KEYINPUT45), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT44), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n638), .A2(new_n700), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n701), .B1(new_n472), .B2(new_n482), .ZN(new_n702));
  NOR3_X1   g501(.A1(new_n552), .A2(new_n597), .A3(new_n663), .ZN(new_n703));
  NOR3_X1   g502(.A1(new_n479), .A2(new_n469), .A3(new_n470), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT35), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n477), .A2(new_n475), .A3(new_n476), .ZN(new_n706));
  INV_X1    g505(.A(new_n481), .ZN(new_n707));
  OAI22_X1  g506(.A1(new_n704), .A2(new_n705), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n418), .A2(new_n687), .A3(new_n471), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n638), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  OAI211_X1 g509(.A(new_n702), .B(new_n703), .C1(new_n710), .C2(KEYINPUT44), .ZN(new_n711));
  OAI21_X1  g510(.A(G29gat), .B1(new_n711), .B2(new_n474), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n699), .A2(new_n712), .ZN(G1328gat));
  OAI21_X1  g512(.A(G36gat), .B1(new_n711), .B2(new_n476), .ZN(new_n714));
  NAND4_X1  g513(.A1(new_n553), .A2(new_n497), .A3(new_n470), .A4(new_n697), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT104), .ZN(new_n716));
  AND3_X1   g515(.A1(new_n715), .A2(new_n716), .A3(KEYINPUT46), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n716), .B1(new_n715), .B2(KEYINPUT46), .ZN(new_n718));
  OAI221_X1 g517(.A(new_n714), .B1(KEYINPUT46), .B2(new_n715), .C1(new_n717), .C2(new_n718), .ZN(G1329gat));
  INV_X1    g518(.A(KEYINPUT105), .ZN(new_n720));
  OAI21_X1  g519(.A(G43gat), .B1(new_n711), .B2(new_n687), .ZN(new_n721));
  NAND4_X1  g520(.A1(new_n553), .A2(new_n421), .A3(new_n475), .A4(new_n697), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n720), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT47), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n723), .B(new_n724), .ZN(G1330gat));
  OAI21_X1  g524(.A(G50gat), .B1(new_n711), .B2(new_n477), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT107), .ZN(new_n727));
  AOI21_X1  g526(.A(KEYINPUT48), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n553), .A2(new_n697), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n463), .A2(new_n508), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(KEYINPUT106), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n726), .B1(new_n729), .B2(new_n731), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n728), .B(new_n732), .ZN(G1331gat));
  NAND4_X1  g532(.A1(new_n552), .A2(new_n597), .A3(new_n638), .A4(new_n663), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n734), .B1(new_n708), .B2(new_n709), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(new_n469), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(G57gat), .ZN(G1332gat));
  INV_X1    g536(.A(new_n735), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n738), .A2(new_n476), .ZN(new_n739));
  NOR2_X1   g538(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n740));
  AND2_X1   g539(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n739), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n742), .B1(new_n739), .B2(new_n740), .ZN(G1333gat));
  NAND4_X1  g542(.A1(new_n735), .A2(G71gat), .A3(new_n686), .A4(new_n683), .ZN(new_n744));
  AND2_X1   g543(.A1(new_n735), .A2(new_n475), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n744), .B1(new_n745), .B2(G71gat), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g546(.A1(new_n735), .A2(new_n463), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g548(.A1(new_n694), .A2(new_n552), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(KEYINPUT108), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n751), .A2(new_n664), .ZN(new_n752));
  OAI211_X1 g551(.A(new_n702), .B(new_n752), .C1(new_n710), .C2(KEYINPUT44), .ZN(new_n753));
  NOR3_X1   g552(.A1(new_n753), .A2(new_n278), .A3(new_n474), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n708), .A2(new_n709), .ZN(new_n755));
  INV_X1    g554(.A(new_n751), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n755), .A2(new_n695), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(KEYINPUT51), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT51), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n710), .A2(new_n759), .A3(new_n756), .ZN(new_n760));
  AND2_X1   g559(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n761), .A2(new_n469), .A3(new_n663), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n754), .B1(new_n762), .B2(new_n278), .ZN(G1336gat));
  NOR3_X1   g562(.A1(new_n476), .A2(new_n664), .A3(G92gat), .ZN(new_n764));
  AOI21_X1  g563(.A(KEYINPUT52), .B1(new_n761), .B2(new_n764), .ZN(new_n765));
  OAI21_X1  g564(.A(KEYINPUT110), .B1(new_n753), .B2(new_n476), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(G92gat), .ZN(new_n767));
  NOR3_X1   g566(.A1(new_n753), .A2(KEYINPUT110), .A3(new_n476), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n765), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n757), .A2(KEYINPUT109), .A3(KEYINPUT51), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT109), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n771), .B1(new_n710), .B2(new_n756), .ZN(new_n772));
  OAI211_X1 g571(.A(new_n770), .B(new_n764), .C1(KEYINPUT51), .C2(new_n772), .ZN(new_n773));
  OAI21_X1  g572(.A(G92gat), .B1(new_n753), .B2(new_n476), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(KEYINPUT52), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n769), .A2(new_n776), .ZN(G1337gat));
  INV_X1    g576(.A(G99gat), .ZN(new_n778));
  NOR3_X1   g577(.A1(new_n753), .A2(new_n778), .A3(new_n687), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n761), .A2(new_n475), .A3(new_n663), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n779), .B1(new_n780), .B2(new_n778), .ZN(G1338gat));
  INV_X1    g580(.A(KEYINPUT111), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n477), .A2(G106gat), .A3(new_n664), .ZN(new_n783));
  OAI211_X1 g582(.A(new_n770), .B(new_n783), .C1(new_n772), .C2(KEYINPUT51), .ZN(new_n784));
  OAI21_X1  g583(.A(G106gat), .B1(new_n753), .B2(new_n477), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n782), .B1(new_n786), .B2(KEYINPUT53), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT53), .ZN(new_n788));
  AOI211_X1 g587(.A(KEYINPUT111), .B(new_n788), .C1(new_n784), .C2(new_n785), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT112), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n755), .A2(new_n695), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(new_n700), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n792), .A2(new_n463), .A3(new_n702), .A4(new_n752), .ZN(new_n793));
  AOI21_X1  g592(.A(KEYINPUT53), .B1(new_n793), .B2(G106gat), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n477), .A2(G106gat), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n758), .A2(new_n663), .A3(new_n760), .A4(new_n795), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n790), .B1(new_n794), .B2(new_n796), .ZN(new_n797));
  AND4_X1   g596(.A1(new_n790), .A2(new_n785), .A3(new_n788), .A4(new_n796), .ZN(new_n798));
  OAI22_X1  g597(.A1(new_n787), .A2(new_n789), .B1(new_n797), .B2(new_n798), .ZN(G1339gat));
  AOI21_X1  g598(.A(KEYINPUT18), .B1(new_n543), .B2(new_n525), .ZN(new_n800));
  INV_X1    g599(.A(new_n525), .ZN(new_n801));
  NOR4_X1   g600(.A1(new_n542), .A2(new_n540), .A3(new_n801), .A4(new_n523), .ZN(new_n802));
  NOR3_X1   g601(.A1(new_n800), .A2(new_n802), .A3(new_n527), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n490), .B1(new_n803), .B2(KEYINPUT90), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n652), .A2(new_n653), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(new_n655), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n652), .A2(new_n643), .A3(new_n653), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n806), .A2(new_n807), .A3(KEYINPUT54), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT54), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n660), .B1(new_n654), .B2(new_n809), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n808), .A2(KEYINPUT55), .A3(new_n810), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n811), .B1(new_n661), .B2(new_n662), .ZN(new_n812));
  INV_X1    g611(.A(new_n812), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n548), .A2(new_n549), .A3(new_n489), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT55), .ZN(new_n815));
  AND3_X1   g614(.A1(new_n652), .A2(new_n643), .A3(new_n653), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n816), .A2(new_n654), .A3(new_n809), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n805), .A2(new_n809), .A3(new_n655), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(new_n641), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n815), .B1(new_n817), .B2(new_n819), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n804), .A2(new_n813), .A3(new_n814), .A4(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n541), .A2(new_n544), .A3(new_n489), .ZN(new_n822));
  INV_X1    g621(.A(new_n488), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n543), .A2(new_n525), .ZN(new_n824));
  AND2_X1   g623(.A1(new_n524), .A2(new_n526), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n823), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  AND3_X1   g625(.A1(new_n663), .A2(new_n822), .A3(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n695), .B1(new_n821), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n820), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n822), .A2(new_n826), .ZN(new_n831));
  NOR3_X1   g630(.A1(new_n830), .A2(new_n638), .A3(new_n831), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n694), .B1(new_n829), .B2(new_n832), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n552), .A2(new_n597), .A3(new_n638), .A4(new_n664), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n474), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(new_n480), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n836), .A2(new_n552), .ZN(new_n837));
  XNOR2_X1  g636(.A(new_n837), .B(new_n285), .ZN(G1340gat));
  NOR2_X1   g637(.A1(new_n836), .A2(new_n664), .ZN(new_n839));
  XNOR2_X1  g638(.A(new_n839), .B(new_n283), .ZN(G1341gat));
  INV_X1    g639(.A(new_n836), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(new_n597), .ZN(new_n842));
  XNOR2_X1  g641(.A(new_n842), .B(G127gat), .ZN(G1342gat));
  NAND2_X1  g642(.A1(new_n841), .A2(new_n695), .ZN(new_n844));
  OR3_X1    g643(.A1(new_n844), .A2(KEYINPUT56), .A3(G134gat), .ZN(new_n845));
  OAI21_X1  g644(.A(KEYINPUT56), .B1(new_n844), .B2(G134gat), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n844), .A2(G134gat), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n845), .A2(new_n846), .A3(new_n847), .ZN(G1343gat));
  AOI21_X1  g647(.A(new_n477), .B1(new_n683), .B2(new_n686), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT116), .ZN(new_n850));
  OR2_X1    g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n470), .B1(new_n849), .B2(new_n850), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n851), .A2(new_n835), .A3(new_n852), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n853), .A2(G141gat), .A3(new_n552), .ZN(new_n854));
  INV_X1    g653(.A(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT58), .ZN(new_n856));
  AOI211_X1 g655(.A(new_n350), .B(new_n470), .C1(new_n466), .C2(new_n468), .ZN(new_n857));
  NOR3_X1   g656(.A1(new_n458), .A2(new_n459), .A3(new_n682), .ZN(new_n858));
  AOI21_X1  g657(.A(KEYINPUT102), .B1(new_n685), .B2(new_n457), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n857), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT57), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n477), .B1(new_n833), .B2(new_n834), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n860), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(new_n832), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT113), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n820), .A2(new_n865), .ZN(new_n866));
  OAI211_X1 g665(.A(KEYINPUT113), .B(new_n815), .C1(new_n817), .C2(new_n819), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n868), .A2(new_n804), .A3(new_n814), .A4(new_n813), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n695), .B1(new_n869), .B2(new_n828), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT114), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n864), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n812), .B1(new_n866), .B2(new_n867), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n827), .B1(new_n551), .B2(new_n873), .ZN(new_n874));
  NOR3_X1   g673(.A1(new_n874), .A2(KEYINPUT114), .A3(new_n695), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n694), .B1(new_n872), .B2(new_n875), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n477), .B1(new_n876), .B2(new_n834), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n863), .B1(new_n877), .B2(new_n861), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n295), .B1(new_n878), .B2(new_n552), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n855), .A2(new_n856), .A3(new_n879), .ZN(new_n880));
  INV_X1    g679(.A(new_n834), .ZN(new_n881));
  OAI21_X1  g680(.A(KEYINPUT114), .B1(new_n874), .B2(new_n695), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n869), .A2(new_n828), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n883), .A2(new_n871), .A3(new_n638), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n882), .A2(new_n884), .A3(new_n864), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n881), .B1(new_n885), .B2(new_n694), .ZN(new_n886));
  OAI21_X1  g685(.A(KEYINPUT57), .B1(new_n886), .B2(new_n477), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT115), .ZN(new_n888));
  AND3_X1   g687(.A1(new_n887), .A2(new_n888), .A3(new_n863), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n888), .B1(new_n887), .B2(new_n863), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n551), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n854), .B1(new_n891), .B2(new_n295), .ZN(new_n892));
  NOR3_X1   g691(.A1(new_n892), .A2(KEYINPUT117), .A3(new_n856), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT117), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n878), .A2(KEYINPUT115), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n887), .A2(new_n888), .A3(new_n863), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n552), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(new_n295), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n855), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n894), .B1(new_n899), .B2(KEYINPUT58), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n880), .B1(new_n893), .B2(new_n900), .ZN(G1344gat));
  INV_X1    g700(.A(KEYINPUT121), .ZN(new_n902));
  NOR3_X1   g701(.A1(new_n870), .A2(new_n902), .A3(new_n832), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n883), .A2(new_n638), .ZN(new_n904));
  AOI21_X1  g703(.A(KEYINPUT121), .B1(new_n904), .B2(new_n864), .ZN(new_n905));
  NOR3_X1   g704(.A1(new_n903), .A2(new_n597), .A3(new_n905), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n667), .A2(new_n552), .A3(new_n668), .ZN(new_n907));
  XNOR2_X1  g706(.A(new_n907), .B(KEYINPUT120), .ZN(new_n908));
  OAI211_X1 g707(.A(new_n861), .B(new_n463), .C1(new_n906), .C2(new_n908), .ZN(new_n909));
  INV_X1    g708(.A(new_n862), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(KEYINPUT57), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n860), .A2(new_n664), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n909), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT122), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(G148gat), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n913), .A2(new_n914), .ZN(new_n917));
  OAI21_X1  g716(.A(KEYINPUT59), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n664), .B1(new_n895), .B2(new_n896), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n296), .A2(KEYINPUT59), .ZN(new_n920));
  INV_X1    g719(.A(new_n920), .ZN(new_n921));
  OR3_X1    g720(.A1(new_n919), .A2(KEYINPUT119), .A3(new_n921), .ZN(new_n922));
  OAI21_X1  g721(.A(KEYINPUT119), .B1(new_n919), .B2(new_n921), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n918), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  NOR3_X1   g723(.A1(new_n853), .A2(G148gat), .A3(new_n664), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n925), .B(KEYINPUT118), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n924), .A2(new_n926), .ZN(G1345gat));
  INV_X1    g726(.A(new_n853), .ZN(new_n928));
  AOI21_X1  g727(.A(G155gat), .B1(new_n928), .B2(new_n597), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n895), .A2(new_n896), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n694), .A2(new_n299), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n929), .B1(new_n930), .B2(new_n931), .ZN(G1346gat));
  NAND2_X1  g731(.A1(new_n930), .A2(new_n695), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n933), .A2(G162gat), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT123), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n928), .A2(new_n300), .A3(new_n695), .ZN(new_n936));
  AND3_X1   g735(.A1(new_n934), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n935), .B1(new_n934), .B2(new_n936), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n937), .A2(new_n938), .ZN(G1347gat));
  NAND2_X1  g738(.A1(new_n833), .A2(new_n834), .ZN(new_n940));
  NOR3_X1   g739(.A1(new_n479), .A2(new_n469), .A3(new_n476), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g741(.A(new_n942), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n943), .A2(new_n551), .ZN(new_n944));
  XNOR2_X1  g743(.A(new_n944), .B(G169gat), .ZN(G1348gat));
  NAND2_X1  g744(.A1(new_n943), .A2(new_n663), .ZN(new_n946));
  XNOR2_X1  g745(.A(new_n946), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g746(.A1(new_n943), .A2(new_n597), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n948), .A2(new_n237), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n949), .B1(G183gat), .B2(new_n948), .ZN(new_n950));
  NAND2_X1  g749(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n951));
  XNOR2_X1  g750(.A(new_n950), .B(new_n951), .ZN(G1350gat));
  OAI21_X1  g751(.A(G190gat), .B1(new_n942), .B2(new_n638), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n953), .A2(KEYINPUT61), .ZN(new_n954));
  AND2_X1   g753(.A1(new_n953), .A2(KEYINPUT61), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n943), .A2(new_n241), .A3(new_n695), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n954), .B1(new_n955), .B2(new_n956), .ZN(G1351gat));
  NAND3_X1  g756(.A1(new_n687), .A2(new_n474), .A3(new_n470), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n910), .A2(new_n958), .ZN(new_n959));
  INV_X1    g758(.A(G197gat), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n959), .A2(new_n960), .A3(new_n551), .ZN(new_n961));
  XNOR2_X1  g760(.A(new_n958), .B(KEYINPUT125), .ZN(new_n962));
  AND3_X1   g761(.A1(new_n909), .A2(new_n962), .A3(new_n911), .ZN(new_n963));
  AND2_X1   g762(.A1(new_n963), .A2(new_n551), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n961), .B1(new_n964), .B2(new_n960), .ZN(G1352gat));
  INV_X1    g764(.A(G204gat), .ZN(new_n966));
  AOI21_X1  g765(.A(new_n966), .B1(new_n963), .B2(new_n663), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT62), .ZN(new_n968));
  NOR2_X1   g767(.A1(new_n664), .A2(G204gat), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n959), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  OR2_X1    g769(.A1(new_n970), .A2(KEYINPUT126), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n959), .A2(new_n969), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n972), .A2(KEYINPUT62), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n970), .A2(KEYINPUT126), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n971), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  INV_X1    g774(.A(KEYINPUT127), .ZN(new_n976));
  OR3_X1    g775(.A1(new_n967), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  OAI21_X1  g776(.A(new_n976), .B1(new_n967), .B2(new_n975), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n977), .A2(new_n978), .ZN(G1353gat));
  NAND3_X1  g778(.A1(new_n959), .A2(new_n204), .A3(new_n597), .ZN(new_n980));
  NOR2_X1   g779(.A1(new_n958), .A2(new_n694), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n909), .A2(new_n911), .A3(new_n981), .ZN(new_n982));
  AND3_X1   g781(.A1(new_n982), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n983));
  AOI21_X1  g782(.A(KEYINPUT63), .B1(new_n982), .B2(G211gat), .ZN(new_n984));
  OAI21_X1  g783(.A(new_n980), .B1(new_n983), .B2(new_n984), .ZN(G1354gat));
  AOI21_X1  g784(.A(G218gat), .B1(new_n959), .B2(new_n695), .ZN(new_n986));
  NOR2_X1   g785(.A1(new_n638), .A2(new_n203), .ZN(new_n987));
  AOI21_X1  g786(.A(new_n986), .B1(new_n963), .B2(new_n987), .ZN(G1355gat));
endmodule


