//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 0 0 1 0 1 1 0 0 0 1 0 1 1 1 0 1 1 0 1 1 1 1 0 0 1 0 1 0 0 0 0 0 1 1 0 1 1 1 0 1 0 1 0 0 0 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:56 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n554, new_n555, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n574, new_n575,
    new_n576, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n613, new_n614, new_n617, new_n619,
    new_n620, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT64), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT65), .ZN(new_n451));
  INV_X1    g026(.A(KEYINPUT2), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT66), .Z(G319));
  XNOR2_X1  g034(.A(KEYINPUT3), .B(G2104), .ZN(new_n460));
  AND2_X1   g035(.A1(new_n460), .A2(G125), .ZN(new_n461));
  AND2_X1   g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  XNOR2_X1  g037(.A(new_n462), .B(KEYINPUT67), .ZN(new_n463));
  OAI21_X1  g038(.A(G2105), .B1(new_n461), .B2(new_n463), .ZN(new_n464));
  OR2_X1    g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(G2105), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n469), .A2(KEYINPUT68), .A3(G101), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n471), .A2(G101), .A3(G2104), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT68), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AOI22_X1  g049(.A1(G137), .A2(new_n467), .B1(new_n470), .B2(new_n474), .ZN(new_n475));
  AND2_X1   g050(.A1(new_n464), .A2(new_n475), .ZN(G160));
  NAND2_X1  g051(.A1(new_n460), .A2(G2105), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  XOR2_X1   g054(.A(new_n479), .B(KEYINPUT69), .Z(new_n480));
  OR2_X1    g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  INV_X1    g056(.A(G112), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n468), .B1(new_n482), .B2(G2105), .ZN(new_n483));
  AOI22_X1  g058(.A1(new_n467), .A2(G136), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n480), .A2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  AND2_X1   g061(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n487));
  NOR2_X1   g062(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n488));
  OAI211_X1 g063(.A(G138), .B(new_n471), .C1(new_n487), .C2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n460), .A2(KEYINPUT4), .A3(G138), .A4(new_n471), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT71), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n460), .A2(G126), .A3(G2105), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(new_n496));
  OAI21_X1  g071(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT70), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n498), .B1(new_n471), .B2(G114), .ZN(new_n499));
  INV_X1    g074(.A(G114), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n500), .A2(KEYINPUT70), .A3(G2105), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n497), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n494), .B1(new_n496), .B2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n502), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n504), .A2(new_n495), .A3(KEYINPUT71), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n493), .B1(new_n503), .B2(new_n505), .ZN(G164));
  INV_X1    g081(.A(G651), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT73), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT5), .ZN(new_n509));
  OAI21_X1  g084(.A(G543), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n508), .B1(new_n509), .B2(KEYINPUT72), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  OAI211_X1 g087(.A(new_n508), .B(G543), .C1(new_n509), .C2(KEYINPUT72), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n512), .A2(G62), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(G75), .A2(G543), .ZN(new_n515));
  XNOR2_X1  g090(.A(new_n515), .B(KEYINPUT74), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n507), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  XNOR2_X1  g092(.A(KEYINPUT6), .B(G651), .ZN(new_n518));
  NAND4_X1  g093(.A1(new_n512), .A2(new_n518), .A3(new_n513), .A4(G88), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n518), .A2(G50), .A3(G543), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n517), .A2(new_n521), .ZN(G166));
  AND3_X1   g097(.A1(new_n512), .A2(new_n518), .A3(new_n513), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G89), .ZN(new_n524));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n525), .B(KEYINPUT7), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n518), .A2(G543), .ZN(new_n527));
  INV_X1    g102(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G51), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n524), .A2(new_n526), .A3(new_n529), .ZN(new_n530));
  NAND4_X1  g105(.A1(new_n512), .A2(new_n513), .A3(G63), .A4(G651), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n531), .B(KEYINPUT75), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n530), .A2(new_n532), .ZN(G168));
  NAND2_X1  g108(.A1(G77), .A2(G543), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n512), .A2(new_n513), .ZN(new_n535));
  INV_X1    g110(.A(G64), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G651), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n523), .A2(G90), .B1(new_n528), .B2(G52), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n538), .A2(new_n539), .ZN(G301));
  INV_X1    g115(.A(G301), .ZN(G171));
  NAND2_X1  g116(.A1(G68), .A2(G543), .ZN(new_n542));
  INV_X1    g117(.A(G56), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n542), .B1(new_n535), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G651), .ZN(new_n545));
  INV_X1    g120(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n528), .A2(G43), .ZN(new_n547));
  INV_X1    g122(.A(new_n523), .ZN(new_n548));
  INV_X1    g123(.A(G81), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n546), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  NAND4_X1  g127(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT8), .ZN(new_n555));
  NAND4_X1  g130(.A1(G319), .A2(G483), .A3(G661), .A4(new_n555), .ZN(G188));
  INV_X1    g131(.A(KEYINPUT9), .ZN(new_n557));
  OAI211_X1 g132(.A(new_n528), .B(G53), .C1(KEYINPUT76), .C2(new_n557), .ZN(new_n558));
  XOR2_X1   g133(.A(KEYINPUT76), .B(KEYINPUT9), .Z(new_n559));
  INV_X1    g134(.A(G53), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n559), .B1(new_n527), .B2(new_n560), .ZN(new_n561));
  AOI22_X1  g136(.A1(new_n558), .A2(new_n561), .B1(G91), .B2(new_n523), .ZN(new_n562));
  NAND2_X1  g137(.A1(G78), .A2(G543), .ZN(new_n563));
  XOR2_X1   g138(.A(new_n563), .B(KEYINPUT77), .Z(new_n564));
  INV_X1    g139(.A(G65), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n564), .B1(new_n535), .B2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT78), .ZN(new_n567));
  AOI21_X1  g142(.A(new_n507), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  OAI211_X1 g143(.A(KEYINPUT78), .B(new_n564), .C1(new_n535), .C2(new_n565), .ZN(new_n569));
  AND3_X1   g144(.A1(new_n568), .A2(KEYINPUT79), .A3(new_n569), .ZN(new_n570));
  AOI21_X1  g145(.A(KEYINPUT79), .B1(new_n568), .B2(new_n569), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n562), .B1(new_n570), .B2(new_n571), .ZN(G299));
  INV_X1    g147(.A(G168), .ZN(G286));
  NAND2_X1  g148(.A1(G166), .A2(KEYINPUT80), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT80), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n575), .B1(new_n517), .B2(new_n521), .ZN(new_n576));
  AND2_X1   g151(.A1(new_n574), .A2(new_n576), .ZN(G303));
  AOI22_X1  g152(.A1(new_n523), .A2(G87), .B1(new_n528), .B2(G49), .ZN(new_n578));
  AND2_X1   g153(.A1(new_n512), .A2(new_n513), .ZN(new_n579));
  OAI21_X1  g154(.A(G651), .B1(new_n579), .B2(G74), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(new_n582));
  OR2_X1    g157(.A1(new_n582), .A2(KEYINPUT81), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(KEYINPUT81), .ZN(new_n584));
  AND2_X1   g159(.A1(new_n583), .A2(new_n584), .ZN(G288));
  NAND2_X1  g160(.A1(G73), .A2(G543), .ZN(new_n586));
  INV_X1    g161(.A(G61), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n535), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n588), .A2(G651), .ZN(new_n589));
  AND2_X1   g164(.A1(G48), .A2(G543), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n518), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT82), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n518), .A2(KEYINPUT82), .A3(new_n590), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n523), .A2(G86), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n589), .A2(new_n595), .ZN(G305));
  AOI22_X1  g171(.A1(new_n579), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n597));
  OR2_X1    g172(.A1(new_n597), .A2(new_n507), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n523), .A2(G85), .B1(new_n528), .B2(G47), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(G290));
  NAND2_X1  g175(.A1(G301), .A2(G868), .ZN(new_n601));
  AND3_X1   g176(.A1(new_n523), .A2(KEYINPUT10), .A3(G92), .ZN(new_n602));
  AOI21_X1  g177(.A(KEYINPUT10), .B1(new_n523), .B2(G92), .ZN(new_n603));
  OR2_X1    g178(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(G79), .A2(G543), .ZN(new_n605));
  INV_X1    g180(.A(G66), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n535), .B2(new_n606), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n607), .A2(G651), .B1(G54), .B2(new_n528), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n601), .B1(new_n610), .B2(G868), .ZN(G284));
  XOR2_X1   g186(.A(G284), .B(KEYINPUT83), .Z(G321));
  NAND2_X1  g187(.A1(G286), .A2(G868), .ZN(new_n613));
  INV_X1    g188(.A(G299), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n613), .B1(new_n614), .B2(G868), .ZN(G297));
  OAI21_X1  g190(.A(new_n613), .B1(new_n614), .B2(G868), .ZN(G280));
  INV_X1    g191(.A(G559), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n610), .B1(new_n617), .B2(G860), .ZN(G148));
  NAND2_X1  g193(.A1(new_n610), .A2(new_n617), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n619), .A2(G868), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n620), .B1(G868), .B2(new_n551), .ZN(G323));
  XNOR2_X1  g196(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g197(.A1(new_n460), .A2(new_n469), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT12), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT13), .ZN(new_n625));
  INV_X1    g200(.A(G2100), .ZN(new_n626));
  OR2_X1    g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n625), .A2(new_n626), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n467), .A2(G135), .ZN(new_n629));
  NOR2_X1   g204(.A1(G99), .A2(G2105), .ZN(new_n630));
  OAI21_X1  g205(.A(G2104), .B1(new_n471), .B2(G111), .ZN(new_n631));
  INV_X1    g206(.A(G123), .ZN(new_n632));
  OAI221_X1 g207(.A(new_n629), .B1(new_n630), .B2(new_n631), .C1(new_n632), .C2(new_n477), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(G2096), .Z(new_n634));
  NAND3_X1  g209(.A1(new_n627), .A2(new_n628), .A3(new_n634), .ZN(G156));
  XOR2_X1   g210(.A(G2451), .B(G2454), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT16), .ZN(new_n637));
  XNOR2_X1  g212(.A(G1341), .B(G1348), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2443), .B(G2446), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2427), .B(G2438), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2430), .ZN(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT15), .B(G2435), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n643), .A2(new_n644), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n645), .A2(new_n646), .A3(KEYINPUT14), .ZN(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(new_n648));
  OR2_X1    g223(.A1(new_n641), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n641), .A2(new_n648), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n649), .A2(new_n650), .A3(G14), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT84), .ZN(G401));
  XNOR2_X1  g227(.A(G2072), .B(G2078), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2084), .B(G2090), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT85), .ZN(new_n655));
  XOR2_X1   g230(.A(G2067), .B(G2678), .Z(new_n656));
  NOR2_X1   g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(KEYINPUT86), .B(KEYINPUT18), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n653), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  INV_X1    g234(.A(new_n658), .ZN(new_n660));
  INV_X1    g235(.A(KEYINPUT17), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n657), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n655), .A2(new_n656), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n660), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  MUX2_X1   g239(.A(new_n659), .B(new_n653), .S(new_n664), .Z(new_n665));
  XOR2_X1   g240(.A(G2096), .B(G2100), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(G227));
  XNOR2_X1  g242(.A(G1971), .B(G1976), .ZN(new_n668));
  INV_X1    g243(.A(KEYINPUT19), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1956), .B(G2474), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1961), .B(G1966), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT20), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n670), .A2(new_n671), .A3(new_n672), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n671), .B(new_n672), .ZN(new_n677));
  AOI21_X1  g252(.A(new_n670), .B1(new_n677), .B2(KEYINPUT87), .ZN(new_n678));
  OAI21_X1  g253(.A(new_n678), .B1(KEYINPUT87), .B2(new_n677), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n675), .A2(new_n676), .A3(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(G1986), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n683));
  AND2_X1   g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n682), .A2(new_n683), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1991), .B(G1996), .ZN(new_n687));
  INV_X1    g262(.A(G1981), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  AND2_X1   g264(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n686), .A2(new_n689), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n690), .A2(new_n691), .ZN(G229));
  INV_X1    g267(.A(KEYINPUT36), .ZN(new_n693));
  INV_X1    g268(.A(G16), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(G6), .ZN(new_n695));
  INV_X1    g270(.A(G305), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n695), .B1(new_n696), .B2(new_n694), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT32), .ZN(new_n698));
  OR2_X1    g273(.A1(new_n698), .A2(G1981), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n698), .A2(G1981), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n694), .A2(G22), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n701), .B1(G166), .B2(new_n694), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n702), .A2(G1971), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n702), .A2(G1971), .ZN(new_n704));
  AND2_X1   g279(.A1(new_n694), .A2(G23), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n705), .B1(new_n581), .B2(G16), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT33), .B(G1976), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n704), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  AOI211_X1 g283(.A(new_n703), .B(new_n708), .C1(new_n706), .C2(new_n707), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n699), .A2(new_n700), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(KEYINPUT34), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n467), .A2(G131), .ZN(new_n712));
  OR2_X1    g287(.A1(G95), .A2(G2105), .ZN(new_n713));
  OAI211_X1 g288(.A(new_n713), .B(G2104), .C1(G107), .C2(new_n471), .ZN(new_n714));
  INV_X1    g289(.A(G119), .ZN(new_n715));
  OAI211_X1 g290(.A(new_n712), .B(new_n714), .C1(new_n715), .C2(new_n477), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT88), .ZN(new_n717));
  MUX2_X1   g292(.A(G25), .B(new_n717), .S(G29), .Z(new_n718));
  XOR2_X1   g293(.A(KEYINPUT35), .B(G1991), .Z(new_n719));
  INV_X1    g294(.A(new_n719), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n718), .B(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n721), .A2(KEYINPUT89), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n721), .A2(KEYINPUT89), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n694), .A2(G24), .ZN(new_n724));
  INV_X1    g299(.A(G290), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n724), .B1(new_n725), .B2(new_n694), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(G1986), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n723), .A2(new_n727), .ZN(new_n728));
  AND3_X1   g303(.A1(new_n711), .A2(new_n722), .A3(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(KEYINPUT90), .ZN(new_n730));
  OR2_X1    g305(.A1(new_n710), .A2(KEYINPUT34), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n729), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(new_n732), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n730), .B1(new_n729), .B2(new_n731), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n693), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  INV_X1    g310(.A(new_n734), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n736), .A2(KEYINPUT36), .A3(new_n732), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n694), .A2(G21), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(G168), .B2(new_n694), .ZN(new_n740));
  OR2_X1    g315(.A1(new_n740), .A2(G1966), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n740), .A2(G1966), .ZN(new_n742));
  INV_X1    g317(.A(G29), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n743), .A2(G27), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G164), .B2(new_n743), .ZN(new_n745));
  INV_X1    g320(.A(G2078), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n741), .A2(new_n742), .A3(new_n747), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n743), .B1(KEYINPUT24), .B2(G34), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(KEYINPUT24), .B2(G34), .ZN(new_n750));
  INV_X1    g325(.A(G160), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n750), .B1(new_n751), .B2(G29), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(KEYINPUT92), .Z(new_n753));
  NAND2_X1  g328(.A1(new_n753), .A2(G2084), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT93), .ZN(new_n755));
  NOR2_X1   g330(.A1(G5), .A2(G16), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(KEYINPUT95), .Z(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(G301), .B2(new_n694), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(KEYINPUT96), .Z(new_n759));
  AOI211_X1 g334(.A(new_n748), .B(new_n755), .C1(G1961), .C2(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n743), .A2(G35), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(G162), .B2(new_n743), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(KEYINPUT98), .Z(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT29), .ZN(new_n764));
  OR2_X1    g339(.A1(new_n764), .A2(G2090), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n694), .A2(G4), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(new_n610), .B2(new_n694), .ZN(new_n767));
  INV_X1    g342(.A(G1348), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n767), .B(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n743), .A2(G33), .ZN(new_n770));
  NAND3_X1  g345(.A1(new_n471), .A2(G103), .A3(G2104), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT25), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n460), .A2(G127), .ZN(new_n773));
  NAND2_X1  g348(.A1(G115), .A2(G2104), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n471), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  AOI211_X1 g350(.A(new_n772), .B(new_n775), .C1(G139), .C2(new_n467), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n770), .B1(new_n776), .B2(new_n743), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n777), .A2(G2072), .ZN(new_n778));
  XNOR2_X1  g353(.A(KEYINPUT31), .B(G11), .ZN(new_n779));
  XNOR2_X1  g354(.A(KEYINPUT94), .B(G28), .ZN(new_n780));
  INV_X1    g355(.A(KEYINPUT30), .ZN(new_n781));
  AOI21_X1  g356(.A(G29), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(new_n781), .B2(new_n780), .ZN(new_n783));
  OAI211_X1 g358(.A(new_n779), .B(new_n783), .C1(new_n633), .C2(new_n743), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n778), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n478), .A2(G129), .ZN(new_n786));
  AOI22_X1  g361(.A1(new_n467), .A2(G141), .B1(G105), .B2(new_n469), .ZN(new_n787));
  NAND3_X1  g362(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(KEYINPUT26), .Z(new_n789));
  NAND3_X1  g364(.A1(new_n786), .A2(new_n787), .A3(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n791), .A2(new_n743), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(new_n743), .B2(G32), .ZN(new_n793));
  XNOR2_X1  g368(.A(KEYINPUT27), .B(G1996), .ZN(new_n794));
  AOI22_X1  g369(.A1(new_n793), .A2(new_n794), .B1(G2072), .B2(new_n777), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n467), .A2(G140), .ZN(new_n796));
  NOR2_X1   g371(.A1(G104), .A2(G2105), .ZN(new_n797));
  OAI21_X1  g372(.A(G2104), .B1(new_n471), .B2(G116), .ZN(new_n798));
  INV_X1    g373(.A(G128), .ZN(new_n799));
  OAI221_X1 g374(.A(new_n796), .B1(new_n797), .B2(new_n798), .C1(new_n799), .C2(new_n477), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n800), .A2(G29), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n743), .A2(G26), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT28), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(G2067), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  AND3_X1   g381(.A1(new_n785), .A2(new_n795), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n694), .A2(G19), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(new_n551), .B2(new_n694), .ZN(new_n809));
  XOR2_X1   g384(.A(KEYINPUT91), .B(G1341), .Z(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  NAND3_X1  g386(.A1(new_n769), .A2(new_n807), .A3(new_n811), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(new_n764), .B2(G2090), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n760), .A2(new_n765), .A3(new_n813), .ZN(new_n814));
  OR2_X1    g389(.A1(new_n793), .A2(new_n794), .ZN(new_n815));
  OAI221_X1 g390(.A(new_n815), .B1(new_n759), .B2(G1961), .C1(G2084), .C2(new_n753), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT97), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n694), .A2(G20), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT23), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n819), .B1(new_n614), .B2(new_n694), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT100), .ZN(new_n821));
  XOR2_X1   g396(.A(KEYINPUT99), .B(G1956), .Z(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  NOR3_X1   g398(.A1(new_n814), .A2(new_n817), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n738), .A2(new_n824), .ZN(G150));
  INV_X1    g400(.A(G150), .ZN(G311));
  NAND2_X1  g401(.A1(G80), .A2(G543), .ZN(new_n827));
  INV_X1    g402(.A(G67), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n827), .B1(new_n535), .B2(new_n828), .ZN(new_n829));
  AND2_X1   g404(.A1(new_n829), .A2(G651), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n523), .A2(G93), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n528), .A2(G55), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n830), .A2(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(G860), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT37), .ZN(new_n837));
  OAI22_X1  g412(.A1(new_n546), .A2(new_n550), .B1(new_n830), .B2(new_n833), .ZN(new_n838));
  AND2_X1   g413(.A1(new_n831), .A2(new_n832), .ZN(new_n839));
  AOI22_X1  g414(.A1(new_n523), .A2(G81), .B1(new_n528), .B2(G43), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n829), .A2(G651), .ZN(new_n841));
  NAND4_X1  g416(.A1(new_n839), .A2(new_n545), .A3(new_n840), .A4(new_n841), .ZN(new_n842));
  AND2_X1   g417(.A1(new_n838), .A2(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT38), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n609), .A2(new_n617), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n844), .B(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n847), .A2(KEYINPUT39), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT101), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n835), .B1(new_n847), .B2(KEYINPUT39), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n837), .B1(new_n849), .B2(new_n850), .ZN(G145));
  XNOR2_X1  g426(.A(new_n717), .B(new_n790), .ZN(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n496), .A2(new_n502), .ZN(new_n854));
  AND3_X1   g429(.A1(new_n491), .A2(new_n492), .A3(KEYINPUT102), .ZN(new_n855));
  AOI21_X1  g430(.A(KEYINPUT102), .B1(new_n491), .B2(new_n492), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n854), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(new_n800), .ZN(new_n858));
  OR2_X1    g433(.A1(new_n858), .A2(new_n776), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n776), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n467), .A2(G142), .ZN(new_n861));
  NOR2_X1   g436(.A1(G106), .A2(G2105), .ZN(new_n862));
  OAI21_X1  g437(.A(G2104), .B1(new_n471), .B2(G118), .ZN(new_n863));
  INV_X1    g438(.A(G130), .ZN(new_n864));
  OAI221_X1 g439(.A(new_n861), .B1(new_n862), .B2(new_n863), .C1(new_n864), .C2(new_n477), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(new_n624), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n859), .A2(new_n860), .A3(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n867), .B1(new_n859), .B2(new_n860), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n853), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n485), .B(new_n633), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(G160), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n858), .B(new_n776), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n874), .A2(new_n866), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n875), .A2(new_n852), .A3(new_n868), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n871), .A2(new_n873), .A3(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT103), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND4_X1  g454(.A1(new_n871), .A2(KEYINPUT103), .A3(new_n873), .A4(new_n876), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n873), .B1(new_n871), .B2(new_n876), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n882), .A2(G37), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g460(.A1(new_n838), .A2(new_n842), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(KEYINPUT104), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(new_n619), .ZN(new_n888));
  NAND2_X1  g463(.A1(G299), .A2(new_n610), .ZN(new_n889));
  OAI211_X1 g464(.A(new_n609), .B(new_n562), .C1(new_n571), .C2(new_n570), .ZN(new_n890));
  AOI21_X1  g465(.A(KEYINPUT41), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n889), .A2(KEYINPUT41), .A3(new_n890), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n888), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n889), .A2(new_n890), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n895), .B1(new_n897), .B2(new_n888), .ZN(new_n898));
  XNOR2_X1  g473(.A(G290), .B(new_n696), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n581), .B(G166), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n899), .B(new_n900), .ZN(new_n901));
  XOR2_X1   g476(.A(new_n901), .B(KEYINPUT42), .Z(new_n902));
  XNOR2_X1  g477(.A(new_n898), .B(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n903), .A2(G868), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n904), .B1(G868), .B2(new_n834), .ZN(G295));
  OAI21_X1  g480(.A(new_n904), .B1(G868), .B2(new_n834), .ZN(G331));
  AND3_X1   g481(.A1(new_n524), .A2(new_n526), .A3(new_n529), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT75), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n531), .B(new_n908), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n907), .A2(new_n909), .A3(new_n538), .A4(new_n539), .ZN(new_n910));
  OAI21_X1  g485(.A(G301), .B1(new_n532), .B2(new_n530), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(new_n886), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT106), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n912), .A2(new_n886), .A3(KEYINPUT106), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND4_X1  g492(.A1(new_n843), .A2(KEYINPUT107), .A3(new_n911), .A4(new_n910), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n910), .A2(new_n838), .A3(new_n911), .A4(new_n842), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT107), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n918), .A2(new_n921), .ZN(new_n922));
  AND2_X1   g497(.A1(new_n917), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n923), .A2(new_n896), .ZN(new_n924));
  INV_X1    g499(.A(new_n893), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT109), .ZN(new_n926));
  NOR3_X1   g501(.A1(new_n925), .A2(new_n926), .A3(new_n891), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n891), .A2(new_n926), .ZN(new_n928));
  NAND4_X1  g503(.A1(new_n843), .A2(KEYINPUT108), .A3(new_n911), .A4(new_n910), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT108), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n919), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n929), .A2(new_n913), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n928), .A2(new_n932), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n924), .B1(new_n927), .B2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(new_n901), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n932), .A2(new_n897), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n917), .A2(new_n922), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n937), .B1(new_n894), .B2(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(G37), .B1(new_n939), .B2(new_n901), .ZN(new_n940));
  XNOR2_X1  g515(.A(KEYINPUT105), .B(KEYINPUT43), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n936), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  AOI22_X1  g517(.A1(new_n892), .A2(new_n893), .B1(new_n917), .B2(new_n922), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n935), .B1(new_n943), .B2(new_n937), .ZN(new_n944));
  OR2_X1    g519(.A1(new_n932), .A2(new_n897), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n925), .A2(new_n891), .ZN(new_n946));
  OAI211_X1 g521(.A(new_n945), .B(new_n901), .C1(new_n946), .C2(new_n923), .ZN(new_n947));
  INV_X1    g522(.A(G37), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n944), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(new_n941), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n942), .A2(new_n951), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n952), .A2(KEYINPUT44), .ZN(new_n953));
  OAI211_X1 g528(.A(new_n928), .B(new_n932), .C1(new_n894), .C2(new_n926), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n901), .B1(new_n954), .B2(new_n924), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n947), .A2(new_n948), .ZN(new_n956));
  OAI21_X1  g531(.A(KEYINPUT43), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n957), .B1(new_n950), .B2(new_n949), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n953), .B1(KEYINPUT44), .B2(new_n958), .ZN(G397));
  INV_X1    g534(.A(G1384), .ZN(new_n960));
  AOI21_X1  g535(.A(KEYINPUT45), .B1(new_n857), .B2(new_n960), .ZN(new_n961));
  AND3_X1   g536(.A1(new_n464), .A2(G40), .A3(new_n475), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  XNOR2_X1  g538(.A(new_n963), .B(KEYINPUT110), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n964), .A2(G1996), .A3(new_n790), .ZN(new_n965));
  XNOR2_X1  g540(.A(new_n965), .B(KEYINPUT111), .ZN(new_n966));
  XNOR2_X1  g541(.A(new_n800), .B(G2067), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n963), .A2(G1996), .ZN(new_n968));
  AOI22_X1  g543(.A1(new_n964), .A2(new_n967), .B1(new_n791), .B2(new_n968), .ZN(new_n969));
  AND2_X1   g544(.A1(new_n966), .A2(new_n969), .ZN(new_n970));
  AND2_X1   g545(.A1(new_n717), .A2(new_n720), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n717), .A2(new_n720), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n964), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n970), .A2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(new_n963), .ZN(new_n975));
  XNOR2_X1  g550(.A(G290), .B(G1986), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n974), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT120), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n574), .A2(G8), .A3(new_n576), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT55), .ZN(new_n980));
  XNOR2_X1  g555(.A(new_n979), .B(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(G8), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n857), .A2(KEYINPUT45), .A3(new_n960), .ZN(new_n983));
  NOR2_X1   g558(.A1(G164), .A2(G1384), .ZN(new_n984));
  OAI211_X1 g559(.A(new_n983), .B(new_n962), .C1(new_n984), .C2(KEYINPUT45), .ZN(new_n985));
  INV_X1    g560(.A(G1971), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT50), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n984), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n857), .A2(new_n960), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(KEYINPUT50), .ZN(new_n991));
  XOR2_X1   g566(.A(KEYINPUT112), .B(G2090), .Z(new_n992));
  NAND4_X1  g567(.A1(new_n989), .A2(new_n991), .A3(new_n962), .A4(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n987), .A2(new_n993), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n982), .B1(new_n994), .B2(KEYINPUT116), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT116), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n987), .A2(new_n996), .A3(new_n993), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n981), .B1(new_n995), .B2(new_n997), .ZN(new_n998));
  AND2_X1   g573(.A1(new_n985), .A2(new_n986), .ZN(new_n999));
  OAI21_X1  g574(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n857), .A2(new_n988), .A3(new_n960), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n1000), .A2(new_n962), .A3(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(new_n992), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  OAI211_X1 g579(.A(G8), .B(new_n981), .C1(new_n999), .C2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n962), .A2(new_n857), .A3(new_n960), .ZN(new_n1006));
  AOI21_X1  g581(.A(KEYINPUT113), .B1(new_n1006), .B2(G8), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1006), .A2(KEYINPUT113), .A3(G8), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n589), .A2(KEYINPUT114), .ZN(new_n1011));
  NAND3_X1  g586(.A1(G305), .A2(new_n1011), .A3(G1981), .ZN(new_n1012));
  OAI211_X1 g587(.A(new_n589), .B(new_n595), .C1(KEYINPUT114), .C2(new_n688), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1012), .A2(KEYINPUT49), .A3(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(KEYINPUT49), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT115), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  AOI211_X1 g592(.A(KEYINPUT115), .B(KEYINPUT49), .C1(new_n1012), .C2(new_n1013), .ZN(new_n1018));
  OAI211_X1 g593(.A(new_n1010), .B(new_n1014), .C1(new_n1017), .C2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n582), .A2(G1976), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1009), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1020), .B1(new_n1021), .B2(new_n1007), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(KEYINPUT52), .ZN(new_n1023));
  INV_X1    g598(.A(G1976), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n583), .A2(new_n1024), .A3(new_n584), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT52), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n1010), .A2(new_n1025), .A3(new_n1026), .A4(new_n1020), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n1005), .A2(new_n1019), .A3(new_n1023), .A4(new_n1027), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n998), .A2(new_n1028), .ZN(new_n1029));
  NOR2_X1   g604(.A1(G286), .A2(new_n982), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1030), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1002), .A2(G2084), .ZN(new_n1032));
  INV_X1    g607(.A(new_n962), .ZN(new_n1033));
  OAI21_X1  g608(.A(KEYINPUT117), .B1(new_n961), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT117), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT102), .ZN(new_n1036));
  AOI21_X1  g611(.A(KEYINPUT4), .B1(new_n467), .B2(G138), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n489), .A2(new_n490), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1036), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n491), .A2(new_n492), .A3(KEYINPUT102), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(G1384), .B1(new_n1041), .B2(new_n854), .ZN(new_n1042));
  OAI211_X1 g617(.A(new_n1035), .B(new_n962), .C1(new_n1042), .C2(KEYINPUT45), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n984), .A2(KEYINPUT45), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1034), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(G1966), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1032), .B1(new_n1047), .B2(KEYINPUT118), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT118), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1045), .A2(new_n1049), .A3(new_n1046), .ZN(new_n1050));
  AOI211_X1 g625(.A(KEYINPUT119), .B(new_n1031), .C1(new_n1048), .C2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT119), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1047), .A2(KEYINPUT118), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1032), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1053), .A2(new_n1050), .A3(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1052), .B1(new_n1055), .B2(new_n1030), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1029), .B1(new_n1051), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT63), .ZN(new_n1058));
  AND3_X1   g633(.A1(new_n1045), .A2(new_n1049), .A3(new_n1046), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1049), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1060));
  NOR3_X1   g635(.A1(new_n1059), .A2(new_n1060), .A3(new_n1032), .ZN(new_n1061));
  OAI21_X1  g636(.A(KEYINPUT119), .B1(new_n1061), .B2(new_n1031), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1055), .A2(new_n1052), .A3(new_n1030), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n999), .A2(new_n1004), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1065), .A2(new_n982), .ZN(new_n1066));
  OAI21_X1  g641(.A(KEYINPUT63), .B1(new_n1066), .B2(new_n981), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1067), .A2(new_n1028), .ZN(new_n1068));
  AOI22_X1  g643(.A1(new_n1057), .A2(new_n1058), .B1(new_n1064), .B2(new_n1068), .ZN(new_n1069));
  NOR2_X1   g644(.A1(G288), .A2(G1976), .ZN(new_n1070));
  AOI22_X1  g645(.A1(new_n1019), .A2(new_n1070), .B1(new_n688), .B2(new_n696), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1010), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1005), .ZN(new_n1074));
  AND3_X1   g649(.A1(new_n1019), .A2(new_n1023), .A3(new_n1027), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1073), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1076), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n978), .B1(new_n1069), .B2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g653(.A(KEYINPUT63), .B1(new_n1064), .B2(new_n1029), .ZN(new_n1079));
  AOI211_X1 g654(.A(new_n1028), .B(new_n1067), .C1(new_n1062), .C2(new_n1063), .ZN(new_n1080));
  OAI211_X1 g655(.A(KEYINPUT120), .B(new_n1076), .C1(new_n1079), .C2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1078), .A2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1029), .ZN(new_n1083));
  NOR2_X1   g658(.A1(KEYINPUT124), .A2(KEYINPUT51), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1084), .B1(new_n1055), .B2(G286), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1053), .A2(G168), .A3(new_n1050), .A4(new_n1054), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(G8), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1088));
  AND2_X1   g663(.A1(KEYINPUT124), .A2(KEYINPUT51), .ZN(new_n1089));
  AOI211_X1 g664(.A(new_n1084), .B(new_n1089), .C1(new_n1086), .C2(G8), .ZN(new_n1090));
  OAI21_X1  g665(.A(KEYINPUT62), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1089), .A2(new_n1084), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1087), .A2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT62), .ZN(new_n1094));
  OAI211_X1 g669(.A(new_n1093), .B(new_n1094), .C1(new_n1087), .C2(new_n1085), .ZN(new_n1095));
  OR2_X1    g670(.A1(G164), .A2(G1384), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT45), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1033), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1098), .A2(new_n746), .A3(new_n983), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT53), .ZN(new_n1100));
  INV_X1    g675(.A(G1961), .ZN(new_n1101));
  AOI22_X1  g676(.A1(new_n1099), .A2(new_n1100), .B1(new_n1101), .B2(new_n1002), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1100), .A2(G2078), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1034), .A2(new_n1043), .A3(new_n1044), .A4(new_n1103), .ZN(new_n1104));
  AND2_X1   g679(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1105), .A2(G301), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1091), .A2(new_n1095), .A3(new_n1106), .ZN(new_n1107));
  XNOR2_X1  g682(.A(G301), .B(KEYINPUT54), .ZN(new_n1108));
  INV_X1    g683(.A(new_n961), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1109), .A2(new_n983), .A3(new_n962), .A4(new_n1103), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1108), .B1(new_n1102), .B2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1111), .B1(new_n1108), .B2(new_n1105), .ZN(new_n1112));
  NAND2_X1  g687(.A1(KEYINPUT122), .A2(KEYINPUT61), .ZN(new_n1113));
  XNOR2_X1  g688(.A(KEYINPUT56), .B(G2072), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1098), .A2(new_n983), .A3(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n989), .A2(new_n962), .A3(new_n991), .ZN(new_n1116));
  INV_X1    g691(.A(G1956), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1115), .A2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(KEYINPUT121), .B1(new_n558), .B2(new_n561), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1120), .A2(KEYINPUT57), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1121), .ZN(new_n1122));
  XNOR2_X1  g697(.A(G299), .B(new_n1122), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1113), .B1(new_n1119), .B2(new_n1123), .ZN(new_n1124));
  XNOR2_X1  g699(.A(G299), .B(new_n1121), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1113), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1125), .A2(new_n1118), .A3(new_n1115), .A4(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1119), .A2(new_n1123), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1124), .A2(new_n1127), .A3(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1006), .ZN(new_n1130));
  XNOR2_X1  g705(.A(KEYINPUT58), .B(G1341), .ZN(new_n1131));
  OAI22_X1  g706(.A1(new_n985), .A2(G1996), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1132), .A2(new_n551), .ZN(new_n1133));
  XNOR2_X1  g708(.A(new_n1133), .B(KEYINPUT59), .ZN(new_n1134));
  AOI22_X1  g709(.A1(new_n1002), .A2(new_n768), .B1(new_n805), .B2(new_n1130), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1135), .A2(KEYINPUT60), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1136), .A2(KEYINPUT123), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1137), .A2(new_n610), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1136), .A2(KEYINPUT123), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  OAI22_X1  g715(.A1(new_n1137), .A2(new_n610), .B1(KEYINPUT60), .B2(new_n1135), .ZN(new_n1141));
  OAI211_X1 g716(.A(new_n1129), .B(new_n1134), .C1(new_n1140), .C2(new_n1141), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1135), .A2(new_n609), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1143), .B1(new_n1119), .B2(new_n1123), .ZN(new_n1144));
  AND2_X1   g719(.A1(new_n1144), .A2(new_n1128), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1112), .B1(new_n1142), .B2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1093), .B1(new_n1087), .B2(new_n1085), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1083), .B1(new_n1107), .B2(new_n1148), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n977), .B1(new_n1082), .B2(new_n1149), .ZN(new_n1150));
  XOR2_X1   g725(.A(new_n968), .B(KEYINPUT46), .Z(new_n1151));
  OAI21_X1  g726(.A(new_n964), .B1(new_n790), .B2(new_n967), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  XOR2_X1   g728(.A(KEYINPUT125), .B(KEYINPUT47), .Z(new_n1154));
  XNOR2_X1  g729(.A(new_n1153), .B(new_n1154), .ZN(new_n1155));
  NOR3_X1   g730(.A1(new_n963), .A2(G1986), .A3(G290), .ZN(new_n1156));
  XNOR2_X1  g731(.A(new_n1156), .B(KEYINPUT48), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1155), .B1(new_n974), .B2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n970), .A2(new_n972), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1159), .B1(G2067), .B2(new_n800), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1158), .B1(new_n964), .B2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1150), .A2(new_n1161), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g737(.A(KEYINPUT127), .ZN(new_n1164));
  INV_X1    g738(.A(KEYINPUT126), .ZN(new_n1165));
  NAND2_X1  g739(.A1(G319), .A2(new_n651), .ZN(new_n1166));
  NOR2_X1   g740(.A1(new_n1166), .A2(G227), .ZN(new_n1167));
  OAI21_X1  g741(.A(new_n1167), .B1(new_n690), .B2(new_n691), .ZN(new_n1168));
  AOI21_X1  g742(.A(new_n1168), .B1(new_n881), .B2(new_n883), .ZN(new_n1169));
  AND3_X1   g743(.A1(new_n952), .A2(new_n1165), .A3(new_n1169), .ZN(new_n1170));
  AOI21_X1  g744(.A(new_n1165), .B1(new_n952), .B2(new_n1169), .ZN(new_n1171));
  OAI21_X1  g745(.A(new_n1164), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g746(.A1(new_n952), .A2(new_n1169), .ZN(new_n1173));
  NAND2_X1  g747(.A1(new_n1173), .A2(KEYINPUT126), .ZN(new_n1174));
  NAND3_X1  g748(.A1(new_n952), .A2(new_n1165), .A3(new_n1169), .ZN(new_n1175));
  NAND3_X1  g749(.A1(new_n1174), .A2(KEYINPUT127), .A3(new_n1175), .ZN(new_n1176));
  NAND2_X1  g750(.A1(new_n1172), .A2(new_n1176), .ZN(G308));
  NAND2_X1  g751(.A1(new_n1174), .A2(new_n1175), .ZN(G225));
endmodule


