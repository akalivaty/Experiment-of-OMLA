//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 0 1 1 1 1 0 1 1 1 0 1 1 0 0 0 0 0 1 0 1 0 1 1 0 1 1 0 0 1 0 1 0 1 0 1 1 1 0 0 0 1 0 1 1 1 0 0 0 1 0 1 0 1 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n708, new_n709, new_n710,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n742,
    new_n743, new_n744, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n753, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n782,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n840, new_n841,
    new_n843, new_n844, new_n846, new_n847, new_n848, new_n849, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n915, new_n916,
    new_n917, new_n919, new_n920, new_n921, new_n922, new_n923, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n990, new_n991;
  INV_X1    g000(.A(KEYINPUT91), .ZN(new_n202));
  NAND2_X1  g001(.A1(G229gat), .A2(G233gat), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(G43gat), .B(G50gat), .ZN(new_n205));
  OAI21_X1  g004(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  NOR3_X1   g006(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n208));
  OAI22_X1  g007(.A1(new_n205), .A2(KEYINPUT15), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  AND2_X1   g008(.A1(new_n205), .A2(KEYINPUT15), .ZN(new_n210));
  INV_X1    g009(.A(G29gat), .ZN(new_n211));
  INV_X1    g010(.A(G36gat), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NOR3_X1   g012(.A1(new_n209), .A2(new_n210), .A3(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n206), .A2(KEYINPUT86), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT86), .ZN(new_n216));
  OAI211_X1 g015(.A(new_n216), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(new_n208), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n213), .B1(new_n220), .B2(KEYINPUT87), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n208), .B1(new_n215), .B2(new_n217), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT87), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n221), .A2(new_n224), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n214), .B1(new_n225), .B2(new_n210), .ZN(new_n226));
  XNOR2_X1  g025(.A(G15gat), .B(G22gat), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n227), .A2(G1gat), .ZN(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT16), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n227), .B1(new_n230), .B2(G1gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  OAI21_X1  g031(.A(G8gat), .B1(new_n228), .B2(KEYINPUT88), .ZN(new_n233));
  XNOR2_X1  g032(.A(new_n232), .B(new_n233), .ZN(new_n234));
  OAI21_X1  g033(.A(KEYINPUT90), .B1(new_n226), .B2(new_n234), .ZN(new_n235));
  OAI22_X1  g034(.A1(new_n222), .A2(new_n223), .B1(new_n211), .B2(new_n212), .ZN(new_n236));
  AND2_X1   g035(.A1(new_n222), .A2(new_n223), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n210), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(new_n214), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT90), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n233), .A2(new_n229), .A3(new_n231), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n233), .B1(new_n229), .B2(new_n231), .ZN(new_n244));
  OAI211_X1 g043(.A(new_n240), .B(new_n241), .C1(new_n243), .C2(new_n244), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n204), .B1(new_n235), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n240), .A2(KEYINPUT17), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT17), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n238), .A2(new_n248), .A3(new_n239), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(KEYINPUT89), .B1(new_n250), .B2(new_n234), .ZN(new_n251));
  AND3_X1   g050(.A1(new_n238), .A2(new_n248), .A3(new_n239), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n248), .B1(new_n238), .B2(new_n239), .ZN(new_n253));
  OAI211_X1 g052(.A(KEYINPUT89), .B(new_n234), .C1(new_n252), .C2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n246), .B1(new_n251), .B2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT18), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n234), .B1(new_n252), .B2(new_n253), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT89), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(new_n254), .ZN(new_n262));
  AOI211_X1 g061(.A(new_n257), .B(new_n204), .C1(new_n235), .C2(new_n245), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n235), .A2(new_n245), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n226), .A2(new_n234), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  XOR2_X1   g065(.A(new_n203), .B(KEYINPUT13), .Z(new_n267));
  AOI22_X1  g066(.A1(new_n262), .A2(new_n263), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  XNOR2_X1  g067(.A(G113gat), .B(G141gat), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n269), .B(G197gat), .ZN(new_n270));
  XOR2_X1   g069(.A(KEYINPUT11), .B(G169gat), .Z(new_n271));
  XNOR2_X1  g070(.A(new_n270), .B(new_n271), .ZN(new_n272));
  XOR2_X1   g071(.A(new_n272), .B(KEYINPUT12), .Z(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  AND3_X1   g073(.A1(new_n258), .A2(new_n268), .A3(new_n274), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n274), .B1(new_n258), .B2(new_n268), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n202), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n258), .A2(new_n268), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(new_n273), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n258), .A2(new_n268), .A3(new_n274), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n279), .A2(new_n280), .A3(KEYINPUT91), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n277), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  XNOR2_X1  g082(.A(G190gat), .B(G218gat), .ZN(new_n284));
  XNOR2_X1  g083(.A(KEYINPUT99), .B(KEYINPUT100), .ZN(new_n285));
  XOR2_X1   g084(.A(new_n284), .B(new_n285), .Z(new_n286));
  INV_X1    g085(.A(G85gat), .ZN(new_n287));
  INV_X1    g086(.A(G92gat), .ZN(new_n288));
  OAI211_X1 g087(.A(KEYINPUT97), .B(KEYINPUT7), .C1(new_n287), .C2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(KEYINPUT97), .A2(KEYINPUT7), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n290), .A2(G85gat), .A3(G92gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(G99gat), .A2(G106gat), .ZN(new_n293));
  AOI22_X1  g092(.A1(KEYINPUT8), .A2(new_n293), .B1(new_n287), .B2(new_n288), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  XOR2_X1   g094(.A(G99gat), .B(G106gat), .Z(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n296), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n298), .A2(new_n292), .A3(new_n294), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT98), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n297), .A2(KEYINPUT98), .A3(new_n299), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n250), .A2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n304), .ZN(new_n306));
  AND2_X1   g105(.A1(G232gat), .A2(G233gat), .ZN(new_n307));
  AOI22_X1  g106(.A1(new_n306), .A2(new_n240), .B1(KEYINPUT41), .B2(new_n307), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n286), .B1(new_n305), .B2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT101), .ZN(new_n310));
  XOR2_X1   g109(.A(G134gat), .B(G162gat), .Z(new_n311));
  NOR2_X1   g110(.A1(new_n307), .A2(KEYINPUT41), .ZN(new_n312));
  XNOR2_X1  g111(.A(new_n311), .B(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n309), .B1(new_n310), .B2(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n305), .A2(new_n308), .A3(new_n286), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n313), .A2(KEYINPUT101), .ZN(new_n317));
  XOR2_X1   g116(.A(new_n317), .B(KEYINPUT102), .Z(new_n318));
  AND3_X1   g117(.A1(new_n315), .A2(new_n316), .A3(new_n318), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n318), .B1(new_n315), .B2(new_n316), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(G71gat), .A2(G78gat), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT93), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  OR2_X1    g124(.A1(G71gat), .A2(G78gat), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT92), .ZN(new_n327));
  NAND3_X1  g126(.A1(KEYINPUT93), .A2(G71gat), .A3(G78gat), .ZN(new_n328));
  NAND4_X1  g127(.A1(new_n325), .A2(new_n326), .A3(new_n327), .A4(new_n328), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n327), .B1(G71gat), .B2(G78gat), .ZN(new_n330));
  AND3_X1   g129(.A1(KEYINPUT93), .A2(G71gat), .A3(G78gat), .ZN(new_n331));
  AOI21_X1  g130(.A(KEYINPUT93), .B1(G71gat), .B2(G78gat), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n330), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n329), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(G57gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(G64gat), .ZN(new_n336));
  INV_X1    g135(.A(G64gat), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(G57gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT9), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n323), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n334), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n326), .A2(new_n323), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT94), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n326), .A2(KEYINPUT94), .A3(new_n323), .ZN(new_n347));
  NAND4_X1  g146(.A1(new_n346), .A2(new_n341), .A3(new_n339), .A4(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n343), .A2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT21), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(G231gat), .A2(G233gat), .ZN(new_n352));
  XNOR2_X1  g151(.A(new_n351), .B(new_n352), .ZN(new_n353));
  XNOR2_X1  g152(.A(G127gat), .B(G155gat), .ZN(new_n354));
  XNOR2_X1  g153(.A(new_n354), .B(KEYINPUT20), .ZN(new_n355));
  XNOR2_X1  g154(.A(new_n353), .B(new_n355), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n234), .B1(new_n350), .B2(new_n349), .ZN(new_n357));
  XNOR2_X1  g156(.A(new_n357), .B(KEYINPUT96), .ZN(new_n358));
  XNOR2_X1  g157(.A(new_n356), .B(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(G183gat), .B(G211gat), .ZN(new_n360));
  XNOR2_X1  g159(.A(KEYINPUT95), .B(KEYINPUT19), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n360), .B(new_n361), .ZN(new_n362));
  AND2_X1   g161(.A1(new_n359), .A2(new_n362), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n359), .A2(new_n362), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n322), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(G230gat), .A2(G233gat), .ZN(new_n367));
  AOI21_X1  g166(.A(KEYINPUT94), .B1(new_n326), .B2(new_n323), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n342), .A2(new_n368), .ZN(new_n369));
  AOI22_X1  g168(.A1(new_n369), .A2(new_n347), .B1(new_n334), .B2(new_n342), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n298), .A2(KEYINPUT103), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n370), .A2(new_n299), .A3(new_n297), .A4(new_n372), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n300), .B1(new_n349), .B2(new_n371), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n367), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  OR2_X1    g174(.A1(new_n375), .A2(KEYINPUT104), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n373), .A2(new_n374), .ZN(new_n377));
  INV_X1    g176(.A(new_n367), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n377), .A2(KEYINPUT104), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n376), .A2(new_n379), .ZN(new_n380));
  OR2_X1    g179(.A1(new_n380), .A2(KEYINPUT105), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT10), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n373), .A2(new_n374), .A3(new_n382), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n302), .A2(KEYINPUT10), .A3(new_n370), .A4(new_n303), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(new_n367), .ZN(new_n386));
  XNOR2_X1  g185(.A(G120gat), .B(G148gat), .ZN(new_n387));
  XNOR2_X1  g186(.A(G176gat), .B(G204gat), .ZN(new_n388));
  XOR2_X1   g187(.A(new_n387), .B(new_n388), .Z(new_n389));
  NAND2_X1  g188(.A1(new_n380), .A2(KEYINPUT105), .ZN(new_n390));
  NAND4_X1  g189(.A1(new_n381), .A2(new_n386), .A3(new_n389), .A4(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(new_n389), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n378), .B1(new_n383), .B2(new_n384), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n392), .B1(new_n380), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n391), .A2(new_n394), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n366), .A2(new_n395), .ZN(new_n396));
  XNOR2_X1  g195(.A(G211gat), .B(G218gat), .ZN(new_n397));
  XNOR2_X1  g196(.A(new_n397), .B(KEYINPUT77), .ZN(new_n398));
  XNOR2_X1  g197(.A(G197gat), .B(G204gat), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT22), .ZN(new_n400));
  INV_X1    g199(.A(G211gat), .ZN(new_n401));
  INV_X1    g200(.A(G218gat), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n400), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n399), .A2(new_n403), .ZN(new_n404));
  OR2_X1    g203(.A1(new_n398), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n398), .A2(new_n404), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NOR2_X1   g206(.A1(G169gat), .A2(G176gat), .ZN(new_n408));
  XNOR2_X1  g207(.A(new_n408), .B(KEYINPUT26), .ZN(new_n409));
  NAND2_X1  g208(.A1(G169gat), .A2(G176gat), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT66), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(KEYINPUT66), .A2(G169gat), .A3(G176gat), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n409), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(G183gat), .A2(G190gat), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT71), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT70), .ZN(new_n419));
  INV_X1    g218(.A(G183gat), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(KEYINPUT27), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT27), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(G183gat), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n419), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n419), .B1(new_n422), .B2(G183gat), .ZN(new_n425));
  INV_X1    g224(.A(G190gat), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n418), .B1(new_n424), .B2(new_n427), .ZN(new_n428));
  AOI21_X1  g227(.A(G190gat), .B1(new_n421), .B2(new_n419), .ZN(new_n429));
  XNOR2_X1  g228(.A(KEYINPUT27), .B(G183gat), .ZN(new_n430));
  OAI211_X1 g229(.A(new_n429), .B(KEYINPUT71), .C1(new_n419), .C2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT28), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n428), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n430), .A2(KEYINPUT28), .A3(new_n426), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT72), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n417), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n433), .A2(KEYINPUT72), .A3(new_n434), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT25), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n408), .A2(KEYINPUT23), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT65), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  OR2_X1    g242(.A1(new_n408), .A2(KEYINPUT23), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n408), .A2(KEYINPUT65), .A3(KEYINPUT23), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n443), .A2(new_n444), .A3(new_n414), .A4(new_n445), .ZN(new_n446));
  AND2_X1   g245(.A1(new_n446), .A2(KEYINPUT67), .ZN(new_n447));
  OAI211_X1 g246(.A(KEYINPUT64), .B(KEYINPUT24), .C1(G183gat), .C2(G190gat), .ZN(new_n448));
  INV_X1    g247(.A(new_n416), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NOR2_X1   g249(.A1(KEYINPUT64), .A2(KEYINPUT24), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n451), .A2(new_n416), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n450), .B1(new_n448), .B2(new_n452), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n453), .B1(new_n446), .B2(KEYINPUT67), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n440), .B1(new_n447), .B2(new_n454), .ZN(new_n455));
  XNOR2_X1  g254(.A(new_n414), .B(KEYINPUT68), .ZN(new_n456));
  NOR3_X1   g255(.A1(new_n416), .A2(KEYINPUT69), .A3(KEYINPUT24), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n457), .B1(KEYINPUT23), .B2(new_n408), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n420), .A2(new_n426), .ZN(new_n459));
  OAI211_X1 g258(.A(new_n459), .B(new_n416), .C1(KEYINPUT69), .C2(KEYINPUT24), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n458), .A2(new_n460), .A3(KEYINPUT25), .A4(new_n444), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n455), .B1(new_n456), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(G226gat), .A2(G233gat), .ZN(new_n463));
  AND3_X1   g262(.A1(new_n439), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT29), .ZN(new_n465));
  AOI22_X1  g264(.A1(new_n439), .A2(new_n462), .B1(new_n465), .B2(new_n463), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n407), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n463), .A2(new_n465), .ZN(new_n468));
  AND3_X1   g267(.A1(new_n433), .A2(KEYINPUT72), .A3(new_n434), .ZN(new_n469));
  AOI21_X1  g268(.A(KEYINPUT72), .B1(new_n433), .B2(new_n434), .ZN(new_n470));
  NOR3_X1   g269(.A1(new_n469), .A2(new_n470), .A3(new_n417), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n461), .A2(new_n456), .ZN(new_n472));
  OR2_X1    g271(.A1(new_n446), .A2(KEYINPUT67), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n446), .A2(KEYINPUT67), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n473), .A2(new_n474), .A3(new_n453), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n472), .B1(new_n475), .B2(new_n440), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n468), .B1(new_n471), .B2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(new_n407), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n439), .A2(new_n462), .A3(new_n463), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n477), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT78), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n467), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n477), .A2(new_n479), .A3(KEYINPUT78), .A4(new_n478), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  XNOR2_X1  g283(.A(G8gat), .B(G36gat), .ZN(new_n485));
  XNOR2_X1  g284(.A(G64gat), .B(G92gat), .ZN(new_n486));
  XOR2_X1   g285(.A(new_n485), .B(new_n486), .Z(new_n487));
  NAND2_X1  g286(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  XOR2_X1   g287(.A(new_n487), .B(KEYINPUT79), .Z(new_n489));
  NAND3_X1  g288(.A1(new_n482), .A2(new_n489), .A3(new_n483), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(KEYINPUT30), .ZN(new_n492));
  INV_X1    g291(.A(new_n487), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n493), .B1(new_n482), .B2(new_n483), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n494), .A2(KEYINPUT30), .ZN(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n492), .A2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(G113gat), .ZN(new_n498));
  INV_X1    g297(.A(G120gat), .ZN(new_n499));
  AOI21_X1  g298(.A(KEYINPUT1), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  XNOR2_X1  g299(.A(G127gat), .B(G134gat), .ZN(new_n501));
  OAI221_X1 g300(.A(new_n500), .B1(new_n498), .B2(new_n499), .C1(new_n501), .C2(KEYINPUT73), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(KEYINPUT73), .ZN(new_n503));
  XOR2_X1   g302(.A(new_n502), .B(new_n503), .Z(new_n504));
  XOR2_X1   g303(.A(G141gat), .B(G148gat), .Z(new_n505));
  XNOR2_X1  g304(.A(G155gat), .B(G162gat), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT2), .ZN(new_n508));
  XNOR2_X1  g307(.A(KEYINPUT80), .B(G155gat), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n508), .B1(new_n509), .B2(G162gat), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n506), .B1(new_n505), .B2(new_n508), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n504), .A2(KEYINPUT4), .A3(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT4), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n502), .B(new_n503), .ZN(new_n516));
  OR2_X1    g315(.A1(new_n511), .A2(new_n512), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  AND2_X1   g317(.A1(new_n514), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(G225gat), .A2(G233gat), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n517), .A2(KEYINPUT3), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT3), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n513), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n521), .A2(new_n523), .A3(new_n516), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n519), .A2(KEYINPUT5), .A3(new_n520), .A4(new_n524), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n524), .A2(new_n514), .A3(new_n518), .ZN(new_n526));
  INV_X1    g325(.A(new_n520), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT5), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n516), .B(new_n517), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n529), .B1(new_n530), .B2(new_n527), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n525), .B1(new_n528), .B2(new_n531), .ZN(new_n532));
  XNOR2_X1  g331(.A(G1gat), .B(G29gat), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n533), .B(KEYINPUT0), .ZN(new_n534));
  XNOR2_X1  g333(.A(G57gat), .B(G85gat), .ZN(new_n535));
  XOR2_X1   g334(.A(new_n534), .B(new_n535), .Z(new_n536));
  NAND2_X1  g335(.A1(new_n532), .A2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(new_n536), .ZN(new_n538));
  OAI211_X1 g337(.A(new_n525), .B(new_n538), .C1(new_n528), .C2(new_n531), .ZN(new_n539));
  XNOR2_X1  g338(.A(KEYINPUT81), .B(KEYINPUT6), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n537), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  OR2_X1    g340(.A1(new_n539), .A2(new_n540), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n497), .A2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT35), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT34), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n504), .B1(new_n471), .B2(new_n476), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n439), .A2(new_n516), .A3(new_n462), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(G227gat), .ZN(new_n551));
  INV_X1    g350(.A(G233gat), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n547), .B1(new_n550), .B2(new_n554), .ZN(new_n555));
  AOI211_X1 g354(.A(KEYINPUT34), .B(new_n553), .C1(new_n548), .C2(new_n549), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n548), .A2(new_n553), .A3(new_n549), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n558), .A2(KEYINPUT32), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT33), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  XOR2_X1   g360(.A(G15gat), .B(G43gat), .Z(new_n562));
  XNOR2_X1  g361(.A(G71gat), .B(G99gat), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n562), .B(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n559), .A2(new_n561), .A3(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n564), .ZN(new_n566));
  OAI211_X1 g365(.A(new_n558), .B(KEYINPUT32), .C1(new_n560), .C2(new_n566), .ZN(new_n567));
  AND3_X1   g366(.A1(new_n557), .A2(new_n565), .A3(new_n567), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n557), .B1(new_n565), .B2(new_n567), .ZN(new_n569));
  OR2_X1    g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(KEYINPUT31), .B(G50gat), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n405), .A2(new_n406), .A3(new_n465), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n513), .B1(new_n573), .B2(new_n522), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  AOI21_X1  g374(.A(KEYINPUT29), .B1(new_n513), .B2(new_n522), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n575), .B1(new_n478), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n577), .A2(G228gat), .A3(G233gat), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n575), .A2(KEYINPUT82), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT82), .ZN(new_n580));
  AOI22_X1  g379(.A1(new_n574), .A2(new_n580), .B1(G228gat), .B2(G233gat), .ZN(new_n581));
  OAI21_X1  g380(.A(KEYINPUT83), .B1(new_n478), .B2(new_n576), .ZN(new_n582));
  OR3_X1    g381(.A1(new_n478), .A2(new_n576), .A3(KEYINPUT83), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n579), .A2(new_n581), .A3(new_n582), .A4(new_n583), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n572), .B1(new_n578), .B2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(G78gat), .B(G106gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n587), .B(G22gat), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n578), .A2(new_n584), .A3(new_n572), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n586), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n588), .ZN(new_n591));
  INV_X1    g390(.A(new_n589), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n591), .B1(new_n592), .B2(new_n585), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n570), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n545), .A2(new_n546), .A3(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n594), .A2(new_n568), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT75), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n565), .A2(new_n567), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n600), .A2(KEYINPUT74), .ZN(new_n601));
  INV_X1    g400(.A(new_n557), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT74), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n565), .A2(new_n603), .A3(new_n567), .ZN(new_n604));
  AND4_X1   g403(.A1(new_n599), .A2(new_n601), .A3(new_n602), .A4(new_n604), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n557), .B1(new_n600), .B2(KEYINPUT74), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n599), .B1(new_n606), .B2(new_n604), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n598), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT85), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  OAI211_X1 g409(.A(KEYINPUT85), .B(new_n598), .C1(new_n605), .C2(new_n607), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n610), .A2(new_n545), .A3(new_n611), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n597), .B1(new_n612), .B2(KEYINPUT35), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT36), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n568), .A2(new_n614), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n615), .B1(new_n605), .B2(new_n607), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n614), .B1(new_n568), .B2(new_n569), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n617), .A2(KEYINPUT76), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT76), .ZN(new_n619));
  OAI211_X1 g418(.A(new_n619), .B(new_n614), .C1(new_n568), .C2(new_n569), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  AND2_X1   g420(.A1(new_n616), .A2(new_n621), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n543), .A2(new_n494), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT37), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n484), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n482), .A2(KEYINPUT37), .A3(new_n483), .ZN(new_n626));
  AND2_X1   g425(.A1(new_n493), .A2(KEYINPUT38), .ZN(new_n627));
  AND3_X1   g426(.A1(new_n625), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n489), .ZN(new_n629));
  INV_X1    g428(.A(new_n480), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n624), .B1(new_n630), .B2(KEYINPUT84), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT84), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n467), .A2(new_n480), .A3(new_n632), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n629), .B1(new_n631), .B2(new_n633), .ZN(new_n634));
  AOI21_X1  g433(.A(KEYINPUT38), .B1(new_n625), .B2(new_n634), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n623), .B1(new_n628), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n526), .A2(new_n527), .ZN(new_n637));
  OR2_X1    g436(.A1(new_n637), .A2(KEYINPUT39), .ZN(new_n638));
  OAI211_X1 g437(.A(new_n637), .B(KEYINPUT39), .C1(new_n527), .C2(new_n530), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n638), .A2(new_n639), .A3(new_n536), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT40), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n539), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n642), .B1(new_n641), .B2(new_n640), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT30), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n644), .B1(new_n488), .B2(new_n490), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n643), .B1(new_n645), .B2(new_n495), .ZN(new_n646));
  INV_X1    g445(.A(new_n594), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n636), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n594), .B1(new_n497), .B2(new_n544), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n622), .A2(new_n650), .ZN(new_n651));
  OAI211_X1 g450(.A(new_n283), .B(new_n396), .C1(new_n613), .C2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n653), .A2(new_n544), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(G1gat), .ZN(G1324gat));
  INV_X1    g454(.A(new_n497), .ZN(new_n656));
  OR3_X1    g455(.A1(new_n652), .A2(KEYINPUT106), .A3(new_n656), .ZN(new_n657));
  OAI21_X1  g456(.A(KEYINPUT106), .B1(new_n652), .B2(new_n656), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n657), .A2(G8gat), .A3(new_n658), .ZN(new_n659));
  XOR2_X1   g458(.A(KEYINPUT16), .B(G8gat), .Z(new_n660));
  NAND4_X1  g459(.A1(new_n653), .A2(KEYINPUT42), .A3(new_n497), .A4(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n660), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n662), .B1(new_n657), .B2(new_n658), .ZN(new_n663));
  OAI211_X1 g462(.A(new_n659), .B(new_n661), .C1(new_n663), .C2(KEYINPUT42), .ZN(G1325gat));
  INV_X1    g463(.A(KEYINPUT108), .ZN(new_n665));
  AND3_X1   g464(.A1(new_n616), .A2(new_n621), .A3(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n665), .B1(new_n616), .B2(new_n621), .ZN(new_n667));
  OR2_X1    g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n653), .A2(G15gat), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n612), .A2(KEYINPUT35), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n670), .A2(new_n596), .ZN(new_n671));
  INV_X1    g470(.A(new_n651), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n570), .ZN(new_n674));
  NAND4_X1  g473(.A1(new_n673), .A2(new_n674), .A3(new_n283), .A4(new_n396), .ZN(new_n675));
  INV_X1    g474(.A(G15gat), .ZN(new_n676));
  AOI21_X1  g475(.A(KEYINPUT107), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  OAI211_X1 g476(.A(KEYINPUT107), .B(new_n676), .C1(new_n652), .C2(new_n570), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n669), .B1(new_n677), .B2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT109), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  OAI211_X1 g481(.A(KEYINPUT109), .B(new_n669), .C1(new_n677), .C2(new_n679), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(G1326gat));
  NOR2_X1   g483(.A1(new_n652), .A2(new_n647), .ZN(new_n685));
  XOR2_X1   g484(.A(KEYINPUT43), .B(G22gat), .Z(new_n686));
  XNOR2_X1  g485(.A(new_n685), .B(new_n686), .ZN(G1327gat));
  NOR3_X1   g486(.A1(new_n666), .A2(new_n667), .A3(new_n650), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n321), .B1(new_n613), .B2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT44), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  OAI211_X1 g490(.A(KEYINPUT44), .B(new_n321), .C1(new_n613), .C2(new_n651), .ZN(new_n692));
  AND2_X1   g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n365), .ZN(new_n694));
  INV_X1    g493(.A(new_n395), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n279), .A2(new_n280), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n693), .A2(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(G29gat), .B1(new_n700), .B2(new_n543), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n696), .A2(new_n322), .ZN(new_n702));
  OAI211_X1 g501(.A(new_n283), .B(new_n702), .C1(new_n613), .C2(new_n651), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n704), .A2(new_n211), .A3(new_n544), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(KEYINPUT45), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n701), .A2(new_n706), .ZN(G1328gat));
  OAI21_X1  g506(.A(G36gat), .B1(new_n700), .B2(new_n656), .ZN(new_n708));
  NOR3_X1   g507(.A1(new_n703), .A2(G36gat), .A3(new_n656), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(KEYINPUT46), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n708), .A2(new_n710), .ZN(G1329gat));
  INV_X1    g510(.A(KEYINPUT47), .ZN(new_n712));
  NAND4_X1  g511(.A1(new_n691), .A2(new_n668), .A3(new_n692), .A4(new_n699), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(G43gat), .ZN(new_n714));
  NOR3_X1   g513(.A1(new_n703), .A2(G43gat), .A3(new_n570), .ZN(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n712), .B1(new_n714), .B2(new_n716), .ZN(new_n717));
  AOI211_X1 g516(.A(KEYINPUT47), .B(new_n715), .C1(new_n713), .C2(G43gat), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n717), .A2(new_n718), .ZN(G1330gat));
  NAND4_X1  g518(.A1(new_n691), .A2(new_n594), .A3(new_n692), .A4(new_n699), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(G50gat), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n647), .A2(G50gat), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n704), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n721), .A2(KEYINPUT48), .A3(new_n723), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n282), .B1(new_n671), .B2(new_n672), .ZN(new_n725));
  NAND4_X1  g524(.A1(new_n725), .A2(KEYINPUT111), .A3(new_n702), .A4(new_n722), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT111), .ZN(new_n727));
  INV_X1    g526(.A(new_n722), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n727), .B1(new_n703), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n726), .A2(new_n729), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n730), .B1(G50gat), .B2(new_n720), .ZN(new_n731));
  XOR2_X1   g530(.A(KEYINPUT110), .B(KEYINPUT48), .Z(new_n732));
  OAI21_X1  g531(.A(new_n724), .B1(new_n731), .B2(new_n732), .ZN(G1331gat));
  NOR2_X1   g532(.A1(new_n666), .A2(new_n667), .ZN(new_n734));
  INV_X1    g533(.A(new_n650), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n671), .A2(new_n736), .ZN(new_n737));
  NOR3_X1   g536(.A1(new_n366), .A2(new_n697), .A3(new_n695), .ZN(new_n738));
  AND2_X1   g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(new_n544), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g540(.A1(new_n739), .A2(new_n497), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n742), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n743));
  XOR2_X1   g542(.A(KEYINPUT49), .B(G64gat), .Z(new_n744));
  OAI21_X1  g543(.A(new_n743), .B1(new_n742), .B2(new_n744), .ZN(G1333gat));
  INV_X1    g544(.A(G71gat), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n739), .A2(new_n746), .A3(new_n674), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n737), .A2(new_n738), .ZN(new_n748));
  OAI21_X1  g547(.A(G71gat), .B1(new_n748), .B2(new_n734), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT50), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n750), .B(new_n751), .ZN(G1334gat));
  NAND2_X1  g551(.A1(new_n739), .A2(new_n594), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g553(.A1(new_n365), .A2(new_n697), .ZN(new_n755));
  OAI211_X1 g554(.A(new_n321), .B(new_n755), .C1(new_n613), .C2(new_n688), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT112), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT51), .ZN(new_n758));
  NOR3_X1   g557(.A1(new_n756), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  AND2_X1   g558(.A1(new_n756), .A2(new_n758), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND4_X1  g560(.A1(new_n737), .A2(KEYINPUT51), .A3(new_n321), .A4(new_n755), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(new_n757), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  NOR3_X1   g563(.A1(new_n695), .A2(new_n543), .A3(G85gat), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NOR3_X1   g565(.A1(new_n365), .A2(new_n697), .A3(new_n695), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n693), .A2(new_n767), .ZN(new_n768));
  OAI21_X1  g567(.A(G85gat), .B1(new_n768), .B2(new_n543), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n766), .A2(new_n769), .ZN(G1336gat));
  NOR3_X1   g569(.A1(new_n656), .A2(G92gat), .A3(new_n695), .ZN(new_n771));
  INV_X1    g570(.A(new_n771), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n772), .B1(new_n761), .B2(new_n763), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n691), .A2(new_n497), .A3(new_n692), .A4(new_n767), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(G92gat), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT52), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n756), .A2(new_n758), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n778), .ZN(new_n779));
  AOI22_X1  g578(.A1(G92gat), .A2(new_n774), .B1(new_n779), .B2(new_n771), .ZN(new_n780));
  OAI22_X1  g579(.A1(new_n773), .A2(new_n777), .B1(new_n780), .B2(new_n776), .ZN(G1337gat));
  NOR3_X1   g580(.A1(new_n570), .A2(G99gat), .A3(new_n695), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n764), .A2(new_n782), .ZN(new_n783));
  OAI21_X1  g582(.A(G99gat), .B1(new_n768), .B2(new_n734), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(G1338gat));
  NOR3_X1   g584(.A1(new_n647), .A2(G106gat), .A3(new_n695), .ZN(new_n786));
  INV_X1    g585(.A(new_n786), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n787), .B1(new_n761), .B2(new_n763), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n691), .A2(new_n594), .A3(new_n692), .A4(new_n767), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(G106gat), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT53), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  AOI22_X1  g591(.A1(G106gat), .A2(new_n789), .B1(new_n779), .B2(new_n786), .ZN(new_n793));
  OAI22_X1  g592(.A1(new_n788), .A2(new_n792), .B1(new_n793), .B2(new_n791), .ZN(G1339gat));
  INV_X1    g593(.A(new_n595), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n383), .A2(new_n378), .A3(new_n384), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n386), .A2(KEYINPUT54), .A3(new_n796), .ZN(new_n797));
  XOR2_X1   g596(.A(KEYINPUT113), .B(KEYINPUT54), .Z(new_n798));
  AOI21_X1  g597(.A(new_n389), .B1(new_n393), .B2(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n797), .A2(KEYINPUT55), .A3(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT114), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n797), .A2(new_n799), .A3(KEYINPUT114), .A4(KEYINPUT55), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  AND2_X1   g603(.A1(new_n804), .A2(new_n391), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT55), .ZN(new_n806));
  AND3_X1   g605(.A1(new_n383), .A2(new_n378), .A3(new_n384), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT54), .ZN(new_n808));
  NOR3_X1   g607(.A1(new_n807), .A2(new_n393), .A3(new_n808), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n385), .A2(new_n367), .A3(new_n798), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(new_n392), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n806), .B1(new_n809), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n805), .A2(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT115), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n805), .A2(KEYINPUT115), .A3(new_n812), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n815), .A2(new_n697), .A3(new_n816), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n266), .A2(new_n267), .ZN(new_n818));
  XOR2_X1   g617(.A(new_n818), .B(KEYINPUT116), .Z(new_n819));
  AOI21_X1  g618(.A(new_n203), .B1(new_n262), .B2(new_n264), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n272), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n821), .A2(new_n280), .A3(new_n395), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n321), .B1(new_n817), .B2(new_n822), .ZN(new_n823));
  AND2_X1   g622(.A1(new_n821), .A2(new_n280), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n824), .A2(new_n815), .A3(new_n321), .A4(new_n816), .ZN(new_n825));
  INV_X1    g624(.A(new_n825), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n694), .B1(new_n823), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n396), .A2(new_n698), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n795), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n497), .A2(new_n543), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NOR3_X1   g630(.A1(new_n831), .A2(new_n498), .A3(new_n282), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n543), .B1(new_n827), .B2(new_n828), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n610), .A2(new_n611), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n834), .A2(new_n497), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(new_n697), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n832), .B1(new_n498), .B2(new_n838), .ZN(G1340gat));
  NOR3_X1   g638(.A1(new_n831), .A2(new_n499), .A3(new_n695), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n837), .A2(new_n395), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n840), .B1(new_n499), .B2(new_n841), .ZN(G1341gat));
  OAI21_X1  g641(.A(G127gat), .B1(new_n831), .B2(new_n694), .ZN(new_n843));
  OR2_X1    g642(.A1(new_n694), .A2(G127gat), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n843), .B1(new_n836), .B2(new_n844), .ZN(G1342gat));
  OR3_X1    g644(.A1(new_n836), .A2(G134gat), .A3(new_n322), .ZN(new_n846));
  OR2_X1    g645(.A1(new_n846), .A2(KEYINPUT56), .ZN(new_n847));
  OAI21_X1  g646(.A(G134gat), .B1(new_n831), .B2(new_n322), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n846), .A2(KEYINPUT56), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n847), .A2(new_n848), .A3(new_n849), .ZN(G1343gat));
  NAND2_X1  g649(.A1(new_n734), .A2(new_n594), .ZN(new_n851));
  INV_X1    g650(.A(new_n851), .ZN(new_n852));
  AND3_X1   g651(.A1(new_n852), .A2(new_n656), .A3(new_n833), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n282), .A2(G141gat), .ZN(new_n854));
  AND2_X1   g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n734), .A2(new_n830), .ZN(new_n856));
  INV_X1    g655(.A(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT57), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n647), .A2(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT120), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT117), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n862), .B1(new_n809), .B2(new_n811), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n797), .A2(KEYINPUT117), .A3(new_n799), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n863), .A2(new_n806), .A3(new_n864), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n804), .A2(new_n391), .A3(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT118), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n804), .A2(new_n865), .A3(new_n391), .A4(KEYINPUT118), .ZN(new_n869));
  NAND4_X1  g668(.A1(new_n868), .A2(new_n281), .A3(new_n277), .A4(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n321), .B1(new_n870), .B2(new_n822), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n825), .B1(new_n871), .B2(KEYINPUT119), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT119), .ZN(new_n873));
  AOI211_X1 g672(.A(new_n873), .B(new_n321), .C1(new_n870), .C2(new_n822), .ZN(new_n874));
  OAI211_X1 g673(.A(new_n861), .B(new_n694), .C1(new_n872), .C2(new_n874), .ZN(new_n875));
  AND2_X1   g674(.A1(new_n875), .A2(new_n828), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n694), .B1(new_n872), .B2(new_n874), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(KEYINPUT120), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n860), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n827), .A2(new_n828), .ZN(new_n880));
  AOI21_X1  g679(.A(KEYINPUT57), .B1(new_n880), .B2(new_n594), .ZN(new_n881));
  OAI211_X1 g680(.A(new_n697), .B(new_n857), .C1(new_n879), .C2(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n855), .B1(new_n882), .B2(G141gat), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT58), .ZN(new_n884));
  INV_X1    g683(.A(G141gat), .ZN(new_n885));
  INV_X1    g684(.A(new_n878), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n875), .A2(new_n828), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n859), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(new_n881), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n856), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n885), .B1(new_n890), .B2(new_n283), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n853), .A2(new_n854), .ZN(new_n892));
  XOR2_X1   g691(.A(KEYINPUT121), .B(KEYINPUT58), .Z(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  OAI22_X1  g693(.A1(new_n883), .A2(new_n884), .B1(new_n891), .B2(new_n894), .ZN(G1344gat));
  INV_X1    g694(.A(G148gat), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n853), .A2(new_n896), .A3(new_n395), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT59), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(G148gat), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n899), .B1(new_n890), .B2(new_n395), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n880), .A2(new_n594), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(KEYINPUT57), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n594), .A2(new_n858), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT122), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n904), .B1(new_n813), .B2(new_n322), .ZN(new_n905));
  NAND4_X1  g704(.A1(new_n321), .A2(new_n805), .A3(KEYINPUT122), .A4(new_n812), .ZN(new_n906));
  AND3_X1   g705(.A1(new_n905), .A2(new_n906), .A3(new_n824), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n694), .B1(new_n907), .B2(new_n871), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n396), .A2(new_n282), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n903), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(new_n910), .ZN(new_n911));
  NAND4_X1  g710(.A1(new_n902), .A2(new_n395), .A3(new_n857), .A4(new_n911), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n898), .B1(new_n912), .B2(G148gat), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n897), .B1(new_n900), .B2(new_n913), .ZN(G1345gat));
  INV_X1    g713(.A(new_n509), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n853), .A2(new_n915), .A3(new_n365), .ZN(new_n916));
  AND2_X1   g715(.A1(new_n890), .A2(new_n365), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n916), .B1(new_n917), .B2(new_n915), .ZN(G1346gat));
  NOR2_X1   g717(.A1(new_n322), .A2(G162gat), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n853), .A2(new_n919), .ZN(new_n920));
  XNOR2_X1  g719(.A(new_n920), .B(KEYINPUT123), .ZN(new_n921));
  AND2_X1   g720(.A1(new_n890), .A2(new_n321), .ZN(new_n922));
  INV_X1    g721(.A(G162gat), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n921), .B1(new_n922), .B2(new_n923), .ZN(G1347gat));
  AOI21_X1  g723(.A(new_n544), .B1(new_n827), .B2(new_n828), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n834), .A2(new_n656), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  INV_X1    g726(.A(new_n927), .ZN(new_n928));
  AOI21_X1  g727(.A(G169gat), .B1(new_n928), .B2(new_n697), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n656), .A2(new_n544), .ZN(new_n930));
  AND3_X1   g729(.A1(new_n829), .A2(KEYINPUT124), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g730(.A(KEYINPUT124), .B1(new_n829), .B2(new_n930), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  AND2_X1   g732(.A1(new_n283), .A2(G169gat), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n929), .B1(new_n933), .B2(new_n934), .ZN(G1348gat));
  NAND2_X1  g734(.A1(new_n829), .A2(new_n930), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT124), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n829), .A2(KEYINPUT124), .A3(new_n930), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g739(.A(G176gat), .B1(new_n940), .B2(new_n695), .ZN(new_n941));
  OR2_X1    g740(.A1(new_n695), .A2(G176gat), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n941), .B1(new_n927), .B2(new_n942), .ZN(G1349gat));
  AOI21_X1  g742(.A(new_n420), .B1(new_n933), .B2(new_n365), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n928), .A2(new_n430), .A3(new_n365), .ZN(new_n945));
  INV_X1    g744(.A(new_n945), .ZN(new_n946));
  OAI21_X1  g745(.A(KEYINPUT60), .B1(new_n944), .B2(new_n946), .ZN(new_n947));
  OAI21_X1  g746(.A(G183gat), .B1(new_n940), .B2(new_n694), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT60), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n948), .A2(new_n945), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n947), .A2(new_n950), .ZN(G1350gat));
  NAND3_X1  g750(.A1(new_n928), .A2(new_n426), .A3(new_n321), .ZN(new_n952));
  XNOR2_X1  g751(.A(new_n952), .B(KEYINPUT125), .ZN(new_n953));
  OAI21_X1  g752(.A(G190gat), .B1(new_n940), .B2(new_n322), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT61), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  OAI211_X1 g755(.A(KEYINPUT61), .B(G190gat), .C1(new_n940), .C2(new_n322), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n953), .A2(new_n956), .A3(new_n957), .ZN(G1351gat));
  NOR2_X1   g757(.A1(new_n851), .A2(new_n656), .ZN(new_n959));
  AND2_X1   g758(.A1(new_n959), .A2(new_n925), .ZN(new_n960));
  AOI21_X1  g759(.A(G197gat), .B1(new_n960), .B2(new_n697), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n858), .B1(new_n880), .B2(new_n594), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n734), .A2(new_n930), .ZN(new_n963));
  NOR3_X1   g762(.A1(new_n962), .A2(new_n910), .A3(new_n963), .ZN(new_n964));
  AND2_X1   g763(.A1(new_n283), .A2(G197gat), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n961), .B1(new_n964), .B2(new_n965), .ZN(G1352gat));
  NOR2_X1   g765(.A1(new_n695), .A2(G204gat), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n959), .A2(new_n925), .A3(new_n967), .ZN(new_n968));
  XNOR2_X1  g767(.A(new_n968), .B(KEYINPUT62), .ZN(new_n969));
  INV_X1    g768(.A(G204gat), .ZN(new_n970));
  AOI21_X1  g769(.A(new_n970), .B1(new_n964), .B2(new_n395), .ZN(new_n971));
  OAI21_X1  g770(.A(KEYINPUT126), .B1(new_n969), .B2(new_n971), .ZN(new_n972));
  INV_X1    g771(.A(new_n963), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n902), .A2(new_n911), .A3(new_n973), .ZN(new_n974));
  OAI21_X1  g773(.A(G204gat), .B1(new_n974), .B2(new_n695), .ZN(new_n975));
  INV_X1    g774(.A(KEYINPUT126), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n968), .A2(KEYINPUT62), .ZN(new_n977));
  OR2_X1    g776(.A1(new_n968), .A2(KEYINPUT62), .ZN(new_n978));
  NAND4_X1  g777(.A1(new_n975), .A2(new_n976), .A3(new_n977), .A4(new_n978), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n972), .A2(new_n979), .ZN(G1353gat));
  NOR2_X1   g779(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n981));
  NOR4_X1   g780(.A1(new_n962), .A2(new_n694), .A3(new_n910), .A4(new_n963), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n981), .B1(new_n982), .B2(new_n401), .ZN(new_n983));
  INV_X1    g782(.A(new_n981), .ZN(new_n984));
  OAI211_X1 g783(.A(G211gat), .B(new_n984), .C1(new_n974), .C2(new_n694), .ZN(new_n985));
  NAND2_X1  g784(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n986));
  NAND3_X1  g785(.A1(new_n983), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  NAND3_X1  g786(.A1(new_n960), .A2(new_n401), .A3(new_n365), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n987), .A2(new_n988), .ZN(G1354gat));
  OAI21_X1  g788(.A(G218gat), .B1(new_n974), .B2(new_n322), .ZN(new_n990));
  NAND3_X1  g789(.A1(new_n960), .A2(new_n402), .A3(new_n321), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n990), .A2(new_n991), .ZN(G1355gat));
endmodule


