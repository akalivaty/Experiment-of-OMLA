//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 0 1 0 0 0 1 1 0 0 1 1 0 0 1 0 0 1 0 1 1 1 1 0 0 1 1 0 0 0 1 0 0 0 0 0 1 0 1 1 1 1 1 0 1 0 1 0 0 1 0 0 0 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:53 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n450, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n543,
    new_n544, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n593, new_n594, new_n595,
    new_n596, new_n599, new_n601, new_n602, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1105, new_n1106,
    new_n1107;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT64), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT65), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT66), .Z(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT67), .ZN(G217));
  NOR4_X1   g026(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  AND2_X1   g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  OAI21_X1  g035(.A(G137), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g036(.A1(G101), .A2(G2104), .ZN(new_n462));
  AOI21_X1  g037(.A(G2105), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  OAI21_X1  g038(.A(G125), .B1(new_n459), .B2(new_n460), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT68), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  OAI211_X1 g041(.A(KEYINPUT68), .B(G125), .C1(new_n459), .C2(new_n460), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n466), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n463), .B1(new_n469), .B2(G2105), .ZN(G160));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  OAI21_X1  g046(.A(G2104), .B1(new_n471), .B2(G112), .ZN(new_n472));
  INV_X1    g047(.A(G100), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n472), .B1(new_n473), .B2(new_n471), .ZN(new_n474));
  XNOR2_X1  g049(.A(new_n474), .B(KEYINPUT70), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n459), .A2(new_n460), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n476), .A2(new_n471), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n475), .B1(G124), .B2(new_n477), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n476), .A2(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G136), .ZN(new_n480));
  XOR2_X1   g055(.A(new_n480), .B(KEYINPUT69), .Z(new_n481));
  NAND2_X1  g056(.A1(new_n478), .A2(new_n481), .ZN(new_n482));
  XNOR2_X1  g057(.A(new_n482), .B(KEYINPUT71), .ZN(G162));
  NAND2_X1  g058(.A1(KEYINPUT4), .A2(G138), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT3), .ZN(new_n485));
  INV_X1    g060(.A(G2104), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n484), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  AND2_X1   g064(.A1(G102), .A2(G2104), .ZN(new_n490));
  OAI21_X1  g065(.A(new_n471), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(G126), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n492), .B1(new_n487), .B2(new_n488), .ZN(new_n493));
  AND2_X1   g068(.A1(G114), .A2(G2104), .ZN(new_n494));
  OAI21_X1  g069(.A(G2105), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  OAI211_X1 g070(.A(G138), .B(new_n471), .C1(new_n459), .C2(new_n460), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n491), .A2(new_n495), .A3(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  XNOR2_X1  g075(.A(KEYINPUT6), .B(G651), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n501), .A2(G50), .A3(G543), .ZN(new_n502));
  XNOR2_X1  g077(.A(new_n502), .B(KEYINPUT72), .ZN(new_n503));
  OR2_X1    g078(.A1(KEYINPUT5), .A2(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(KEYINPUT5), .A2(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n506), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n506), .A2(new_n501), .ZN(new_n509));
  INV_X1    g084(.A(G88), .ZN(new_n510));
  OAI22_X1  g085(.A1(new_n507), .A2(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n503), .A2(new_n511), .ZN(G166));
  XOR2_X1   g087(.A(KEYINPUT73), .B(KEYINPUT7), .Z(new_n513));
  NAND3_X1  g088(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n514));
  XNOR2_X1  g089(.A(new_n513), .B(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(G51), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n501), .A2(G543), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n506), .A2(G63), .A3(G651), .ZN(new_n519));
  INV_X1    g094(.A(G89), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n519), .B1(new_n509), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n518), .A2(new_n521), .ZN(G168));
  AOI22_X1  g097(.A1(new_n506), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n523), .A2(new_n508), .ZN(new_n524));
  INV_X1    g099(.A(G90), .ZN(new_n525));
  INV_X1    g100(.A(G52), .ZN(new_n526));
  OAI22_X1  g101(.A1(new_n509), .A2(new_n525), .B1(new_n517), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n524), .A2(new_n527), .ZN(G171));
  AND2_X1   g103(.A1(new_n506), .A2(G56), .ZN(new_n529));
  AND2_X1   g104(.A1(G68), .A2(G543), .ZN(new_n530));
  OAI21_X1  g105(.A(G651), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT74), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(G81), .ZN(new_n534));
  INV_X1    g109(.A(G43), .ZN(new_n535));
  OAI22_X1  g110(.A1(new_n509), .A2(new_n534), .B1(new_n517), .B2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n533), .A2(new_n537), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n531), .A2(new_n532), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G860), .ZN(G153));
  NAND4_X1  g116(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g117(.A1(G1), .A2(G3), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT8), .ZN(new_n544));
  NAND4_X1  g119(.A1(G319), .A2(G483), .A3(G661), .A4(new_n544), .ZN(G188));
  INV_X1    g120(.A(new_n517), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G53), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT9), .ZN(new_n548));
  XNOR2_X1  g123(.A(KEYINPUT75), .B(G65), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n506), .A2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(new_n551));
  AND2_X1   g126(.A1(G78), .A2(G543), .ZN(new_n552));
  OAI21_X1  g127(.A(G651), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(G91), .ZN(new_n554));
  OAI211_X1 g129(.A(new_n548), .B(new_n553), .C1(new_n554), .C2(new_n509), .ZN(G299));
  XNOR2_X1  g130(.A(G171), .B(KEYINPUT76), .ZN(G301));
  INV_X1    g131(.A(G168), .ZN(G286));
  INV_X1    g132(.A(G166), .ZN(G303));
  NAND3_X1  g133(.A1(new_n506), .A2(new_n501), .A3(G87), .ZN(new_n559));
  INV_X1    g134(.A(G49), .ZN(new_n560));
  OAI21_X1  g135(.A(G651), .B1(new_n506), .B2(G74), .ZN(new_n561));
  OAI221_X1 g136(.A(new_n559), .B1(new_n517), .B2(new_n560), .C1(new_n561), .C2(KEYINPUT77), .ZN(new_n562));
  AND2_X1   g137(.A1(new_n561), .A2(KEYINPUT77), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(new_n564), .ZN(G288));
  AOI22_X1  g140(.A1(new_n506), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n566));
  OR2_X1    g141(.A1(new_n566), .A2(new_n508), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n506), .A2(new_n501), .A3(G86), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n501), .A2(G48), .A3(G543), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT78), .ZN(G305));
  INV_X1    g146(.A(G85), .ZN(new_n572));
  INV_X1    g147(.A(G47), .ZN(new_n573));
  OAI22_X1  g148(.A1(new_n509), .A2(new_n572), .B1(new_n517), .B2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(KEYINPUT79), .ZN(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n575), .A2(KEYINPUT79), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n506), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n579));
  OAI22_X1  g154(.A1(new_n577), .A2(new_n578), .B1(new_n508), .B2(new_n579), .ZN(G290));
  INV_X1    g155(.A(G868), .ZN(new_n581));
  NOR2_X1   g156(.A1(G301), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n506), .A2(new_n501), .A3(G92), .ZN(new_n583));
  XOR2_X1   g158(.A(new_n583), .B(KEYINPUT10), .Z(new_n584));
  NAND2_X1  g159(.A1(new_n506), .A2(G66), .ZN(new_n585));
  NAND2_X1  g160(.A1(G79), .A2(G543), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n508), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n587), .B1(G54), .B2(new_n546), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n584), .A2(new_n588), .ZN(new_n589));
  XNOR2_X1  g164(.A(new_n589), .B(KEYINPUT80), .ZN(new_n590));
  AOI21_X1  g165(.A(new_n582), .B1(new_n590), .B2(new_n581), .ZN(G321));
  XOR2_X1   g166(.A(G321), .B(KEYINPUT81), .Z(G284));
  NAND2_X1  g167(.A1(G299), .A2(new_n581), .ZN(new_n593));
  NAND3_X1  g168(.A1(G286), .A2(KEYINPUT82), .A3(G868), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT82), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n595), .B1(G168), .B2(new_n581), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n593), .A2(new_n594), .A3(new_n596), .ZN(G297));
  NAND3_X1  g172(.A1(new_n593), .A2(new_n594), .A3(new_n596), .ZN(G280));
  INV_X1    g173(.A(G559), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n590), .B1(new_n599), .B2(G860), .ZN(G148));
  OAI21_X1  g175(.A(new_n581), .B1(new_n538), .B2(new_n539), .ZN(new_n601));
  AND2_X1   g176(.A1(new_n590), .A2(new_n599), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n602), .B2(new_n581), .ZN(G323));
  XNOR2_X1  g178(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g179(.A1(new_n479), .A2(G2104), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n605), .B(KEYINPUT12), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(KEYINPUT13), .ZN(new_n607));
  INV_X1    g182(.A(new_n607), .ZN(new_n608));
  OR2_X1    g183(.A1(new_n608), .A2(G2100), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(G2100), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n479), .A2(G135), .ZN(new_n611));
  NOR2_X1   g186(.A1(G99), .A2(G2105), .ZN(new_n612));
  OAI21_X1  g187(.A(G2104), .B1(new_n471), .B2(G111), .ZN(new_n613));
  AND3_X1   g188(.A1(new_n477), .A2(KEYINPUT83), .A3(G123), .ZN(new_n614));
  AOI21_X1  g189(.A(KEYINPUT83), .B1(new_n477), .B2(G123), .ZN(new_n615));
  OAI221_X1 g190(.A(new_n611), .B1(new_n612), .B2(new_n613), .C1(new_n614), .C2(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(G2096), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n616), .B(new_n617), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n609), .A2(new_n610), .A3(new_n618), .ZN(new_n619));
  XOR2_X1   g194(.A(new_n619), .B(KEYINPUT84), .Z(G156));
  XOR2_X1   g195(.A(KEYINPUT15), .B(G2435), .Z(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(G2438), .ZN(new_n622));
  XNOR2_X1  g197(.A(G2427), .B(G2430), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT86), .ZN(new_n624));
  OR2_X1    g199(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n622), .A2(new_n624), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n625), .A2(KEYINPUT14), .A3(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(G1341), .B(G1348), .Z(new_n628));
  XNOR2_X1  g203(.A(KEYINPUT85), .B(KEYINPUT16), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n627), .B(new_n630), .ZN(new_n631));
  INV_X1    g206(.A(new_n631), .ZN(new_n632));
  XOR2_X1   g207(.A(G2443), .B(G2446), .Z(new_n633));
  XNOR2_X1  g208(.A(G2451), .B(G2454), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  INV_X1    g210(.A(new_n635), .ZN(new_n636));
  OAI21_X1  g211(.A(G14), .B1(new_n632), .B2(new_n636), .ZN(new_n637));
  AOI21_X1  g212(.A(new_n637), .B1(new_n636), .B2(new_n632), .ZN(G401));
  XOR2_X1   g213(.A(G2072), .B(G2078), .Z(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(KEYINPUT17), .Z(new_n640));
  XOR2_X1   g215(.A(G2084), .B(G2090), .Z(new_n641));
  XNOR2_X1  g216(.A(G2067), .B(G2678), .ZN(new_n642));
  OAI21_X1  g217(.A(new_n640), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n641), .A2(new_n642), .ZN(new_n644));
  INV_X1    g219(.A(new_n641), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n645), .A2(new_n639), .ZN(new_n646));
  OAI211_X1 g221(.A(new_n643), .B(new_n644), .C1(new_n642), .C2(new_n646), .ZN(new_n647));
  NOR2_X1   g222(.A1(new_n644), .A2(new_n639), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT18), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(new_n617), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2100), .ZN(G227));
  XOR2_X1   g227(.A(G1971), .B(G1976), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT87), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT19), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1956), .B(G2474), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1961), .B(G1966), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT20), .ZN(new_n660));
  AND2_X1   g235(.A1(new_n656), .A2(new_n657), .ZN(new_n661));
  NOR3_X1   g236(.A1(new_n655), .A2(new_n658), .A3(new_n661), .ZN(new_n662));
  AOI21_X1  g237(.A(new_n662), .B1(new_n655), .B2(new_n661), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(KEYINPUT88), .B(G1986), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1991), .B(G1996), .ZN(new_n669));
  INV_X1    g244(.A(G1981), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n668), .B(new_n671), .ZN(G229));
  INV_X1    g247(.A(G16), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n564), .A2(new_n673), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n674), .B1(new_n673), .B2(G23), .ZN(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT33), .B(G1976), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NOR2_X1   g252(.A1(G166), .A2(new_n673), .ZN(new_n678));
  AOI21_X1  g253(.A(new_n678), .B1(new_n673), .B2(G22), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n677), .B1(new_n680), .B2(G1971), .ZN(new_n681));
  OR2_X1    g256(.A1(G6), .A2(G16), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n682), .B1(G305), .B2(new_n673), .ZN(new_n683));
  XOR2_X1   g258(.A(KEYINPUT32), .B(G1981), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT89), .ZN(new_n685));
  OR2_X1    g260(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n683), .A2(new_n685), .ZN(new_n687));
  INV_X1    g262(.A(G1971), .ZN(new_n688));
  AOI22_X1  g263(.A1(new_n675), .A2(new_n676), .B1(new_n679), .B2(new_n688), .ZN(new_n689));
  NAND4_X1  g264(.A1(new_n681), .A2(new_n686), .A3(new_n687), .A4(new_n689), .ZN(new_n690));
  OR2_X1    g265(.A1(new_n690), .A2(KEYINPUT34), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n690), .A2(KEYINPUT34), .ZN(new_n692));
  OR2_X1    g267(.A1(G16), .A2(G24), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n693), .B1(G290), .B2(new_n673), .ZN(new_n694));
  INV_X1    g269(.A(G1986), .ZN(new_n695));
  AND2_X1   g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n694), .A2(new_n695), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n479), .A2(G131), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n477), .A2(G119), .ZN(new_n699));
  NOR2_X1   g274(.A1(G95), .A2(G2105), .ZN(new_n700));
  OAI21_X1  g275(.A(G2104), .B1(new_n471), .B2(G107), .ZN(new_n701));
  OAI211_X1 g276(.A(new_n698), .B(new_n699), .C1(new_n700), .C2(new_n701), .ZN(new_n702));
  MUX2_X1   g277(.A(G25), .B(new_n702), .S(G29), .Z(new_n703));
  XOR2_X1   g278(.A(KEYINPUT35), .B(G1991), .Z(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n703), .B(new_n705), .ZN(new_n706));
  NOR3_X1   g281(.A1(new_n696), .A2(new_n697), .A3(new_n706), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n691), .A2(new_n692), .A3(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT36), .ZN(new_n709));
  XOR2_X1   g284(.A(KEYINPUT31), .B(G11), .Z(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT97), .B(G28), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n711), .A2(KEYINPUT30), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n712), .A2(G29), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n711), .A2(KEYINPUT30), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n710), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(G29), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n715), .B1(new_n616), .B2(new_n716), .ZN(new_n717));
  NOR2_X1   g292(.A1(G168), .A2(new_n673), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(new_n673), .B2(G21), .ZN(new_n719));
  XNOR2_X1  g294(.A(KEYINPUT96), .B(G1966), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n717), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n673), .A2(G5), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(G171), .B2(new_n673), .ZN(new_n723));
  OAI221_X1 g298(.A(new_n721), .B1(G1961), .B2(new_n723), .C1(new_n719), .C2(new_n720), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n716), .A2(G32), .ZN(new_n725));
  NAND3_X1  g300(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n726));
  XOR2_X1   g301(.A(new_n726), .B(KEYINPUT26), .Z(new_n727));
  NAND2_X1  g302(.A1(new_n479), .A2(G141), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n477), .A2(G129), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n471), .A2(G105), .A3(G2104), .ZN(new_n730));
  AND4_X1   g305(.A1(new_n727), .A2(new_n728), .A3(new_n729), .A4(new_n730), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n725), .B1(new_n731), .B2(new_n716), .ZN(new_n732));
  XNOR2_X1  g307(.A(KEYINPUT27), .B(G1996), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n732), .B(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n716), .A2(G27), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(G164), .B2(new_n716), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n734), .B1(G2078), .B2(new_n736), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n724), .A2(new_n737), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n716), .B1(KEYINPUT24), .B2(G34), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(KEYINPUT24), .B2(G34), .ZN(new_n740));
  INV_X1    g315(.A(G160), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n740), .B1(new_n741), .B2(G29), .ZN(new_n742));
  INV_X1    g317(.A(G2084), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n742), .A2(new_n743), .ZN(new_n745));
  NOR2_X1   g320(.A1(G29), .A2(G33), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT93), .Z(new_n747));
  XNOR2_X1  g322(.A(KEYINPUT94), .B(KEYINPUT25), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n471), .A2(G103), .A3(G2104), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n487), .A2(new_n488), .ZN(new_n751));
  AOI22_X1  g326(.A1(new_n751), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n752));
  NOR3_X1   g327(.A1(new_n752), .A2(KEYINPUT95), .A3(new_n471), .ZN(new_n753));
  AOI211_X1 g328(.A(new_n750), .B(new_n753), .C1(G139), .C2(new_n479), .ZN(new_n754));
  OAI21_X1  g329(.A(KEYINPUT95), .B1(new_n752), .B2(new_n471), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n747), .B1(new_n756), .B2(new_n716), .ZN(new_n757));
  INV_X1    g332(.A(G2072), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n745), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  AOI211_X1 g334(.A(new_n744), .B(new_n759), .C1(new_n758), .C2(new_n757), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n723), .A2(KEYINPUT98), .A3(G1961), .ZN(new_n761));
  AOI21_X1  g336(.A(KEYINPUT98), .B1(new_n723), .B2(G1961), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(G2078), .B2(new_n736), .ZN(new_n763));
  NAND4_X1  g338(.A1(new_n738), .A2(new_n760), .A3(new_n761), .A4(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(KEYINPUT99), .ZN(new_n765));
  OR2_X1    g340(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n716), .A2(G35), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT100), .Z(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G162), .B2(new_n716), .ZN(new_n769));
  XOR2_X1   g344(.A(KEYINPUT29), .B(G2090), .Z(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n673), .A2(G4), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(new_n590), .B2(new_n673), .ZN(new_n773));
  XOR2_X1   g348(.A(KEYINPUT90), .B(G1348), .Z(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n673), .A2(G19), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(new_n540), .B2(new_n673), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(G1341), .Z(new_n778));
  NAND2_X1  g353(.A1(new_n673), .A2(G20), .ZN(new_n779));
  XOR2_X1   g354(.A(new_n779), .B(KEYINPUT23), .Z(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(G299), .B2(G16), .ZN(new_n781));
  INV_X1    g356(.A(G1956), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n479), .A2(G140), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n477), .A2(G128), .ZN(new_n785));
  NOR2_X1   g360(.A1(G104), .A2(G2105), .ZN(new_n786));
  OAI21_X1  g361(.A(G2104), .B1(new_n471), .B2(G116), .ZN(new_n787));
  OAI211_X1 g362(.A(new_n784), .B(new_n785), .C1(new_n786), .C2(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n788), .A2(G29), .ZN(new_n789));
  XOR2_X1   g364(.A(KEYINPUT91), .B(KEYINPUT28), .Z(new_n790));
  NAND2_X1  g365(.A1(new_n716), .A2(G26), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n789), .A2(new_n792), .ZN(new_n793));
  XOR2_X1   g368(.A(KEYINPUT92), .B(G2067), .Z(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n783), .A2(new_n795), .ZN(new_n796));
  NAND4_X1  g371(.A1(new_n771), .A2(new_n775), .A3(new_n778), .A4(new_n796), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(new_n764), .B2(new_n765), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n709), .A2(new_n766), .A3(new_n798), .ZN(G150));
  INV_X1    g374(.A(G150), .ZN(G311));
  NAND2_X1  g375(.A1(new_n506), .A2(G67), .ZN(new_n801));
  NAND2_X1  g376(.A1(G80), .A2(G543), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n508), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(KEYINPUT101), .ZN(new_n804));
  OR2_X1    g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n803), .A2(new_n804), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n546), .A2(G55), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n506), .A2(new_n501), .A3(G93), .ZN(new_n808));
  NAND4_X1  g383(.A1(new_n805), .A2(new_n806), .A3(new_n807), .A4(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n809), .A2(G860), .ZN(new_n810));
  XOR2_X1   g385(.A(new_n810), .B(KEYINPUT37), .Z(new_n811));
  AOI21_X1  g386(.A(new_n809), .B1(new_n540), .B2(KEYINPUT102), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n540), .A2(KEYINPUT102), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n812), .B(new_n813), .Z(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT38), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n590), .A2(G559), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT39), .ZN(new_n818));
  OR2_X1    g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  AOI21_X1  g394(.A(G860), .B1(new_n817), .B2(new_n818), .ZN(new_n820));
  AND3_X1   g395(.A1(new_n819), .A2(KEYINPUT103), .A3(new_n820), .ZN(new_n821));
  AOI21_X1  g396(.A(KEYINPUT103), .B1(new_n819), .B2(new_n820), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n811), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n823), .A2(KEYINPUT104), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT104), .ZN(new_n825));
  OAI211_X1 g400(.A(new_n825), .B(new_n811), .C1(new_n821), .C2(new_n822), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n824), .A2(new_n826), .ZN(G145));
  XNOR2_X1  g402(.A(G164), .B(new_n788), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n756), .B(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n702), .B(KEYINPUT105), .ZN(new_n830));
  XOR2_X1   g405(.A(new_n830), .B(new_n606), .Z(new_n831));
  XNOR2_X1  g406(.A(new_n829), .B(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n479), .A2(G142), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n477), .A2(G130), .ZN(new_n834));
  NOR2_X1   g409(.A1(G106), .A2(G2105), .ZN(new_n835));
  OAI21_X1  g410(.A(G2104), .B1(new_n471), .B2(G118), .ZN(new_n836));
  OAI211_X1 g411(.A(new_n833), .B(new_n834), .C1(new_n835), .C2(new_n836), .ZN(new_n837));
  XOR2_X1   g412(.A(new_n731), .B(new_n837), .Z(new_n838));
  XNOR2_X1  g413(.A(new_n832), .B(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n616), .B(G160), .ZN(new_n840));
  XNOR2_X1  g415(.A(G162), .B(new_n840), .ZN(new_n841));
  XOR2_X1   g416(.A(new_n841), .B(KEYINPUT107), .Z(new_n842));
  NAND2_X1  g417(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT108), .ZN(new_n844));
  INV_X1    g419(.A(G37), .ZN(new_n845));
  AND2_X1   g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(new_n841), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n839), .A2(new_n847), .ZN(new_n848));
  XOR2_X1   g423(.A(new_n848), .B(KEYINPUT106), .Z(new_n849));
  AOI21_X1  g424(.A(KEYINPUT40), .B1(new_n846), .B2(new_n849), .ZN(new_n850));
  AND4_X1   g425(.A1(KEYINPUT40), .A2(new_n849), .A3(new_n845), .A4(new_n844), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n850), .A2(new_n851), .ZN(G395));
  NAND2_X1  g427(.A1(new_n809), .A2(new_n581), .ZN(new_n853));
  INV_X1    g428(.A(new_n589), .ZN(new_n854));
  XNOR2_X1  g429(.A(G299), .B(new_n854), .ZN(new_n855));
  XOR2_X1   g430(.A(new_n855), .B(KEYINPUT41), .Z(new_n856));
  XNOR2_X1  g431(.A(new_n814), .B(new_n602), .ZN(new_n857));
  MUX2_X1   g432(.A(new_n855), .B(new_n856), .S(new_n857), .Z(new_n858));
  XOR2_X1   g433(.A(G305), .B(G290), .Z(new_n859));
  XNOR2_X1  g434(.A(new_n564), .B(G166), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n859), .B(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n861), .A2(KEYINPUT109), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(KEYINPUT42), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n858), .B(new_n863), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n853), .B1(new_n864), .B2(new_n581), .ZN(G295));
  OAI21_X1  g440(.A(new_n853), .B1(new_n864), .B2(new_n581), .ZN(G331));
  INV_X1    g441(.A(KEYINPUT110), .ZN(new_n867));
  INV_X1    g442(.A(G171), .ZN(new_n868));
  NAND2_X1  g443(.A1(G286), .A2(new_n868), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n869), .B1(G286), .B2(G301), .ZN(new_n870));
  XOR2_X1   g445(.A(new_n814), .B(new_n870), .Z(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(new_n855), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n814), .B(new_n870), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n873), .A2(new_n856), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n867), .B1(new_n875), .B2(new_n861), .ZN(new_n876));
  AOI21_X1  g451(.A(G37), .B1(new_n875), .B2(new_n861), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT43), .ZN(new_n878));
  INV_X1    g453(.A(new_n861), .ZN(new_n879));
  NAND4_X1  g454(.A1(new_n872), .A2(KEYINPUT110), .A3(new_n879), .A4(new_n874), .ZN(new_n880));
  NAND4_X1  g455(.A1(new_n876), .A2(new_n877), .A3(new_n878), .A4(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n881), .A2(KEYINPUT111), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(KEYINPUT44), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n876), .A2(new_n877), .A3(new_n880), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n884), .A2(KEYINPUT43), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n885), .A2(new_n881), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n883), .A2(new_n886), .ZN(new_n887));
  NAND4_X1  g462(.A1(new_n882), .A2(new_n885), .A3(KEYINPUT44), .A4(new_n881), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(G397));
  XNOR2_X1  g464(.A(new_n731), .B(G1996), .ZN(new_n890));
  XOR2_X1   g465(.A(new_n788), .B(G2067), .Z(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  OR2_X1    g467(.A1(new_n702), .A2(new_n705), .ZN(new_n893));
  OAI22_X1  g468(.A1(new_n892), .A2(new_n893), .B1(G2067), .B2(new_n788), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n469), .A2(G2105), .ZN(new_n895));
  INV_X1    g470(.A(new_n463), .ZN(new_n896));
  AND4_X1   g471(.A1(KEYINPUT112), .A2(new_n895), .A3(G40), .A4(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(KEYINPUT112), .B1(G160), .B2(G40), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(G1384), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n499), .A2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT45), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n899), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n894), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n702), .A2(new_n705), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n890), .A2(new_n891), .A3(new_n893), .A4(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(new_n904), .ZN(new_n908));
  NOR2_X1   g483(.A1(G290), .A2(G1986), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n904), .A2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n908), .B1(new_n911), .B2(KEYINPUT48), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT48), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n910), .A2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(G1996), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n904), .A2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT46), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n891), .A2(new_n731), .ZN(new_n918));
  AOI22_X1  g493(.A1(new_n916), .A2(new_n917), .B1(new_n904), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n919), .B1(new_n917), .B2(new_n916), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT47), .ZN(new_n921));
  OAI221_X1 g496(.A(new_n905), .B1(new_n912), .B2(new_n914), .C1(new_n920), .C2(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n922), .B1(new_n921), .B2(new_n920), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT127), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n499), .A2(KEYINPUT45), .A3(new_n900), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(KEYINPUT113), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT113), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n499), .A2(new_n927), .A3(KEYINPUT45), .A4(new_n900), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n926), .A2(new_n903), .A3(new_n928), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n688), .B1(new_n899), .B2(new_n929), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n895), .A2(G40), .A3(new_n896), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT112), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(G160), .A2(KEYINPUT112), .A3(G40), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(G2090), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT50), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n937), .B1(new_n499), .B2(new_n900), .ZN(new_n938));
  INV_X1    g513(.A(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n499), .A2(new_n937), .A3(new_n900), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n935), .A2(new_n936), .A3(new_n939), .A4(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n930), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(G8), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT116), .ZN(new_n944));
  OAI21_X1  g519(.A(G8), .B1(new_n503), .B2(new_n511), .ZN(new_n945));
  XNOR2_X1  g520(.A(new_n945), .B(KEYINPUT55), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n943), .A2(new_n944), .A3(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(G8), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n948), .B1(new_n930), .B2(new_n941), .ZN(new_n949));
  INV_X1    g524(.A(new_n946), .ZN(new_n950));
  OAI21_X1  g525(.A(KEYINPUT116), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n940), .A2(KEYINPUT114), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n952), .A2(new_n938), .ZN(new_n953));
  AND2_X1   g528(.A1(new_n499), .A2(new_n900), .ZN(new_n954));
  NOR3_X1   g529(.A1(new_n954), .A2(KEYINPUT114), .A3(new_n937), .ZN(new_n955));
  OAI211_X1 g530(.A(new_n936), .B(new_n935), .C1(new_n953), .C2(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n948), .B1(new_n930), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(new_n950), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n954), .B1(new_n897), .B2(new_n898), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n564), .A2(G1976), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n959), .A2(G8), .A3(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(KEYINPUT52), .ZN(new_n962));
  XNOR2_X1  g537(.A(KEYINPUT115), .B(G86), .ZN(new_n963));
  OAI221_X1 g538(.A(new_n569), .B1(new_n509), .B2(new_n963), .C1(new_n566), .C2(new_n508), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(G1981), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n567), .A2(new_n568), .A3(new_n569), .A4(new_n670), .ZN(new_n966));
  AND3_X1   g541(.A1(new_n965), .A2(new_n966), .A3(KEYINPUT49), .ZN(new_n967));
  AOI21_X1  g542(.A(KEYINPUT49), .B1(new_n965), .B2(new_n966), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n969), .A2(G8), .A3(new_n959), .ZN(new_n970));
  INV_X1    g545(.A(G1976), .ZN(new_n971));
  AOI21_X1  g546(.A(KEYINPUT52), .B1(G288), .B2(new_n971), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n972), .A2(new_n959), .A3(G8), .A4(new_n960), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n962), .A2(new_n970), .A3(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(new_n974), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n947), .A2(new_n951), .A3(new_n958), .A4(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(KEYINPUT125), .ZN(new_n977));
  AOI211_X1 g552(.A(new_n948), .B(new_n946), .C1(new_n930), .C2(new_n956), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n978), .A2(new_n974), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT125), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n979), .A2(new_n980), .A3(new_n947), .A4(new_n951), .ZN(new_n981));
  AND2_X1   g556(.A1(new_n977), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(G1961), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n935), .B1(new_n953), .B2(new_n955), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n903), .A2(new_n925), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n899), .A2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT53), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n987), .A2(G2078), .ZN(new_n988));
  AOI22_X1  g563(.A1(new_n983), .A2(new_n984), .B1(new_n986), .B2(new_n988), .ZN(new_n989));
  AOI21_X1  g564(.A(KEYINPUT45), .B1(new_n499), .B2(new_n900), .ZN(new_n990));
  AND3_X1   g565(.A1(new_n499), .A2(KEYINPUT45), .A3(new_n900), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n990), .B1(new_n991), .B2(new_n927), .ZN(new_n992));
  INV_X1    g567(.A(G2078), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n935), .A2(new_n992), .A3(new_n993), .A4(new_n926), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(new_n987), .ZN(new_n995));
  AOI21_X1  g570(.A(G301), .B1(new_n989), .B2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT123), .ZN(new_n997));
  XOR2_X1   g572(.A(KEYINPUT117), .B(G2084), .Z(new_n998));
  OAI211_X1 g573(.A(new_n935), .B(new_n998), .C1(new_n953), .C2(new_n955), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n720), .B1(new_n899), .B2(new_n985), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n999), .A2(new_n1000), .A3(G168), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(G8), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(KEYINPUT51), .ZN(new_n1003));
  AOI21_X1  g578(.A(G168), .B1(new_n999), .B2(new_n1000), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT51), .ZN(new_n1005));
  OAI211_X1 g580(.A(G8), .B(new_n1001), .C1(new_n1004), .C2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n997), .B1(new_n1003), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1003), .A2(new_n1006), .A3(new_n997), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1008), .A2(KEYINPUT62), .A3(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT62), .ZN(new_n1011));
  AND3_X1   g586(.A1(new_n1003), .A2(new_n1006), .A3(new_n997), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1011), .B1(new_n1012), .B2(new_n1007), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n982), .A2(new_n996), .A3(new_n1010), .A4(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT63), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n999), .A2(new_n1000), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1016), .A2(G8), .A3(G168), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1015), .B1(new_n976), .B2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(KEYINPUT118), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT118), .ZN(new_n1020));
  OAI211_X1 g595(.A(new_n1020), .B(new_n1015), .C1(new_n976), .C2(new_n1017), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1017), .A2(new_n1015), .ZN(new_n1022));
  OAI211_X1 g597(.A(new_n979), .B(new_n1022), .C1(new_n957), .C2(new_n950), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1019), .A2(new_n1021), .A3(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n959), .A2(G8), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n970), .A2(new_n971), .A3(new_n564), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1025), .B1(new_n1026), .B2(new_n966), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1027), .B1(new_n978), .B2(new_n975), .ZN(new_n1028));
  AND3_X1   g603(.A1(new_n1014), .A2(new_n1024), .A3(new_n1028), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1012), .A2(new_n1007), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT124), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n984), .A2(new_n983), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n986), .A2(new_n988), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1032), .A2(new_n995), .A3(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(G301), .ZN(new_n1035));
  INV_X1    g610(.A(new_n929), .ZN(new_n1036));
  NOR3_X1   g611(.A1(new_n931), .A2(new_n987), .A3(G2078), .ZN(new_n1037));
  AOI22_X1  g612(.A1(new_n994), .A2(new_n987), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1035), .B1(new_n984), .B2(new_n983), .ZN(new_n1039));
  AOI22_X1  g614(.A1(new_n1034), .A2(new_n1035), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1031), .B1(new_n1040), .B2(KEYINPUT54), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT54), .ZN(new_n1042));
  AND2_X1   g617(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1043));
  OAI211_X1 g618(.A(KEYINPUT124), .B(new_n1042), .C1(new_n996), .C2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1041), .A2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g620(.A(KEYINPUT54), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n868), .B1(new_n1038), .B2(new_n1032), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1048), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1030), .A2(new_n1045), .A3(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n977), .A2(new_n981), .ZN(new_n1051));
  OAI21_X1  g626(.A(KEYINPUT126), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  NOR3_X1   g627(.A1(new_n1012), .A2(new_n1007), .A3(new_n1048), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT126), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n982), .A2(new_n1053), .A3(new_n1054), .A4(new_n1045), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n899), .A2(new_n929), .ZN(new_n1056));
  XNOR2_X1  g631(.A(KEYINPUT56), .B(G2072), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n935), .A2(new_n939), .A3(new_n940), .ZN(new_n1059));
  AND3_X1   g634(.A1(new_n1059), .A2(KEYINPUT119), .A3(new_n782), .ZN(new_n1060));
  AOI21_X1  g635(.A(KEYINPUT119), .B1(new_n1059), .B2(new_n782), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1058), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  XNOR2_X1  g637(.A(G299), .B(KEYINPUT57), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n959), .A2(G2067), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1065), .B1(new_n774), .B2(new_n984), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1064), .B1(new_n589), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1063), .ZN(new_n1068));
  OAI211_X1 g643(.A(new_n1068), .B(new_n1058), .C1(new_n1060), .C2(new_n1061), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(KEYINPUT120), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT120), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1067), .A2(new_n1072), .A3(new_n1069), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT61), .ZN(new_n1074));
  AND3_X1   g649(.A1(new_n1064), .A2(new_n1069), .A3(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1074), .B1(new_n1064), .B2(new_n1069), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  AND2_X1   g652(.A1(new_n540), .A2(KEYINPUT122), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1056), .A2(new_n915), .ZN(new_n1079));
  XOR2_X1   g654(.A(KEYINPUT58), .B(G1341), .Z(new_n1080));
  NAND2_X1  g655(.A1(new_n959), .A2(new_n1080), .ZN(new_n1081));
  AND3_X1   g656(.A1(new_n1079), .A2(KEYINPUT121), .A3(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(KEYINPUT121), .B1(new_n1079), .B2(new_n1081), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1078), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT59), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1066), .A2(new_n589), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1087), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1066), .A2(new_n589), .ZN(new_n1089));
  OAI21_X1  g664(.A(KEYINPUT60), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  OAI211_X1 g665(.A(KEYINPUT59), .B(new_n1078), .C1(new_n1082), .C2(new_n1083), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1066), .ZN(new_n1092));
  OR3_X1    g667(.A1(new_n1092), .A2(KEYINPUT60), .A3(new_n589), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1086), .A2(new_n1090), .A3(new_n1091), .A4(new_n1093), .ZN(new_n1094));
  OAI211_X1 g669(.A(new_n1071), .B(new_n1073), .C1(new_n1077), .C2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1052), .A2(new_n1055), .A3(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1029), .A2(new_n1096), .ZN(new_n1097));
  XNOR2_X1  g672(.A(G290), .B(G1986), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n904), .B1(new_n1098), .B2(new_n907), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n924), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1099), .ZN(new_n1101));
  AOI211_X1 g676(.A(KEYINPUT127), .B(new_n1101), .C1(new_n1029), .C2(new_n1096), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n923), .B1(new_n1100), .B2(new_n1102), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g678(.A1(new_n846), .A2(new_n849), .ZN(new_n1105));
  INV_X1    g679(.A(G319), .ZN(new_n1106));
  NOR4_X1   g680(.A1(G229), .A2(new_n1106), .A3(G401), .A4(G227), .ZN(new_n1107));
  NAND3_X1  g681(.A1(new_n1105), .A2(new_n886), .A3(new_n1107), .ZN(G225));
  INV_X1    g682(.A(G225), .ZN(G308));
endmodule


