//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 1 0 0 0 1 1 1 1 1 1 1 0 0 0 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 0 0 1 0 1 1 1 1 0 1 0 0 1 1 1 1 1 1 1 1 0 0 1 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:14 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n749, new_n751, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n790, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n990, new_n991, new_n992, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1013, new_n1014, new_n1015, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  NAND2_X1  g004(.A1(KEYINPUT81), .A2(KEYINPUT25), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G140), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G125), .ZN(new_n194));
  INV_X1    g008(.A(G125), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G140), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n194), .A2(new_n196), .A3(KEYINPUT76), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n193), .A2(G125), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT76), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n197), .A2(new_n200), .A3(KEYINPUT16), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n195), .A2(G140), .ZN(new_n202));
  OR2_X1    g016(.A1(new_n202), .A2(KEYINPUT16), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n201), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G146), .ZN(new_n205));
  NAND2_X1  g019(.A1(KEYINPUT23), .A2(G119), .ZN(new_n206));
  OAI21_X1  g020(.A(KEYINPUT74), .B1(new_n206), .B2(G128), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT74), .ZN(new_n208));
  INV_X1    g022(.A(G128), .ZN(new_n209));
  NAND4_X1  g023(.A1(new_n208), .A2(new_n209), .A3(KEYINPUT23), .A4(G119), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n207), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G110), .ZN(new_n212));
  OAI211_X1 g026(.A(KEYINPUT75), .B(KEYINPUT23), .C1(new_n209), .C2(G119), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n209), .A2(G119), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G119), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G128), .ZN(new_n217));
  AOI21_X1  g031(.A(KEYINPUT75), .B1(new_n217), .B2(KEYINPUT23), .ZN(new_n218));
  OAI211_X1 g032(.A(new_n211), .B(new_n212), .C1(new_n215), .C2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT73), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n217), .A2(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n216), .A2(KEYINPUT73), .A3(G128), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n221), .A2(new_n222), .A3(new_n214), .ZN(new_n223));
  XNOR2_X1  g037(.A(KEYINPUT24), .B(G110), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n219), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g040(.A(KEYINPUT77), .B1(new_n202), .B2(new_n198), .ZN(new_n227));
  INV_X1    g041(.A(G146), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT77), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n194), .A2(new_n196), .A3(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n227), .A2(new_n228), .A3(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n205), .A2(new_n226), .A3(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(KEYINPUT78), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n228), .B1(new_n201), .B2(new_n203), .ZN(new_n234));
  INV_X1    g048(.A(new_n231), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT78), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n236), .A2(new_n237), .A3(new_n226), .ZN(new_n238));
  XNOR2_X1  g052(.A(new_n204), .B(G146), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n223), .A2(new_n224), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n211), .B1(new_n215), .B2(new_n218), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n240), .B1(new_n241), .B2(G110), .ZN(new_n242));
  AOI22_X1  g056(.A1(new_n233), .A2(new_n238), .B1(new_n239), .B2(new_n242), .ZN(new_n243));
  XNOR2_X1  g057(.A(KEYINPUT22), .B(G137), .ZN(new_n244));
  INV_X1    g058(.A(G953), .ZN(new_n245));
  AND3_X1   g059(.A1(new_n245), .A2(G221), .A3(G234), .ZN(new_n246));
  XOR2_X1   g060(.A(new_n244), .B(new_n246), .Z(new_n247));
  OAI21_X1  g061(.A(KEYINPUT79), .B1(new_n243), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n239), .A2(new_n242), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n232), .A2(KEYINPUT78), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n237), .B1(new_n236), .B2(new_n226), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n249), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT79), .ZN(new_n253));
  INV_X1    g067(.A(new_n247), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n252), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n248), .A2(new_n255), .ZN(new_n256));
  OAI211_X1 g070(.A(new_n249), .B(new_n247), .C1(new_n250), .C2(new_n251), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT80), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n243), .A2(KEYINPUT80), .A3(new_n247), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n256), .A2(new_n261), .A3(new_n188), .ZN(new_n262));
  NOR2_X1   g076(.A1(KEYINPUT81), .A2(KEYINPUT25), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n192), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(new_n263), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n256), .A2(new_n261), .A3(new_n188), .A4(new_n265), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n190), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  AND2_X1   g081(.A1(new_n256), .A2(new_n261), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n190), .A2(new_n188), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n269), .B(KEYINPUT82), .ZN(new_n270));
  AND2_X1   g084(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n267), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g086(.A(KEYINPUT2), .B(G113), .ZN(new_n273));
  INV_X1    g087(.A(G116), .ZN(new_n274));
  OAI21_X1  g088(.A(KEYINPUT69), .B1(new_n274), .B2(G119), .ZN(new_n275));
  XNOR2_X1  g089(.A(KEYINPUT68), .B(G116), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n275), .B1(new_n276), .B2(G119), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT69), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n274), .A2(KEYINPUT68), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT68), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(G116), .ZN(new_n281));
  AND4_X1   g095(.A1(new_n278), .A2(new_n279), .A3(new_n281), .A4(G119), .ZN(new_n282));
  NOR3_X1   g096(.A1(new_n277), .A2(new_n282), .A3(KEYINPUT70), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT70), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n279), .A2(new_n281), .A3(G119), .ZN(new_n285));
  INV_X1    g099(.A(new_n275), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n276), .A2(new_n278), .A3(G119), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n284), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n273), .B1(new_n283), .B2(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n273), .B1(new_n287), .B2(new_n288), .ZN(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n228), .A2(G143), .ZN(new_n293));
  INV_X1    g107(.A(G143), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(G146), .ZN(new_n295));
  AND2_X1   g109(.A1(KEYINPUT0), .A2(G128), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n293), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(KEYINPUT65), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT65), .ZN(new_n299));
  NAND4_X1  g113(.A1(new_n293), .A2(new_n295), .A3(new_n296), .A4(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT0), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n301), .A2(new_n209), .A3(KEYINPUT64), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT64), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n303), .B1(KEYINPUT0), .B2(G128), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n296), .B1(new_n293), .B2(new_n295), .ZN(new_n306));
  AOI22_X1  g120(.A1(new_n298), .A2(new_n300), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT66), .ZN(new_n308));
  INV_X1    g122(.A(G134), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n308), .B1(new_n309), .B2(G137), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(KEYINPUT11), .ZN(new_n311));
  INV_X1    g125(.A(G131), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT11), .ZN(new_n313));
  OAI211_X1 g127(.A(new_n308), .B(new_n313), .C1(new_n309), .C2(G137), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n309), .A2(G137), .ZN(new_n315));
  NAND4_X1  g129(.A1(new_n311), .A2(new_n312), .A3(new_n314), .A4(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(G137), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n318), .A2(G134), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n319), .B1(new_n310), .B2(KEYINPUT11), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n312), .B1(new_n320), .B2(new_n314), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n307), .B1(new_n317), .B2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT1), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n293), .A2(new_n295), .A3(new_n323), .A4(G128), .ZN(new_n324));
  OAI211_X1 g138(.A(new_n294), .B(G146), .C1(new_n209), .C2(KEYINPUT1), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n209), .A2(new_n228), .A3(G143), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n324), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n309), .A2(G137), .ZN(new_n328));
  OAI21_X1  g142(.A(G131), .B1(new_n328), .B2(new_n319), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n316), .A2(new_n327), .A3(new_n329), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n290), .A2(new_n292), .A3(new_n322), .A4(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(KEYINPUT28), .ZN(new_n332));
  INV_X1    g146(.A(new_n273), .ZN(new_n333));
  OAI21_X1  g147(.A(KEYINPUT70), .B1(new_n277), .B2(new_n282), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n287), .A2(new_n288), .A3(new_n284), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n333), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n336), .A2(new_n291), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT28), .ZN(new_n338));
  NAND4_X1  g152(.A1(new_n337), .A2(new_n338), .A3(new_n322), .A4(new_n330), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n332), .A2(new_n339), .ZN(new_n340));
  OR2_X1    g154(.A1(KEYINPUT71), .A2(G237), .ZN(new_n341));
  NAND2_X1  g155(.A1(KEYINPUT71), .A2(G237), .ZN(new_n342));
  AOI21_X1  g156(.A(G953), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(G210), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n344), .B(KEYINPUT27), .ZN(new_n345));
  XOR2_X1   g159(.A(KEYINPUT26), .B(G101), .Z(new_n346));
  XNOR2_X1  g160(.A(new_n345), .B(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n290), .A2(new_n292), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n322), .A2(new_n330), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n340), .A2(KEYINPUT29), .A3(new_n348), .A4(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(G902), .B1(new_n352), .B2(KEYINPUT72), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n353), .B1(KEYINPUT72), .B2(new_n352), .ZN(new_n354));
  AND3_X1   g168(.A1(new_n324), .A2(new_n325), .A3(new_n326), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n316), .A2(new_n329), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT67), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n355), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n316), .A2(KEYINPUT67), .A3(new_n329), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n320), .A2(new_n314), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(G131), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(new_n316), .ZN(new_n362));
  AOI22_X1  g176(.A1(new_n358), .A2(new_n359), .B1(new_n362), .B2(new_n307), .ZN(new_n363));
  OR2_X1    g177(.A1(new_n363), .A2(new_n337), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n340), .A2(new_n364), .A3(new_n348), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT29), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(new_n331), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n356), .A2(new_n357), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n369), .A2(new_n359), .A3(new_n327), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT30), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n370), .A2(new_n371), .A3(new_n322), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n350), .A2(KEYINPUT30), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n368), .B1(new_n374), .B2(new_n349), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n375), .A2(new_n348), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n367), .A2(new_n376), .ZN(new_n377));
  OAI21_X1  g191(.A(G472), .B1(new_n354), .B2(new_n377), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n348), .B1(new_n340), .B2(new_n364), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  AOI21_X1  g194(.A(KEYINPUT31), .B1(new_n375), .B2(new_n348), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n337), .B1(new_n372), .B2(new_n373), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT31), .ZN(new_n383));
  NOR4_X1   g197(.A1(new_n382), .A2(new_n383), .A3(new_n368), .A4(new_n347), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n380), .B1(new_n381), .B2(new_n384), .ZN(new_n385));
  NOR2_X1   g199(.A1(G472), .A2(G902), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n385), .A2(KEYINPUT32), .A3(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT32), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n371), .B1(new_n322), .B2(new_n330), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n389), .B1(new_n363), .B2(new_n371), .ZN(new_n390));
  OAI211_X1 g204(.A(new_n331), .B(new_n348), .C1(new_n390), .C2(new_n337), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(new_n383), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n375), .A2(KEYINPUT31), .A3(new_n348), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n379), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(new_n386), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n388), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n378), .A2(new_n387), .A3(new_n396), .ZN(new_n397));
  AND2_X1   g211(.A1(new_n272), .A2(new_n397), .ZN(new_n398));
  OAI21_X1  g212(.A(G210), .B1(G237), .B2(G902), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n355), .A2(new_n195), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n401), .B1(new_n195), .B2(new_n307), .ZN(new_n402));
  INV_X1    g216(.A(G224), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n403), .A2(G953), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n402), .B(new_n404), .ZN(new_n405));
  AND2_X1   g219(.A1(KEYINPUT83), .A2(G101), .ZN(new_n406));
  NOR2_X1   g220(.A1(KEYINPUT83), .A2(G101), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(G104), .ZN(new_n409));
  OAI21_X1  g223(.A(KEYINPUT3), .B1(new_n409), .B2(G107), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT3), .ZN(new_n411));
  INV_X1    g225(.A(G107), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n411), .A2(new_n412), .A3(G104), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n409), .A2(G107), .ZN(new_n414));
  NAND4_X1  g228(.A1(new_n408), .A2(new_n410), .A3(new_n413), .A4(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n410), .A2(new_n413), .A3(new_n414), .ZN(new_n416));
  AOI22_X1  g230(.A1(new_n415), .A2(KEYINPUT4), .B1(new_n416), .B2(G101), .ZN(new_n417));
  AND3_X1   g231(.A1(new_n416), .A2(KEYINPUT4), .A3(G101), .ZN(new_n418));
  OR2_X1    g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n419), .B1(new_n336), .B2(new_n291), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n334), .A2(KEYINPUT5), .A3(new_n335), .ZN(new_n421));
  INV_X1    g235(.A(G113), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n274), .A2(G119), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT5), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n422), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n421), .A2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT84), .ZN(new_n427));
  XNOR2_X1  g241(.A(G104), .B(G107), .ZN(new_n428));
  INV_X1    g242(.A(G101), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n427), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n412), .A2(G104), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(new_n414), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n432), .A2(KEYINPUT84), .A3(G101), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n415), .A2(new_n430), .A3(new_n433), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n291), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n426), .A2(new_n435), .ZN(new_n436));
  XNOR2_X1  g250(.A(G110), .B(G122), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n420), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n420), .A2(new_n436), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n437), .A2(KEYINPUT89), .ZN(new_n440));
  AOI22_X1  g254(.A1(new_n438), .A2(KEYINPUT6), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  AOI22_X1  g255(.A1(new_n349), .A2(new_n419), .B1(new_n426), .B2(new_n435), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT6), .ZN(new_n443));
  INV_X1    g257(.A(new_n440), .ZN(new_n444));
  NOR3_X1   g258(.A1(new_n442), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  OAI211_X1 g259(.A(KEYINPUT90), .B(new_n405), .C1(new_n441), .C2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n404), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(KEYINPUT7), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT92), .ZN(new_n449));
  OAI211_X1 g263(.A(new_n402), .B(new_n448), .C1(new_n449), .C2(new_n404), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n402), .B1(new_n449), .B2(new_n404), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n451), .A2(KEYINPUT7), .A3(new_n447), .ZN(new_n452));
  AND3_X1   g266(.A1(new_n438), .A2(new_n450), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n426), .A2(new_n292), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(new_n434), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n424), .B1(new_n287), .B2(new_n288), .ZN(new_n456));
  INV_X1    g270(.A(new_n425), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n435), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n455), .A2(new_n458), .ZN(new_n459));
  XNOR2_X1  g273(.A(KEYINPUT91), .B(KEYINPUT8), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n437), .B(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(G902), .B1(new_n453), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n446), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n439), .A2(KEYINPUT6), .A3(new_n440), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n443), .B1(new_n442), .B2(new_n437), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n442), .A2(new_n444), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  AOI21_X1  g282(.A(KEYINPUT90), .B1(new_n468), .B2(new_n405), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n400), .B1(new_n464), .B2(new_n469), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n405), .B1(new_n441), .B2(new_n445), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT90), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n473), .A2(new_n399), .A3(new_n446), .A4(new_n463), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n470), .A2(KEYINPUT93), .A3(new_n474), .ZN(new_n475));
  OAI21_X1  g289(.A(G214), .B1(G237), .B2(G902), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n464), .A2(new_n469), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT93), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n477), .A2(new_n478), .A3(new_n399), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n475), .A2(new_n476), .A3(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(G475), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n204), .A2(G146), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n483), .A2(new_n234), .ZN(new_n484));
  AND2_X1   g298(.A1(KEYINPUT71), .A2(G237), .ZN(new_n485));
  NOR2_X1   g299(.A1(KEYINPUT71), .A2(G237), .ZN(new_n486));
  OAI211_X1 g300(.A(G214), .B(new_n245), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(new_n294), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n341), .A2(new_n342), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n489), .A2(G143), .A3(G214), .A4(new_n245), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n491), .A2(KEYINPUT17), .A3(G131), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(G131), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n488), .A2(new_n490), .A3(new_n312), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  OAI211_X1 g309(.A(new_n484), .B(new_n492), .C1(KEYINPUT17), .C2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT94), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n197), .A2(new_n200), .A3(G146), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n231), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(KEYINPUT18), .A2(G131), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n488), .A2(new_n490), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n500), .B1(new_n488), .B2(new_n490), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n497), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n503), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n505), .A2(KEYINPUT94), .A3(new_n499), .A4(new_n501), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  XNOR2_X1  g321(.A(G113), .B(G122), .ZN(new_n508));
  XNOR2_X1  g322(.A(KEYINPUT96), .B(G104), .ZN(new_n509));
  XOR2_X1   g323(.A(new_n508), .B(new_n509), .Z(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n496), .A2(new_n507), .A3(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n511), .B1(new_n496), .B2(new_n507), .ZN(new_n514));
  OR2_X1    g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n482), .B1(new_n515), .B2(new_n188), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT19), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n227), .A2(new_n518), .A3(new_n230), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n197), .A2(new_n200), .A3(KEYINPUT19), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n519), .A2(new_n228), .A3(new_n520), .ZN(new_n521));
  AND2_X1   g335(.A1(new_n205), .A2(new_n521), .ZN(new_n522));
  AOI22_X1  g336(.A1(new_n504), .A2(new_n506), .B1(new_n522), .B2(new_n495), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n510), .B1(new_n523), .B2(KEYINPUT95), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n522), .A2(new_n495), .ZN(new_n525));
  AND3_X1   g339(.A1(new_n507), .A2(KEYINPUT95), .A3(new_n525), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n512), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT20), .ZN(new_n528));
  NOR2_X1   g342(.A1(G475), .A2(G902), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n527), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(KEYINPUT97), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT97), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n527), .A2(new_n532), .A3(new_n528), .A4(new_n529), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n527), .A2(new_n529), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(KEYINPUT20), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n531), .A2(new_n533), .A3(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(G952), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n537), .A2(G953), .ZN(new_n538));
  INV_X1    g352(.A(G234), .ZN(new_n539));
  INV_X1    g353(.A(G237), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  AOI211_X1 g356(.A(new_n188), .B(new_n245), .C1(G234), .C2(G237), .ZN(new_n543));
  XNOR2_X1  g357(.A(KEYINPUT21), .B(G898), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  XNOR2_X1  g360(.A(KEYINPUT9), .B(G234), .ZN(new_n547));
  NOR3_X1   g361(.A1(new_n547), .A2(new_n187), .A3(G953), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  XNOR2_X1  g363(.A(G128), .B(G143), .ZN(new_n550));
  OR2_X1    g364(.A1(new_n550), .A2(G134), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n279), .A2(new_n281), .A3(G122), .ZN(new_n552));
  INV_X1    g366(.A(G122), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(G116), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n552), .A2(new_n412), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n550), .A2(G134), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n551), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT14), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n554), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n552), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(KEYINPUT98), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT98), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n552), .A2(new_n562), .A3(new_n559), .ZN(new_n563));
  INV_X1    g377(.A(new_n552), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(new_n558), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n561), .A2(new_n563), .A3(new_n565), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n557), .B1(new_n566), .B2(G107), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n552), .A2(new_n554), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(G107), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(new_n555), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n209), .A2(G143), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT13), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n309), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n573), .B(new_n550), .ZN(new_n574));
  AND2_X1   g388(.A1(new_n570), .A2(new_n574), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n549), .B1(new_n567), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n570), .A2(new_n574), .ZN(new_n577));
  AOI22_X1  g391(.A1(new_n560), .A2(KEYINPUT98), .B1(new_n564), .B2(new_n558), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n412), .B1(new_n578), .B2(new_n563), .ZN(new_n579));
  OAI211_X1 g393(.A(new_n577), .B(new_n548), .C1(new_n579), .C2(new_n557), .ZN(new_n580));
  AOI21_X1  g394(.A(G902), .B1(new_n576), .B2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(G478), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n582), .A2(KEYINPUT15), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n581), .B(new_n583), .ZN(new_n584));
  AND4_X1   g398(.A1(new_n517), .A2(new_n536), .A3(new_n546), .A4(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT87), .ZN(new_n586));
  XNOR2_X1  g400(.A(G110), .B(G140), .ZN(new_n587));
  INV_X1    g401(.A(G227), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n588), .A2(G953), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n587), .B(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n434), .A2(new_n355), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n325), .A2(KEYINPUT85), .A3(new_n326), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(new_n324), .ZN(new_n595));
  AOI21_X1  g409(.A(KEYINPUT85), .B1(new_n325), .B2(new_n326), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n597), .A2(new_n434), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n362), .B1(new_n593), .B2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT12), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n592), .B1(new_n434), .B2(new_n597), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n602), .A2(KEYINPUT12), .A3(new_n362), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n362), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT10), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n606), .B1(new_n597), .B2(new_n434), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n307), .B1(new_n417), .B2(new_n418), .ZN(new_n608));
  AND2_X1   g422(.A1(new_n430), .A2(new_n433), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n609), .A2(KEYINPUT10), .A3(new_n327), .A4(new_n415), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n605), .A2(new_n607), .A3(new_n608), .A4(new_n610), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n591), .B1(new_n604), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n591), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n607), .A2(new_n608), .A3(new_n610), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT86), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n605), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n607), .A2(new_n608), .A3(new_n610), .A4(KEYINPUT86), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n613), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n586), .B1(new_n612), .B2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n603), .ZN(new_n620));
  AOI21_X1  g434(.A(KEYINPUT12), .B1(new_n602), .B2(new_n362), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n611), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(new_n590), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n616), .A2(new_n617), .ZN(new_n624));
  INV_X1    g438(.A(new_n613), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n623), .A2(new_n626), .A3(KEYINPUT87), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n619), .A2(new_n627), .A3(G469), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n625), .A2(new_n604), .ZN(new_n629));
  INV_X1    g443(.A(new_n611), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n630), .B1(new_n616), .B2(new_n617), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n629), .B1(new_n631), .B2(new_n591), .ZN(new_n632));
  INV_X1    g446(.A(G469), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n632), .A2(new_n633), .A3(new_n188), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n633), .A2(new_n188), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n628), .A2(new_n634), .A3(new_n636), .ZN(new_n637));
  OAI21_X1  g451(.A(G221), .B1(new_n547), .B2(G902), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT88), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n637), .A2(KEYINPUT88), .A3(new_n638), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  AND4_X1   g457(.A1(new_n398), .A2(new_n481), .A3(new_n585), .A4(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(new_n408), .ZN(G3));
  OR2_X1    g459(.A1(new_n267), .A2(new_n271), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n394), .A2(G902), .ZN(new_n647));
  INV_X1    g461(.A(G472), .ZN(new_n648));
  OR2_X1    g462(.A1(new_n648), .A2(KEYINPUT99), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n647), .B(new_n649), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n646), .A2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT100), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n582), .A2(G902), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT33), .ZN(new_n654));
  AND3_X1   g468(.A1(new_n576), .A2(new_n580), .A3(new_n654), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n654), .B1(new_n576), .B2(new_n580), .ZN(new_n656));
  OAI211_X1 g470(.A(new_n652), .B(new_n653), .C1(new_n655), .C2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n653), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n576), .A2(new_n580), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(KEYINPUT33), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n576), .A2(new_n580), .A3(new_n654), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n658), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  OAI21_X1  g476(.A(KEYINPUT100), .B1(new_n581), .B2(G478), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n657), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(KEYINPUT101), .ZN(new_n665));
  INV_X1    g479(.A(KEYINPUT101), .ZN(new_n666));
  OAI211_X1 g480(.A(new_n657), .B(new_n666), .C1(new_n662), .C2(new_n663), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n669), .B1(new_n517), .B2(new_n536), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n470), .A2(new_n474), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(new_n476), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n672), .A2(new_n545), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n651), .A2(new_n643), .A3(new_n670), .A4(new_n673), .ZN(new_n674));
  XOR2_X1   g488(.A(KEYINPUT34), .B(G104), .Z(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G6));
  NAND2_X1  g490(.A1(new_n385), .A2(new_n188), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(new_n649), .ZN(new_n678));
  AND3_X1   g492(.A1(new_n637), .A2(KEYINPUT88), .A3(new_n638), .ZN(new_n679));
  AOI21_X1  g493(.A(KEYINPUT88), .B1(new_n637), .B2(new_n638), .ZN(new_n680));
  OAI211_X1 g494(.A(new_n272), .B(new_n678), .C1(new_n679), .C2(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(new_n476), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n682), .B1(new_n470), .B2(new_n474), .ZN(new_n683));
  AOI211_X1 g497(.A(new_n584), .B(new_n516), .C1(new_n535), .C2(new_n530), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n683), .A2(new_n684), .A3(new_n546), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n681), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(KEYINPUT35), .B(G107), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(G9));
  NOR2_X1   g502(.A1(new_n254), .A2(KEYINPUT36), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n252), .B(new_n689), .ZN(new_n690));
  AND2_X1   g504(.A1(new_n690), .A2(new_n270), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n262), .A2(new_n263), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n692), .A2(new_n266), .A3(new_n191), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n691), .B1(new_n693), .B2(new_n189), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n650), .A2(new_n694), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n481), .A2(new_n695), .A3(new_n585), .A4(new_n643), .ZN(new_n696));
  XOR2_X1   g510(.A(KEYINPUT37), .B(G110), .Z(new_n697));
  XNOR2_X1  g511(.A(new_n696), .B(new_n697), .ZN(G12));
  NOR2_X1   g512(.A1(new_n672), .A2(new_n694), .ZN(new_n699));
  INV_X1    g513(.A(new_n535), .ZN(new_n700));
  INV_X1    g514(.A(new_n530), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n517), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(G900), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n543), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(new_n541), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  NOR3_X1   g520(.A1(new_n702), .A2(new_n584), .A3(new_n706), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n699), .A2(new_n643), .A3(new_n397), .A4(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G128), .ZN(G30));
  XNOR2_X1  g523(.A(new_n705), .B(KEYINPUT39), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n643), .A2(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT40), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n643), .A2(KEYINPUT40), .A3(new_n710), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(new_n584), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(new_n476), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n717), .B1(new_n536), .B2(new_n517), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(new_n694), .ZN(new_n719));
  XOR2_X1   g533(.A(new_n719), .B(KEYINPUT103), .Z(new_n720));
  NOR2_X1   g534(.A1(new_n348), .A2(new_n368), .ZN(new_n721));
  AOI21_X1  g535(.A(G902), .B1(new_n721), .B2(new_n351), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n348), .B1(new_n382), .B2(new_n368), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n648), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n396), .A2(new_n387), .A3(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(KEYINPUT102), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n392), .A2(new_n393), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n395), .B1(new_n728), .B2(new_n380), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n724), .B1(new_n729), .B2(KEYINPUT32), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT102), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n730), .A2(new_n731), .A3(new_n396), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n727), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n475), .A2(new_n479), .ZN(new_n734));
  XOR2_X1   g548(.A(new_n734), .B(KEYINPUT38), .Z(new_n735));
  NAND4_X1  g549(.A1(new_n715), .A2(new_n720), .A3(new_n733), .A4(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G143), .ZN(G45));
  AOI221_X4 g551(.A(new_n706), .B1(new_n665), .B2(new_n667), .C1(new_n536), .C2(new_n517), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n699), .A2(new_n643), .A3(new_n397), .A4(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G146), .ZN(G48));
  NAND2_X1  g554(.A1(new_n632), .A2(new_n188), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(G469), .ZN(new_n742));
  AND3_X1   g556(.A1(new_n742), .A2(new_n638), .A3(new_n634), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n398), .A2(new_n673), .A3(new_n670), .A4(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(KEYINPUT41), .B(G113), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n744), .B(new_n745), .ZN(G15));
  NAND2_X1  g560(.A1(new_n272), .A2(new_n397), .ZN(new_n747));
  INV_X1    g561(.A(new_n743), .ZN(new_n748));
  NOR3_X1   g562(.A1(new_n747), .A2(new_n685), .A3(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(new_n274), .ZN(G18));
  NAND4_X1  g564(.A1(new_n699), .A2(new_n397), .A3(new_n585), .A4(new_n743), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G119), .ZN(G21));
  XNOR2_X1  g566(.A(KEYINPUT104), .B(G472), .ZN(new_n753));
  AND2_X1   g567(.A1(new_n340), .A2(new_n351), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n728), .B1(new_n348), .B2(new_n754), .ZN(new_n755));
  AOI22_X1  g569(.A1(new_n677), .A2(new_n753), .B1(new_n755), .B2(new_n386), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n272), .A2(new_n546), .A3(new_n743), .A4(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n718), .A2(new_n671), .ZN(new_n758));
  OR2_X1    g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G122), .ZN(G24));
  NOR2_X1   g574(.A1(new_n672), .A2(new_n748), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n693), .A2(new_n189), .ZN(new_n762));
  INV_X1    g576(.A(new_n691), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n761), .A2(new_n764), .A3(new_n738), .A4(new_n756), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G125), .ZN(G27));
  INV_X1    g580(.A(new_n738), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n767), .A2(KEYINPUT42), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n682), .B1(new_n475), .B2(new_n479), .ZN(new_n769));
  INV_X1    g583(.A(new_n638), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n612), .A2(new_n618), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n635), .B1(new_n771), .B2(G469), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n770), .B1(new_n772), .B2(new_n634), .ZN(new_n773));
  AND3_X1   g587(.A1(new_n769), .A2(KEYINPUT105), .A3(new_n773), .ZN(new_n774));
  AOI21_X1  g588(.A(KEYINPUT105), .B1(new_n769), .B2(new_n773), .ZN(new_n775));
  OAI211_X1 g589(.A(new_n768), .B(new_n398), .C1(new_n774), .C2(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n387), .A2(KEYINPUT106), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT106), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n729), .A2(new_n778), .A3(KEYINPUT32), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n777), .A2(new_n378), .A3(new_n779), .A4(new_n396), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n738), .A2(new_n272), .A3(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n734), .A2(new_n476), .A3(new_n773), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT105), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n769), .A2(KEYINPUT105), .A3(new_n773), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n781), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT42), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n776), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(new_n312), .ZN(G33));
  OAI211_X1 g603(.A(new_n398), .B(new_n707), .C1(new_n774), .C2(new_n775), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G134), .ZN(G36));
  INV_X1    g605(.A(KEYINPUT111), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n650), .A2(new_n764), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n536), .A2(new_n668), .A3(new_n517), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(KEYINPUT110), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n795), .A2(KEYINPUT43), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT43), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n794), .A2(KEYINPUT110), .A3(new_n797), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n793), .B1(new_n796), .B2(new_n798), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n792), .B1(new_n799), .B2(KEYINPUT44), .ZN(new_n800));
  INV_X1    g614(.A(new_n769), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n801), .B1(new_n799), .B2(KEYINPUT44), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT112), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n678), .A2(new_n694), .ZN(new_n804));
  AND3_X1   g618(.A1(new_n794), .A2(KEYINPUT110), .A3(new_n797), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n797), .B1(new_n794), .B2(KEYINPUT110), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n804), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT44), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n807), .A2(KEYINPUT111), .A3(new_n808), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n800), .A2(new_n802), .A3(new_n803), .A4(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT108), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT46), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT45), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n612), .A2(new_n618), .A3(new_n586), .ZN(new_n814));
  AOI21_X1  g628(.A(KEYINPUT87), .B1(new_n623), .B2(new_n626), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n813), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT107), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n633), .B1(new_n771), .B2(KEYINPUT45), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n816), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  AOI21_X1  g633(.A(KEYINPUT45), .B1(new_n619), .B2(new_n627), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n623), .A2(new_n626), .ZN(new_n821));
  OAI21_X1  g635(.A(G469), .B1(new_n821), .B2(new_n813), .ZN(new_n822));
  OAI21_X1  g636(.A(KEYINPUT107), .B1(new_n820), .B2(new_n822), .ZN(new_n823));
  AOI211_X1 g637(.A(new_n812), .B(new_n635), .C1(new_n819), .C2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(new_n634), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n811), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n635), .B1(new_n819), .B2(new_n823), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n827), .A2(KEYINPUT46), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n828), .A2(KEYINPUT108), .A3(new_n634), .ZN(new_n829));
  OR3_X1    g643(.A1(new_n827), .A2(KEYINPUT109), .A3(KEYINPUT46), .ZN(new_n830));
  OAI21_X1  g644(.A(KEYINPUT109), .B1(new_n827), .B2(KEYINPUT46), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n826), .A2(new_n829), .A3(new_n830), .A4(new_n831), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n832), .A2(new_n638), .A3(new_n710), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n810), .A2(new_n833), .ZN(new_n834));
  AOI21_X1  g648(.A(KEYINPUT111), .B1(new_n807), .B2(new_n808), .ZN(new_n835));
  OAI211_X1 g649(.A(KEYINPUT44), .B(new_n804), .C1(new_n805), .C2(new_n806), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(new_n769), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n803), .B1(new_n838), .B2(new_n809), .ZN(new_n839));
  OR2_X1    g653(.A1(new_n834), .A2(new_n839), .ZN(new_n840));
  XNOR2_X1  g654(.A(new_n840), .B(G137), .ZN(G39));
  NAND2_X1  g655(.A1(new_n832), .A2(new_n638), .ZN(new_n842));
  XNOR2_X1  g656(.A(KEYINPUT113), .B(KEYINPUT47), .ZN(new_n843));
  INV_X1    g657(.A(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n832), .A2(new_n638), .A3(new_n843), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NOR4_X1   g661(.A1(new_n801), .A2(new_n767), .A3(new_n272), .A4(new_n397), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  XNOR2_X1  g663(.A(new_n849), .B(G140), .ZN(G42));
  NAND2_X1  g664(.A1(new_n537), .A2(new_n245), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n541), .B1(new_n796), .B2(new_n798), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n852), .A2(new_n743), .A3(new_n769), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n764), .A2(new_n756), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n646), .A2(new_n541), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n731), .B1(new_n730), .B2(new_n396), .ZN(new_n856));
  AND4_X1   g670(.A1(new_n731), .A2(new_n396), .A3(new_n387), .A4(new_n725), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n855), .A2(new_n858), .A3(new_n743), .A4(new_n769), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n536), .A2(new_n517), .ZN(new_n860));
  INV_X1    g674(.A(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(new_n669), .ZN(new_n862));
  OAI22_X1  g676(.A1(new_n853), .A2(new_n854), .B1(new_n859), .B2(new_n862), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n735), .A2(new_n476), .A3(new_n748), .ZN(new_n864));
  AND2_X1   g678(.A1(new_n272), .A2(new_n756), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n852), .A2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n864), .A2(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT50), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n864), .A2(KEYINPUT50), .A3(new_n867), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n863), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  AND2_X1   g686(.A1(new_n742), .A2(new_n634), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n847), .B1(new_n770), .B2(new_n873), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n866), .A2(new_n801), .ZN(new_n875));
  INV_X1    g689(.A(new_n875), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n872), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT51), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(new_n670), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n538), .B1(new_n859), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n780), .A2(new_n272), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n853), .A2(new_n882), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n883), .B(KEYINPUT48), .ZN(new_n884));
  AOI211_X1 g698(.A(new_n881), .B(new_n884), .C1(new_n761), .C2(new_n867), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n874), .A2(KEYINPUT117), .ZN(new_n886));
  INV_X1    g700(.A(new_n846), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n843), .B1(new_n832), .B2(new_n638), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(new_n873), .ZN(new_n890));
  OAI211_X1 g704(.A(new_n889), .B(KEYINPUT117), .C1(new_n638), .C2(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n891), .A2(new_n875), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n886), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n872), .A2(KEYINPUT51), .ZN(new_n894));
  OAI211_X1 g708(.A(new_n879), .B(new_n885), .C1(new_n893), .C2(new_n894), .ZN(new_n895));
  AND3_X1   g709(.A1(new_n378), .A2(new_n387), .A3(new_n396), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n896), .B1(new_n641), .B2(new_n642), .ZN(new_n897));
  NOR4_X1   g711(.A1(new_n694), .A2(new_n702), .A3(new_n716), .A4(new_n706), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n897), .A2(new_n769), .A3(new_n898), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n767), .A2(new_n854), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n900), .B1(new_n774), .B2(new_n775), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n790), .A2(new_n899), .A3(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(new_n781), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n904), .B1(new_n774), .B2(new_n775), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n747), .B1(new_n784), .B2(new_n785), .ZN(new_n906));
  AOI22_X1  g720(.A1(KEYINPUT42), .A2(new_n905), .B1(new_n906), .B2(new_n768), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n480), .A2(new_n545), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n536), .A2(new_n517), .A3(new_n716), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n909), .B1(new_n861), .B2(new_n669), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n908), .A2(new_n651), .A3(new_n643), .A4(new_n910), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n398), .A2(new_n673), .A3(new_n684), .A4(new_n743), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n911), .A2(new_n696), .A3(new_n744), .A4(new_n912), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n398), .A2(new_n481), .A3(new_n585), .A4(new_n643), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n759), .A2(new_n914), .A3(new_n751), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n903), .A2(new_n907), .A3(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT52), .ZN(new_n918));
  AOI211_X1 g732(.A(new_n770), .B(new_n706), .C1(new_n772), .C2(new_n634), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n718), .A2(new_n694), .A3(new_n671), .A4(new_n919), .ZN(new_n920));
  OAI21_X1  g734(.A(KEYINPUT114), .B1(new_n858), .B2(new_n920), .ZN(new_n921));
  AND2_X1   g735(.A1(new_n718), .A2(new_n671), .ZN(new_n922));
  AND2_X1   g736(.A1(new_n694), .A2(new_n919), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT114), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n922), .A2(new_n733), .A3(new_n923), .A4(new_n924), .ZN(new_n925));
  AND2_X1   g739(.A1(new_n921), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n708), .A2(new_n739), .A3(new_n765), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n918), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n921), .A2(new_n925), .ZN(new_n929));
  OAI211_X1 g743(.A(new_n897), .B(new_n699), .C1(new_n707), .C2(new_n738), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n929), .A2(new_n930), .A3(KEYINPUT52), .A4(new_n765), .ZN(new_n931));
  AND2_X1   g745(.A1(new_n928), .A2(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT53), .ZN(new_n933));
  NOR3_X1   g747(.A1(new_n917), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n585), .A2(new_n683), .A3(new_n764), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n397), .A2(new_n743), .ZN(new_n936));
  OAI22_X1  g750(.A1(new_n935), .A2(new_n936), .B1(new_n757), .B2(new_n758), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n644), .A2(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(new_n909), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n670), .A2(new_n939), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n940), .A2(new_n681), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n749), .B1(new_n941), .B2(new_n908), .ZN(new_n942));
  AND2_X1   g756(.A1(new_n744), .A2(new_n696), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n938), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  NOR3_X1   g758(.A1(new_n944), .A2(new_n788), .A3(new_n902), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT115), .ZN(new_n946));
  AND3_X1   g760(.A1(new_n928), .A2(new_n946), .A3(new_n931), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n946), .B1(new_n928), .B2(new_n931), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n945), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n934), .B1(new_n933), .B2(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT54), .ZN(new_n951));
  XOR2_X1   g765(.A(KEYINPUT116), .B(KEYINPUT54), .Z(new_n952));
  INV_X1    g766(.A(new_n952), .ZN(new_n953));
  OAI211_X1 g767(.A(KEYINPUT53), .B(new_n945), .C1(new_n947), .C2(new_n948), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n933), .B1(new_n917), .B2(new_n932), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  OAI22_X1  g770(.A1(new_n950), .A2(new_n951), .B1(new_n953), .B2(new_n956), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n851), .B1(new_n895), .B2(new_n957), .ZN(new_n958));
  OR2_X1    g772(.A1(new_n890), .A2(KEYINPUT49), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n890), .A2(KEYINPUT49), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n959), .A2(new_n476), .A3(new_n638), .A4(new_n960), .ZN(new_n961));
  NOR3_X1   g775(.A1(new_n961), .A2(new_n646), .A3(new_n794), .ZN(new_n962));
  INV_X1    g776(.A(new_n735), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n962), .A2(new_n963), .A3(new_n858), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n958), .A2(new_n964), .ZN(G75));
  NOR2_X1   g779(.A1(new_n245), .A2(G952), .ZN(new_n966));
  INV_X1    g780(.A(new_n966), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n188), .B1(new_n954), .B2(new_n955), .ZN(new_n968));
  AOI21_X1  g782(.A(KEYINPUT56), .B1(new_n968), .B2(G210), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n468), .B(KEYINPUT118), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n970), .B(KEYINPUT55), .Z(new_n971));
  XNOR2_X1  g785(.A(new_n971), .B(new_n405), .ZN(new_n972));
  XNOR2_X1  g786(.A(KEYINPUT119), .B(KEYINPUT120), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n972), .B(new_n973), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n967), .B1(new_n969), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n968), .A2(G210), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT56), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n976), .A2(new_n977), .A3(new_n974), .ZN(new_n978));
  INV_X1    g792(.A(KEYINPUT121), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n969), .A2(KEYINPUT121), .A3(new_n974), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n975), .B1(new_n980), .B2(new_n981), .ZN(G51));
  XNOR2_X1  g796(.A(new_n635), .B(KEYINPUT57), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n956), .A2(new_n953), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n952), .B1(new_n954), .B2(new_n955), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n983), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n986), .A2(new_n632), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n968), .A2(new_n819), .A3(new_n823), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n966), .B1(new_n987), .B2(new_n988), .ZN(G54));
  AND2_X1   g803(.A1(KEYINPUT58), .A2(G475), .ZN(new_n990));
  AND3_X1   g804(.A1(new_n968), .A2(new_n527), .A3(new_n990), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n527), .B1(new_n968), .B2(new_n990), .ZN(new_n992));
  NOR3_X1   g806(.A1(new_n991), .A2(new_n992), .A3(new_n966), .ZN(G60));
  NAND2_X1  g807(.A1(new_n660), .A2(new_n661), .ZN(new_n994));
  NAND2_X1  g808(.A1(G478), .A2(G902), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n995), .B(KEYINPUT59), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n994), .B1(new_n957), .B2(new_n996), .ZN(new_n997));
  AND2_X1   g811(.A1(new_n994), .A2(new_n996), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n998), .B1(new_n984), .B2(new_n985), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n999), .A2(new_n967), .ZN(new_n1000));
  NOR2_X1   g814(.A1(new_n997), .A2(new_n1000), .ZN(G63));
  INV_X1    g815(.A(KEYINPUT61), .ZN(new_n1002));
  NAND2_X1  g816(.A1(G217), .A2(G902), .ZN(new_n1003));
  XNOR2_X1  g817(.A(new_n1003), .B(KEYINPUT60), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n1004), .B1(new_n954), .B2(new_n955), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1005), .A2(new_n690), .ZN(new_n1006));
  INV_X1    g820(.A(new_n1006), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n967), .B1(new_n1005), .B2(new_n268), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n1002), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  OR2_X1    g823(.A1(new_n1005), .A2(new_n268), .ZN(new_n1010));
  NAND4_X1  g824(.A1(new_n1010), .A2(KEYINPUT61), .A3(new_n967), .A4(new_n1006), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1009), .A2(new_n1011), .ZN(G66));
  OAI21_X1  g826(.A(G953), .B1(new_n544), .B2(new_n403), .ZN(new_n1013));
  OAI21_X1  g827(.A(new_n1013), .B1(new_n916), .B2(G953), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n970), .B1(G898), .B2(new_n245), .ZN(new_n1015));
  XNOR2_X1  g829(.A(new_n1014), .B(new_n1015), .ZN(G69));
  NAND2_X1  g830(.A1(new_n519), .A2(new_n520), .ZN(new_n1017));
  XNOR2_X1  g831(.A(new_n374), .B(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g832(.A(new_n1018), .B(KEYINPUT122), .ZN(new_n1019));
  INV_X1    g833(.A(new_n848), .ZN(new_n1020));
  INV_X1    g834(.A(new_n927), .ZN(new_n1021));
  AND3_X1   g835(.A1(new_n736), .A2(KEYINPUT62), .A3(new_n1021), .ZN(new_n1022));
  AOI21_X1  g836(.A(KEYINPUT62), .B1(new_n736), .B2(new_n1021), .ZN(new_n1023));
  OAI22_X1  g837(.A1(new_n889), .A2(new_n1020), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  OR4_X1    g838(.A1(new_n747), .A2(new_n711), .A3(new_n940), .A4(new_n801), .ZN(new_n1025));
  OAI21_X1  g839(.A(new_n1025), .B1(new_n834), .B2(new_n839), .ZN(new_n1026));
  INV_X1    g840(.A(KEYINPUT123), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  OAI211_X1 g842(.A(KEYINPUT123), .B(new_n1025), .C1(new_n834), .C2(new_n839), .ZN(new_n1029));
  AOI21_X1  g843(.A(new_n1024), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g844(.A(new_n1019), .B1(new_n1030), .B2(G953), .ZN(new_n1031));
  AOI21_X1  g845(.A(new_n1018), .B1(G900), .B2(G953), .ZN(new_n1032));
  NAND3_X1  g846(.A1(new_n907), .A2(new_n790), .A3(new_n1021), .ZN(new_n1033));
  AOI21_X1  g847(.A(new_n1033), .B1(new_n847), .B2(new_n848), .ZN(new_n1034));
  NOR2_X1   g848(.A1(new_n882), .A2(new_n758), .ZN(new_n1035));
  NAND4_X1  g849(.A1(new_n832), .A2(new_n638), .A3(new_n710), .A4(new_n1035), .ZN(new_n1036));
  XNOR2_X1  g850(.A(new_n1036), .B(KEYINPUT124), .ZN(new_n1037));
  NAND3_X1  g851(.A1(new_n1034), .A2(new_n840), .A3(new_n1037), .ZN(new_n1038));
  OAI21_X1  g852(.A(new_n1032), .B1(new_n1038), .B2(G953), .ZN(new_n1039));
  AOI21_X1  g853(.A(new_n245), .B1(G227), .B2(G900), .ZN(new_n1040));
  XNOR2_X1  g854(.A(new_n1040), .B(KEYINPUT125), .ZN(new_n1041));
  AND3_X1   g855(.A1(new_n1031), .A2(new_n1039), .A3(new_n1041), .ZN(new_n1042));
  AOI21_X1  g856(.A(new_n1041), .B1(new_n1031), .B2(new_n1039), .ZN(new_n1043));
  NOR2_X1   g857(.A1(new_n1042), .A2(new_n1043), .ZN(G72));
  NAND4_X1  g858(.A1(new_n1034), .A2(new_n840), .A3(new_n916), .A4(new_n1037), .ZN(new_n1045));
  INV_X1    g859(.A(KEYINPUT126), .ZN(new_n1046));
  NAND2_X1  g860(.A1(G472), .A2(G902), .ZN(new_n1047));
  XOR2_X1   g861(.A(new_n1047), .B(KEYINPUT63), .Z(new_n1048));
  AND3_X1   g862(.A1(new_n1045), .A2(new_n1046), .A3(new_n1048), .ZN(new_n1049));
  AOI21_X1  g863(.A(new_n1046), .B1(new_n1045), .B2(new_n1048), .ZN(new_n1050));
  NAND2_X1  g864(.A1(new_n375), .A2(new_n347), .ZN(new_n1051));
  NOR3_X1   g865(.A1(new_n1049), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  NAND2_X1  g866(.A1(new_n1030), .A2(new_n916), .ZN(new_n1053));
  AOI21_X1  g867(.A(new_n723), .B1(new_n1053), .B2(new_n1048), .ZN(new_n1054));
  NAND3_X1  g868(.A1(new_n1051), .A2(new_n723), .A3(new_n1048), .ZN(new_n1055));
  XOR2_X1   g869(.A(new_n1055), .B(KEYINPUT127), .Z(new_n1056));
  OAI21_X1  g870(.A(new_n967), .B1(new_n950), .B2(new_n1056), .ZN(new_n1057));
  NOR3_X1   g871(.A1(new_n1052), .A2(new_n1054), .A3(new_n1057), .ZN(G57));
endmodule


