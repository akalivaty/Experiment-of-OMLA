//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 0 1 1 0 0 0 1 0 1 0 1 1 1 1 0 1 1 1 0 1 0 0 0 1 0 0 1 1 1 1 1 1 0 1 0 1 1 1 0 1 1 0 0 0 0 1 1 0 1 0 0 0 1 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:34 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1201, new_n1202, new_n1203, new_n1205, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1266, new_n1267, new_n1268, new_n1269;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XOR2_X1   g0011(.A(new_n211), .B(KEYINPUT0), .Z(new_n212));
  AND2_X1   g0012(.A1(G116), .A2(G270), .ZN(new_n213));
  INV_X1    g0013(.A(G77), .ZN(new_n214));
  INV_X1    g0014(.A(G244), .ZN(new_n215));
  INV_X1    g0015(.A(G97), .ZN(new_n216));
  INV_X1    g0016(.A(G257), .ZN(new_n217));
  OAI22_X1  g0017(.A1(new_n214), .A2(new_n215), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  AOI211_X1 g0018(.A(new_n213), .B(new_n218), .C1(G87), .C2(G250), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G50), .A2(G226), .ZN(new_n220));
  AND2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(G58), .ZN(new_n222));
  INV_X1    g0022(.A(G232), .ZN(new_n223));
  INV_X1    g0023(.A(G107), .ZN(new_n224));
  INV_X1    g0024(.A(G264), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n221), .B1(new_n222), .B2(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  AND2_X1   g0026(.A1(G68), .A2(G238), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n209), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT1), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n230), .A2(new_n207), .ZN(new_n231));
  OAI21_X1  g0031(.A(G50), .B1(G58), .B2(G68), .ZN(new_n232));
  INV_X1    g0032(.A(new_n232), .ZN(new_n233));
  AOI211_X1 g0033(.A(new_n212), .B(new_n229), .C1(new_n231), .C2(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G250), .B(G257), .Z(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XNOR2_X1  g0042(.A(G50), .B(G58), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(KEYINPUT64), .ZN(new_n244));
  XOR2_X1   g0044(.A(G68), .B(G77), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G87), .B(G97), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(G116), .ZN(new_n248));
  XNOR2_X1  g0048(.A(KEYINPUT65), .B(G107), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n246), .B(new_n250), .ZN(G351));
  INV_X1    g0051(.A(KEYINPUT14), .ZN(new_n252));
  OAI21_X1  g0052(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n253));
  INV_X1    g0053(.A(G274), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G33), .ZN(new_n256));
  INV_X1    g0056(.A(G41), .ZN(new_n257));
  OAI211_X1 g0057(.A(G1), .B(G13), .C1(new_n256), .C2(new_n257), .ZN(new_n258));
  AND2_X1   g0058(.A1(new_n258), .A2(new_n253), .ZN(new_n259));
  XNOR2_X1  g0059(.A(new_n259), .B(KEYINPUT66), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n255), .B1(new_n260), .B2(G238), .ZN(new_n261));
  NAND2_X1  g0061(.A1(G33), .A2(G97), .ZN(new_n262));
  XNOR2_X1  g0062(.A(KEYINPUT3), .B(G33), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n223), .A2(G1698), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n265), .B1(G226), .B2(G1698), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n262), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  OR2_X1    g0067(.A1(new_n267), .A2(KEYINPUT71), .ZN(new_n268));
  INV_X1    g0068(.A(new_n258), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n267), .A2(KEYINPUT71), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n268), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n261), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(KEYINPUT13), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT13), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n261), .A2(new_n274), .A3(new_n271), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n252), .B1(new_n276), .B2(G169), .ZN(new_n277));
  INV_X1    g0077(.A(G169), .ZN(new_n278));
  AOI211_X1 g0078(.A(KEYINPUT14), .B(new_n278), .C1(new_n273), .C2(new_n275), .ZN(new_n279));
  INV_X1    g0079(.A(G179), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n276), .A2(new_n280), .ZN(new_n281));
  NOR3_X1   g0081(.A1(new_n277), .A2(new_n279), .A3(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(new_n230), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n207), .A2(new_n256), .ZN(new_n286));
  OAI22_X1  g0086(.A1(new_n286), .A2(new_n202), .B1(new_n207), .B2(G68), .ZN(new_n287));
  NOR3_X1   g0087(.A1(new_n256), .A2(new_n214), .A3(G20), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n285), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  XNOR2_X1  g0089(.A(new_n289), .B(KEYINPUT11), .ZN(new_n290));
  INV_X1    g0090(.A(G68), .ZN(new_n291));
  INV_X1    g0091(.A(new_n285), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n292), .B1(G1), .B2(new_n207), .ZN(new_n293));
  INV_X1    g0093(.A(G13), .ZN(new_n294));
  NOR3_X1   g0094(.A1(new_n294), .A2(new_n207), .A3(G1), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(new_n291), .ZN(new_n296));
  AND2_X1   g0096(.A1(new_n296), .A2(KEYINPUT12), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n296), .A2(KEYINPUT12), .ZN(new_n298));
  OAI221_X1 g0098(.A(new_n290), .B1(new_n291), .B2(new_n293), .C1(new_n297), .C2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n283), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n276), .A2(G200), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(KEYINPUT72), .ZN(new_n302));
  INV_X1    g0102(.A(new_n299), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n273), .A2(G190), .A3(new_n275), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT72), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n276), .A2(new_n305), .A3(G200), .ZN(new_n306));
  NAND4_X1  g0106(.A1(new_n302), .A2(new_n303), .A3(new_n304), .A4(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n300), .A2(new_n307), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n295), .A2(G50), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n309), .B1(new_n293), .B2(G50), .ZN(new_n310));
  XNOR2_X1  g0110(.A(new_n310), .B(KEYINPUT68), .ZN(new_n311));
  OR3_X1    g0111(.A1(new_n222), .A2(KEYINPUT67), .A3(KEYINPUT8), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n222), .A2(KEYINPUT8), .ZN(new_n313));
  AOI21_X1  g0113(.A(KEYINPUT67), .B1(new_n222), .B2(KEYINPUT8), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n312), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n256), .A2(G20), .ZN(new_n316));
  INV_X1    g0116(.A(new_n286), .ZN(new_n317));
  AOI22_X1  g0117(.A1(new_n315), .A2(new_n316), .B1(G150), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n203), .A2(G20), .ZN(new_n319));
  AND2_X1   g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n311), .B1(new_n292), .B2(new_n320), .ZN(new_n321));
  XNOR2_X1  g0121(.A(new_n321), .B(KEYINPUT9), .ZN(new_n322));
  NOR2_X1   g0122(.A1(G222), .A2(G1698), .ZN(new_n323));
  INV_X1    g0123(.A(G1698), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n324), .A2(G223), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n263), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  OAI211_X1 g0126(.A(new_n326), .B(new_n269), .C1(G77), .C2(new_n263), .ZN(new_n327));
  INV_X1    g0127(.A(new_n255), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n329), .B1(new_n260), .B2(G226), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(G190), .ZN(new_n331));
  INV_X1    g0131(.A(G200), .ZN(new_n332));
  OAI211_X1 g0132(.A(new_n322), .B(new_n331), .C1(new_n332), .C2(new_n330), .ZN(new_n333));
  XNOR2_X1  g0133(.A(new_n333), .B(KEYINPUT10), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n330), .A2(new_n280), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n321), .B(new_n335), .C1(G169), .C2(new_n330), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(G58), .A2(G68), .ZN(new_n338));
  XNOR2_X1  g0138(.A(new_n338), .B(KEYINPUT75), .ZN(new_n339));
  OAI21_X1  g0139(.A(G20), .B1(new_n339), .B2(new_n201), .ZN(new_n340));
  INV_X1    g0140(.A(G159), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n340), .B1(new_n341), .B2(new_n286), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n256), .A2(KEYINPUT3), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT3), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(G33), .ZN(new_n345));
  AOI21_X1  g0145(.A(G20), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  OAI21_X1  g0146(.A(KEYINPUT76), .B1(new_n346), .B2(KEYINPUT7), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT76), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT7), .ZN(new_n349));
  OAI211_X1 g0149(.A(new_n348), .B(new_n349), .C1(new_n263), .C2(G20), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n347), .A2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT73), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(new_n344), .ZN(new_n353));
  NAND2_X1  g0153(.A1(KEYINPUT73), .A2(KEYINPUT3), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n353), .A2(new_n256), .A3(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(G20), .B1(new_n355), .B2(new_n345), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(KEYINPUT7), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n351), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n342), .B1(new_n358), .B2(G68), .ZN(new_n359));
  OAI21_X1  g0159(.A(KEYINPUT77), .B1(new_n359), .B2(KEYINPUT16), .ZN(new_n360));
  AND2_X1   g0160(.A1(KEYINPUT73), .A2(KEYINPUT3), .ZN(new_n361));
  NOR2_X1   g0161(.A1(KEYINPUT73), .A2(KEYINPUT3), .ZN(new_n362));
  OAI21_X1  g0162(.A(G33), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT74), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n364), .B1(KEYINPUT3), .B2(new_n256), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  OAI211_X1 g0166(.A(new_n364), .B(G33), .C1(new_n361), .C2(new_n362), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n366), .A2(new_n349), .A3(new_n207), .A4(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n256), .B1(new_n353), .B2(new_n354), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n343), .A2(KEYINPUT74), .ZN(new_n370));
  OAI211_X1 g0170(.A(new_n367), .B(new_n207), .C1(new_n369), .C2(new_n370), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n291), .B1(new_n371), .B2(KEYINPUT7), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n342), .B1(new_n368), .B2(new_n372), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n292), .B1(new_n373), .B2(KEYINPUT16), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT77), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT16), .ZN(new_n376));
  AOI22_X1  g0176(.A1(new_n347), .A2(new_n350), .B1(new_n356), .B2(KEYINPUT7), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n377), .A2(new_n291), .ZN(new_n378));
  OAI211_X1 g0178(.A(new_n375), .B(new_n376), .C1(new_n378), .C2(new_n342), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n360), .A2(new_n374), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n293), .A2(new_n315), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n381), .B1(new_n295), .B2(new_n315), .ZN(new_n382));
  XOR2_X1   g0182(.A(new_n382), .B(KEYINPUT78), .Z(new_n383));
  INV_X1    g0183(.A(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT79), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n255), .B1(new_n259), .B2(G232), .ZN(new_n386));
  INV_X1    g0186(.A(G223), .ZN(new_n387));
  AOI22_X1  g0187(.A1(new_n366), .A2(new_n367), .B1(new_n387), .B2(new_n324), .ZN(new_n388));
  OR2_X1    g0188(.A1(new_n324), .A2(G226), .ZN(new_n389));
  AOI22_X1  g0189(.A1(new_n388), .A2(new_n389), .B1(G33), .B2(G87), .ZN(new_n390));
  OAI211_X1 g0190(.A(new_n385), .B(new_n386), .C1(new_n390), .C2(new_n258), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n367), .B1(new_n369), .B2(new_n370), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n387), .A2(new_n324), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n392), .A2(new_n393), .A3(new_n389), .ZN(new_n394));
  NAND2_X1  g0194(.A1(G33), .A2(G87), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n258), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(new_n386), .ZN(new_n397));
  OAI21_X1  g0197(.A(KEYINPUT79), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  AOI21_X1  g0198(.A(G200), .B1(new_n391), .B2(new_n398), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n396), .A2(new_n397), .ZN(new_n400));
  INV_X1    g0200(.A(G190), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n380), .B(new_n384), .C1(new_n399), .C2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT17), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n391), .A2(new_n398), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(new_n332), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(new_n402), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n409), .A2(KEYINPUT17), .A3(new_n384), .A4(new_n380), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n380), .A2(new_n384), .ZN(new_n411));
  AOI22_X1  g0211(.A1(new_n407), .A2(new_n278), .B1(new_n280), .B2(new_n400), .ZN(new_n412));
  AND3_X1   g0212(.A1(new_n411), .A2(KEYINPUT18), .A3(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(KEYINPUT18), .B1(new_n411), .B2(new_n412), .ZN(new_n414));
  OAI211_X1 g0214(.A(new_n406), .B(new_n410), .C1(new_n413), .C2(new_n414), .ZN(new_n415));
  XOR2_X1   g0215(.A(KEYINPUT15), .B(G87), .Z(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(new_n316), .ZN(new_n417));
  XNOR2_X1  g0217(.A(new_n417), .B(KEYINPUT70), .ZN(new_n418));
  XNOR2_X1  g0218(.A(KEYINPUT8), .B(G58), .ZN(new_n419));
  OAI221_X1 g0219(.A(new_n418), .B1(new_n207), .B2(new_n214), .C1(new_n286), .C2(new_n419), .ZN(new_n420));
  AOI22_X1  g0220(.A1(new_n420), .A2(new_n285), .B1(new_n214), .B2(new_n295), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n421), .B1(new_n214), .B2(new_n293), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n260), .A2(G244), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n263), .A2(G232), .A3(new_n324), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n263), .A2(G238), .A3(G1698), .ZN(new_n425));
  XNOR2_X1  g0225(.A(KEYINPUT69), .B(G107), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  OAI211_X1 g0227(.A(new_n424), .B(new_n425), .C1(new_n263), .C2(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n255), .B1(new_n428), .B2(new_n269), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n423), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(new_n278), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n423), .A2(new_n280), .A3(new_n429), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n422), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  OR2_X1    g0234(.A1(new_n415), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n422), .B1(G200), .B2(new_n430), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n423), .A2(G190), .A3(new_n429), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  NOR4_X1   g0239(.A1(new_n308), .A2(new_n337), .A3(new_n435), .A4(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n217), .A2(G1698), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n392), .B(new_n441), .C1(G250), .C2(G1698), .ZN(new_n442));
  NAND2_X1  g0242(.A1(G33), .A2(G294), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n258), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(G45), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n445), .A2(G1), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n257), .A2(KEYINPUT5), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT5), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(G41), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n446), .A2(new_n447), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(new_n258), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n451), .A2(new_n225), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n446), .A2(new_n447), .A3(new_n449), .A4(G274), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  NOR3_X1   g0254(.A1(new_n444), .A2(new_n452), .A3(new_n454), .ZN(new_n455));
  OAI21_X1  g0255(.A(KEYINPUT88), .B1(new_n455), .B2(G200), .ZN(new_n456));
  INV_X1    g0256(.A(new_n452), .ZN(new_n457));
  AND2_X1   g0257(.A1(new_n442), .A2(new_n443), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n457), .B(new_n453), .C1(new_n458), .C2(new_n258), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT88), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n459), .A2(new_n460), .A3(new_n332), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n455), .A2(new_n401), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n456), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n295), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n206), .A2(G33), .ZN(new_n465));
  AND3_X1   g0265(.A1(new_n464), .A2(new_n292), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(G107), .ZN(new_n467));
  XOR2_X1   g0267(.A(KEYINPUT86), .B(KEYINPUT22), .Z(new_n468));
  INV_X1    g0268(.A(G87), .ZN(new_n469));
  NOR4_X1   g0269(.A1(new_n264), .A2(new_n468), .A3(G20), .A4(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n392), .A2(new_n207), .A3(G87), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n470), .B1(new_n471), .B2(KEYINPUT22), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT23), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n473), .A2(new_n224), .A3(G20), .ZN(new_n474));
  NAND2_X1  g0274(.A1(G33), .A2(G116), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n426), .A2(new_n207), .ZN(new_n476));
  OAI221_X1 g0276(.A(new_n474), .B1(G20), .B2(new_n475), .C1(new_n476), .C2(new_n473), .ZN(new_n477));
  OAI21_X1  g0277(.A(KEYINPUT87), .B1(new_n472), .B2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT87), .ZN(new_n479));
  INV_X1    g0279(.A(new_n477), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT22), .ZN(new_n481));
  AOI21_X1  g0281(.A(G20), .B1(new_n366), .B2(new_n367), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n481), .B1(new_n482), .B2(G87), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n479), .B(new_n480), .C1(new_n483), .C2(new_n470), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n478), .A2(KEYINPUT24), .A3(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT24), .ZN(new_n486));
  OAI211_X1 g0286(.A(KEYINPUT87), .B(new_n486), .C1(new_n472), .C2(new_n477), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n485), .A2(new_n285), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n295), .A2(new_n224), .ZN(new_n489));
  XOR2_X1   g0289(.A(new_n489), .B(KEYINPUT25), .Z(new_n490));
  NAND4_X1  g0290(.A1(new_n463), .A2(new_n467), .A3(new_n488), .A4(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n488), .A2(new_n467), .A3(new_n490), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n455), .A2(G169), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n493), .B1(new_n280), .B2(new_n455), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  AND2_X1   g0295(.A1(new_n491), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n317), .A2(G77), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n224), .A2(KEYINPUT6), .A3(G97), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n216), .A2(new_n224), .ZN(new_n499));
  NOR2_X1   g0299(.A1(G97), .A2(G107), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n498), .B1(new_n501), .B2(KEYINPUT6), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(G20), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n497), .B(new_n503), .C1(new_n377), .C2(new_n427), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(new_n285), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n295), .A2(new_n216), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n466), .A2(G97), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n505), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n450), .A2(G257), .A3(new_n258), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT80), .ZN(new_n510));
  AND3_X1   g0310(.A1(new_n509), .A2(new_n510), .A3(new_n453), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n510), .B1(new_n509), .B2(new_n453), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n263), .A2(KEYINPUT4), .A3(G244), .A4(new_n324), .ZN(new_n514));
  NAND2_X1  g0314(.A1(G33), .A2(G283), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n263), .A2(G250), .A3(G1698), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n392), .A2(G244), .A3(new_n324), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT4), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n513), .B1(new_n520), .B2(new_n258), .ZN(new_n521));
  INV_X1    g0321(.A(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n508), .B1(G190), .B2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT81), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n521), .A2(new_n524), .ZN(new_n525));
  OAI211_X1 g0325(.A(KEYINPUT81), .B(new_n513), .C1(new_n520), .C2(new_n258), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n525), .A2(G200), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(KEYINPUT82), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT82), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n525), .A2(new_n529), .A3(G200), .A4(new_n526), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n523), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n450), .A2(G270), .A3(new_n258), .ZN(new_n532));
  INV_X1    g0332(.A(G303), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n263), .A2(new_n533), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n366), .A2(new_n367), .B1(new_n217), .B2(new_n324), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n225), .A2(G1698), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n453), .B(new_n532), .C1(new_n537), .C2(new_n258), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n538), .A2(new_n280), .ZN(new_n539));
  INV_X1    g0339(.A(G116), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n295), .A2(new_n540), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n464), .A2(G116), .A3(new_n292), .A4(new_n465), .ZN(new_n542));
  AOI22_X1  g0342(.A1(new_n284), .A2(new_n230), .B1(G20), .B2(new_n540), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n515), .B(new_n207), .C1(G33), .C2(new_n216), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n543), .A2(KEYINPUT20), .A3(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(new_n545), .ZN(new_n546));
  AOI21_X1  g0346(.A(KEYINPUT20), .B1(new_n543), .B2(new_n544), .ZN(new_n547));
  OAI211_X1 g0347(.A(new_n541), .B(new_n542), .C1(new_n546), .C2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(KEYINPUT85), .ZN(new_n549));
  INV_X1    g0349(.A(new_n547), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n545), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT85), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n551), .A2(new_n552), .A3(new_n541), .A4(new_n542), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n549), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n539), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n538), .A2(new_n554), .A3(G169), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT21), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n538), .A2(G200), .ZN(new_n559));
  INV_X1    g0359(.A(new_n554), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n217), .A2(new_n324), .ZN(new_n561));
  AND3_X1   g0361(.A1(new_n392), .A2(new_n561), .A3(new_n536), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n269), .B1(new_n562), .B2(new_n534), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n563), .A2(G190), .A3(new_n453), .A4(new_n532), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n559), .A2(new_n560), .A3(new_n564), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n538), .A2(new_n554), .A3(KEYINPUT21), .A4(G169), .ZN(new_n566));
  AND4_X1   g0366(.A1(new_n555), .A2(new_n558), .A3(new_n565), .A4(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n521), .A2(new_n278), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n280), .B(new_n513), .C1(new_n520), .C2(new_n258), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n508), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n466), .A2(G87), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n464), .A2(new_n416), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n482), .A2(G68), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n224), .A2(KEYINPUT69), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT69), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(G107), .ZN(new_n576));
  AOI21_X1  g0376(.A(G97), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n469), .A2(KEYINPUT84), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT84), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(G87), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n207), .B1(new_n577), .B2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT19), .ZN(new_n583));
  INV_X1    g0383(.A(new_n262), .ZN(new_n584));
  NOR3_X1   g0384(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  NOR3_X1   g0385(.A1(new_n262), .A2(KEYINPUT19), .A3(G20), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n573), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n572), .B1(new_n587), .B2(new_n285), .ZN(new_n588));
  NOR2_X1   g0388(.A1(G238), .A2(G1698), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n324), .A2(G244), .ZN(new_n590));
  AOI211_X1 g0390(.A(new_n589), .B(new_n590), .C1(new_n366), .C2(new_n367), .ZN(new_n591));
  INV_X1    g0391(.A(new_n475), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n269), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n446), .A2(G274), .ZN(new_n594));
  XNOR2_X1  g0394(.A(new_n594), .B(KEYINPUT83), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n258), .B(G250), .C1(G1), .C2(new_n445), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(new_n597), .ZN(new_n598));
  AOI21_X1  g0398(.A(G200), .B1(new_n593), .B2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(new_n589), .ZN(new_n600));
  INV_X1    g0400(.A(new_n590), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n392), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n258), .B1(new_n602), .B2(new_n475), .ZN(new_n603));
  NOR3_X1   g0403(.A1(new_n603), .A2(G190), .A3(new_n597), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n571), .B(new_n588), .C1(new_n599), .C2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(new_n572), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n466), .A2(new_n416), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n575), .A2(G107), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n224), .A2(KEYINPUT69), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n216), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  AND2_X1   g0410(.A1(new_n578), .A2(new_n580), .ZN(new_n611));
  OAI21_X1  g0411(.A(G20), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n612), .A2(KEYINPUT19), .A3(new_n262), .ZN(new_n613));
  INV_X1    g0413(.A(new_n586), .ZN(new_n614));
  AOI22_X1  g0414(.A1(new_n613), .A2(new_n614), .B1(G68), .B2(new_n482), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n606), .B(new_n607), .C1(new_n615), .C2(new_n292), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n593), .A2(new_n280), .A3(new_n598), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n278), .B1(new_n603), .B2(new_n597), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n616), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n605), .A2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  AND4_X1   g0421(.A1(new_n531), .A2(new_n567), .A3(new_n570), .A4(new_n621), .ZN(new_n622));
  AND3_X1   g0422(.A1(new_n440), .A2(new_n496), .A3(new_n622), .ZN(G372));
  NOR2_X1   g0423(.A1(new_n413), .A2(new_n414), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n307), .A2(new_n434), .ZN(new_n626));
  AND2_X1   g0426(.A1(new_n300), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n406), .A2(new_n410), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n625), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  OR2_X1    g0429(.A1(new_n629), .A2(KEYINPUT93), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(KEYINPUT93), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n630), .A2(new_n334), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(new_n336), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n440), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT91), .ZN(new_n636));
  XNOR2_X1  g0436(.A(new_n570), .B(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n620), .A2(KEYINPUT89), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT89), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n605), .A2(new_n619), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(KEYINPUT26), .B1(new_n637), .B2(new_n641), .ZN(new_n642));
  AOI22_X1  g0442(.A1(new_n504), .A2(new_n285), .B1(new_n216), .B2(new_n295), .ZN(new_n643));
  AOI22_X1  g0443(.A1(new_n643), .A2(new_n507), .B1(new_n278), .B2(new_n521), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n644), .A2(new_n569), .A3(new_n605), .A4(new_n619), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT26), .ZN(new_n646));
  OAI21_X1  g0446(.A(KEYINPUT92), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT92), .ZN(new_n648));
  INV_X1    g0448(.A(new_n570), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n621), .A2(new_n648), .A3(KEYINPUT26), .A4(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n619), .B1(new_n642), .B2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT90), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n641), .A2(new_n491), .A3(new_n531), .A4(new_n570), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n558), .A2(new_n555), .A3(new_n566), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n655), .B1(new_n492), .B2(new_n494), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n653), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  AND3_X1   g0457(.A1(new_n605), .A2(new_n639), .A3(new_n619), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n639), .B1(new_n605), .B2(new_n619), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n570), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  AND3_X1   g0460(.A1(new_n523), .A2(new_n528), .A3(new_n530), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n656), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n662), .A2(KEYINPUT90), .A3(new_n491), .A4(new_n663), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n652), .B1(new_n657), .B2(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n634), .B1(new_n635), .B2(new_n665), .ZN(G369));
  NOR2_X1   g0466(.A1(new_n294), .A2(G20), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(new_n206), .ZN(new_n668));
  OR2_X1    g0468(.A1(new_n668), .A2(KEYINPUT27), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(KEYINPUT27), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n669), .A2(G213), .A3(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(G343), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n492), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n496), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n673), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n675), .B1(new_n495), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n554), .A2(new_n673), .ZN(new_n678));
  XNOR2_X1  g0478(.A(new_n678), .B(KEYINPUT94), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n567), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n655), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n680), .B1(new_n681), .B2(new_n679), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(G330), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n677), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n681), .A2(new_n673), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n496), .A2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n495), .A2(new_n673), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n685), .A2(new_n690), .ZN(G399));
  NAND2_X1  g0491(.A1(new_n210), .A2(new_n257), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(G1), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n577), .A2(new_n540), .A3(new_n581), .ZN(new_n694));
  OAI22_X1  g0494(.A1(new_n693), .A2(new_n694), .B1(new_n232), .B2(new_n692), .ZN(new_n695));
  XNOR2_X1  g0495(.A(new_n695), .B(KEYINPUT28), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT96), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n664), .A2(new_n657), .ZN(new_n698));
  INV_X1    g0498(.A(new_n619), .ZN(new_n699));
  INV_X1    g0499(.A(new_n651), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n658), .A2(new_n659), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n644), .A2(new_n636), .A3(new_n569), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n570), .A2(KEYINPUT91), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n646), .B1(new_n701), .B2(new_n704), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n699), .B1(new_n700), .B2(new_n705), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n673), .B1(new_n698), .B2(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n697), .B1(new_n707), .B2(KEYINPUT29), .ZN(new_n708));
  OAI21_X1  g0508(.A(KEYINPUT26), .B1(new_n701), .B2(new_n704), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n645), .A2(KEYINPUT26), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n710), .A2(new_n699), .ZN(new_n711));
  OAI211_X1 g0511(.A(new_n709), .B(new_n711), .C1(new_n654), .C2(new_n656), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n712), .A2(KEYINPUT29), .A3(new_n676), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT29), .ZN(new_n714));
  OAI211_X1 g0514(.A(KEYINPUT96), .B(new_n714), .C1(new_n665), .C2(new_n673), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n708), .A2(new_n713), .A3(new_n715), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n622), .A2(new_n496), .A3(new_n676), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n444), .A2(new_n452), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n603), .A2(new_n597), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  OR2_X1    g0520(.A1(new_n720), .A2(KEYINPUT95), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n521), .B1(new_n720), .B2(KEYINPUT95), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n721), .A2(new_n539), .A3(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT30), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n721), .A2(new_n722), .A3(KEYINPUT30), .A4(new_n539), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n522), .A2(G179), .ZN(new_n727));
  INV_X1    g0527(.A(new_n719), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n727), .A2(new_n459), .A3(new_n728), .A4(new_n538), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n725), .A2(new_n726), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(new_n673), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n717), .A2(KEYINPUT31), .A3(new_n731), .ZN(new_n732));
  OR2_X1    g0532(.A1(new_n731), .A2(KEYINPUT31), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(G330), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n716), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n696), .B1(new_n739), .B2(G1), .ZN(G364));
  AOI21_X1  g0540(.A(new_n693), .B1(G45), .B2(new_n667), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n684), .A2(new_n741), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n742), .B1(G330), .B2(new_n682), .ZN(new_n743));
  NOR2_X1   g0543(.A1(G13), .A2(G33), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(G20), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  OR2_X1    g0547(.A1(new_n682), .A2(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n230), .B1(G20), .B2(new_n278), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n207), .A2(new_n401), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n280), .A2(new_n332), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(G326), .ZN(new_n753));
  NOR2_X1   g0553(.A1(G179), .A2(G200), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n207), .B1(new_n754), .B2(G190), .ZN(new_n755));
  INV_X1    g0555(.A(G294), .ZN(new_n756));
  OAI22_X1  g0556(.A1(new_n752), .A2(new_n753), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  XNOR2_X1  g0557(.A(new_n757), .B(KEYINPUT98), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n207), .A2(G190), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n280), .A2(G200), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(G311), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n759), .A2(new_n754), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  AOI211_X1 g0565(.A(new_n263), .B(new_n763), .C1(G329), .C2(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n751), .A2(new_n759), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  XNOR2_X1  g0568(.A(KEYINPUT33), .B(G317), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n750), .A2(new_n760), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  AOI22_X1  g0571(.A1(new_n768), .A2(new_n769), .B1(new_n771), .B2(G322), .ZN(new_n772));
  INV_X1    g0572(.A(G283), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n759), .A2(new_n280), .A3(G200), .ZN(new_n774));
  OR2_X1    g0574(.A1(new_n774), .A2(KEYINPUT97), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n774), .A2(KEYINPUT97), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  OAI211_X1 g0577(.A(new_n766), .B(new_n772), .C1(new_n773), .C2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n750), .ZN(new_n779));
  NOR3_X1   g0579(.A1(new_n779), .A2(new_n332), .A3(G179), .ZN(new_n780));
  AOI211_X1 g0580(.A(new_n758), .B(new_n778), .C1(G303), .C2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n777), .ZN(new_n782));
  AOI22_X1  g0582(.A1(new_n782), .A2(G107), .B1(G68), .B2(new_n768), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n783), .B1(new_n202), .B2(new_n752), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n755), .A2(new_n216), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n764), .A2(new_n341), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(KEYINPUT32), .ZN(new_n788));
  INV_X1    g0588(.A(new_n761), .ZN(new_n789));
  AOI22_X1  g0589(.A1(G58), .A2(new_n771), .B1(new_n789), .B2(G77), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n788), .A2(new_n790), .A3(new_n263), .ZN(new_n791));
  INV_X1    g0591(.A(new_n780), .ZN(new_n792));
  OAI22_X1  g0592(.A1(new_n792), .A2(new_n581), .B1(new_n787), .B2(KEYINPUT32), .ZN(new_n793));
  NOR4_X1   g0593(.A1(new_n784), .A2(new_n785), .A3(new_n791), .A4(new_n793), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n749), .B1(new_n781), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n233), .A2(new_n445), .ZN(new_n796));
  INV_X1    g0596(.A(new_n392), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n797), .A2(new_n210), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  OAI211_X1 g0599(.A(new_n796), .B(new_n799), .C1(new_n246), .C2(new_n445), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n210), .A2(G355), .A3(new_n263), .ZN(new_n801));
  OAI211_X1 g0601(.A(new_n800), .B(new_n801), .C1(G116), .C2(new_n210), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n746), .A2(new_n749), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND4_X1  g0604(.A1(new_n748), .A2(new_n795), .A3(new_n804), .A4(new_n741), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n743), .A2(new_n805), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n806), .B(KEYINPUT99), .ZN(G396));
  NOR2_X1   g0607(.A1(new_n433), .A2(new_n673), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n422), .A2(new_n673), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n438), .A2(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n808), .B1(new_n810), .B2(new_n433), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n707), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n810), .A2(new_n433), .ZN(new_n813));
  INV_X1    g0613(.A(new_n808), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  AOI211_X1 g0615(.A(new_n673), .B(new_n815), .C1(new_n698), .C2(new_n706), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n812), .A2(new_n816), .ZN(new_n817));
  XNOR2_X1  g0617(.A(new_n817), .B(new_n736), .ZN(new_n818));
  OR2_X1    g0618(.A1(new_n818), .A2(new_n741), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n815), .A2(new_n744), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n777), .A2(new_n469), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n821), .A2(new_n263), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n771), .A2(G294), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n785), .B1(G283), .B2(new_n768), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n761), .A2(new_n540), .ZN(new_n825));
  OAI22_X1  g0625(.A1(new_n752), .A2(new_n533), .B1(new_n764), .B2(new_n762), .ZN(new_n826));
  AOI211_X1 g0626(.A(new_n825), .B(new_n826), .C1(G107), .C2(new_n780), .ZN(new_n827));
  NAND4_X1  g0627(.A1(new_n822), .A2(new_n823), .A3(new_n824), .A4(new_n827), .ZN(new_n828));
  XOR2_X1   g0628(.A(KEYINPUT100), .B(G143), .Z(new_n829));
  AOI22_X1  g0629(.A1(new_n771), .A2(new_n829), .B1(new_n789), .B2(G159), .ZN(new_n830));
  INV_X1    g0630(.A(G137), .ZN(new_n831));
  INV_X1    g0631(.A(G150), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n830), .B1(new_n831), .B2(new_n752), .C1(new_n832), .C2(new_n767), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT34), .ZN(new_n834));
  OR2_X1    g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n780), .A2(G50), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n755), .A2(new_n222), .ZN(new_n837));
  AOI211_X1 g0637(.A(new_n837), .B(new_n797), .C1(G132), .C2(new_n765), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n782), .A2(G68), .ZN(new_n839));
  NAND4_X1  g0639(.A1(new_n835), .A2(new_n836), .A3(new_n838), .A4(new_n839), .ZN(new_n840));
  AND2_X1   g0640(.A1(new_n833), .A2(new_n834), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n828), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(new_n749), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n749), .A2(new_n744), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(new_n214), .ZN(new_n845));
  NAND4_X1  g0645(.A1(new_n820), .A2(new_n741), .A3(new_n843), .A4(new_n845), .ZN(new_n846));
  AND2_X1   g0646(.A1(new_n819), .A2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(G384));
  AOI21_X1  g0648(.A(new_n540), .B1(new_n502), .B2(KEYINPUT35), .ZN(new_n849));
  OAI211_X1 g0649(.A(new_n849), .B(new_n231), .C1(KEYINPUT35), .C2(new_n502), .ZN(new_n850));
  XNOR2_X1  g0650(.A(new_n850), .B(KEYINPUT36), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n233), .A2(G77), .ZN(new_n852));
  OAI22_X1  g0652(.A1(new_n339), .A2(new_n852), .B1(G50), .B2(new_n291), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n853), .A2(G1), .A3(new_n294), .ZN(new_n854));
  NAND4_X1  g0654(.A1(new_n708), .A2(new_n440), .A3(new_n713), .A4(new_n715), .ZN(new_n855));
  OR2_X1    g0655(.A1(new_n855), .A2(KEYINPUT103), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n855), .A2(KEYINPUT103), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n633), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n671), .ZN(new_n859));
  OR2_X1    g0659(.A1(new_n373), .A2(KEYINPUT16), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n383), .B1(new_n860), .B2(new_n374), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n415), .A2(new_n859), .A3(new_n862), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n412), .A2(new_n859), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n404), .B1(new_n864), .B2(new_n861), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(KEYINPUT37), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n411), .A2(new_n412), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n411), .A2(new_n859), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT37), .ZN(new_n869));
  NAND4_X1  g0669(.A1(new_n867), .A2(new_n868), .A3(new_n869), .A4(new_n404), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n866), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n863), .A2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT38), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n863), .A2(new_n871), .A3(KEYINPUT38), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n283), .A2(new_n299), .A3(new_n673), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n299), .A2(new_n673), .ZN(new_n878));
  OAI211_X1 g0678(.A(new_n307), .B(new_n878), .C1(new_n282), .C2(new_n303), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  OAI211_X1 g0680(.A(new_n876), .B(new_n880), .C1(new_n816), .C2(new_n808), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n625), .A2(new_n859), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT39), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n884), .B1(new_n874), .B2(new_n875), .ZN(new_n885));
  AND3_X1   g0685(.A1(new_n863), .A2(new_n871), .A3(KEYINPUT38), .ZN(new_n886));
  INV_X1    g0686(.A(new_n868), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n887), .B1(new_n624), .B2(new_n628), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(KEYINPUT102), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT102), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n415), .A2(new_n890), .A3(new_n887), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n867), .A2(new_n868), .A3(new_n404), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(KEYINPUT37), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n893), .A2(KEYINPUT101), .A3(new_n870), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT101), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n892), .A2(new_n895), .A3(KEYINPUT37), .ZN(new_n896));
  NAND4_X1  g0696(.A1(new_n889), .A2(new_n891), .A3(new_n894), .A4(new_n896), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n886), .B1(new_n897), .B2(new_n873), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n885), .B1(new_n898), .B2(new_n884), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n300), .A2(new_n673), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n881), .B(new_n883), .C1(new_n899), .C2(new_n901), .ZN(new_n902));
  XOR2_X1   g0702(.A(new_n858), .B(new_n902), .Z(new_n903));
  INV_X1    g0703(.A(new_n734), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT40), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n894), .A2(new_n896), .ZN(new_n906));
  AND3_X1   g0706(.A1(new_n415), .A2(new_n890), .A3(new_n887), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n890), .B1(new_n415), .B2(new_n887), .ZN(new_n908));
  NOR3_X1   g0708(.A1(new_n906), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n875), .B1(new_n909), .B2(KEYINPUT38), .ZN(new_n910));
  NAND4_X1  g0710(.A1(new_n732), .A2(new_n733), .A3(new_n811), .A4(new_n880), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(KEYINPUT104), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n905), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(KEYINPUT38), .B1(new_n863), .B2(new_n871), .ZN(new_n914));
  NOR3_X1   g0714(.A1(new_n886), .A2(new_n914), .A3(KEYINPUT40), .ZN(new_n915));
  NAND2_X1  g0715(.A1(KEYINPUT104), .A2(KEYINPUT40), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  NOR3_X1   g0717(.A1(new_n915), .A2(new_n911), .A3(new_n917), .ZN(new_n918));
  OAI211_X1 g0718(.A(new_n440), .B(new_n904), .C1(new_n913), .C2(new_n918), .ZN(new_n919));
  AND2_X1   g0719(.A1(new_n911), .A2(KEYINPUT104), .ZN(new_n920));
  OAI21_X1  g0720(.A(KEYINPUT40), .B1(new_n920), .B2(new_n898), .ZN(new_n921));
  OR3_X1    g0721(.A1(new_n915), .A2(new_n911), .A3(new_n917), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n735), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n736), .A2(new_n440), .ZN(new_n924));
  INV_X1    g0724(.A(new_n924), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n919), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  OAI22_X1  g0726(.A1(new_n903), .A2(new_n926), .B1(new_n206), .B2(new_n667), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n927), .B(KEYINPUT105), .ZN(new_n928));
  AND2_X1   g0728(.A1(new_n903), .A2(new_n926), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n851), .B(new_n854), .C1(new_n928), .C2(new_n929), .ZN(G367));
  AOI21_X1  g0730(.A(new_n206), .B1(new_n667), .B2(G45), .ZN(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n508), .A2(new_n673), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n531), .A2(new_n570), .A3(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n934), .B1(new_n570), .B2(new_n676), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n690), .A2(new_n935), .ZN(new_n936));
  XOR2_X1   g0736(.A(new_n936), .B(KEYINPUT45), .Z(new_n937));
  NOR2_X1   g0737(.A1(new_n690), .A2(new_n935), .ZN(new_n938));
  XNOR2_X1  g0738(.A(KEYINPUT107), .B(KEYINPUT44), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n938), .B(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n937), .A2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n685), .ZN(new_n942));
  AOI21_X1  g0742(.A(KEYINPUT108), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n941), .B(new_n942), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n943), .B1(new_n944), .B2(KEYINPUT108), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n687), .B1(new_n677), .B2(new_n686), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n946), .B(new_n683), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n738), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n945), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n949), .A2(new_n739), .ZN(new_n950));
  XOR2_X1   g0750(.A(new_n692), .B(KEYINPUT41), .Z(new_n951));
  AOI21_X1  g0751(.A(new_n932), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n688), .A2(new_n935), .ZN(new_n953));
  XOR2_X1   g0753(.A(new_n953), .B(KEYINPUT42), .Z(new_n954));
  OAI21_X1  g0754(.A(new_n570), .B1(new_n934), .B2(new_n495), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n955), .A2(new_n676), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n588), .A2(new_n571), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n958), .A2(new_n673), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n641), .A2(new_n959), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n699), .A2(new_n958), .A3(new_n673), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n957), .A2(KEYINPUT43), .A3(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(KEYINPUT43), .B2(new_n962), .ZN(new_n964));
  AOI21_X1  g0764(.A(KEYINPUT106), .B1(new_n954), .B2(new_n956), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n964), .B(new_n965), .Z(new_n966));
  NAND2_X1  g0766(.A1(new_n942), .A2(new_n935), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n966), .B(new_n967), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n962), .A2(new_n747), .ZN(new_n969));
  INV_X1    g0769(.A(new_n752), .ZN(new_n970));
  AOI22_X1  g0770(.A1(G311), .A2(new_n970), .B1(new_n771), .B2(G303), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n971), .B1(new_n756), .B2(new_n767), .ZN(new_n972));
  AOI211_X1 g0772(.A(new_n392), .B(new_n972), .C1(G97), .C2(new_n782), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n765), .A2(G317), .ZN(new_n974));
  OAI22_X1  g0774(.A1(new_n427), .A2(new_n755), .B1(new_n761), .B2(new_n773), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n975), .B(KEYINPUT109), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n780), .A2(G116), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(KEYINPUT46), .ZN(new_n978));
  NAND4_X1  g0778(.A1(new_n973), .A2(new_n974), .A3(new_n976), .A4(new_n978), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n764), .A2(new_n831), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n777), .A2(new_n214), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n981), .A2(new_n264), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n982), .A2(KEYINPUT110), .ZN(new_n983));
  AOI211_X1 g0783(.A(new_n980), .B(new_n983), .C1(G159), .C2(new_n768), .ZN(new_n984));
  OAI22_X1  g0784(.A1(new_n792), .A2(new_n222), .B1(new_n832), .B2(new_n770), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n985), .B1(new_n982), .B2(KEYINPUT110), .ZN(new_n986));
  AOI22_X1  g0786(.A1(new_n970), .A2(new_n829), .B1(new_n789), .B2(G50), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n984), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n755), .A2(new_n291), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n979), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  XOR2_X1   g0790(.A(new_n990), .B(KEYINPUT111), .Z(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT47), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n992), .A2(new_n749), .ZN(new_n993));
  INV_X1    g0793(.A(new_n416), .ZN(new_n994));
  OAI221_X1 g0794(.A(new_n803), .B1(new_n210), .B2(new_n994), .C1(new_n798), .C2(new_n241), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n993), .A2(new_n741), .A3(new_n995), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n952), .A2(new_n968), .B1(new_n969), .B2(new_n996), .ZN(G387));
  OR2_X1    g0797(.A1(new_n677), .A2(new_n747), .ZN(new_n998));
  AOI22_X1  g0798(.A1(new_n782), .A2(G97), .B1(new_n315), .B2(new_n768), .ZN(new_n999));
  OAI221_X1 g0799(.A(new_n999), .B1(new_n202), .B2(new_n770), .C1(new_n291), .C2(new_n761), .ZN(new_n1000));
  AOI211_X1 g0800(.A(new_n797), .B(new_n1000), .C1(G150), .C2(new_n765), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT112), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n1002), .B1(new_n970), .B2(G159), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1003), .B1(G77), .B2(new_n780), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n970), .A2(new_n1002), .A3(G159), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n755), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1006), .A2(new_n416), .ZN(new_n1007));
  NAND4_X1  g0807(.A1(new_n1001), .A2(new_n1004), .A3(new_n1005), .A4(new_n1007), .ZN(new_n1008));
  XOR2_X1   g0808(.A(new_n1008), .B(KEYINPUT113), .Z(new_n1009));
  OAI21_X1  g0809(.A(new_n797), .B1(new_n753), .B2(new_n764), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(G322), .A2(new_n970), .B1(new_n768), .B2(G311), .ZN(new_n1011));
  INV_X1    g0811(.A(G317), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n1011), .B1(new_n533), .B2(new_n761), .C1(new_n1012), .C2(new_n770), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT48), .ZN(new_n1014));
  OR2_X1    g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n780), .A2(G294), .B1(G283), .B2(new_n1006), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1017), .B(KEYINPUT114), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1015), .A2(new_n1016), .A3(new_n1018), .ZN(new_n1019));
  XOR2_X1   g0819(.A(new_n1019), .B(KEYINPUT49), .Z(new_n1020));
  AOI211_X1 g0820(.A(new_n1010), .B(new_n1020), .C1(G116), .C2(new_n782), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n749), .B1(new_n1009), .B2(new_n1021), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n419), .A2(G50), .ZN(new_n1023));
  XOR2_X1   g0823(.A(new_n1023), .B(KEYINPUT50), .Z(new_n1024));
  NOR2_X1   g0824(.A1(new_n291), .A2(new_n214), .ZN(new_n1025));
  NOR4_X1   g0825(.A1(new_n1024), .A2(G45), .A3(new_n1025), .A4(new_n694), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n799), .B1(new_n238), .B2(new_n445), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n694), .A2(new_n210), .A3(new_n263), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1026), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n210), .A2(G107), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n803), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n998), .A2(new_n1022), .A3(new_n741), .A4(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n692), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n947), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1033), .B1(new_n739), .B2(new_n1034), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n1032), .B1(new_n931), .B2(new_n947), .C1(new_n1035), .C2(new_n948), .ZN(G393));
  OAI21_X1  g0836(.A(new_n944), .B1(new_n738), .B2(new_n947), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n949), .A2(new_n1033), .A3(new_n1037), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n944), .A2(new_n931), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n777), .A2(new_n224), .B1(new_n756), .B2(new_n761), .ZN(new_n1040));
  AOI211_X1 g0840(.A(new_n263), .B(new_n1040), .C1(G303), .C2(new_n768), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n765), .A2(G322), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n752), .A2(new_n1012), .B1(new_n770), .B2(new_n762), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT52), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n780), .A2(G283), .B1(G116), .B2(new_n1006), .ZN(new_n1045));
  NAND4_X1  g0845(.A1(new_n1041), .A2(new_n1042), .A3(new_n1044), .A4(new_n1045), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n767), .A2(new_n202), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n821), .B1(G68), .B2(new_n780), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n752), .A2(new_n832), .B1(new_n770), .B2(new_n341), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT51), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1006), .A2(G77), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n761), .A2(new_n419), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n1052), .B(new_n797), .C1(new_n765), .C2(new_n829), .ZN(new_n1053));
  NAND4_X1  g0853(.A1(new_n1048), .A2(new_n1050), .A3(new_n1051), .A4(new_n1053), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1046), .B1(new_n1047), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1055), .A2(new_n749), .ZN(new_n1056));
  OR2_X1    g0856(.A1(new_n935), .A2(new_n747), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n803), .B1(new_n216), .B2(new_n210), .C1(new_n250), .C2(new_n798), .ZN(new_n1058));
  AND3_X1   g0858(.A1(new_n1057), .A2(new_n741), .A3(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1039), .B1(new_n1056), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1038), .A2(new_n1060), .ZN(G390));
  NAND4_X1  g0861(.A1(new_n732), .A2(new_n733), .A3(G330), .A4(new_n811), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n880), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n712), .A2(new_n676), .A3(new_n813), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1063), .B1(new_n1065), .B2(new_n814), .ZN(new_n1066));
  NOR3_X1   g0866(.A1(new_n898), .A2(new_n1066), .A3(new_n900), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n808), .B1(new_n707), .B2(new_n811), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n901), .B1(new_n1068), .B2(new_n1063), .ZN(new_n1069));
  AOI211_X1 g0869(.A(new_n1064), .B(new_n1067), .C1(new_n1069), .C2(new_n899), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n1064), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n698), .A2(new_n706), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1072), .A2(new_n676), .A3(new_n811), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1063), .B1(new_n1073), .B2(new_n814), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n899), .B1(new_n1074), .B2(new_n900), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1067), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1071), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n1070), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n899), .A2(new_n744), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n782), .A2(G50), .B1(G125), .B2(new_n765), .ZN(new_n1080));
  XOR2_X1   g0880(.A(KEYINPUT54), .B(G143), .Z(new_n1081));
  NAND2_X1  g0881(.A1(new_n789), .A2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1080), .A2(new_n263), .A3(new_n1082), .ZN(new_n1083));
  AND2_X1   g0883(.A1(new_n970), .A2(G128), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n780), .A2(G150), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1085), .B(KEYINPUT53), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(G132), .A2(new_n771), .B1(new_n768), .B2(G137), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1087), .B1(new_n341), .B2(new_n755), .ZN(new_n1088));
  NOR4_X1   g0888(.A1(new_n1083), .A2(new_n1084), .A3(new_n1086), .A4(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n839), .A2(new_n1051), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n752), .A2(new_n773), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n263), .B1(new_n768), .B2(new_n426), .ZN(new_n1092));
  OAI221_X1 g0892(.A(new_n1092), .B1(new_n216), .B2(new_n761), .C1(new_n792), .C2(new_n469), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n770), .A2(new_n540), .B1(new_n764), .B2(new_n756), .ZN(new_n1094));
  NOR4_X1   g0894(.A1(new_n1090), .A2(new_n1091), .A3(new_n1093), .A4(new_n1094), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n749), .B1(new_n1089), .B2(new_n1095), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n844), .B(new_n312), .C1(new_n313), .C2(new_n314), .ZN(new_n1097));
  AND3_X1   g0897(.A1(new_n1079), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n1078), .A2(new_n932), .B1(new_n741), .B2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n880), .B1(KEYINPUT115), .B2(new_n811), .ZN(new_n1100));
  XOR2_X1   g0900(.A(new_n1062), .B(new_n1100), .Z(new_n1101));
  NAND3_X1  g0901(.A1(new_n1101), .A2(new_n814), .A3(new_n1065), .ZN(new_n1102));
  AND2_X1   g0902(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n1103), .A2(new_n1064), .B1(new_n808), .B2(new_n816), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1105));
  NAND4_X1  g0905(.A1(new_n1078), .A2(new_n858), .A3(new_n924), .A4(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1106), .A2(new_n1033), .ZN(new_n1107));
  AND2_X1   g0907(.A1(new_n855), .A2(KEYINPUT103), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n855), .A2(KEYINPUT103), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n634), .B(new_n924), .C1(new_n1108), .C2(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1078), .B1(new_n1111), .B2(new_n1105), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1099), .B1(new_n1107), .B2(new_n1112), .ZN(G378));
  NAND2_X1  g0913(.A1(new_n923), .A2(new_n902), .ZN(new_n1114));
  OAI21_X1  g0914(.A(G330), .B1(new_n913), .B2(new_n918), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n910), .A2(KEYINPUT39), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n900), .B1(new_n1116), .B2(new_n885), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n882), .B1(new_n1074), .B2(new_n876), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1115), .A2(new_n1117), .A3(new_n1118), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(new_n337), .B(KEYINPUT119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n321), .A2(new_n859), .ZN(new_n1121));
  OR2_X1    g0921(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1124));
  AND3_X1   g0924(.A1(new_n1122), .A2(new_n1123), .A3(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1124), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1114), .A2(new_n1119), .A3(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1114), .A2(new_n1119), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1127), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n1106), .A2(new_n1111), .B1(new_n1128), .B2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n692), .B1(new_n1132), .B2(KEYINPUT57), .ZN(new_n1133));
  INV_X1    g0933(.A(KEYINPUT57), .ZN(new_n1134));
  AND3_X1   g0934(.A1(new_n1114), .A2(new_n1119), .A3(new_n1127), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1127), .B1(new_n1114), .B2(new_n1119), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1110), .B1(new_n1078), .B2(new_n1105), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1134), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT120), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  OAI211_X1 g0941(.A(KEYINPUT120), .B(new_n1134), .C1(new_n1137), .C2(new_n1138), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1133), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1127), .A2(new_n744), .ZN(new_n1144));
  OAI22_X1  g0944(.A1(new_n994), .A2(new_n761), .B1(new_n216), .B2(new_n767), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(new_n1145), .B(KEYINPUT116), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n797), .A2(new_n257), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1147), .B1(G283), .B2(new_n765), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n782), .A2(G58), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  AOI211_X1 g0950(.A(new_n1146), .B(new_n1150), .C1(G77), .C2(new_n780), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n989), .B1(G116), .B2(new_n970), .ZN(new_n1152));
  XOR2_X1   g0952(.A(new_n1152), .B(KEYINPUT117), .Z(new_n1153));
  OAI211_X1 g0953(.A(new_n1151), .B(new_n1153), .C1(new_n224), .C2(new_n770), .ZN(new_n1154));
  XOR2_X1   g0954(.A(new_n1154), .B(KEYINPUT58), .Z(new_n1155));
  OAI211_X1 g0955(.A(new_n1147), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(G132), .A2(new_n768), .B1(new_n789), .B2(G137), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(new_n970), .A2(G125), .B1(new_n1006), .B2(G150), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n780), .A2(new_n1081), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n771), .A2(G128), .ZN(new_n1160));
  NAND4_X1  g0960(.A1(new_n1157), .A2(new_n1158), .A3(new_n1159), .A4(new_n1160), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(new_n1161), .B(KEYINPUT59), .ZN(new_n1162));
  AOI211_X1 g0962(.A(G33), .B(G41), .C1(new_n765), .C2(G124), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1163), .B1(new_n777), .B2(new_n341), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1156), .B1(new_n1162), .B2(new_n1164), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n749), .B1(new_n1155), .B2(new_n1165), .ZN(new_n1166));
  XOR2_X1   g0966(.A(new_n1166), .B(KEYINPUT118), .Z(new_n1167));
  NAND3_X1  g0967(.A1(new_n1144), .A2(new_n741), .A3(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1168), .B1(new_n202), .B2(new_n844), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1137), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1169), .B1(new_n1170), .B2(new_n932), .ZN(new_n1171));
  AND2_X1   g0971(.A1(new_n1143), .A2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(G375));
  NAND2_X1  g0973(.A1(new_n1111), .A2(new_n1105), .ZN(new_n1174));
  AND2_X1   g0974(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1110), .A2(new_n1175), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1174), .A2(new_n951), .A3(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1105), .A2(new_n932), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1063), .A2(new_n744), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n780), .A2(G97), .B1(G303), .B2(new_n765), .ZN(new_n1180));
  XNOR2_X1  g0980(.A(new_n1180), .B(KEYINPUT121), .ZN(new_n1181));
  AOI211_X1 g0981(.A(new_n981), .B(new_n1181), .C1(G294), .C2(new_n970), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n1182), .B(new_n264), .C1(new_n427), .C2(new_n761), .ZN(new_n1183));
  OAI221_X1 g0983(.A(new_n1007), .B1(new_n540), .B2(new_n767), .C1(new_n773), .C2(new_n770), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n755), .A2(new_n202), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n789), .A2(G150), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n765), .A2(G128), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n768), .A2(new_n1081), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n1149), .A2(new_n1186), .A3(new_n1187), .A4(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1189), .B1(G159), .B2(new_n780), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(G132), .A2(new_n970), .B1(new_n771), .B2(G137), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1190), .A2(new_n392), .A3(new_n1191), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n1183), .A2(new_n1184), .B1(new_n1185), .B2(new_n1192), .ZN(new_n1193));
  XOR2_X1   g0993(.A(new_n1193), .B(KEYINPUT122), .Z(new_n1194));
  NAND2_X1  g0994(.A1(new_n1194), .A2(new_n749), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n844), .A2(new_n291), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n1179), .A2(new_n1195), .A3(new_n741), .A4(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1178), .A2(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1177), .A2(new_n1199), .ZN(G381));
  NOR2_X1   g1000(.A1(G375), .A2(G378), .ZN(new_n1201));
  OR2_X1    g1001(.A1(G393), .A2(G396), .ZN(new_n1202));
  NOR4_X1   g1002(.A1(G387), .A2(G384), .A3(G390), .A4(new_n1202), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1201), .A2(new_n1199), .A3(new_n1177), .A4(new_n1203), .ZN(G407));
  NAND2_X1  g1004(.A1(new_n1201), .A2(new_n672), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(G407), .A2(G213), .A3(new_n1205), .ZN(G409));
  NAND3_X1  g1006(.A1(new_n1143), .A2(G378), .A3(new_n1171), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1207), .A2(KEYINPUT123), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT123), .ZN(new_n1209));
  NAND4_X1  g1009(.A1(new_n1143), .A2(G378), .A3(new_n1209), .A4(new_n1171), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1208), .A2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(G378), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1171), .ZN(new_n1213));
  AND2_X1   g1013(.A1(new_n1132), .A2(new_n951), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1212), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1211), .A2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n672), .A2(G213), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  OAI21_X1  g1018(.A(KEYINPUT60), .B1(new_n1110), .B2(new_n1175), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1219), .A2(new_n1176), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1110), .A2(KEYINPUT60), .A3(new_n1175), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1220), .A2(new_n1033), .A3(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1222), .A2(KEYINPUT124), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT124), .ZN(new_n1224));
  NAND4_X1  g1024(.A1(new_n1220), .A2(new_n1224), .A3(new_n1033), .A4(new_n1221), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1223), .A2(new_n1225), .ZN(new_n1226));
  AOI21_X1  g1026(.A(G384), .B1(new_n1226), .B2(new_n1199), .ZN(new_n1227));
  AOI211_X1 g1027(.A(new_n847), .B(new_n1198), .C1(new_n1223), .C2(new_n1225), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT125), .ZN(new_n1229));
  NOR3_X1   g1029(.A1(new_n1227), .A2(new_n1228), .A3(new_n1229), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1229), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1231));
  INV_X1    g1031(.A(G2897), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1217), .A2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1231), .A2(new_n1233), .ZN(new_n1234));
  OAI221_X1 g1034(.A(new_n1229), .B1(new_n1232), .B2(new_n1217), .C1(new_n1227), .C2(new_n1228), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1230), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(KEYINPUT61), .B1(new_n1218), .B2(new_n1236), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n1211), .A2(new_n1215), .B1(G213), .B2(new_n672), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT62), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1238), .A2(new_n1239), .A3(new_n1240), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1216), .A2(new_n1217), .A3(new_n1240), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(KEYINPUT62), .ZN(new_n1243));
  AND3_X1   g1043(.A1(new_n1237), .A2(new_n1241), .A3(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(G390), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(G387), .A2(new_n1245), .ZN(new_n1246));
  OR2_X1    g1046(.A1(G387), .A2(new_n1245), .ZN(new_n1247));
  XOR2_X1   g1047(.A(G393), .B(G396), .Z(new_n1248));
  INV_X1    g1048(.A(new_n1248), .ZN(new_n1249));
  OR2_X1    g1049(.A1(new_n1249), .A2(KEYINPUT126), .ZN(new_n1250));
  AND2_X1   g1050(.A1(new_n1247), .A2(new_n1250), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(new_n1247), .A2(new_n1249), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1246), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  OR2_X1    g1053(.A1(new_n1246), .A2(new_n1250), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(KEYINPUT61), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT63), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1257), .B1(new_n1218), .B2(new_n1236), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1242), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1256), .B1(new_n1258), .B2(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT127), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1261), .B1(new_n1242), .B2(new_n1257), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1238), .A2(KEYINPUT127), .A3(KEYINPUT63), .A4(new_n1240), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  OAI22_X1  g1064(.A1(new_n1244), .A2(new_n1255), .B1(new_n1260), .B2(new_n1264), .ZN(G405));
  NAND2_X1  g1065(.A1(G375), .A2(new_n1212), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1266), .A2(new_n1211), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1240), .ZN(new_n1268));
  XNOR2_X1  g1068(.A(new_n1267), .B(new_n1268), .ZN(new_n1269));
  XNOR2_X1  g1069(.A(new_n1269), .B(new_n1255), .ZN(G402));
endmodule


