//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 0 0 1 0 0 0 0 0 0 0 0 1 1 0 1 1 0 0 0 1 1 1 0 1 0 1 0 1 0 1 0 0 1 0 0 1 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:54 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n566, new_n567, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n578, new_n579, new_n580,
    new_n581, new_n585, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n630,
    new_n633, new_n635, new_n636, new_n637, new_n638, new_n639, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT65), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT66), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n455), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n453), .A2(G2106), .ZN(new_n459));
  INV_X1    g034(.A(KEYINPUT67), .ZN(new_n460));
  OAI21_X1  g035(.A(new_n458), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  AOI21_X1  g036(.A(new_n461), .B1(new_n460), .B2(new_n459), .ZN(G319));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G125), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n463), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n464), .A2(G2105), .ZN(new_n471));
  AOI22_X1  g046(.A1(new_n470), .A2(G2105), .B1(G101), .B2(new_n471), .ZN(new_n472));
  OAI21_X1  g047(.A(KEYINPUT68), .B1(new_n466), .B2(G2104), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT68), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n474), .A2(new_n464), .A3(KEYINPUT3), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n473), .A2(new_n475), .A3(new_n467), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n476), .A2(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G137), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n472), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G160));
  NAND2_X1  g055(.A1(new_n477), .A2(G136), .ZN(new_n481));
  INV_X1    g056(.A(G2105), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n482), .A2(G112), .ZN(new_n483));
  OAI21_X1  g058(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n481), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND4_X1  g060(.A1(new_n473), .A2(new_n475), .A3(G2105), .A4(new_n467), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(KEYINPUT69), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT69), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n486), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n485), .B1(new_n492), .B2(G124), .ZN(new_n493));
  XOR2_X1   g068(.A(new_n493), .B(KEYINPUT70), .Z(G162));
  OAI21_X1  g069(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT71), .ZN(new_n497));
  INV_X1    g072(.A(G114), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n497), .B1(new_n498), .B2(G2105), .ZN(new_n499));
  NOR3_X1   g074(.A1(new_n482), .A2(KEYINPUT71), .A3(G114), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n496), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(G126), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n501), .B1(new_n486), .B2(new_n502), .ZN(new_n503));
  AND2_X1   g078(.A1(new_n475), .A2(new_n467), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT72), .ZN(new_n505));
  INV_X1    g080(.A(G138), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n506), .A2(G2105), .ZN(new_n507));
  NAND4_X1  g082(.A1(new_n504), .A2(new_n505), .A3(new_n473), .A4(new_n507), .ZN(new_n508));
  NAND4_X1  g083(.A1(new_n473), .A2(new_n475), .A3(new_n467), .A4(new_n507), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(KEYINPUT72), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n508), .A2(KEYINPUT4), .A3(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT4), .ZN(new_n512));
  NAND4_X1  g087(.A1(new_n507), .A2(new_n465), .A3(new_n467), .A4(new_n512), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n503), .B1(new_n511), .B2(new_n513), .ZN(G164));
  INV_X1    g089(.A(G543), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT6), .ZN(new_n516));
  INV_X1    g091(.A(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(KEYINPUT6), .A2(G651), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n515), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G50), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT5), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(new_n515), .ZN(new_n523));
  NAND2_X1  g098(.A1(KEYINPUT5), .A2(G543), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n518), .A2(new_n519), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(G88), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n521), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n525), .A2(G62), .ZN(new_n530));
  NAND2_X1  g105(.A1(G75), .A2(G543), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n517), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n529), .A2(new_n532), .ZN(G166));
  XNOR2_X1  g108(.A(new_n520), .B(KEYINPUT73), .ZN(new_n534));
  INV_X1    g109(.A(G51), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  XNOR2_X1  g111(.A(KEYINPUT74), .B(KEYINPUT7), .ZN(new_n537));
  AND3_X1   g112(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n537), .B(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n526), .A2(G89), .ZN(new_n540));
  NAND2_X1  g115(.A1(G63), .A2(G651), .ZN(new_n541));
  AND2_X1   g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(new_n525), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n539), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n536), .A2(new_n544), .ZN(G168));
  INV_X1    g120(.A(KEYINPUT73), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n520), .B(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G52), .ZN(new_n548));
  NAND2_X1  g123(.A1(G77), .A2(G543), .ZN(new_n549));
  INV_X1    g124(.A(G64), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n549), .B1(new_n543), .B2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(new_n527), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n551), .A2(G651), .B1(new_n552), .B2(G90), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n548), .A2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(G171));
  NAND2_X1  g130(.A1(new_n547), .A2(G43), .ZN(new_n556));
  NAND2_X1  g131(.A1(G68), .A2(G543), .ZN(new_n557));
  INV_X1    g132(.A(G56), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n557), .B1(new_n543), .B2(new_n558), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n559), .A2(G651), .B1(new_n552), .B2(G81), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n556), .A2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(G860), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT75), .ZN(G153));
  NAND4_X1  g139(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g140(.A1(G1), .A2(G3), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT8), .ZN(new_n567));
  NAND4_X1  g142(.A1(G319), .A2(G483), .A3(G661), .A4(new_n567), .ZN(G188));
  NAND2_X1  g143(.A1(new_n552), .A2(G91), .ZN(new_n569));
  XNOR2_X1  g144(.A(KEYINPUT76), .B(G65), .ZN(new_n570));
  NOR2_X1   g145(.A1(new_n543), .A2(new_n570), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n571), .B1(G78), .B2(G543), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n569), .B1(new_n572), .B2(new_n517), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n520), .A2(G53), .ZN(new_n574));
  XOR2_X1   g149(.A(new_n574), .B(KEYINPUT9), .Z(new_n575));
  NOR2_X1   g150(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(G299));
  INV_X1    g152(.A(KEYINPUT77), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n548), .A2(new_n553), .A3(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(new_n579), .ZN(new_n580));
  AOI21_X1  g155(.A(new_n578), .B1(new_n548), .B2(new_n553), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n580), .A2(new_n581), .ZN(G301));
  OR2_X1    g157(.A1(new_n536), .A2(new_n544), .ZN(G286));
  INV_X1    g158(.A(G166), .ZN(G303));
  NAND2_X1  g159(.A1(new_n552), .A2(G87), .ZN(new_n585));
  INV_X1    g160(.A(G74), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n523), .A2(new_n586), .A3(new_n524), .ZN(new_n587));
  AOI22_X1  g162(.A1(G49), .A2(new_n520), .B1(new_n587), .B2(G651), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n585), .A2(new_n588), .ZN(G288));
  INV_X1    g164(.A(KEYINPUT78), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n525), .A2(new_n590), .A3(G61), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(G73), .A2(G543), .ZN(new_n593));
  INV_X1    g168(.A(G61), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n594), .B1(new_n523), .B2(new_n524), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n593), .B1(new_n595), .B2(new_n590), .ZN(new_n596));
  OAI21_X1  g171(.A(G651), .B1(new_n592), .B2(new_n596), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n552), .A2(G86), .B1(G48), .B2(new_n520), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n597), .A2(new_n598), .ZN(G305));
  AND2_X1   g174(.A1(new_n547), .A2(G47), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n525), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n601));
  INV_X1    g176(.A(G85), .ZN(new_n602));
  OAI22_X1  g177(.A1(new_n601), .A2(new_n517), .B1(new_n527), .B2(new_n602), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(G290));
  INV_X1    g180(.A(KEYINPUT10), .ZN(new_n606));
  INV_X1    g181(.A(G92), .ZN(new_n607));
  OAI21_X1  g182(.A(KEYINPUT79), .B1(new_n527), .B2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(new_n609));
  NOR3_X1   g184(.A1(new_n527), .A2(KEYINPUT79), .A3(new_n607), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n606), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(new_n610), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n612), .A2(KEYINPUT10), .A3(new_n608), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  AND2_X1   g189(.A1(new_n525), .A2(G66), .ZN(new_n615));
  NAND2_X1  g190(.A1(G79), .A2(G543), .ZN(new_n616));
  XOR2_X1   g191(.A(new_n616), .B(KEYINPUT80), .Z(new_n617));
  OAI21_X1  g192(.A(G651), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(G54), .ZN(new_n619));
  OAI211_X1 g194(.A(new_n618), .B(KEYINPUT81), .C1(new_n534), .C2(new_n619), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n618), .B1(new_n534), .B2(new_n619), .ZN(new_n621));
  INV_X1    g196(.A(KEYINPUT81), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  AOI21_X1  g198(.A(new_n614), .B1(new_n620), .B2(new_n623), .ZN(new_n624));
  INV_X1    g199(.A(G868), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n626), .B1(new_n625), .B2(G301), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT82), .ZN(G284));
  INV_X1    g203(.A(new_n627), .ZN(G321));
  NAND2_X1  g204(.A1(G286), .A2(G868), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n630), .B1(G868), .B2(new_n576), .ZN(G297));
  OAI21_X1  g206(.A(new_n630), .B1(G868), .B2(new_n576), .ZN(G280));
  INV_X1    g207(.A(G559), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n624), .B1(new_n633), .B2(G860), .ZN(G148));
  NOR2_X1   g209(.A1(new_n561), .A2(G868), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n623), .A2(new_n620), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n636), .A2(new_n613), .A3(new_n611), .ZN(new_n637));
  NOR2_X1   g212(.A1(new_n637), .A2(G559), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT83), .ZN(new_n639));
  AOI21_X1  g214(.A(new_n635), .B1(new_n639), .B2(G868), .ZN(G323));
  XNOR2_X1  g215(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g216(.A1(new_n477), .A2(G135), .ZN(new_n642));
  OAI21_X1  g217(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n643));
  INV_X1    g218(.A(KEYINPUT85), .ZN(new_n644));
  INV_X1    g219(.A(G111), .ZN(new_n645));
  AOI22_X1  g220(.A1(new_n643), .A2(new_n644), .B1(new_n645), .B2(G2105), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n646), .B1(new_n644), .B2(new_n643), .ZN(new_n647));
  INV_X1    g222(.A(G123), .ZN(new_n648));
  OAI211_X1 g223(.A(new_n642), .B(new_n647), .C1(new_n491), .C2(new_n648), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n649), .A2(G2096), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n649), .A2(G2096), .ZN(new_n651));
  XNOR2_X1  g226(.A(KEYINPUT84), .B(KEYINPUT12), .ZN(new_n652));
  NOR3_X1   g227(.A1(new_n466), .A2(new_n464), .A3(G2105), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n652), .B(new_n653), .Z(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT13), .B(G2100), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n650), .A2(new_n651), .A3(new_n656), .ZN(G156));
  XNOR2_X1  g232(.A(KEYINPUT15), .B(G2435), .ZN(new_n658));
  XNOR2_X1  g233(.A(KEYINPUT87), .B(G2438), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n658), .B(new_n659), .Z(new_n660));
  XNOR2_X1  g235(.A(G2427), .B(G2430), .ZN(new_n661));
  OR2_X1    g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n660), .A2(new_n661), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n662), .A2(KEYINPUT14), .A3(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1341), .B(G1348), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2443), .B(G2446), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n664), .B(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(G2451), .B(G2454), .Z(new_n669));
  XNOR2_X1  g244(.A(KEYINPUT86), .B(KEYINPUT16), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n672), .A2(G14), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n668), .A2(new_n671), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n673), .A2(new_n674), .ZN(G401));
  XOR2_X1   g250(.A(KEYINPUT88), .B(KEYINPUT18), .Z(new_n676));
  XOR2_X1   g251(.A(G2084), .B(G2090), .Z(new_n677));
  XNOR2_X1  g252(.A(G2067), .B(G2678), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n679), .A2(KEYINPUT17), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n677), .A2(new_n678), .ZN(new_n681));
  OAI21_X1  g256(.A(new_n676), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT89), .ZN(new_n683));
  XOR2_X1   g258(.A(G2072), .B(G2078), .Z(new_n684));
  INV_X1    g259(.A(new_n676), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n684), .B1(new_n679), .B2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n683), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(G2096), .B(G2100), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(G227));
  XNOR2_X1  g264(.A(G1971), .B(G1976), .ZN(new_n690));
  INV_X1    g265(.A(KEYINPUT19), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XOR2_X1   g267(.A(G1956), .B(G2474), .Z(new_n693));
  XOR2_X1   g268(.A(G1961), .B(G1966), .Z(new_n694));
  AND2_X1   g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n692), .A2(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(KEYINPUT20), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n693), .A2(new_n694), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n695), .A2(new_n699), .ZN(new_n700));
  MUX2_X1   g275(.A(new_n700), .B(new_n699), .S(new_n692), .Z(new_n701));
  NOR2_X1   g276(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(G1981), .ZN(new_n703));
  INV_X1    g278(.A(G1986), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  XOR2_X1   g280(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT90), .ZN(new_n707));
  AND2_X1   g282(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n705), .A2(new_n707), .ZN(new_n709));
  XNOR2_X1  g284(.A(G1991), .B(G1996), .ZN(new_n710));
  INV_X1    g285(.A(new_n710), .ZN(new_n711));
  OR3_X1    g286(.A1(new_n708), .A2(new_n709), .A3(new_n711), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n711), .B1(new_n708), .B2(new_n709), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n712), .A2(new_n713), .ZN(G229));
  INV_X1    g289(.A(G16), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n715), .A2(G21), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(G168), .B2(new_n715), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(KEYINPUT102), .Z(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(G1966), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(KEYINPUT103), .Z(new_n720));
  INV_X1    g295(.A(G29), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n721), .A2(G27), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(G164), .B2(new_n721), .ZN(new_n723));
  INV_X1    g298(.A(G2078), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  AND2_X1   g300(.A1(new_n720), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n721), .A2(G35), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(G162), .B2(new_n721), .ZN(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(new_n729));
  XOR2_X1   g304(.A(KEYINPUT29), .B(G2090), .Z(new_n730));
  OR2_X1    g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n715), .A2(G4), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(new_n624), .B2(new_n715), .ZN(new_n733));
  INV_X1    g308(.A(G1348), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n733), .B(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n729), .A2(new_n730), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n731), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n721), .A2(G32), .ZN(new_n739));
  NAND3_X1  g314(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n740));
  INV_X1    g315(.A(KEYINPUT26), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n740), .A2(new_n741), .ZN(new_n743));
  AOI22_X1  g318(.A1(new_n742), .A2(new_n743), .B1(G105), .B2(new_n471), .ZN(new_n744));
  INV_X1    g319(.A(new_n477), .ZN(new_n745));
  INV_X1    g320(.A(G141), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n744), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n492), .A2(KEYINPUT100), .A3(G129), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT100), .ZN(new_n749));
  INV_X1    g324(.A(G129), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n749), .B1(new_n491), .B2(new_n750), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n747), .B1(new_n748), .B2(new_n751), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n739), .B1(new_n752), .B2(new_n721), .ZN(new_n753));
  XNOR2_X1  g328(.A(KEYINPUT27), .B(G1996), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT101), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n753), .B(new_n755), .Z(new_n756));
  INV_X1    g331(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n718), .A2(G1966), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n715), .A2(G20), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT23), .Z(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(G299), .B2(G16), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(G1956), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n721), .A2(G26), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT28), .Z(new_n764));
  NAND2_X1  g339(.A1(new_n492), .A2(G128), .ZN(new_n765));
  OAI21_X1  g340(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n766));
  INV_X1    g341(.A(G116), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n766), .B1(new_n767), .B2(G2105), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(new_n477), .B2(G140), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n765), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n764), .B1(new_n770), .B2(G29), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(G2067), .ZN(new_n772));
  INV_X1    g347(.A(G19), .ZN(new_n773));
  OR3_X1    g348(.A1(new_n773), .A2(KEYINPUT97), .A3(G16), .ZN(new_n774));
  OAI21_X1  g349(.A(KEYINPUT97), .B1(new_n773), .B2(G16), .ZN(new_n775));
  INV_X1    g350(.A(new_n561), .ZN(new_n776));
  OAI211_X1 g351(.A(new_n774), .B(new_n775), .C1(new_n776), .C2(new_n715), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(G1341), .Z(new_n778));
  NAND2_X1  g353(.A1(new_n721), .A2(G33), .ZN(new_n779));
  NAND2_X1  g354(.A1(G115), .A2(G2104), .ZN(new_n780));
  INV_X1    g355(.A(G127), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n780), .B1(new_n468), .B2(new_n781), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n482), .B1(new_n782), .B2(KEYINPUT99), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(KEYINPUT99), .B2(new_n782), .ZN(new_n784));
  XNOR2_X1  g359(.A(KEYINPUT98), .B(KEYINPUT25), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n482), .A2(G103), .A3(G2104), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(G139), .B2(new_n477), .ZN(new_n788));
  AND2_X1   g363(.A1(new_n784), .A2(new_n788), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n779), .B1(new_n789), .B2(new_n721), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n790), .A2(G2072), .ZN(new_n791));
  NAND4_X1  g366(.A1(new_n762), .A2(new_n772), .A3(new_n778), .A4(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n715), .A2(G5), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G171), .B2(new_n715), .ZN(new_n794));
  AND2_X1   g369(.A1(new_n794), .A2(G1961), .ZN(new_n795));
  INV_X1    g370(.A(G34), .ZN(new_n796));
  AND2_X1   g371(.A1(new_n796), .A2(KEYINPUT24), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n796), .A2(KEYINPUT24), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n721), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(G160), .B2(new_n721), .ZN(new_n800));
  AND2_X1   g375(.A1(new_n800), .A2(G2084), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n795), .A2(new_n801), .ZN(new_n802));
  OAI221_X1 g377(.A(new_n802), .B1(new_n721), .B2(new_n649), .C1(G2084), .C2(new_n800), .ZN(new_n803));
  XOR2_X1   g378(.A(KEYINPUT31), .B(G11), .Z(new_n804));
  XOR2_X1   g379(.A(KEYINPUT104), .B(G28), .Z(new_n805));
  AOI21_X1  g380(.A(G29), .B1(new_n805), .B2(KEYINPUT30), .ZN(new_n806));
  INV_X1    g381(.A(KEYINPUT105), .ZN(new_n807));
  OR2_X1    g382(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n805), .A2(KEYINPUT30), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(new_n806), .B2(new_n807), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n804), .B1(new_n808), .B2(new_n810), .ZN(new_n811));
  OAI221_X1 g386(.A(new_n811), .B1(new_n794), .B2(G1961), .C1(G2072), .C2(new_n790), .ZN(new_n812));
  NOR4_X1   g387(.A1(new_n758), .A2(new_n792), .A3(new_n803), .A4(new_n812), .ZN(new_n813));
  NAND4_X1  g388(.A1(new_n726), .A2(new_n738), .A3(new_n757), .A4(new_n813), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n492), .A2(KEYINPUT91), .A3(G119), .ZN(new_n815));
  INV_X1    g390(.A(KEYINPUT91), .ZN(new_n816));
  INV_X1    g391(.A(G119), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n816), .B1(new_n491), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n815), .A2(new_n818), .ZN(new_n819));
  OAI21_X1  g394(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n820));
  INV_X1    g395(.A(G107), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n820), .B1(new_n821), .B2(G2105), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n822), .B1(new_n477), .B2(G131), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n819), .A2(new_n823), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT92), .ZN(new_n825));
  MUX2_X1   g400(.A(G25), .B(new_n825), .S(G29), .Z(new_n826));
  XNOR2_X1  g401(.A(KEYINPUT35), .B(G1991), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n827), .B(KEYINPUT93), .Z(new_n828));
  INV_X1    g403(.A(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n826), .B(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(KEYINPUT96), .A2(KEYINPUT36), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n715), .A2(G22), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n832), .B1(G166), .B2(new_n715), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT95), .ZN(new_n834));
  INV_X1    g409(.A(G1971), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n598), .A2(new_n597), .A3(G16), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n836), .B1(G6), .B2(G16), .ZN(new_n837));
  XNOR2_X1  g412(.A(KEYINPUT32), .B(G1981), .ZN(new_n838));
  INV_X1    g413(.A(new_n838), .ZN(new_n839));
  AOI22_X1  g414(.A1(new_n834), .A2(new_n835), .B1(new_n837), .B2(new_n839), .ZN(new_n840));
  AND2_X1   g415(.A1(new_n715), .A2(G23), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n841), .B1(G288), .B2(G16), .ZN(new_n842));
  XNOR2_X1  g417(.A(KEYINPUT33), .B(G1976), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n842), .B(new_n843), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n837), .A2(new_n839), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  OAI211_X1 g421(.A(new_n840), .B(new_n846), .C1(new_n835), .C2(new_n834), .ZN(new_n847));
  XNOR2_X1  g422(.A(KEYINPUT94), .B(KEYINPUT34), .ZN(new_n848));
  OR2_X1    g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n847), .A2(new_n848), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n715), .A2(G24), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n851), .B1(new_n604), .B2(new_n715), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(new_n704), .ZN(new_n853));
  AND3_X1   g428(.A1(new_n849), .A2(new_n850), .A3(new_n853), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n830), .A2(new_n831), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n830), .A2(new_n854), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n856), .A2(KEYINPUT96), .A3(KEYINPUT36), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n814), .B1(new_n855), .B2(new_n857), .ZN(G311));
  INV_X1    g433(.A(G311), .ZN(G150));
  NAND2_X1  g434(.A1(new_n624), .A2(G559), .ZN(new_n860));
  XOR2_X1   g435(.A(KEYINPUT106), .B(KEYINPUT38), .Z(new_n861));
  XNOR2_X1  g436(.A(new_n860), .B(new_n861), .ZN(new_n862));
  AOI22_X1  g437(.A1(new_n525), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n863), .A2(new_n517), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n864), .A2(KEYINPUT107), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n552), .A2(G93), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(G55), .ZN(new_n868));
  OAI22_X1  g443(.A1(new_n534), .A2(new_n868), .B1(new_n864), .B2(KEYINPUT107), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n870), .A2(new_n776), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n561), .B1(new_n867), .B2(new_n869), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n862), .B(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT39), .ZN(new_n876));
  AOI21_X1  g451(.A(G860), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n877), .B1(new_n876), .B2(new_n875), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n870), .A2(new_n562), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(KEYINPUT37), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n878), .A2(new_n880), .ZN(G145));
  OAI21_X1  g456(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n882));
  INV_X1    g457(.A(G118), .ZN(new_n883));
  AOI22_X1  g458(.A1(new_n882), .A2(KEYINPUT109), .B1(new_n883), .B2(G2105), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n884), .B1(KEYINPUT109), .B2(new_n882), .ZN(new_n885));
  INV_X1    g460(.A(G142), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n885), .B1(new_n745), .B2(new_n886), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n887), .B1(new_n492), .B2(G130), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n824), .A2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n888), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n819), .A2(new_n890), .A3(new_n823), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n892), .A2(new_n654), .ZN(new_n893));
  INV_X1    g468(.A(new_n654), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n889), .A2(new_n894), .A3(new_n891), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT108), .ZN(new_n897));
  AND2_X1   g472(.A1(new_n509), .A2(KEYINPUT72), .ZN(new_n898));
  OAI21_X1  g473(.A(KEYINPUT4), .B1(new_n509), .B2(KEYINPUT72), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n513), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n503), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n770), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n765), .A2(G164), .A3(new_n769), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(new_n752), .ZN(new_n906));
  AND2_X1   g481(.A1(new_n748), .A2(new_n751), .ZN(new_n907));
  OAI211_X1 g482(.A(new_n903), .B(new_n904), .C1(new_n907), .C2(new_n747), .ZN(new_n908));
  AOI211_X1 g483(.A(new_n897), .B(new_n789), .C1(new_n906), .C2(new_n908), .ZN(new_n909));
  OR2_X1    g484(.A1(new_n789), .A2(new_n897), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n789), .A2(new_n897), .ZN(new_n911));
  NAND4_X1  g486(.A1(new_n906), .A2(new_n910), .A3(new_n908), .A4(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n896), .B1(new_n909), .B2(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n906), .A2(new_n911), .A3(new_n908), .ZN(new_n915));
  INV_X1    g490(.A(new_n910), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND4_X1  g492(.A1(new_n917), .A2(new_n893), .A3(new_n895), .A4(new_n912), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n914), .A2(new_n918), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n649), .B(new_n479), .ZN(new_n920));
  XNOR2_X1  g495(.A(G162), .B(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n919), .A2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT110), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n919), .A2(KEYINPUT110), .A3(new_n922), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n914), .A2(new_n918), .A3(new_n921), .ZN(new_n928));
  INV_X1    g503(.A(G37), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(KEYINPUT40), .B1(new_n927), .B2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT40), .ZN(new_n933));
  AOI211_X1 g508(.A(new_n933), .B(new_n930), .C1(new_n925), .C2(new_n926), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n932), .A2(new_n934), .ZN(G395));
  XNOR2_X1  g510(.A(new_n639), .B(new_n873), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT111), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n937), .B1(new_n624), .B2(G299), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n637), .A2(KEYINPUT111), .A3(new_n576), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n624), .A2(G299), .ZN(new_n940));
  XOR2_X1   g515(.A(KEYINPUT112), .B(KEYINPUT41), .Z(new_n941));
  INV_X1    g516(.A(new_n941), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n938), .A2(new_n939), .A3(new_n940), .A4(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  AND2_X1   g519(.A1(new_n939), .A2(new_n940), .ZN(new_n945));
  AOI21_X1  g520(.A(KEYINPUT41), .B1(new_n945), .B2(new_n938), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n936), .B1(new_n944), .B2(new_n946), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n639), .B(new_n874), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n945), .A2(new_n938), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  XNOR2_X1  g525(.A(new_n604), .B(G305), .ZN(new_n951));
  XNOR2_X1  g526(.A(G166), .B(G288), .ZN(new_n952));
  XOR2_X1   g527(.A(new_n951), .B(new_n952), .Z(new_n953));
  XOR2_X1   g528(.A(new_n953), .B(KEYINPUT42), .Z(new_n954));
  AND3_X1   g529(.A1(new_n947), .A2(new_n950), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n954), .B1(new_n947), .B2(new_n950), .ZN(new_n956));
  OAI21_X1  g531(.A(G868), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n957), .B1(G868), .B2(new_n870), .ZN(G295));
  OAI21_X1  g533(.A(new_n957), .B1(G868), .B2(new_n870), .ZN(G331));
  INV_X1    g534(.A(new_n581), .ZN(new_n960));
  AOI21_X1  g535(.A(G286), .B1(new_n960), .B2(new_n579), .ZN(new_n961));
  NOR2_X1   g536(.A1(G171), .A2(G168), .ZN(new_n962));
  OAI211_X1 g537(.A(new_n872), .B(new_n871), .C1(new_n961), .C2(new_n962), .ZN(new_n963));
  OAI21_X1  g538(.A(G168), .B1(new_n580), .B2(new_n581), .ZN(new_n964));
  INV_X1    g539(.A(new_n962), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n873), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  AND2_X1   g541(.A1(new_n963), .A2(new_n966), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n967), .B1(new_n946), .B2(new_n944), .ZN(new_n968));
  INV_X1    g543(.A(new_n953), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n963), .A2(new_n966), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n949), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n968), .A2(new_n969), .A3(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT41), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n939), .A2(new_n940), .ZN(new_n974));
  AOI21_X1  g549(.A(KEYINPUT111), .B1(new_n637), .B2(new_n576), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n973), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n970), .B1(new_n976), .B2(new_n943), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n967), .B1(new_n938), .B2(new_n945), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n953), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n972), .A2(new_n979), .A3(new_n929), .ZN(new_n980));
  XOR2_X1   g555(.A(KEYINPUT113), .B(KEYINPUT43), .Z(new_n981));
  INV_X1    g556(.A(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT44), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n938), .A2(new_n939), .A3(new_n973), .A4(new_n940), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n967), .A2(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n941), .B1(new_n945), .B2(new_n938), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n971), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n988), .A2(new_n953), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n989), .A2(new_n972), .A3(new_n929), .A4(new_n981), .ZN(new_n990));
  AND3_X1   g565(.A1(new_n983), .A2(new_n984), .A3(new_n990), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n989), .A2(new_n972), .A3(new_n929), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(KEYINPUT43), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n972), .A2(new_n979), .A3(new_n929), .A4(new_n981), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n984), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n991), .A2(new_n995), .ZN(G397));
  INV_X1    g571(.A(KEYINPUT45), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n997), .B1(G164), .B2(G1384), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n472), .A2(new_n478), .A3(G40), .ZN(new_n999));
  OR2_X1    g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(G2067), .ZN(new_n1001));
  XNOR2_X1  g576(.A(new_n770), .B(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g577(.A(new_n1002), .B(KEYINPUT115), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n1000), .B1(new_n1003), .B2(new_n752), .ZN(new_n1004));
  INV_X1    g579(.A(G1996), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1000), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(new_n1005), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  AOI22_X1  g584(.A1(new_n1004), .A2(new_n1006), .B1(new_n752), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n604), .A2(new_n704), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1000), .A2(new_n1011), .ZN(new_n1012));
  XOR2_X1   g587(.A(new_n1012), .B(KEYINPUT127), .Z(new_n1013));
  XOR2_X1   g588(.A(KEYINPUT126), .B(KEYINPUT48), .Z(new_n1014));
  OR2_X1    g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  XNOR2_X1  g590(.A(new_n824), .B(new_n828), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(new_n1007), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1010), .A2(new_n1015), .A3(new_n1017), .A4(new_n1018), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1009), .A2(KEYINPUT46), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n1004), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT46), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1008), .A2(new_n1022), .ZN(new_n1023));
  XNOR2_X1  g598(.A(new_n1023), .B(KEYINPUT125), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT47), .ZN(new_n1025));
  AND3_X1   g600(.A1(new_n1021), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1025), .B1(new_n1021), .B2(new_n1024), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1019), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n825), .A2(new_n828), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1010), .A2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n765), .A2(new_n1001), .A3(new_n769), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1000), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1028), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(G8), .ZN(new_n1034));
  AOI21_X1  g609(.A(G1384), .B1(new_n900), .B2(new_n901), .ZN(new_n1035));
  INV_X1    g610(.A(new_n999), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1034), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(G1976), .ZN(new_n1038));
  INV_X1    g613(.A(G1981), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1039), .B1(new_n597), .B2(new_n598), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n597), .A2(new_n1039), .A3(new_n598), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1041), .A2(KEYINPUT49), .A3(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT49), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1042), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1044), .B1(new_n1045), .B2(new_n1040), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1043), .A2(new_n1046), .A3(new_n1037), .ZN(new_n1047));
  AND4_X1   g622(.A1(new_n1038), .A2(new_n1047), .A3(new_n585), .A4(new_n588), .ZN(new_n1048));
  XNOR2_X1  g623(.A(new_n1042), .B(KEYINPUT120), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1037), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1035), .A2(KEYINPUT45), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1051), .A2(new_n998), .A3(new_n1036), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(new_n835), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT50), .ZN(new_n1054));
  OAI21_X1  g629(.A(KEYINPUT116), .B1(new_n1035), .B2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n999), .B1(new_n1035), .B2(new_n1054), .ZN(new_n1056));
  INV_X1    g631(.A(G2090), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT116), .ZN(new_n1058));
  OAI211_X1 g633(.A(new_n1058), .B(KEYINPUT50), .C1(G164), .C2(G1384), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1055), .A2(new_n1056), .A3(new_n1057), .A4(new_n1059), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1034), .B1(new_n1053), .B2(new_n1060), .ZN(new_n1061));
  NOR2_X1   g636(.A1(G166), .A2(new_n1034), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT55), .ZN(new_n1063));
  XNOR2_X1  g638(.A(new_n1062), .B(new_n1063), .ZN(new_n1064));
  XNOR2_X1  g639(.A(new_n1064), .B(KEYINPUT117), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1061), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1067));
  INV_X1    g642(.A(G87), .ZN(new_n1068));
  OAI211_X1 g643(.A(new_n588), .B(G1976), .C1(new_n1068), .C2(new_n527), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT118), .ZN(new_n1070));
  XNOR2_X1  g645(.A(new_n1069), .B(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(KEYINPUT52), .B1(G288), .B2(new_n1038), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1067), .A2(new_n1071), .A3(G8), .A4(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT119), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1067), .A2(new_n1071), .A3(G8), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(KEYINPUT52), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1037), .A2(KEYINPUT119), .A3(new_n1071), .A4(new_n1072), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1075), .A2(new_n1077), .A3(new_n1078), .A4(new_n1047), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1050), .B1(new_n1066), .B2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT63), .ZN(new_n1081));
  OAI21_X1  g656(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1082));
  INV_X1    g657(.A(G1384), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n902), .A2(new_n1054), .A3(new_n1083), .ZN(new_n1084));
  AND3_X1   g659(.A1(new_n1082), .A2(new_n1084), .A3(new_n1036), .ZN(new_n1085));
  AOI22_X1  g660(.A1(new_n1085), .A2(new_n1057), .B1(new_n1052), .B2(new_n835), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1064), .B1(new_n1086), .B2(new_n1034), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1079), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1066), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT121), .ZN(new_n1090));
  INV_X1    g665(.A(G2084), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1055), .A2(new_n1056), .A3(new_n1091), .A4(new_n1059), .ZN(new_n1092));
  INV_X1    g667(.A(G1966), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1036), .B1(new_n1035), .B2(KEYINPUT45), .ZN(new_n1094));
  NOR3_X1   g669(.A1(G164), .A2(new_n997), .A3(G1384), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1093), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1092), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(G168), .A2(G8), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1090), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1100));
  AOI211_X1 g675(.A(KEYINPUT121), .B(new_n1098), .C1(new_n1092), .C2(new_n1096), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1081), .B1(new_n1089), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1053), .A2(new_n1060), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(G8), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1081), .B1(new_n1105), .B2(new_n1064), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1079), .B1(new_n1061), .B2(new_n1065), .ZN(new_n1107));
  OAI211_X1 g682(.A(new_n1106), .B(new_n1107), .C1(new_n1101), .C2(new_n1100), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1080), .B1(new_n1103), .B2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1092), .A2(new_n1096), .A3(G168), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(G8), .ZN(new_n1111));
  AOI21_X1  g686(.A(G168), .B1(new_n1092), .B2(new_n1096), .ZN(new_n1112));
  OAI21_X1  g687(.A(KEYINPUT51), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT51), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1110), .A2(new_n1114), .A3(G8), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(KEYINPUT62), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT62), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1113), .A2(new_n1118), .A3(new_n1115), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1055), .A2(new_n1056), .A3(new_n1059), .ZN(new_n1120));
  INV_X1    g695(.A(G1961), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1051), .A2(new_n998), .A3(new_n724), .A4(new_n1036), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT53), .ZN(new_n1123));
  AOI22_X1  g698(.A1(new_n1120), .A2(new_n1121), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1125), .A2(KEYINPUT53), .A3(new_n724), .ZN(new_n1126));
  AOI21_X1  g701(.A(G301), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1127));
  AND3_X1   g702(.A1(new_n1107), .A2(new_n1127), .A3(new_n1087), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1117), .A2(new_n1119), .A3(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1109), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT54), .ZN(new_n1131));
  XNOR2_X1  g706(.A(KEYINPUT123), .B(G2078), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1125), .A2(KEYINPUT53), .A3(new_n1132), .ZN(new_n1133));
  AND3_X1   g708(.A1(new_n1124), .A2(G301), .A3(new_n1133), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1131), .B1(new_n1134), .B2(new_n1127), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1124), .A2(new_n1126), .A3(G301), .ZN(new_n1136));
  AND2_X1   g711(.A1(new_n1124), .A2(new_n1133), .ZN(new_n1137));
  OAI211_X1 g712(.A(KEYINPUT54), .B(new_n1136), .C1(new_n1137), .C2(new_n554), .ZN(new_n1138));
  AND3_X1   g713(.A1(new_n1066), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1135), .A2(new_n1138), .A3(new_n1116), .A4(new_n1139), .ZN(new_n1140));
  OR2_X1    g715(.A1(new_n1140), .A2(KEYINPUT124), .ZN(new_n1141));
  XOR2_X1   g716(.A(KEYINPUT58), .B(G1341), .Z(new_n1142));
  NAND2_X1  g717(.A1(new_n1067), .A2(new_n1142), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1143), .B1(new_n1052), .B2(G1996), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1144), .A2(new_n776), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT59), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n1067), .A2(G2067), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1148), .B1(new_n1120), .B2(new_n734), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1149), .A2(KEYINPUT60), .A3(new_n637), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1144), .A2(KEYINPUT59), .A3(new_n776), .ZN(new_n1151));
  AND3_X1   g726(.A1(new_n1147), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT61), .ZN(new_n1153));
  XNOR2_X1  g728(.A(KEYINPUT56), .B(G2072), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1125), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1056), .A2(new_n1082), .ZN(new_n1156));
  INV_X1    g731(.A(G1956), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  XNOR2_X1  g733(.A(new_n576), .B(KEYINPUT57), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1155), .A2(new_n1158), .A3(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(new_n1160), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1159), .B1(new_n1155), .B2(new_n1158), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1153), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n637), .B1(new_n1149), .B2(KEYINPUT60), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1164), .B1(KEYINPUT60), .B2(new_n1149), .ZN(new_n1165));
  INV_X1    g740(.A(new_n1162), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1166), .A2(KEYINPUT61), .A3(new_n1160), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1152), .A2(new_n1163), .A3(new_n1165), .A4(new_n1167), .ZN(new_n1168));
  OAI21_X1  g743(.A(KEYINPUT122), .B1(new_n1149), .B2(new_n637), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1166), .A2(new_n1169), .ZN(new_n1170));
  NOR3_X1   g745(.A1(new_n1149), .A2(KEYINPUT122), .A3(new_n637), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1160), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  AOI22_X1  g747(.A1(new_n1140), .A2(KEYINPUT124), .B1(new_n1168), .B2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1130), .B1(new_n1141), .B2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1011), .A2(KEYINPUT114), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n604), .A2(new_n704), .ZN(new_n1176));
  XNOR2_X1  g751(.A(new_n1175), .B(new_n1176), .ZN(new_n1177));
  OAI211_X1 g752(.A(new_n1010), .B(new_n1017), .C1(new_n1000), .C2(new_n1177), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1033), .B1(new_n1174), .B2(new_n1178), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g754(.A1(new_n927), .A2(new_n931), .ZN(new_n1181));
  OAI21_X1  g755(.A(G319), .B1(new_n673), .B2(new_n674), .ZN(new_n1182));
  NOR2_X1   g756(.A1(new_n1182), .A2(G227), .ZN(new_n1183));
  AND3_X1   g757(.A1(new_n712), .A2(new_n713), .A3(new_n1183), .ZN(new_n1184));
  NAND2_X1  g758(.A1(new_n983), .A2(new_n990), .ZN(new_n1185));
  AND3_X1   g759(.A1(new_n1181), .A2(new_n1184), .A3(new_n1185), .ZN(G308));
  NAND3_X1  g760(.A1(new_n1181), .A2(new_n1184), .A3(new_n1185), .ZN(G225));
endmodule


