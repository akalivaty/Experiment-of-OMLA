//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 1 0 1 1 1 1 0 1 1 0 0 0 1 1 1 1 0 0 0 0 0 1 1 1 0 0 1 1 0 1 1 0 1 1 0 1 1 1 0 0 0 1 0 0 0 1 1 0 1 0 0 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:57 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n758, new_n759, new_n761, new_n762,
    new_n763, new_n765, new_n766, new_n768, new_n769, new_n770, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n795, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n976, new_n977, new_n978, new_n979, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057;
  XNOR2_X1  g000(.A(G104), .B(G107), .ZN(new_n187));
  INV_X1    g001(.A(G101), .ZN(new_n188));
  OAI21_X1  g002(.A(KEYINPUT76), .B1(new_n187), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G107), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G104), .ZN(new_n191));
  INV_X1    g005(.A(G104), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G107), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT76), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n194), .A2(new_n195), .A3(G101), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n189), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT1), .ZN(new_n198));
  INV_X1    g012(.A(G146), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n198), .B1(G143), .B2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G128), .ZN(new_n201));
  INV_X1    g015(.A(G143), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n202), .A2(G146), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n199), .A2(G143), .ZN(new_n204));
  OAI22_X1  g018(.A1(new_n200), .A2(new_n201), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n199), .A2(G143), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n202), .A2(G146), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n206), .A2(new_n207), .A3(new_n198), .A4(G128), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n205), .A2(new_n208), .ZN(new_n209));
  OAI21_X1  g023(.A(KEYINPUT3), .B1(new_n192), .B2(G107), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT3), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n211), .A2(new_n190), .A3(G104), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n210), .A2(new_n212), .A3(new_n188), .A4(new_n193), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n197), .A2(new_n209), .A3(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT77), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT10), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n197), .A2(new_n209), .A3(KEYINPUT77), .A4(new_n213), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n210), .A2(new_n212), .A3(new_n193), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G101), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n221), .A2(KEYINPUT4), .A3(new_n213), .ZN(new_n222));
  NOR2_X1   g036(.A1(KEYINPUT0), .A2(G128), .ZN(new_n223));
  XNOR2_X1  g037(.A(G143), .B(G146), .ZN(new_n224));
  NAND2_X1  g038(.A1(KEYINPUT0), .A2(G128), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n223), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n206), .A2(new_n207), .ZN(new_n227));
  INV_X1    g041(.A(new_n225), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n226), .A2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT4), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n220), .A2(new_n231), .A3(G101), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n222), .A2(new_n230), .A3(new_n232), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n197), .A2(new_n209), .A3(KEYINPUT10), .A4(new_n213), .ZN(new_n234));
  AND2_X1   g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  OR2_X1    g049(.A1(KEYINPUT65), .A2(G137), .ZN(new_n236));
  NAND2_X1  g050(.A1(KEYINPUT65), .A2(G137), .ZN(new_n237));
  AND2_X1   g051(.A1(KEYINPUT11), .A2(G134), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n236), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(G137), .ZN(new_n240));
  AOI21_X1  g054(.A(KEYINPUT11), .B1(new_n240), .B2(G134), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(G134), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G137), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n239), .A2(new_n242), .A3(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(G131), .ZN(new_n246));
  AOI21_X1  g060(.A(G131), .B1(new_n243), .B2(G137), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n239), .A2(new_n242), .A3(new_n247), .ZN(new_n248));
  AND3_X1   g062(.A1(new_n246), .A2(KEYINPUT78), .A3(new_n248), .ZN(new_n249));
  AOI21_X1  g063(.A(KEYINPUT78), .B1(new_n246), .B2(new_n248), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n219), .A2(new_n235), .A3(new_n251), .ZN(new_n252));
  NOR3_X1   g066(.A1(new_n187), .A2(KEYINPUT76), .A3(new_n188), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n195), .B1(new_n194), .B2(G101), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n213), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n255), .A2(new_n208), .A3(new_n205), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n216), .A2(new_n256), .A3(new_n218), .ZN(new_n257));
  AND2_X1   g071(.A1(KEYINPUT65), .A2(G137), .ZN(new_n258));
  NOR2_X1   g072(.A1(KEYINPUT65), .A2(G137), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n241), .B1(new_n260), .B2(new_n238), .ZN(new_n261));
  AOI22_X1  g075(.A1(G131), .A2(new_n245), .B1(new_n261), .B2(new_n247), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  AND3_X1   g077(.A1(new_n257), .A2(KEYINPUT12), .A3(new_n263), .ZN(new_n264));
  AOI21_X1  g078(.A(KEYINPUT12), .B1(new_n257), .B2(new_n263), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n252), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  XNOR2_X1  g080(.A(G110), .B(G140), .ZN(new_n267));
  INV_X1    g081(.A(G227), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n268), .A2(G953), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n267), .B(new_n269), .ZN(new_n270));
  AND3_X1   g084(.A1(new_n219), .A2(new_n235), .A3(new_n251), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n271), .A2(new_n270), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n219), .A2(new_n235), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(new_n263), .ZN(new_n274));
  AOI22_X1  g088(.A1(new_n266), .A2(new_n270), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  OAI21_X1  g089(.A(G469), .B1(new_n275), .B2(G902), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(KEYINPUT79), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT79), .ZN(new_n278));
  OAI211_X1 g092(.A(new_n278), .B(G469), .C1(new_n275), .C2(G902), .ZN(new_n279));
  INV_X1    g093(.A(G469), .ZN(new_n280));
  INV_X1    g094(.A(G902), .ZN(new_n281));
  INV_X1    g095(.A(new_n270), .ZN(new_n282));
  OAI211_X1 g096(.A(new_n252), .B(new_n282), .C1(new_n264), .C2(new_n265), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n282), .B1(new_n274), .B2(new_n252), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT80), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n283), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n262), .B1(new_n219), .B2(new_n235), .ZN(new_n287));
  OAI211_X1 g101(.A(new_n285), .B(new_n270), .C1(new_n271), .C2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  OAI211_X1 g103(.A(new_n280), .B(new_n281), .C1(new_n286), .C2(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n277), .A2(new_n279), .A3(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(G119), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(G116), .ZN(new_n293));
  INV_X1    g107(.A(G116), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(G119), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT66), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  XNOR2_X1  g112(.A(KEYINPUT2), .B(G113), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n293), .A2(new_n295), .A3(KEYINPUT66), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n298), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT67), .ZN(new_n302));
  NOR3_X1   g116(.A1(new_n296), .A2(new_n299), .A3(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(G113), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(KEYINPUT2), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT2), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(G113), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  XNOR2_X1  g122(.A(G116), .B(G119), .ZN(new_n309));
  AOI21_X1  g123(.A(KEYINPUT67), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n301), .B1(new_n303), .B2(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n311), .A2(new_n222), .A3(new_n232), .ZN(new_n312));
  AND3_X1   g126(.A1(new_n293), .A2(new_n295), .A3(KEYINPUT66), .ZN(new_n313));
  AOI21_X1  g127(.A(KEYINPUT66), .B1(new_n293), .B2(new_n295), .ZN(new_n314));
  OAI21_X1  g128(.A(KEYINPUT5), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT81), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n316), .B1(new_n293), .B2(KEYINPUT5), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT5), .ZN(new_n318));
  NAND4_X1  g132(.A1(new_n318), .A2(new_n292), .A3(KEYINPUT81), .A4(G116), .ZN(new_n319));
  AND3_X1   g133(.A1(new_n317), .A2(G113), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n315), .A2(new_n320), .ZN(new_n321));
  AND3_X1   g135(.A1(new_n210), .A2(new_n212), .A3(new_n193), .ZN(new_n322));
  AOI22_X1  g136(.A1(new_n189), .A2(new_n196), .B1(new_n322), .B2(new_n188), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n302), .B1(new_n296), .B2(new_n299), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n308), .A2(new_n309), .A3(KEYINPUT67), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n321), .A2(new_n323), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n312), .A2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT82), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT6), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n312), .A2(new_n327), .A3(KEYINPUT82), .ZN(new_n332));
  XNOR2_X1  g146(.A(G110), .B(G122), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  NAND4_X1  g148(.A1(new_n330), .A2(new_n331), .A3(new_n332), .A4(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(G125), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n336), .B1(new_n226), .B2(new_n229), .ZN(new_n337));
  AOI21_X1  g151(.A(G125), .B1(new_n205), .B2(new_n208), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(G953), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(G224), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  XNOR2_X1  g156(.A(new_n339), .B(new_n342), .ZN(new_n343));
  AND3_X1   g157(.A1(new_n312), .A2(KEYINPUT82), .A3(new_n327), .ZN(new_n344));
  AOI21_X1  g158(.A(KEYINPUT82), .B1(new_n312), .B2(new_n327), .ZN(new_n345));
  NOR3_X1   g159(.A1(new_n344), .A2(new_n345), .A3(new_n333), .ZN(new_n346));
  OAI21_X1  g160(.A(KEYINPUT6), .B1(new_n328), .B2(new_n334), .ZN(new_n347));
  OAI211_X1 g161(.A(new_n335), .B(new_n343), .C1(new_n346), .C2(new_n347), .ZN(new_n348));
  AND3_X1   g162(.A1(new_n312), .A2(new_n327), .A3(new_n333), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n321), .A2(new_n255), .A3(new_n326), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n317), .A2(G113), .A3(new_n319), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n296), .A2(new_n318), .ZN(new_n352));
  OAI22_X1  g166(.A1(new_n303), .A2(new_n310), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(new_n323), .ZN(new_n354));
  XNOR2_X1  g168(.A(new_n333), .B(KEYINPUT8), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n350), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n209), .A2(new_n336), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT7), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n342), .A2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(new_n223), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n360), .B1(new_n227), .B2(new_n228), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n224), .A2(new_n225), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  OAI211_X1 g177(.A(new_n357), .B(new_n359), .C1(new_n336), .C2(new_n363), .ZN(new_n364));
  OAI22_X1  g178(.A1(new_n337), .A2(new_n338), .B1(new_n358), .B2(new_n342), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n356), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n349), .B1(new_n367), .B2(KEYINPUT83), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT83), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n356), .A2(new_n366), .A3(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(G902), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  OAI21_X1  g185(.A(G210), .B1(G237), .B2(G902), .ZN(new_n372));
  AND3_X1   g186(.A1(new_n348), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  XOR2_X1   g187(.A(new_n372), .B(KEYINPUT84), .Z(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n375), .B1(new_n348), .B2(new_n371), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n373), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(G221), .ZN(new_n378));
  XNOR2_X1  g192(.A(KEYINPUT9), .B(G234), .ZN(new_n379));
  XNOR2_X1  g193(.A(new_n379), .B(KEYINPUT75), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n378), .B1(new_n380), .B2(new_n281), .ZN(new_n381));
  OAI21_X1  g195(.A(G214), .B1(G237), .B2(G902), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  NOR3_X1   g197(.A1(new_n377), .A2(new_n381), .A3(new_n383), .ZN(new_n384));
  AND2_X1   g198(.A1(new_n291), .A2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(G475), .ZN(new_n386));
  INV_X1    g200(.A(G140), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(G125), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n336), .A2(G140), .ZN(new_n389));
  AND2_X1   g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  XNOR2_X1  g204(.A(new_n390), .B(new_n199), .ZN(new_n391));
  INV_X1    g205(.A(G237), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n392), .A2(new_n340), .A3(G214), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(new_n202), .ZN(new_n394));
  NOR2_X1   g208(.A1(G237), .A2(G953), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n395), .A2(G143), .A3(G214), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n397), .A2(KEYINPUT18), .A3(G131), .ZN(new_n398));
  NAND2_X1  g212(.A1(KEYINPUT18), .A2(G131), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n394), .A2(new_n396), .A3(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n391), .A2(new_n398), .A3(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT87), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT17), .ZN(new_n403));
  AND3_X1   g217(.A1(new_n395), .A2(G143), .A3(G214), .ZN(new_n404));
  AOI21_X1  g218(.A(G143), .B1(new_n395), .B2(G214), .ZN(new_n405));
  OAI21_X1  g219(.A(G131), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(KEYINPUT85), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT85), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n397), .A2(new_n408), .A3(G131), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n403), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n388), .A2(new_n389), .A3(KEYINPUT16), .ZN(new_n411));
  OR3_X1    g225(.A1(new_n336), .A2(KEYINPUT16), .A3(G140), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(new_n199), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n411), .A2(new_n412), .A3(G146), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n402), .B1(new_n410), .B2(new_n416), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n408), .B1(new_n397), .B2(G131), .ZN(new_n418));
  INV_X1    g232(.A(G131), .ZN(new_n419));
  AOI211_X1 g233(.A(KEYINPUT85), .B(new_n419), .C1(new_n394), .C2(new_n396), .ZN(new_n420));
  OAI21_X1  g234(.A(KEYINPUT17), .B1(new_n418), .B2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n416), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n421), .A2(KEYINPUT87), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n417), .A2(new_n423), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n418), .A2(new_n420), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT88), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n394), .A2(new_n419), .A3(new_n396), .ZN(new_n427));
  NAND4_X1  g241(.A1(new_n425), .A2(new_n426), .A3(new_n403), .A4(new_n427), .ZN(new_n428));
  NAND4_X1  g242(.A1(new_n407), .A2(new_n409), .A3(new_n403), .A4(new_n427), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(KEYINPUT88), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n401), .B1(new_n424), .B2(new_n431), .ZN(new_n432));
  XNOR2_X1  g246(.A(G113), .B(G122), .ZN(new_n433));
  XNOR2_X1  g247(.A(new_n433), .B(new_n192), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n432), .A2(new_n435), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n434), .B(new_n401), .C1(new_n424), .C2(new_n431), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n386), .B1(new_n438), .B2(new_n281), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT20), .ZN(new_n441));
  AND3_X1   g255(.A1(new_n407), .A2(new_n409), .A3(new_n427), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT73), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n415), .A2(new_n443), .ZN(new_n444));
  NAND4_X1  g258(.A1(new_n411), .A2(new_n412), .A3(KEYINPUT73), .A4(G146), .ZN(new_n445));
  AND3_X1   g259(.A1(new_n388), .A2(new_n389), .A3(KEYINPUT19), .ZN(new_n446));
  AOI21_X1  g260(.A(KEYINPUT19), .B1(new_n388), .B2(new_n389), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  OAI211_X1 g262(.A(new_n444), .B(new_n445), .C1(G146), .C2(new_n448), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n401), .B1(new_n442), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(KEYINPUT86), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT86), .ZN(new_n452));
  OAI211_X1 g266(.A(new_n452), .B(new_n401), .C1(new_n442), .C2(new_n449), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n451), .A2(new_n435), .A3(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT89), .ZN(new_n455));
  AND3_X1   g269(.A1(new_n437), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n455), .B1(new_n437), .B2(new_n454), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NOR2_X1   g272(.A1(G475), .A2(G902), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n441), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n437), .A2(new_n454), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n461), .A2(new_n441), .A3(new_n459), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n440), .B1(new_n460), .B2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(G952), .ZN(new_n465));
  AOI211_X1 g279(.A(G953), .B(new_n465), .C1(G234), .C2(G237), .ZN(new_n466));
  AOI211_X1 g280(.A(new_n281), .B(new_n340), .C1(G234), .C2(G237), .ZN(new_n467));
  XNOR2_X1  g281(.A(KEYINPUT21), .B(G898), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n466), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT90), .ZN(new_n470));
  INV_X1    g284(.A(G122), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(G116), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n294), .A2(G122), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n472), .A2(new_n473), .A3(new_n190), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n190), .B1(new_n472), .B2(new_n473), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n470), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n202), .A2(G128), .ZN(new_n478));
  OAI21_X1  g292(.A(G134), .B1(new_n478), .B2(KEYINPUT13), .ZN(new_n479));
  XNOR2_X1  g293(.A(G128), .B(G143), .ZN(new_n480));
  OR2_X1    g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n294), .A2(G122), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n471), .A2(G116), .ZN(new_n483));
  OAI21_X1  g297(.A(G107), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n484), .A2(KEYINPUT90), .A3(new_n474), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n479), .A2(new_n480), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n477), .A2(new_n481), .A3(new_n485), .A4(new_n486), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n472), .B1(new_n473), .B2(KEYINPUT14), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT14), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n483), .A2(new_n489), .ZN(new_n490));
  OAI21_X1  g304(.A(G107), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n480), .A2(G134), .ZN(new_n492));
  OR2_X1    g306(.A1(new_n480), .A2(G134), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n491), .A2(new_n474), .A3(new_n492), .A4(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n487), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n380), .A2(G217), .A3(new_n340), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n496), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n498), .A2(new_n487), .A3(new_n494), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n497), .A2(KEYINPUT91), .A3(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT91), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n498), .A2(new_n487), .A3(new_n501), .A4(new_n494), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n500), .A2(new_n281), .A3(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(G478), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n504), .A2(KEYINPUT15), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(new_n505), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n500), .A2(new_n281), .A3(new_n502), .A4(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  NOR3_X1   g323(.A1(new_n464), .A2(new_n469), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n292), .A2(G128), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n201), .A2(KEYINPUT23), .A3(G119), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n292), .A2(G128), .ZN(new_n513));
  OAI211_X1 g327(.A(new_n511), .B(new_n512), .C1(new_n513), .C2(KEYINPUT23), .ZN(new_n514));
  XOR2_X1   g328(.A(KEYINPUT24), .B(G110), .Z(new_n515));
  XNOR2_X1  g329(.A(G119), .B(G128), .ZN(new_n516));
  AOI22_X1  g330(.A1(new_n514), .A2(G110), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n416), .A2(new_n517), .ZN(new_n518));
  XNOR2_X1  g332(.A(KEYINPUT72), .B(G110), .ZN(new_n519));
  OAI22_X1  g333(.A1(new_n514), .A2(new_n519), .B1(new_n515), .B2(new_n516), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n390), .A2(new_n199), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n444), .A2(new_n520), .A3(new_n445), .A4(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n518), .A2(new_n522), .ZN(new_n523));
  XNOR2_X1  g337(.A(KEYINPUT22), .B(G137), .ZN(new_n524));
  AND3_X1   g338(.A1(new_n340), .A2(G221), .A3(G234), .ZN(new_n525));
  XOR2_X1   g339(.A(new_n524), .B(new_n525), .Z(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n523), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n518), .A2(new_n522), .A3(new_n526), .ZN(new_n529));
  AND2_X1   g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  AOI21_X1  g344(.A(KEYINPUT25), .B1(new_n530), .B2(new_n281), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n530), .A2(KEYINPUT25), .A3(new_n281), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n532), .A2(KEYINPUT74), .A3(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(G217), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n535), .B1(G234), .B2(new_n281), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT74), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n537), .B1(new_n531), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n536), .A2(G902), .ZN(new_n540));
  AOI22_X1  g354(.A1(new_n534), .A2(new_n539), .B1(new_n530), .B2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(G472), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n395), .A2(G210), .ZN(new_n544));
  XNOR2_X1  g358(.A(new_n544), .B(KEYINPUT27), .ZN(new_n545));
  XNOR2_X1  g359(.A(KEYINPUT26), .B(G101), .ZN(new_n546));
  XNOR2_X1  g360(.A(new_n545), .B(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT28), .ZN(new_n549));
  AOI22_X1  g363(.A1(new_n246), .A2(new_n248), .B1(new_n229), .B2(new_n226), .ZN(new_n550));
  AOI21_X1  g364(.A(G134), .B1(new_n236), .B2(new_n237), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n240), .A2(G134), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  OAI21_X1  g367(.A(G131), .B1(new_n551), .B2(new_n553), .ZN(new_n554));
  AND3_X1   g368(.A1(new_n209), .A2(new_n248), .A3(new_n554), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n311), .B1(new_n550), .B2(new_n555), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n313), .A2(new_n314), .ZN(new_n557));
  AOI22_X1  g371(.A1(new_n557), .A2(new_n299), .B1(new_n324), .B2(new_n325), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n209), .A2(new_n248), .A3(new_n554), .ZN(new_n559));
  OAI211_X1 g373(.A(new_n558), .B(new_n559), .C1(new_n262), .C2(new_n363), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n549), .B1(new_n556), .B2(new_n560), .ZN(new_n561));
  AND2_X1   g375(.A1(new_n560), .A2(new_n549), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n548), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n560), .A2(new_n547), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n419), .B1(new_n261), .B2(new_n244), .ZN(new_n565));
  INV_X1    g379(.A(new_n248), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n230), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT68), .ZN(new_n568));
  NAND4_X1  g382(.A1(new_n567), .A2(new_n568), .A3(KEYINPUT30), .A4(new_n559), .ZN(new_n569));
  INV_X1    g383(.A(new_n208), .ZN(new_n570));
  OAI21_X1  g384(.A(KEYINPUT1), .B1(new_n202), .B2(G146), .ZN(new_n571));
  AOI22_X1  g385(.A1(new_n571), .A2(G128), .B1(new_n206), .B2(new_n207), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n248), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n243), .B1(new_n258), .B2(new_n259), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n419), .B1(new_n574), .B2(new_n552), .ZN(new_n575));
  OAI21_X1  g389(.A(KEYINPUT30), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(KEYINPUT68), .B1(new_n576), .B2(new_n550), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n569), .A2(new_n577), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n559), .B1(new_n262), .B2(new_n363), .ZN(new_n579));
  XNOR2_X1  g393(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n558), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n564), .B1(new_n578), .B2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT31), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n563), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  AOI211_X1 g398(.A(KEYINPUT31), .B(new_n564), .C1(new_n578), .C2(new_n581), .ZN(new_n585));
  OAI211_X1 g399(.A(new_n543), .B(new_n281), .C1(new_n584), .C2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT32), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NOR3_X1   g402(.A1(new_n587), .A2(G472), .A3(G902), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n589), .B1(new_n584), .B2(new_n585), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT71), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  OAI211_X1 g406(.A(KEYINPUT71), .B(new_n589), .C1(new_n584), .C2(new_n585), .ZN(new_n593));
  AND3_X1   g407(.A1(new_n588), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT29), .ZN(new_n595));
  INV_X1    g409(.A(new_n560), .ZN(new_n596));
  AOI211_X1 g410(.A(new_n596), .B(new_n547), .C1(new_n578), .C2(new_n581), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n558), .B1(new_n567), .B2(new_n559), .ZN(new_n598));
  OAI21_X1  g412(.A(KEYINPUT28), .B1(new_n596), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n560), .A2(new_n549), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n548), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  OAI211_X1 g415(.A(KEYINPUT69), .B(new_n595), .C1(new_n597), .C2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT70), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n547), .A2(KEYINPUT29), .ZN(new_n604));
  NOR3_X1   g418(.A1(new_n561), .A2(new_n562), .A3(new_n604), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n603), .B1(new_n605), .B2(G902), .ZN(new_n606));
  INV_X1    g420(.A(new_n604), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n599), .A2(new_n600), .A3(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n608), .A2(KEYINPUT70), .A3(new_n281), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n602), .A2(new_n606), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n578), .A2(new_n581), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n611), .A2(new_n560), .A3(new_n548), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n547), .B1(new_n561), .B2(new_n562), .ZN(new_n613));
  AOI21_X1  g427(.A(KEYINPUT29), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n614), .A2(KEYINPUT69), .ZN(new_n615));
  OAI21_X1  g429(.A(G472), .B1(new_n610), .B2(new_n615), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n542), .B1(new_n594), .B2(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n385), .A2(new_n510), .A3(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(G101), .ZN(G3));
  OAI21_X1  g433(.A(new_n270), .B1(new_n271), .B2(new_n287), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n257), .A2(new_n263), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT12), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n257), .A2(KEYINPUT12), .A3(new_n263), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  AOI22_X1  g439(.A1(KEYINPUT80), .A2(new_n620), .B1(new_n272), .B2(new_n625), .ZN(new_n626));
  AOI21_X1  g440(.A(G902), .B1(new_n626), .B2(new_n288), .ZN(new_n627));
  AOI22_X1  g441(.A1(new_n280), .A2(new_n627), .B1(new_n276), .B2(KEYINPUT79), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n381), .B1(new_n628), .B2(new_n279), .ZN(new_n629));
  INV_X1    g443(.A(new_n564), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n611), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(KEYINPUT31), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n582), .A2(new_n583), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n632), .A2(new_n633), .A3(new_n563), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(new_n281), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(G472), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(new_n586), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n637), .A2(new_n542), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n629), .A2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n469), .ZN(new_n640));
  XOR2_X1   g454(.A(KEYINPUT92), .B(KEYINPUT33), .Z(new_n641));
  NAND3_X1  g455(.A1(new_n500), .A2(new_n502), .A3(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT93), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(new_n644));
  AND2_X1   g458(.A1(new_n499), .A2(KEYINPUT33), .ZN(new_n645));
  AND3_X1   g459(.A1(new_n495), .A2(KEYINPUT94), .A3(new_n496), .ZN(new_n646));
  AOI21_X1  g460(.A(KEYINPUT94), .B1(new_n495), .B2(new_n496), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n645), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(KEYINPUT95), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT95), .ZN(new_n650));
  OAI211_X1 g464(.A(new_n645), .B(new_n650), .C1(new_n647), .C2(new_n646), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n504), .A2(G902), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n644), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n503), .A2(new_n504), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(KEYINPUT96), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n372), .B1(new_n348), .B2(new_n371), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n348), .A2(new_n371), .A3(new_n372), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n383), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n464), .A2(new_n640), .A3(new_n657), .A4(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n639), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(KEYINPUT34), .B(G104), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G6));
  XNOR2_X1  g479(.A(new_n469), .B(KEYINPUT97), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n661), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n461), .A2(KEYINPUT89), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n437), .A2(new_n454), .A3(new_n455), .ZN(new_n669));
  AND4_X1   g483(.A1(new_n441), .A2(new_n668), .A3(new_n459), .A4(new_n669), .ZN(new_n670));
  OAI211_X1 g484(.A(new_n440), .B(new_n509), .C1(new_n460), .C2(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n667), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n672), .A2(new_n629), .A3(new_n638), .ZN(new_n673));
  XOR2_X1   g487(.A(KEYINPUT35), .B(G107), .Z(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(G9));
  NAND2_X1  g489(.A1(new_n534), .A2(new_n539), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n527), .A2(KEYINPUT36), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n523), .B(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(new_n540), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n680), .A2(new_n636), .A3(new_n586), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n385), .A2(new_n510), .A3(new_n682), .ZN(new_n683));
  XOR2_X1   g497(.A(KEYINPUT37), .B(G110), .Z(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(G12));
  INV_X1    g499(.A(new_n680), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n686), .B1(new_n594), .B2(new_n616), .ZN(new_n687));
  XOR2_X1   g501(.A(new_n466), .B(KEYINPUT98), .Z(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(G900), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n689), .B1(new_n690), .B2(new_n467), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n671), .A2(new_n691), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n687), .A2(new_n692), .A3(new_n629), .A4(new_n661), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G128), .ZN(G30));
  XOR2_X1   g508(.A(new_n691), .B(KEYINPUT39), .Z(new_n695));
  NAND2_X1  g509(.A1(new_n629), .A2(new_n695), .ZN(new_n696));
  XOR2_X1   g510(.A(new_n696), .B(KEYINPUT40), .Z(new_n697));
  NAND3_X1  g511(.A1(new_n588), .A2(new_n592), .A3(new_n593), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT101), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n547), .B1(new_n556), .B2(new_n560), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(KEYINPUT100), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n701), .A2(G472), .A3(new_n631), .ZN(new_n702));
  NAND2_X1  g516(.A1(G472), .A2(G902), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n699), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  AND3_X1   g518(.A1(new_n702), .A2(new_n699), .A3(new_n703), .ZN(new_n705));
  NOR3_X1   g519(.A1(new_n698), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  XOR2_X1   g521(.A(KEYINPUT99), .B(KEYINPUT38), .Z(new_n708));
  XNOR2_X1  g522(.A(new_n377), .B(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n668), .A2(new_n459), .A3(new_n669), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n463), .B1(new_n711), .B2(KEYINPUT20), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n712), .A2(new_n439), .ZN(new_n713));
  INV_X1    g527(.A(new_n509), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n715), .A2(new_n382), .A3(new_n686), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n710), .B1(KEYINPUT102), .B2(new_n716), .ZN(new_n717));
  OAI211_X1 g531(.A(new_n697), .B(new_n717), .C1(KEYINPUT102), .C2(new_n716), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G143), .ZN(G45));
  INV_X1    g533(.A(new_n691), .ZN(new_n720));
  OAI211_X1 g534(.A(new_n657), .B(new_n720), .C1(new_n712), .C2(new_n439), .ZN(new_n721));
  INV_X1    g535(.A(new_n721), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n687), .A2(new_n629), .A3(new_n722), .A4(new_n661), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT103), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT69), .ZN(new_n726));
  AOI211_X1 g540(.A(new_n726), .B(KEYINPUT29), .C1(new_n612), .C2(new_n613), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n606), .A2(new_n609), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(new_n615), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n543), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n680), .B1(new_n731), .B2(new_n698), .ZN(new_n732));
  INV_X1    g546(.A(new_n381), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n291), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n735), .A2(KEYINPUT103), .A3(new_n661), .A4(new_n722), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n725), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G146), .ZN(G48));
  AOI21_X1  g552(.A(KEYINPUT71), .B1(new_n634), .B2(new_n589), .ZN(new_n739));
  INV_X1    g553(.A(new_n593), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n741), .A2(new_n616), .A3(new_n588), .ZN(new_n742));
  INV_X1    g556(.A(new_n290), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n620), .A2(KEYINPUT80), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n744), .A2(new_n288), .A3(new_n283), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n280), .B1(new_n745), .B2(new_n281), .ZN(new_n746));
  NOR3_X1   g560(.A1(new_n743), .A2(new_n746), .A3(new_n381), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n742), .A2(new_n541), .A3(new_n747), .ZN(new_n748));
  OAI21_X1  g562(.A(KEYINPUT104), .B1(new_n748), .B2(new_n662), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n661), .A2(new_n640), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n657), .B1(new_n712), .B2(new_n439), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT104), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n752), .A2(new_n617), .A3(new_n753), .A4(new_n747), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n749), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(KEYINPUT41), .B(G113), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n755), .B(new_n756), .ZN(G15));
  NAND3_X1  g571(.A1(new_n672), .A2(new_n617), .A3(new_n747), .ZN(new_n758));
  XNOR2_X1  g572(.A(KEYINPUT105), .B(G116), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n758), .B(new_n759), .ZN(G18));
  OAI21_X1  g574(.A(new_n382), .B1(new_n373), .B2(new_n658), .ZN(new_n761));
  NOR4_X1   g575(.A1(new_n761), .A2(new_n743), .A3(new_n746), .A4(new_n381), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n510), .A2(new_n687), .A3(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G119), .ZN(G21));
  AND4_X1   g578(.A1(new_n586), .A2(new_n636), .A3(new_n541), .A4(new_n666), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n762), .A2(new_n715), .A3(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G122), .ZN(G24));
  NOR2_X1   g581(.A1(new_n721), .A2(new_n681), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(new_n762), .ZN(new_n769));
  XNOR2_X1  g583(.A(KEYINPUT106), .B(G125), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n769), .B(new_n770), .ZN(G27));
  AOI21_X1  g585(.A(KEYINPUT108), .B1(new_n377), .B2(new_n382), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n348), .A2(new_n371), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(new_n374), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n774), .A2(KEYINPUT108), .A3(new_n382), .A4(new_n660), .ZN(new_n775));
  INV_X1    g589(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n772), .A2(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT107), .ZN(new_n778));
  AND3_X1   g592(.A1(new_n290), .A2(new_n276), .A3(new_n778), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n778), .B1(new_n290), .B2(new_n276), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n777), .A2(new_n781), .A3(new_n733), .ZN(new_n782));
  AOI22_X1  g596(.A1(new_n586), .A2(new_n587), .B1(new_n634), .B2(new_n589), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n542), .B1(new_n616), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n722), .A2(new_n784), .ZN(new_n785));
  OAI21_X1  g599(.A(KEYINPUT42), .B1(new_n782), .B2(new_n785), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n721), .A2(KEYINPUT42), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n774), .A2(new_n382), .A3(new_n660), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT108), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  AND3_X1   g604(.A1(new_n790), .A2(new_n733), .A3(new_n775), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n787), .A2(new_n791), .A3(new_n617), .A4(new_n781), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n786), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(new_n419), .ZN(G33));
  NAND4_X1  g608(.A1(new_n617), .A2(new_n791), .A3(new_n692), .A4(new_n781), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(G134), .ZN(G36));
  NAND2_X1  g610(.A1(new_n713), .A2(new_n657), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(KEYINPUT43), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT43), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n713), .A2(new_n799), .A3(new_n657), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n801), .A2(new_n637), .A3(new_n680), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT44), .ZN(new_n803));
  OR2_X1    g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n802), .A2(new_n803), .ZN(new_n805));
  NAND2_X1  g619(.A1(G469), .A2(G902), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n275), .A2(KEYINPUT45), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  OAI21_X1  g622(.A(G469), .B1(new_n275), .B2(KEYINPUT45), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n806), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT46), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n743), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n812), .B1(new_n811), .B2(new_n810), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n813), .A2(new_n733), .ZN(new_n814));
  INV_X1    g628(.A(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(new_n695), .ZN(new_n816));
  INV_X1    g630(.A(new_n816), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n804), .A2(new_n777), .A3(new_n805), .A4(new_n817), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(G137), .ZN(G39));
  NAND2_X1  g633(.A1(new_n815), .A2(KEYINPUT47), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT47), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n814), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(new_n777), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n824), .A2(new_n742), .A3(new_n541), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n823), .A2(new_n722), .A3(new_n825), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n826), .B(G140), .ZN(G42));
  INV_X1    g641(.A(KEYINPUT54), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n713), .A2(new_n714), .A3(new_n761), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT111), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n733), .B1(new_n691), .B2(new_n830), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n831), .B1(new_n830), .B2(new_n691), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n676), .A2(new_n679), .A3(new_n832), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n705), .A2(new_n704), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n833), .B1(new_n594), .B2(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n829), .A2(new_n835), .A3(new_n781), .ZN(new_n836));
  AND3_X1   g650(.A1(new_n693), .A2(new_n836), .A3(new_n769), .ZN(new_n837));
  AND3_X1   g651(.A1(new_n737), .A2(new_n837), .A3(KEYINPUT52), .ZN(new_n838));
  AOI21_X1  g652(.A(KEYINPUT52), .B1(new_n737), .B2(new_n837), .ZN(new_n839));
  OAI21_X1  g653(.A(KEYINPUT53), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n506), .A2(KEYINPUT110), .A3(new_n508), .ZN(new_n841));
  AOI21_X1  g655(.A(KEYINPUT110), .B1(new_n506), .B2(new_n508), .ZN(new_n842));
  OR2_X1    g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n751), .B1(new_n464), .B2(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n385), .A2(new_n844), .A3(new_n765), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n845), .A2(new_n618), .A3(new_n683), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n440), .B1(new_n460), .B2(new_n670), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n720), .B1(new_n841), .B2(new_n842), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n687), .A2(new_n629), .A3(new_n777), .A4(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n768), .A2(new_n791), .A3(new_n781), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n795), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n793), .A2(new_n846), .A3(new_n852), .ZN(new_n853));
  AND3_X1   g667(.A1(new_n758), .A2(new_n763), .A3(new_n766), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n853), .A2(new_n755), .A3(new_n854), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n840), .A2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n737), .A2(new_n837), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT52), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n737), .A2(new_n837), .A3(KEYINPUT52), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n749), .A2(new_n754), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT109), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n758), .A2(new_n763), .A3(new_n766), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  AOI21_X1  g680(.A(KEYINPUT109), .B1(new_n854), .B2(new_n755), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n862), .A2(new_n868), .A3(new_n853), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT53), .ZN(new_n870));
  AOI21_X1  g684(.A(KEYINPUT113), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n838), .A2(new_n839), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n864), .B1(new_n863), .B2(new_n865), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n854), .A2(KEYINPUT109), .A3(new_n755), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n853), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  OAI211_X1 g689(.A(KEYINPUT113), .B(new_n870), .C1(new_n872), .C2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(new_n876), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n828), .B(new_n857), .C1(new_n871), .C2(new_n877), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n870), .B1(new_n872), .B2(new_n875), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n862), .A2(new_n868), .A3(KEYINPUT53), .A4(new_n853), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  AOI21_X1  g695(.A(KEYINPUT112), .B1(new_n881), .B2(KEYINPUT54), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT112), .ZN(new_n883));
  AOI211_X1 g697(.A(new_n883), .B(new_n828), .C1(new_n879), .C2(new_n880), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n878), .B1(new_n882), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(KEYINPUT114), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT114), .ZN(new_n887));
  OAI211_X1 g701(.A(new_n878), .B(new_n887), .C1(new_n882), .C2(new_n884), .ZN(new_n888));
  INV_X1    g702(.A(new_n747), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n824), .A2(new_n889), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n890), .A2(new_n541), .A3(new_n466), .A4(new_n706), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n891), .A2(new_n464), .A3(new_n657), .ZN(new_n892));
  INV_X1    g706(.A(new_n890), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n801), .A2(KEYINPUT115), .A3(new_n689), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n798), .A2(new_n689), .A3(new_n800), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT115), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n893), .B1(new_n894), .B2(new_n897), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n892), .B1(new_n898), .B2(new_n682), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n894), .A2(new_n897), .ZN(new_n900));
  AND2_X1   g714(.A1(new_n900), .A2(new_n638), .ZN(new_n901));
  NOR3_X1   g715(.A1(new_n889), .A2(new_n709), .A3(new_n382), .ZN(new_n902));
  AND3_X1   g716(.A1(new_n901), .A2(KEYINPUT50), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g717(.A(KEYINPUT50), .B1(new_n901), .B2(new_n902), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n899), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT51), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n900), .A2(new_n638), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n907), .A2(new_n824), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n743), .A2(new_n746), .ZN(new_n909));
  INV_X1    g723(.A(new_n909), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n910), .A2(new_n733), .ZN(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n820), .A2(new_n822), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n906), .B1(new_n908), .B2(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(KEYINPUT117), .B1(new_n905), .B2(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(new_n904), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n901), .A2(KEYINPUT50), .A3(new_n902), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT117), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n919), .A2(new_n914), .A3(new_n920), .A4(new_n899), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n916), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n898), .A2(new_n784), .ZN(new_n923));
  XOR2_X1   g737(.A(KEYINPUT119), .B(KEYINPUT48), .Z(new_n924));
  XNOR2_X1  g738(.A(new_n923), .B(new_n924), .ZN(new_n925));
  AND3_X1   g739(.A1(new_n900), .A2(new_n638), .A3(new_n762), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT118), .ZN(new_n927));
  OAI211_X1 g741(.A(G952), .B(new_n340), .C1(new_n891), .C2(new_n751), .ZN(new_n928));
  OR3_X1    g742(.A1(new_n926), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n927), .B1(new_n926), .B2(new_n928), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n925), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT116), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n823), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n933), .A2(new_n912), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n823), .A2(new_n932), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n908), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  OAI211_X1 g750(.A(new_n936), .B(new_n899), .C1(new_n904), .C2(new_n903), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n931), .B1(new_n937), .B2(new_n906), .ZN(new_n938));
  AND2_X1   g752(.A1(new_n922), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n886), .A2(new_n888), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n465), .A2(new_n340), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NOR3_X1   g756(.A1(new_n707), .A2(new_n542), .A3(new_n797), .ZN(new_n943));
  OR2_X1    g757(.A1(new_n910), .A2(KEYINPUT49), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n910), .A2(KEYINPUT49), .ZN(new_n945));
  NOR3_X1   g759(.A1(new_n709), .A2(new_n381), .A3(new_n383), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n943), .A2(new_n944), .A3(new_n945), .A4(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n942), .A2(new_n947), .ZN(G75));
  OAI21_X1  g762(.A(new_n335), .B1(new_n346), .B2(new_n347), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n949), .B(new_n343), .ZN(new_n950));
  XOR2_X1   g764(.A(KEYINPUT120), .B(KEYINPUT55), .Z(new_n951));
  XNOR2_X1  g765(.A(new_n950), .B(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT113), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n879), .A2(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n856), .B1(new_n954), .B2(new_n876), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n955), .A2(new_n281), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n956), .A2(G210), .ZN(new_n957));
  INV_X1    g771(.A(KEYINPUT56), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n952), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n340), .A2(G952), .ZN(new_n960));
  INV_X1    g774(.A(new_n960), .ZN(new_n961));
  NOR3_X1   g775(.A1(new_n955), .A2(new_n281), .A3(new_n375), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n952), .A2(new_n958), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n961), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n959), .A2(new_n964), .ZN(G51));
  NOR2_X1   g779(.A1(new_n808), .A2(new_n809), .ZN(new_n966));
  AND3_X1   g780(.A1(new_n956), .A2(KEYINPUT121), .A3(new_n966), .ZN(new_n967));
  AOI21_X1  g781(.A(KEYINPUT121), .B1(new_n956), .B2(new_n966), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n806), .B(KEYINPUT57), .Z(new_n970));
  INV_X1    g784(.A(new_n878), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n955), .A2(new_n828), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n970), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n973), .A2(new_n745), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n960), .B1(new_n969), .B2(new_n974), .ZN(G54));
  NAND2_X1  g789(.A1(KEYINPUT58), .A2(G475), .ZN(new_n976));
  INV_X1    g790(.A(new_n976), .ZN(new_n977));
  AND3_X1   g791(.A1(new_n956), .A2(new_n458), .A3(new_n977), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n458), .B1(new_n956), .B2(new_n977), .ZN(new_n979));
  NOR3_X1   g793(.A1(new_n978), .A2(new_n979), .A3(new_n960), .ZN(G60));
  AND2_X1   g794(.A1(new_n644), .A2(new_n652), .ZN(new_n981));
  NAND2_X1  g795(.A1(G478), .A2(G902), .ZN(new_n982));
  XOR2_X1   g796(.A(new_n982), .B(KEYINPUT59), .Z(new_n983));
  INV_X1    g797(.A(new_n983), .ZN(new_n984));
  OAI211_X1 g798(.A(new_n981), .B(new_n984), .C1(new_n971), .C2(new_n972), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n985), .A2(new_n961), .ZN(new_n986));
  INV_X1    g800(.A(new_n888), .ZN(new_n987));
  AND3_X1   g801(.A1(new_n853), .A2(new_n873), .A3(new_n874), .ZN(new_n988));
  AOI21_X1  g802(.A(KEYINPUT53), .B1(new_n988), .B2(new_n862), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n840), .A2(new_n875), .ZN(new_n990));
  OAI21_X1  g804(.A(KEYINPUT54), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n991), .A2(new_n883), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n881), .A2(KEYINPUT112), .A3(KEYINPUT54), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n887), .B1(new_n994), .B2(new_n878), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n984), .B1(new_n987), .B2(new_n995), .ZN(new_n996));
  INV_X1    g810(.A(new_n981), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n986), .B1(new_n996), .B2(new_n997), .ZN(G63));
  OAI21_X1  g812(.A(new_n857), .B1(new_n871), .B2(new_n877), .ZN(new_n999));
  NAND2_X1  g813(.A1(G217), .A2(G902), .ZN(new_n1000));
  XNOR2_X1  g814(.A(new_n1000), .B(KEYINPUT122), .ZN(new_n1001));
  XNOR2_X1  g815(.A(new_n1001), .B(KEYINPUT60), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n999), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g817(.A(new_n530), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n960), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n999), .A2(new_n678), .A3(new_n1002), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g821(.A(KEYINPUT61), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g823(.A1(new_n1005), .A2(KEYINPUT61), .A3(new_n1006), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1009), .A2(new_n1010), .ZN(G66));
  OR3_X1    g825(.A1(new_n866), .A2(new_n867), .A3(new_n846), .ZN(new_n1012));
  OR2_X1    g826(.A1(new_n1012), .A2(G953), .ZN(new_n1013));
  INV_X1    g827(.A(new_n468), .ZN(new_n1014));
  NAND3_X1  g828(.A1(new_n1014), .A2(G224), .A3(G953), .ZN(new_n1015));
  NAND3_X1  g829(.A1(new_n1013), .A2(KEYINPUT123), .A3(new_n1015), .ZN(new_n1016));
  INV_X1    g830(.A(new_n1016), .ZN(new_n1017));
  AOI21_X1  g831(.A(KEYINPUT123), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1018));
  OAI21_X1  g832(.A(KEYINPUT124), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g833(.A(new_n1018), .ZN(new_n1020));
  INV_X1    g834(.A(KEYINPUT124), .ZN(new_n1021));
  NAND3_X1  g835(.A1(new_n1020), .A2(new_n1021), .A3(new_n1016), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1019), .A2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g837(.A(new_n949), .B1(G898), .B2(new_n340), .ZN(new_n1024));
  XNOR2_X1  g838(.A(new_n1023), .B(new_n1024), .ZN(G69));
  NAND2_X1  g839(.A1(new_n579), .A2(new_n580), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n578), .A2(new_n1026), .ZN(new_n1027));
  XNOR2_X1  g841(.A(new_n1027), .B(new_n448), .ZN(new_n1028));
  INV_X1    g842(.A(new_n696), .ZN(new_n1029));
  NAND4_X1  g843(.A1(new_n1029), .A2(new_n617), .A3(new_n777), .A4(new_n844), .ZN(new_n1030));
  NAND3_X1  g844(.A1(new_n818), .A2(new_n826), .A3(new_n1030), .ZN(new_n1031));
  AND3_X1   g845(.A1(new_n737), .A2(new_n693), .A3(new_n769), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n718), .A2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g847(.A(new_n1031), .B1(KEYINPUT62), .B2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g848(.A(new_n1034), .B1(KEYINPUT62), .B2(new_n1033), .ZN(new_n1035));
  AOI21_X1  g849(.A(new_n1028), .B1(new_n1035), .B2(new_n340), .ZN(new_n1036));
  INV_X1    g850(.A(new_n795), .ZN(new_n1037));
  AND2_X1   g851(.A1(new_n829), .A2(new_n784), .ZN(new_n1038));
  AOI211_X1 g852(.A(new_n793), .B(new_n1037), .C1(new_n817), .C2(new_n1038), .ZN(new_n1039));
  NAND4_X1  g853(.A1(new_n1039), .A2(new_n818), .A3(new_n826), .A4(new_n1032), .ZN(new_n1040));
  NOR2_X1   g854(.A1(new_n1040), .A2(G953), .ZN(new_n1041));
  OAI21_X1  g855(.A(new_n1028), .B1(new_n690), .B2(new_n340), .ZN(new_n1042));
  OAI21_X1  g856(.A(KEYINPUT125), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NOR2_X1   g857(.A1(new_n1036), .A2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g858(.A(G953), .B1(new_n268), .B2(new_n690), .ZN(new_n1045));
  XNOR2_X1  g859(.A(new_n1044), .B(new_n1045), .ZN(G72));
  XNOR2_X1  g860(.A(new_n703), .B(KEYINPUT63), .ZN(new_n1047));
  INV_X1    g861(.A(new_n1047), .ZN(new_n1048));
  OAI21_X1  g862(.A(new_n1048), .B1(new_n1035), .B2(new_n1012), .ZN(new_n1049));
  AOI21_X1  g863(.A(new_n548), .B1(new_n611), .B2(new_n560), .ZN(new_n1050));
  NAND2_X1  g864(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g865(.A(new_n1048), .B1(new_n1040), .B2(new_n1012), .ZN(new_n1052));
  INV_X1    g866(.A(KEYINPUT126), .ZN(new_n1053));
  AOI21_X1  g867(.A(new_n612), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g868(.A(new_n1054), .B1(new_n1053), .B2(new_n1052), .ZN(new_n1055));
  NOR3_X1   g869(.A1(new_n1050), .A2(new_n597), .A3(new_n1047), .ZN(new_n1056));
  AOI21_X1  g870(.A(new_n960), .B1(new_n881), .B2(new_n1056), .ZN(new_n1057));
  AND3_X1   g871(.A1(new_n1051), .A2(new_n1055), .A3(new_n1057), .ZN(G57));
endmodule


