//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 1 1 0 0 0 0 1 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 1 0 0 0 1 0 1 1 0 0 0 1 1 1 0 0 1 0 1 1 1 1 1 1 1 1 0 1 0 0 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:27 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n685, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n710, new_n711, new_n712, new_n713, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n743, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n765, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n883, new_n884,
    new_n885, new_n886, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  XNOR2_X1  g002(.A(KEYINPUT86), .B(G469), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G134), .ZN(new_n191));
  OAI21_X1  g005(.A(KEYINPUT66), .B1(new_n191), .B2(G137), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(KEYINPUT11), .ZN(new_n193));
  INV_X1    g007(.A(G137), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G134), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT11), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n195), .A2(KEYINPUT66), .A3(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n191), .A2(G137), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n193), .A2(new_n197), .A3(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G131), .ZN(new_n200));
  INV_X1    g014(.A(G131), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n193), .A2(new_n197), .A3(new_n201), .A4(new_n198), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n200), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g017(.A1(KEYINPUT85), .A2(KEYINPUT12), .ZN(new_n204));
  INV_X1    g018(.A(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G104), .ZN(new_n206));
  OAI21_X1  g020(.A(KEYINPUT3), .B1(new_n206), .B2(G107), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT3), .ZN(new_n208));
  INV_X1    g022(.A(G107), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n208), .A2(new_n209), .A3(G104), .ZN(new_n210));
  INV_X1    g024(.A(G101), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n206), .A2(G107), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n207), .A2(new_n210), .A3(new_n211), .A4(new_n212), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n206), .A2(G107), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n209), .A2(G104), .ZN(new_n215));
  OAI21_X1  g029(.A(G101), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n213), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT65), .ZN(new_n218));
  INV_X1    g032(.A(G146), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(KEYINPUT65), .A2(G146), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n220), .A2(G143), .A3(new_n221), .ZN(new_n222));
  AND2_X1   g036(.A1(KEYINPUT69), .A2(KEYINPUT1), .ZN(new_n223));
  NOR2_X1   g037(.A1(KEYINPUT69), .A2(KEYINPUT1), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(G143), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G146), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n222), .A2(new_n225), .A3(G128), .A4(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n217), .A2(new_n228), .ZN(new_n229));
  AND2_X1   g043(.A1(KEYINPUT65), .A2(G146), .ZN(new_n230));
  NOR2_X1   g044(.A1(KEYINPUT65), .A2(G146), .ZN(new_n231));
  NOR3_X1   g045(.A1(new_n230), .A2(new_n231), .A3(new_n226), .ZN(new_n232));
  OAI21_X1  g046(.A(G128), .B1(new_n232), .B2(new_n225), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n226), .A2(G146), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n230), .A2(new_n231), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n235), .B1(new_n236), .B2(G143), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT70), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n233), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(G128), .ZN(new_n240));
  XNOR2_X1  g054(.A(KEYINPUT69), .B(KEYINPUT1), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n240), .B1(new_n222), .B2(new_n241), .ZN(new_n242));
  XNOR2_X1  g056(.A(KEYINPUT65), .B(G146), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n234), .B1(new_n243), .B2(new_n226), .ZN(new_n244));
  OAI21_X1  g058(.A(KEYINPUT70), .B1(new_n242), .B2(new_n244), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n229), .B1(new_n239), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n222), .A2(new_n227), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT1), .ZN(new_n248));
  OAI21_X1  g062(.A(G128), .B1(new_n234), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  AND2_X1   g064(.A1(new_n250), .A2(new_n228), .ZN(new_n251));
  OAI22_X1  g065(.A1(new_n246), .A2(KEYINPUT84), .B1(new_n217), .B2(new_n251), .ZN(new_n252));
  AND2_X1   g066(.A1(new_n246), .A2(KEYINPUT84), .ZN(new_n253));
  OAI211_X1 g067(.A(new_n203), .B(new_n205), .C1(new_n252), .C2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(new_n203), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n217), .B1(new_n250), .B2(new_n228), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n239), .A2(new_n245), .ZN(new_n257));
  INV_X1    g071(.A(new_n229), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT84), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n256), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n246), .A2(KEYINPUT84), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n255), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  AND2_X1   g077(.A1(KEYINPUT85), .A2(KEYINPUT12), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n264), .A2(new_n204), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n254), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(KEYINPUT87), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT87), .ZN(new_n268));
  OAI211_X1 g082(.A(new_n254), .B(new_n268), .C1(new_n263), .C2(new_n265), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n256), .A2(KEYINPUT10), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT83), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n207), .A2(new_n210), .A3(new_n212), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(G101), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n273), .A2(KEYINPUT4), .A3(new_n213), .ZN(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  XOR2_X1   g089(.A(KEYINPUT0), .B(G128), .Z(new_n276));
  AOI21_X1  g090(.A(G143), .B1(new_n220), .B2(new_n221), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n276), .B1(new_n277), .B2(new_n234), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT4), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n272), .A2(new_n279), .A3(G101), .ZN(new_n280));
  NAND4_X1  g094(.A1(new_n222), .A2(KEYINPUT0), .A3(G128), .A4(new_n227), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n278), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n271), .B1(new_n275), .B2(new_n282), .ZN(new_n283));
  AND2_X1   g097(.A1(new_n278), .A2(new_n281), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n284), .A2(new_n274), .A3(KEYINPUT83), .A4(new_n280), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n270), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n238), .B1(new_n233), .B2(new_n237), .ZN(new_n287));
  NOR3_X1   g101(.A1(new_n242), .A2(new_n244), .A3(KEYINPUT70), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n228), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(new_n217), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n289), .A2(KEYINPUT10), .A3(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n286), .A2(new_n255), .A3(new_n291), .ZN(new_n292));
  XNOR2_X1  g106(.A(G110), .B(G140), .ZN(new_n293));
  INV_X1    g107(.A(G953), .ZN(new_n294));
  AND2_X1   g108(.A1(new_n294), .A2(G227), .ZN(new_n295));
  XNOR2_X1  g109(.A(new_n293), .B(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n292), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n267), .A2(new_n269), .A3(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n255), .B1(new_n286), .B2(new_n291), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(new_n292), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(new_n296), .ZN(new_n304));
  AOI211_X1 g118(.A(G902), .B(new_n190), .C1(new_n300), .C2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(G469), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n302), .A2(new_n292), .A3(new_n297), .ZN(new_n307));
  INV_X1    g121(.A(new_n292), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n203), .B1(new_n252), .B2(new_n253), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n309), .B1(new_n264), .B2(new_n204), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n308), .B1(new_n310), .B2(new_n254), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n307), .B1(new_n311), .B2(new_n297), .ZN(new_n312));
  INV_X1    g126(.A(G902), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n306), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n188), .B1(new_n305), .B2(new_n314), .ZN(new_n315));
  XNOR2_X1  g129(.A(G116), .B(G119), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  XNOR2_X1  g131(.A(KEYINPUT2), .B(G113), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(new_n318), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(new_n316), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n274), .A2(new_n322), .A3(new_n280), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n316), .A2(KEYINPUT5), .ZN(new_n324));
  INV_X1    g138(.A(G116), .ZN(new_n325));
  OR3_X1    g139(.A1(new_n325), .A2(KEYINPUT5), .A3(G119), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n324), .A2(G113), .A3(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n290), .A2(new_n321), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n323), .A2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT6), .ZN(new_n330));
  XNOR2_X1  g144(.A(G110), .B(G122), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n329), .A2(new_n330), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n329), .A2(new_n332), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n323), .A2(new_n331), .A3(new_n328), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n334), .A2(KEYINPUT6), .A3(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(new_n228), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n337), .B1(new_n239), .B2(new_n245), .ZN(new_n338));
  INV_X1    g152(.A(G125), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n278), .A2(new_n281), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(G125), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(G224), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n344), .A2(G953), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(new_n345), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n347), .B1(new_n340), .B2(new_n342), .ZN(new_n348));
  OAI211_X1 g162(.A(new_n333), .B(new_n336), .C1(new_n346), .C2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n348), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT7), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n343), .A2(new_n351), .ZN(new_n352));
  XNOR2_X1  g166(.A(new_n331), .B(KEYINPUT8), .ZN(new_n353));
  INV_X1    g167(.A(new_n328), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n290), .B1(new_n321), .B2(new_n327), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n353), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  AND2_X1   g170(.A1(new_n356), .A2(new_n335), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n340), .A2(KEYINPUT7), .A3(new_n347), .A4(new_n342), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n350), .A2(new_n352), .A3(new_n357), .A4(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n349), .A2(new_n313), .A3(new_n359), .ZN(new_n360));
  OAI21_X1  g174(.A(G210), .B1(G237), .B2(G902), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  NAND4_X1  g177(.A1(new_n349), .A2(new_n359), .A3(new_n313), .A4(new_n361), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  OAI21_X1  g179(.A(G214), .B1(G237), .B2(G902), .ZN(new_n366));
  NAND2_X1  g180(.A1(G234), .A2(G237), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n367), .A2(G952), .A3(new_n294), .ZN(new_n368));
  XOR2_X1   g182(.A(KEYINPUT21), .B(G898), .Z(new_n369));
  NAND3_X1  g183(.A1(new_n367), .A2(G902), .A3(G953), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n368), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n365), .A2(new_n366), .A3(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(G237), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n373), .A2(new_n294), .A3(G214), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT88), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n374), .A2(new_n375), .A3(new_n226), .ZN(new_n376));
  NOR2_X1   g190(.A1(G237), .A2(G953), .ZN(new_n377));
  OAI211_X1 g191(.A(new_n377), .B(G214), .C1(KEYINPUT88), .C2(G143), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(G131), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT17), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n376), .A2(new_n201), .A3(new_n378), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n380), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(KEYINPUT89), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT16), .ZN(new_n385));
  INV_X1    g199(.A(G140), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n385), .A2(new_n386), .A3(G125), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(G125), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n339), .A2(G140), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n387), .B1(new_n390), .B2(new_n385), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(new_n219), .ZN(new_n392));
  OAI211_X1 g206(.A(G146), .B(new_n387), .C1(new_n390), .C2(new_n385), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT89), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n380), .A2(new_n396), .A3(new_n381), .A4(new_n382), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n379), .A2(KEYINPUT17), .A3(G131), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n384), .A2(new_n395), .A3(new_n397), .A4(new_n398), .ZN(new_n399));
  XNOR2_X1  g213(.A(G113), .B(G122), .ZN(new_n400));
  XNOR2_X1  g214(.A(new_n400), .B(new_n206), .ZN(new_n401));
  AND2_X1   g215(.A1(KEYINPUT18), .A2(G131), .ZN(new_n402));
  OR2_X1    g216(.A1(new_n379), .A2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n390), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(new_n236), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n405), .B1(new_n219), .B2(new_n404), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n379), .A2(new_n402), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n403), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  AND3_X1   g222(.A1(new_n399), .A2(new_n401), .A3(new_n408), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n401), .B1(new_n399), .B2(new_n408), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n313), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(KEYINPUT90), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT90), .ZN(new_n413));
  OAI211_X1 g227(.A(new_n413), .B(new_n313), .C1(new_n409), .C2(new_n410), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n412), .A2(G475), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n380), .A2(new_n382), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n390), .B(KEYINPUT19), .ZN(new_n417));
  OAI211_X1 g231(.A(new_n416), .B(new_n393), .C1(new_n243), .C2(new_n417), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n401), .B1(new_n418), .B2(new_n408), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n409), .A2(new_n419), .ZN(new_n420));
  NOR2_X1   g234(.A1(G475), .A2(G902), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  OAI21_X1  g236(.A(KEYINPUT20), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT20), .ZN(new_n424));
  OAI211_X1 g238(.A(new_n424), .B(new_n421), .C1(new_n409), .C2(new_n419), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n415), .A2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(KEYINPUT13), .B1(new_n240), .B2(G143), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n429), .A2(new_n191), .ZN(new_n430));
  XNOR2_X1  g244(.A(G128), .B(G143), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n430), .B(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(G122), .ZN(new_n433));
  AND2_X1   g247(.A1(new_n433), .A2(KEYINPUT91), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n433), .A2(KEYINPUT91), .ZN(new_n435));
  OAI21_X1  g249(.A(G116), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n325), .A2(G122), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n436), .A2(new_n209), .A3(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n209), .B1(new_n436), .B2(new_n437), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n432), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(new_n436), .ZN(new_n442));
  XNOR2_X1  g256(.A(new_n437), .B(KEYINPUT14), .ZN(new_n443));
  OAI21_X1  g257(.A(G107), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  XNOR2_X1  g258(.A(new_n431), .B(new_n191), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n444), .A2(new_n438), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n441), .A2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(G217), .ZN(new_n448));
  NOR3_X1   g262(.A1(new_n187), .A2(new_n448), .A3(G953), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n441), .A2(new_n446), .A3(new_n449), .ZN(new_n452));
  AOI21_X1  g266(.A(G902), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(G478), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n454), .A2(KEYINPUT15), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n453), .B(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n428), .A2(new_n456), .ZN(new_n457));
  NOR3_X1   g271(.A1(new_n315), .A2(new_n372), .A3(new_n457), .ZN(new_n458));
  NOR2_X1   g272(.A1(G472), .A2(G902), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT67), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n195), .A2(new_n198), .A3(new_n460), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n191), .A2(KEYINPUT67), .A3(G137), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n461), .A2(G131), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(KEYINPUT68), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT68), .ZN(new_n465));
  NAND4_X1  g279(.A1(new_n461), .A2(new_n465), .A3(G131), .A4(new_n462), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n464), .A2(new_n202), .A3(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n289), .A2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT28), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n203), .A2(new_n284), .ZN(new_n471));
  AND3_X1   g285(.A1(new_n319), .A2(new_n321), .A3(KEYINPUT71), .ZN(new_n472));
  AOI21_X1  g286(.A(KEYINPUT71), .B1(new_n319), .B2(new_n321), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND4_X1  g288(.A1(new_n469), .A2(new_n470), .A3(new_n471), .A4(new_n474), .ZN(new_n475));
  OAI211_X1 g289(.A(new_n471), .B(new_n474), .C1(new_n338), .C2(new_n467), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(KEYINPUT28), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n341), .B1(new_n202), .B2(new_n200), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n478), .B1(new_n289), .B2(new_n468), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  AOI22_X1  g294(.A1(new_n475), .A2(new_n477), .B1(new_n480), .B2(new_n322), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n377), .A2(G210), .ZN(new_n482));
  XNOR2_X1  g296(.A(new_n482), .B(KEYINPUT27), .ZN(new_n483));
  XNOR2_X1  g297(.A(KEYINPUT26), .B(G101), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n483), .B(new_n484), .ZN(new_n485));
  OAI21_X1  g299(.A(KEYINPUT73), .B1(new_n481), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n476), .A2(new_n485), .ZN(new_n487));
  XNOR2_X1  g301(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n467), .B1(new_n257), .B2(new_n228), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n489), .B1(new_n490), .B2(new_n478), .ZN(new_n491));
  INV_X1    g305(.A(new_n322), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT30), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n478), .A2(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n492), .B1(new_n469), .B2(new_n494), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n487), .B1(new_n491), .B2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT31), .ZN(new_n497));
  AOI21_X1  g311(.A(KEYINPUT72), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  OAI211_X1 g312(.A(KEYINPUT30), .B(new_n471), .C1(new_n338), .C2(new_n467), .ZN(new_n499));
  OAI211_X1 g313(.A(new_n322), .B(new_n499), .C1(new_n479), .C2(new_n488), .ZN(new_n500));
  INV_X1    g314(.A(new_n485), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n501), .B1(new_n479), .B2(new_n474), .ZN(new_n502));
  AND4_X1   g316(.A1(KEYINPUT72), .A2(new_n500), .A3(new_n497), .A4(new_n502), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n486), .B1(new_n498), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n475), .A2(new_n477), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n480), .A2(new_n322), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT73), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n507), .A2(new_n508), .A3(new_n501), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n497), .B1(new_n500), .B2(new_n502), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n459), .B1(new_n504), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(KEYINPUT74), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT72), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n500), .A2(new_n502), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n515), .B1(new_n516), .B2(KEYINPUT31), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n496), .A2(KEYINPUT72), .A3(new_n497), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n519), .A2(new_n511), .A3(new_n509), .A4(new_n486), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT74), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n520), .A2(new_n521), .A3(new_n459), .ZN(new_n522));
  XOR2_X1   g336(.A(KEYINPUT75), .B(KEYINPUT32), .Z(new_n523));
  NAND3_X1  g337(.A1(new_n514), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT77), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n479), .A2(new_n474), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n505), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n485), .A2(KEYINPUT29), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n313), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n476), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n531), .B1(new_n495), .B2(new_n491), .ZN(new_n532));
  NOR3_X1   g346(.A1(new_n532), .A2(KEYINPUT76), .A3(new_n485), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT76), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n488), .B1(new_n469), .B2(new_n471), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n471), .A2(KEYINPUT30), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n322), .B1(new_n490), .B2(new_n536), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n476), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n534), .B1(new_n538), .B2(new_n501), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n533), .A2(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(KEYINPUT29), .B1(new_n481), .B2(new_n485), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n530), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(G472), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n525), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n538), .A2(new_n534), .A3(new_n501), .ZN(new_n545));
  OAI21_X1  g359(.A(KEYINPUT76), .B1(new_n532), .B2(new_n485), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n541), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n530), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n549), .A2(KEYINPUT77), .A3(G472), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n544), .A2(new_n550), .ZN(new_n551));
  OAI211_X1 g365(.A(KEYINPUT32), .B(new_n459), .C1(new_n504), .C2(new_n512), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n524), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(G234), .ZN(new_n554));
  OAI21_X1  g368(.A(G217), .B1(new_n554), .B2(G902), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n555), .B(KEYINPUT78), .ZN(new_n556));
  OAI21_X1  g370(.A(KEYINPUT23), .B1(new_n240), .B2(G119), .ZN(new_n557));
  AOI21_X1  g371(.A(KEYINPUT79), .B1(new_n240), .B2(G119), .ZN(new_n558));
  XNOR2_X1  g372(.A(new_n557), .B(new_n558), .ZN(new_n559));
  XNOR2_X1  g373(.A(G119), .B(G128), .ZN(new_n560));
  XOR2_X1   g374(.A(KEYINPUT24), .B(G110), .Z(new_n561));
  AOI22_X1  g375(.A1(new_n559), .A2(G110), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  OAI22_X1  g376(.A1(new_n559), .A2(G110), .B1(new_n560), .B2(new_n561), .ZN(new_n563));
  AND2_X1   g377(.A1(new_n405), .A2(new_n393), .ZN(new_n564));
  AOI22_X1  g378(.A1(new_n394), .A2(new_n562), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  XNOR2_X1  g379(.A(KEYINPUT22), .B(G137), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n294), .A2(G221), .A3(G234), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n566), .B(new_n567), .ZN(new_n568));
  XOR2_X1   g382(.A(new_n568), .B(KEYINPUT80), .Z(new_n569));
  OR2_X1    g383(.A1(new_n565), .A2(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(KEYINPUT81), .B1(new_n565), .B2(new_n568), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n565), .A2(KEYINPUT81), .A3(new_n568), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT82), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT25), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  AND3_X1   g391(.A1(new_n574), .A2(new_n313), .A3(new_n577), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n577), .B1(new_n574), .B2(new_n313), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n556), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n556), .A2(G902), .ZN(new_n581));
  AND2_X1   g395(.A1(new_n574), .A2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n458), .A2(new_n553), .A3(new_n585), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n586), .B(G101), .ZN(G3));
  INV_X1    g401(.A(KEYINPUT92), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n520), .A2(new_n313), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n588), .B1(new_n590), .B2(new_n543), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n589), .A2(KEYINPUT92), .A3(G472), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AND2_X1   g407(.A1(new_n514), .A2(new_n522), .ZN(new_n594));
  AND2_X1   g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n315), .A2(new_n584), .ZN(new_n596));
  AND2_X1   g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT93), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n364), .A2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n366), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n363), .A2(new_n598), .A3(new_n364), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n601), .A2(new_n602), .A3(new_n371), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n451), .A2(new_n452), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(KEYINPUT33), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT33), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n451), .A2(new_n606), .A3(new_n452), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n605), .A2(G478), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n453), .A2(new_n454), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n454), .A2(new_n313), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n608), .A2(new_n609), .A3(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n427), .A2(new_n613), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n603), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n597), .A2(new_n615), .ZN(new_n616));
  XOR2_X1   g430(.A(KEYINPUT34), .B(G104), .Z(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(G6));
  NAND2_X1  g432(.A1(new_n601), .A2(new_n602), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n427), .A2(new_n456), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n371), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(KEYINPUT94), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT94), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n620), .A2(new_n623), .A3(new_n371), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n619), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n597), .A2(new_n625), .ZN(new_n626));
  XOR2_X1   g440(.A(KEYINPUT35), .B(G107), .Z(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(G9));
  INV_X1    g442(.A(KEYINPUT36), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n569), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(new_n565), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(new_n581), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n580), .A2(new_n632), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n593), .A2(new_n458), .A3(new_n594), .A4(new_n633), .ZN(new_n634));
  XOR2_X1   g448(.A(KEYINPUT37), .B(G110), .Z(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G12));
  OR2_X1    g450(.A1(new_n370), .A2(G900), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(new_n368), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  NOR3_X1   g453(.A1(new_n427), .A2(new_n456), .A3(new_n639), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n640), .A2(new_n602), .A3(new_n601), .A4(new_n633), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n641), .A2(new_n315), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n553), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(G128), .ZN(G30));
  INV_X1    g458(.A(new_n524), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n501), .B1(new_n526), .B2(new_n531), .ZN(new_n646));
  AOI21_X1  g460(.A(G902), .B1(new_n516), .B2(new_n646), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n552), .B1(new_n543), .B2(new_n647), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(KEYINPUT96), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n638), .B(KEYINPUT39), .ZN(new_n651));
  OAI211_X1 g465(.A(new_n188), .B(new_n651), .C1(new_n305), .C2(new_n314), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(KEYINPUT40), .ZN(new_n653));
  OR2_X1    g467(.A1(new_n653), .A2(KEYINPUT97), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n653), .A2(KEYINPUT97), .ZN(new_n655));
  XNOR2_X1  g469(.A(KEYINPUT95), .B(KEYINPUT38), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n365), .B(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n456), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n427), .A2(new_n659), .ZN(new_n660));
  NOR4_X1   g474(.A1(new_n658), .A2(new_n600), .A3(new_n633), .A4(new_n660), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n650), .A2(new_n654), .A3(new_n655), .A4(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(KEYINPUT98), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G143), .ZN(G45));
  AOI211_X1 g478(.A(new_n612), .B(new_n639), .C1(new_n415), .C2(new_n426), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n665), .A2(new_n602), .A3(new_n601), .A4(new_n633), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n315), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n553), .A2(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT99), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n553), .A2(new_n667), .A3(KEYINPUT99), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G146), .ZN(G48));
  AOI21_X1  g487(.A(new_n298), .B1(new_n266), .B2(KEYINPUT87), .ZN(new_n674));
  AOI22_X1  g488(.A1(new_n674), .A2(new_n269), .B1(new_n296), .B2(new_n303), .ZN(new_n675));
  OAI21_X1  g489(.A(G469), .B1(new_n675), .B2(G902), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n300), .A2(new_n304), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n677), .A2(new_n313), .A3(new_n189), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n676), .A2(new_n678), .A3(new_n188), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n553), .A2(new_n585), .A3(new_n615), .A4(new_n680), .ZN(new_n681));
  XOR2_X1   g495(.A(KEYINPUT41), .B(G113), .Z(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(KEYINPUT100), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n681), .B(new_n683), .ZN(G15));
  NAND4_X1  g498(.A1(new_n625), .A2(new_n553), .A3(new_n585), .A4(new_n680), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G116), .ZN(G18));
  INV_X1    g500(.A(new_n573), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n687), .B1(new_n570), .B2(new_n571), .ZN(new_n688));
  OAI211_X1 g502(.A(new_n575), .B(new_n576), .C1(new_n688), .C2(G902), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n574), .A2(new_n313), .A3(new_n577), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  AOI22_X1  g505(.A1(new_n691), .A2(new_n556), .B1(new_n581), .B2(new_n631), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n457), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n679), .A2(new_n603), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n553), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G119), .ZN(G21));
  NOR3_X1   g510(.A1(new_n679), .A2(new_n603), .A3(new_n660), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT103), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n584), .B(new_n698), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n485), .B1(new_n505), .B2(new_n527), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT101), .ZN(new_n701));
  OR3_X1    g515(.A1(new_n700), .A2(new_n510), .A3(new_n701), .ZN(new_n702));
  OAI21_X1  g516(.A(new_n701), .B1(new_n700), .B2(new_n510), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n702), .A2(new_n519), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(new_n459), .ZN(new_n705));
  XNOR2_X1  g519(.A(KEYINPUT102), .B(G472), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n589), .A2(new_n706), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n697), .A2(new_n699), .A3(new_n705), .A4(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G122), .ZN(G24));
  AND3_X1   g523(.A1(new_n707), .A2(new_n633), .A3(new_n705), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n665), .A2(new_n602), .A3(new_n601), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n679), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G125), .ZN(G27));
  INV_X1    g528(.A(KEYINPUT32), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n513), .A2(new_n715), .ZN(new_n716));
  AOI21_X1  g530(.A(KEYINPUT77), .B1(new_n549), .B2(G472), .ZN(new_n717));
  AOI211_X1 g531(.A(new_n525), .B(new_n543), .C1(new_n547), .C2(new_n548), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n716), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n552), .A2(KEYINPUT105), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT105), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n520), .A2(new_n721), .A3(KEYINPUT32), .A4(new_n459), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n699), .B1(new_n719), .B2(new_n723), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n363), .A2(new_n188), .A3(new_n364), .A4(new_n366), .ZN(new_n725));
  INV_X1    g539(.A(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT104), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n307), .A2(new_n727), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n302), .A2(KEYINPUT104), .A3(new_n292), .A4(new_n297), .ZN(new_n729));
  OAI211_X1 g543(.A(new_n728), .B(new_n729), .C1(new_n311), .C2(new_n297), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n306), .B1(new_n730), .B2(new_n313), .ZN(new_n731));
  OAI211_X1 g545(.A(new_n726), .B(new_n665), .C1(new_n305), .C2(new_n731), .ZN(new_n732));
  OAI21_X1  g546(.A(KEYINPUT42), .B1(new_n724), .B2(new_n732), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n305), .A2(new_n731), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n734), .A2(new_n725), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n427), .A2(new_n613), .A3(new_n638), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n736), .A2(KEYINPUT42), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n553), .A2(new_n585), .A3(new_n735), .A4(new_n737), .ZN(new_n738));
  AND3_X1   g552(.A1(new_n733), .A2(KEYINPUT106), .A3(new_n738), .ZN(new_n739));
  AOI21_X1  g553(.A(KEYINPUT106), .B1(new_n733), .B2(new_n738), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G131), .ZN(G33));
  NAND4_X1  g556(.A1(new_n553), .A2(new_n585), .A3(new_n640), .A4(new_n735), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G134), .ZN(G36));
  NOR2_X1   g558(.A1(new_n365), .A2(new_n600), .ZN(new_n745));
  INV_X1    g559(.A(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n428), .A2(new_n613), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(KEYINPUT43), .ZN(new_n748));
  OR3_X1    g562(.A1(new_n595), .A2(new_n692), .A3(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT44), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n746), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT45), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n312), .A2(new_n752), .ZN(new_n753));
  OAI211_X1 g567(.A(new_n753), .B(G469), .C1(new_n752), .C2(new_n730), .ZN(new_n754));
  NAND2_X1  g568(.A1(G469), .A2(G902), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT46), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n305), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n758), .B1(new_n757), .B2(new_n756), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(new_n188), .ZN(new_n760));
  INV_X1    g574(.A(new_n760), .ZN(new_n761));
  AND2_X1   g575(.A1(new_n761), .A2(new_n651), .ZN(new_n762));
  OAI211_X1 g576(.A(new_n751), .B(new_n762), .C1(new_n750), .C2(new_n749), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G137), .ZN(G39));
  NOR4_X1   g578(.A1(new_n553), .A2(new_n585), .A3(new_n736), .A4(new_n746), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n761), .A2(KEYINPUT47), .ZN(new_n766));
  AND2_X1   g580(.A1(new_n761), .A2(KEYINPUT47), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n765), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G140), .ZN(G42));
  INV_X1    g583(.A(new_n650), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n676), .A2(new_n678), .ZN(new_n771));
  OR2_X1    g585(.A1(new_n771), .A2(KEYINPUT49), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(KEYINPUT49), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n699), .A2(new_n188), .A3(new_n366), .ZN(new_n774));
  NOR3_X1   g588(.A1(new_n774), .A2(new_n657), .A3(new_n747), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n770), .A2(new_n772), .A3(new_n773), .A4(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT51), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n767), .A2(new_n766), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n778), .B1(new_n188), .B2(new_n771), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n748), .A2(new_n368), .ZN(new_n780));
  AND4_X1   g594(.A1(new_n699), .A2(new_n780), .A3(new_n705), .A4(new_n707), .ZN(new_n781));
  AND3_X1   g595(.A1(new_n779), .A2(new_n745), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n680), .A2(new_n745), .ZN(new_n783));
  NOR3_X1   g597(.A1(new_n783), .A2(new_n584), .A3(new_n368), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n770), .A2(new_n784), .ZN(new_n785));
  NOR3_X1   g599(.A1(new_n785), .A2(new_n427), .A3(new_n613), .ZN(new_n786));
  NOR3_X1   g600(.A1(new_n783), .A2(new_n748), .A3(new_n368), .ZN(new_n787));
  AND2_X1   g601(.A1(new_n787), .A2(new_n710), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT111), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  OAI21_X1  g605(.A(KEYINPUT111), .B1(new_n786), .B2(new_n788), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n781), .A2(new_n680), .ZN(new_n793));
  NOR3_X1   g607(.A1(new_n793), .A2(new_n366), .A3(new_n657), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(KEYINPUT50), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n791), .A2(new_n792), .A3(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT112), .ZN(new_n797));
  OR2_X1    g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n796), .A2(new_n797), .ZN(new_n799));
  AOI211_X1 g613(.A(new_n777), .B(new_n782), .C1(new_n798), .C2(new_n799), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n685), .A2(new_n681), .A3(new_n708), .A4(new_n695), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(KEYINPUT107), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n708), .A2(new_n695), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT107), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n803), .A2(new_n804), .A3(new_n681), .A4(new_n685), .ZN(new_n805));
  NOR3_X1   g619(.A1(new_n315), .A2(new_n639), .A3(new_n746), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n806), .A2(new_n553), .A3(new_n693), .ZN(new_n807));
  INV_X1    g621(.A(new_n732), .ZN(new_n808));
  AOI21_X1  g622(.A(KEYINPUT108), .B1(new_n710), .B2(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n707), .A2(new_n633), .A3(new_n705), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT108), .ZN(new_n811));
  NOR3_X1   g625(.A1(new_n810), .A2(new_n732), .A3(new_n811), .ZN(new_n812));
  OAI211_X1 g626(.A(new_n743), .B(new_n807), .C1(new_n809), .C2(new_n812), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n620), .B1(new_n427), .B2(new_n613), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n814), .A2(new_n372), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n593), .A2(new_n596), .A3(new_n815), .A4(new_n594), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n634), .A2(new_n816), .A3(new_n586), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n813), .A2(new_n817), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n741), .A2(new_n802), .A3(new_n805), .A4(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT53), .ZN(new_n821));
  AOI22_X1  g635(.A1(new_n553), .A2(new_n642), .B1(new_n710), .B2(new_n712), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n692), .A2(new_n188), .A3(new_n638), .ZN(new_n823));
  NOR4_X1   g637(.A1(new_n734), .A2(new_n823), .A3(new_n619), .A4(new_n660), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n824), .B1(new_n645), .B2(new_n648), .ZN(new_n825));
  AND3_X1   g639(.A1(new_n553), .A2(new_n667), .A3(KEYINPUT99), .ZN(new_n826));
  AOI21_X1  g640(.A(KEYINPUT99), .B1(new_n553), .B2(new_n667), .ZN(new_n827));
  OAI211_X1 g641(.A(new_n822), .B(new_n825), .C1(new_n826), .C2(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT109), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT52), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n828), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n828), .A2(new_n830), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n672), .A2(KEYINPUT52), .A3(new_n822), .A4(new_n825), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n832), .A2(new_n833), .A3(KEYINPUT109), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n820), .A2(new_n821), .A3(new_n831), .A4(new_n834), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n832), .A2(new_n833), .ZN(new_n836));
  OAI21_X1  g650(.A(KEYINPUT53), .B1(new_n819), .B2(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n835), .A2(KEYINPUT54), .A3(new_n837), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n821), .B1(new_n819), .B2(new_n836), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n733), .A2(KEYINPUT53), .A3(new_n738), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n801), .A2(new_n840), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n834), .A2(new_n818), .A3(new_n831), .A4(new_n841), .ZN(new_n842));
  XOR2_X1   g656(.A(KEYINPUT110), .B(KEYINPUT54), .Z(new_n843));
  NAND3_X1  g657(.A1(new_n839), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n838), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n795), .A2(new_n789), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n777), .B1(new_n846), .B2(new_n782), .ZN(new_n847));
  INV_X1    g661(.A(new_n724), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n787), .A2(new_n848), .ZN(new_n849));
  XNOR2_X1  g663(.A(new_n849), .B(KEYINPUT48), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n850), .B1(new_n614), .B2(new_n785), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n793), .A2(new_n619), .ZN(new_n852));
  OAI211_X1 g666(.A(G952), .B(new_n294), .C1(new_n852), .C2(KEYINPUT113), .ZN(new_n853));
  AOI211_X1 g667(.A(new_n851), .B(new_n853), .C1(KEYINPUT113), .C2(new_n852), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n847), .A2(new_n854), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n800), .A2(new_n845), .A3(new_n855), .ZN(new_n856));
  NOR2_X1   g670(.A1(G952), .A2(G953), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n776), .B1(new_n856), .B2(new_n857), .ZN(G75));
  NOR2_X1   g672(.A1(new_n294), .A2(G952), .ZN(new_n859));
  XOR2_X1   g673(.A(new_n859), .B(KEYINPUT116), .Z(new_n860));
  NAND2_X1  g674(.A1(new_n839), .A2(new_n842), .ZN(new_n861));
  INV_X1    g675(.A(new_n861), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n862), .A2(new_n313), .ZN(new_n863));
  AOI21_X1  g677(.A(KEYINPUT56), .B1(new_n863), .B2(G210), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n346), .A2(new_n348), .ZN(new_n865));
  XOR2_X1   g679(.A(new_n865), .B(KEYINPUT55), .Z(new_n866));
  NAND2_X1  g680(.A1(new_n336), .A2(new_n333), .ZN(new_n867));
  XNOR2_X1  g681(.A(new_n867), .B(KEYINPUT114), .ZN(new_n868));
  XNOR2_X1  g682(.A(new_n866), .B(new_n868), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n860), .B1(new_n864), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n864), .A2(new_n869), .ZN(new_n871));
  OR2_X1    g685(.A1(new_n871), .A2(KEYINPUT115), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(KEYINPUT115), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n870), .B1(new_n872), .B2(new_n873), .ZN(G51));
  INV_X1    g688(.A(new_n843), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n861), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n876), .A2(new_n844), .ZN(new_n877));
  INV_X1    g691(.A(new_n877), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n755), .B(KEYINPUT57), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n677), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  OR3_X1    g694(.A1(new_n862), .A2(new_n313), .A3(new_n754), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n859), .B1(new_n880), .B2(new_n881), .ZN(G54));
  NAND3_X1  g696(.A1(new_n863), .A2(KEYINPUT58), .A3(G475), .ZN(new_n883));
  OR3_X1    g697(.A1(new_n883), .A2(KEYINPUT117), .A3(new_n420), .ZN(new_n884));
  OAI21_X1  g698(.A(KEYINPUT117), .B1(new_n883), .B2(new_n420), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n859), .B1(new_n883), .B2(new_n420), .ZN(new_n886));
  AND3_X1   g700(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(G60));
  AND2_X1   g701(.A1(new_n605), .A2(new_n607), .ZN(new_n888));
  INV_X1    g702(.A(new_n845), .ZN(new_n889));
  XNOR2_X1  g703(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n611), .B(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(new_n891), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n888), .B1(new_n889), .B2(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(new_n860), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n888), .A2(new_n892), .ZN(new_n895));
  AND3_X1   g709(.A1(new_n839), .A2(new_n842), .A3(new_n843), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n843), .B1(new_n839), .B2(new_n842), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n895), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT119), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  OAI211_X1 g714(.A(KEYINPUT119), .B(new_n895), .C1(new_n896), .C2(new_n897), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n894), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n893), .B1(new_n902), .B2(KEYINPUT120), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT120), .ZN(new_n904));
  AOI211_X1 g718(.A(new_n904), .B(new_n894), .C1(new_n900), .C2(new_n901), .ZN(new_n905));
  OAI21_X1  g719(.A(KEYINPUT121), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(KEYINPUT119), .B1(new_n877), .B2(new_n895), .ZN(new_n907));
  INV_X1    g721(.A(new_n901), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n860), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(new_n904), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n902), .A2(KEYINPUT120), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT121), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n910), .A2(new_n911), .A3(new_n912), .A4(new_n893), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n906), .A2(new_n913), .ZN(G63));
  NAND2_X1  g728(.A1(G217), .A2(G902), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n915), .B(KEYINPUT60), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n916), .B1(new_n839), .B2(new_n842), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n631), .B(KEYINPUT122), .ZN(new_n918));
  AND3_X1   g732(.A1(new_n917), .A2(KEYINPUT123), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(KEYINPUT123), .B1(new_n917), .B2(new_n918), .ZN(new_n920));
  OAI221_X1 g734(.A(new_n860), .B1(new_n574), .B2(new_n917), .C1(new_n919), .C2(new_n920), .ZN(new_n921));
  XOR2_X1   g735(.A(new_n921), .B(KEYINPUT61), .Z(G66));
  AOI21_X1  g736(.A(new_n294), .B1(new_n369), .B2(G224), .ZN(new_n923));
  AND2_X1   g737(.A1(new_n805), .A2(new_n802), .ZN(new_n924));
  INV_X1    g738(.A(new_n817), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n923), .B1(new_n926), .B2(new_n294), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n868), .B1(G898), .B2(new_n294), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n927), .B(new_n928), .Z(G69));
  NOR2_X1   g743(.A1(new_n619), .A2(new_n660), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n762), .A2(new_n848), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n768), .A2(new_n931), .ZN(new_n932));
  AND2_X1   g746(.A1(new_n672), .A2(new_n822), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n763), .A2(new_n933), .ZN(new_n934));
  OR2_X1    g748(.A1(new_n934), .A2(KEYINPUT124), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n934), .A2(KEYINPUT124), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n932), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n741), .A2(new_n743), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(KEYINPUT125), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n937), .A2(new_n294), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n491), .A2(new_n499), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n941), .B(new_n417), .Z(new_n942));
  AOI21_X1  g756(.A(new_n942), .B1(G900), .B2(G953), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n940), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n663), .A2(new_n933), .ZN(new_n945));
  OR2_X1    g759(.A1(new_n945), .A2(KEYINPUT62), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n945), .A2(KEYINPUT62), .ZN(new_n947));
  NOR3_X1   g761(.A1(new_n652), .A2(new_n814), .A3(new_n746), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n948), .A2(new_n553), .A3(new_n585), .ZN(new_n949));
  AND3_X1   g763(.A1(new_n763), .A2(new_n768), .A3(new_n949), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n946), .A2(new_n947), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(new_n294), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(new_n942), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n944), .A2(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n294), .B1(G227), .B2(G900), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n955), .B(KEYINPUT126), .Z(new_n956));
  XNOR2_X1  g770(.A(new_n954), .B(new_n956), .ZN(G72));
  XNOR2_X1  g771(.A(new_n538), .B(KEYINPUT127), .ZN(new_n958));
  NAND4_X1  g772(.A1(new_n937), .A2(new_n924), .A3(new_n925), .A4(new_n939), .ZN(new_n959));
  NAND2_X1  g773(.A1(G472), .A2(G902), .ZN(new_n960));
  XOR2_X1   g774(.A(new_n960), .B(KEYINPUT63), .Z(new_n961));
  AOI211_X1 g775(.A(new_n485), .B(new_n958), .C1(new_n959), .C2(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n958), .A2(new_n485), .ZN(new_n963));
  OR2_X1    g777(.A1(new_n951), .A2(new_n926), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n963), .B1(new_n964), .B2(new_n961), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n540), .A2(new_n516), .ZN(new_n966));
  AND4_X1   g780(.A1(new_n837), .A2(new_n835), .A3(new_n961), .A4(new_n966), .ZN(new_n967));
  NOR4_X1   g781(.A1(new_n962), .A2(new_n965), .A3(new_n859), .A4(new_n967), .ZN(G57));
endmodule


