//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 1 1 1 0 1 1 1 0 1 0 1 1 1 0 0 1 0 0 1 1 1 0 0 1 0 1 0 0 1 1 1 0 1 1 0 1 0 0 0 0 1 0 1 1 0 0 1 1 1 0 1 1 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:44 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1079, new_n1080, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1139,
    new_n1140, new_n1141, new_n1142, new_n1143, new_n1144, new_n1145,
    new_n1146, new_n1147, new_n1148, new_n1149, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1174, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1226, new_n1227,
    new_n1228, new_n1229;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XNOR2_X1  g0003(.A(new_n203), .B(KEYINPUT64), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR3_X1   g0008(.A1(new_n207), .A2(new_n208), .A3(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XOR2_X1   g0010(.A(new_n210), .B(KEYINPUT0), .Z(new_n211));
  AOI22_X1  g0011(.A1(G77), .A2(G244), .B1(G87), .B2(G250), .ZN(new_n212));
  INV_X1    g0012(.A(G116), .ZN(new_n213));
  INV_X1    g0013(.A(G270), .ZN(new_n214));
  OAI21_X1  g0014(.A(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n216));
  INV_X1    g0016(.A(G226), .ZN(new_n217));
  INV_X1    g0017(.A(G68), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n216), .B1(new_n202), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  AOI211_X1 g0020(.A(new_n215), .B(new_n220), .C1(G97), .C2(G257), .ZN(new_n221));
  AOI21_X1  g0021(.A(new_n221), .B1(G1), .B2(G20), .ZN(new_n222));
  XOR2_X1   g0022(.A(new_n222), .B(KEYINPUT1), .Z(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G13), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n224), .A2(new_n208), .ZN(new_n225));
  INV_X1    g0025(.A(new_n201), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n226), .A2(G50), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  AOI211_X1 g0028(.A(new_n211), .B(new_n223), .C1(new_n225), .C2(new_n228), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT2), .B(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT65), .B(G250), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n233), .B(new_n237), .ZN(G358));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XOR2_X1   g0039(.A(G107), .B(G116), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT66), .ZN(new_n242));
  XOR2_X1   g0042(.A(G68), .B(G77), .Z(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G58), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  INV_X1    g0046(.A(G13), .ZN(new_n247));
  NOR3_X1   g0047(.A1(new_n247), .A2(new_n208), .A3(G1), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(new_n202), .ZN(new_n250));
  NAND3_X1  g0050(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(new_n224), .ZN(new_n252));
  AOI21_X1  g0052(.A(new_n252), .B1(new_n207), .B2(G20), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n250), .B1(new_n253), .B2(new_n202), .ZN(new_n254));
  XOR2_X1   g0054(.A(new_n254), .B(KEYINPUT67), .Z(new_n255));
  NAND2_X1  g0055(.A1(new_n204), .A2(G20), .ZN(new_n256));
  INV_X1    g0056(.A(G150), .ZN(new_n257));
  INV_X1    g0057(.A(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n208), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n208), .A2(G33), .ZN(new_n260));
  XNOR2_X1  g0060(.A(KEYINPUT8), .B(G58), .ZN(new_n261));
  OAI221_X1 g0061(.A(new_n256), .B1(new_n257), .B2(new_n259), .C1(new_n260), .C2(new_n261), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n255), .B1(new_n252), .B2(new_n262), .ZN(new_n263));
  AND2_X1   g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  NOR2_X1   g0064(.A1(KEYINPUT3), .A2(G33), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G1698), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n266), .B1(G222), .B2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G223), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n268), .B1(new_n269), .B2(new_n267), .ZN(new_n270));
  INV_X1    g0070(.A(G41), .ZN(new_n271));
  OAI211_X1 g0071(.A(G1), .B(G13), .C1(new_n258), .C2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  XNOR2_X1  g0073(.A(KEYINPUT3), .B(G33), .ZN(new_n274));
  OAI211_X1 g0074(.A(new_n270), .B(new_n273), .C1(G77), .C2(new_n274), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n276));
  INV_X1    g0076(.A(G274), .ZN(new_n277));
  OR2_X1    g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n272), .A2(new_n276), .ZN(new_n279));
  OAI211_X1 g0079(.A(new_n275), .B(new_n278), .C1(new_n217), .C2(new_n279), .ZN(new_n280));
  AOI22_X1  g0080(.A1(new_n263), .A2(KEYINPUT9), .B1(G200), .B2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G190), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n263), .A2(KEYINPUT9), .ZN(new_n283));
  AND2_X1   g0083(.A1(new_n283), .A2(KEYINPUT72), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n283), .A2(KEYINPUT72), .ZN(new_n285));
  OAI221_X1 g0085(.A(new_n281), .B1(new_n282), .B2(new_n280), .C1(new_n284), .C2(new_n285), .ZN(new_n286));
  XNOR2_X1  g0086(.A(new_n286), .B(KEYINPUT10), .ZN(new_n287));
  INV_X1    g0087(.A(G169), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n263), .B1(new_n288), .B2(new_n280), .ZN(new_n289));
  OR2_X1    g0089(.A1(new_n280), .A2(G179), .ZN(new_n290));
  AND2_X1   g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n287), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n253), .A2(G77), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT68), .ZN(new_n295));
  XNOR2_X1  g0095(.A(new_n294), .B(new_n295), .ZN(new_n296));
  XOR2_X1   g0096(.A(KEYINPUT15), .B(G87), .Z(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  OAI22_X1  g0098(.A1(new_n298), .A2(new_n260), .B1(new_n259), .B2(new_n261), .ZN(new_n299));
  INV_X1    g0099(.A(G77), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n208), .A2(new_n300), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n252), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n248), .A2(new_n300), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n296), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(KEYINPUT69), .ZN(new_n305));
  NAND2_X1  g0105(.A1(G238), .A2(G1698), .ZN(new_n306));
  INV_X1    g0106(.A(G232), .ZN(new_n307));
  OAI211_X1 g0107(.A(new_n274), .B(new_n306), .C1(new_n307), .C2(G1698), .ZN(new_n308));
  OAI211_X1 g0108(.A(new_n308), .B(new_n273), .C1(G107), .C2(new_n274), .ZN(new_n309));
  INV_X1    g0109(.A(new_n279), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(G244), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n309), .A2(new_n278), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(G200), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT69), .ZN(new_n314));
  NAND4_X1  g0114(.A1(new_n296), .A2(new_n302), .A3(new_n314), .A4(new_n303), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n305), .A2(new_n313), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(KEYINPUT70), .ZN(new_n317));
  INV_X1    g0117(.A(new_n312), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(G190), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT70), .ZN(new_n320));
  NAND4_X1  g0120(.A1(new_n305), .A2(new_n320), .A3(new_n313), .A4(new_n315), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n317), .A2(new_n319), .A3(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT16), .ZN(new_n324));
  AND2_X1   g0124(.A1(G58), .A2(G68), .ZN(new_n325));
  OAI21_X1  g0125(.A(G20), .B1(new_n325), .B2(new_n201), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n208), .A2(new_n258), .A3(G159), .ZN(new_n327));
  AND3_X1   g0127(.A1(new_n326), .A2(KEYINPUT73), .A3(new_n327), .ZN(new_n328));
  AOI21_X1  g0128(.A(KEYINPUT73), .B1(new_n326), .B2(new_n327), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT7), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n331), .B1(new_n274), .B2(G20), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n266), .A2(KEYINPUT7), .A3(new_n208), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n218), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n324), .B1(new_n330), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n326), .A2(new_n327), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT73), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n326), .A2(KEYINPUT73), .A3(new_n327), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  AOI21_X1  g0140(.A(KEYINPUT7), .B1(new_n266), .B2(new_n208), .ZN(new_n341));
  NOR4_X1   g0141(.A1(new_n264), .A2(new_n265), .A3(new_n331), .A4(G20), .ZN(new_n342));
  OAI21_X1  g0142(.A(G68), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n340), .A2(new_n343), .A3(KEYINPUT16), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n335), .A2(new_n252), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n249), .A2(new_n261), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n346), .B1(new_n253), .B2(new_n261), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n278), .B1(new_n279), .B2(new_n307), .ZN(new_n349));
  OAI211_X1 g0149(.A(G223), .B(new_n267), .C1(new_n264), .C2(new_n265), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT74), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND4_X1  g0152(.A1(new_n274), .A2(KEYINPUT74), .A3(G223), .A4(new_n267), .ZN(new_n353));
  NAND2_X1  g0153(.A1(G33), .A2(G87), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n274), .A2(G226), .A3(G1698), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n352), .A2(new_n353), .A3(new_n354), .A4(new_n355), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n349), .B1(new_n356), .B2(new_n273), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(G179), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n358), .B1(new_n288), .B2(new_n357), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n348), .A2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT18), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n348), .A2(new_n359), .A3(KEYINPUT18), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n362), .A2(KEYINPUT75), .A3(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT17), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n356), .A2(new_n273), .ZN(new_n366));
  INV_X1    g0166(.A(new_n349), .ZN(new_n367));
  AOI21_X1  g0167(.A(G200), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  AOI211_X1 g0168(.A(G190), .B(new_n349), .C1(new_n356), .C2(new_n273), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n365), .B1(new_n348), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n357), .A2(new_n282), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n372), .B1(G200), .B2(new_n357), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n373), .A2(KEYINPUT17), .A3(new_n347), .A4(new_n345), .ZN(new_n374));
  AND2_X1   g0174(.A1(new_n371), .A2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT75), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n360), .A2(new_n376), .A3(new_n361), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n364), .A2(new_n375), .A3(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT13), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n217), .A2(new_n267), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n274), .B(new_n381), .C1(G232), .C2(new_n267), .ZN(new_n382));
  NAND2_X1  g0182(.A1(G33), .A2(G97), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n272), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n278), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n279), .A2(new_n219), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n380), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  NOR4_X1   g0189(.A1(new_n384), .A2(KEYINPUT13), .A3(new_n387), .A4(new_n385), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  OAI21_X1  g0191(.A(KEYINPUT14), .B1(new_n391), .B2(new_n288), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(G179), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT14), .ZN(new_n394));
  OAI211_X1 g0194(.A(new_n394), .B(G169), .C1(new_n389), .C2(new_n390), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n392), .A2(new_n393), .A3(new_n395), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n208), .A2(G68), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n397), .A2(new_n207), .A3(G13), .ZN(new_n398));
  XOR2_X1   g0198(.A(new_n398), .B(KEYINPUT12), .Z(new_n399));
  NAND2_X1  g0199(.A1(new_n253), .A2(G68), .ZN(new_n400));
  OAI22_X1  g0200(.A1(new_n259), .A2(new_n202), .B1(new_n260), .B2(new_n300), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n252), .B1(new_n401), .B2(new_n397), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT11), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n400), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  AOI211_X1 g0204(.A(new_n399), .B(new_n404), .C1(new_n403), .C2(new_n402), .ZN(new_n405));
  INV_X1    g0205(.A(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n396), .A2(new_n406), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n304), .B1(G169), .B2(new_n318), .ZN(new_n408));
  OR2_X1    g0208(.A1(new_n408), .A2(KEYINPUT71), .ZN(new_n409));
  INV_X1    g0209(.A(G179), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n318), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n408), .A2(KEYINPUT71), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n409), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n406), .B1(new_n391), .B2(G190), .ZN(new_n414));
  INV_X1    g0214(.A(G200), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n414), .B1(new_n415), .B2(new_n391), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n379), .A2(new_n407), .A3(new_n413), .A4(new_n416), .ZN(new_n417));
  OAI21_X1  g0217(.A(KEYINPUT23), .B1(new_n208), .B2(G107), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT23), .ZN(new_n419));
  INV_X1    g0219(.A(G107), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n419), .A2(new_n420), .A3(G20), .ZN(new_n421));
  NAND2_X1  g0221(.A1(G33), .A2(G116), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n418), .B(new_n421), .C1(G20), .C2(new_n422), .ZN(new_n423));
  XNOR2_X1  g0223(.A(new_n423), .B(KEYINPUT82), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n274), .A2(new_n208), .A3(G87), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(KEYINPUT81), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT81), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n274), .A2(new_n427), .A3(new_n208), .A4(G87), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n426), .A2(KEYINPUT22), .A3(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT22), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n425), .A2(KEYINPUT81), .A3(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n424), .A2(new_n429), .A3(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT83), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n424), .A2(new_n429), .A3(KEYINPUT83), .A4(new_n431), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n434), .A2(KEYINPUT24), .A3(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT24), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n432), .A2(new_n433), .A3(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n436), .A2(new_n252), .A3(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(G250), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(new_n267), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n274), .B(new_n441), .C1(G257), .C2(new_n267), .ZN(new_n442));
  NAND2_X1  g0242(.A1(G33), .A2(G294), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n272), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT5), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT77), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n445), .B1(new_n446), .B2(G41), .ZN(new_n447));
  INV_X1    g0247(.A(G45), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n448), .A2(G1), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n271), .A2(KEYINPUT77), .A3(KEYINPUT5), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n447), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(new_n272), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n444), .B1(G264), .B2(new_n453), .ZN(new_n454));
  OR2_X1    g0254(.A1(new_n451), .A2(new_n277), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(new_n415), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n457), .B1(G190), .B2(new_n456), .ZN(new_n458));
  NOR4_X1   g0258(.A1(new_n247), .A2(new_n208), .A3(G1), .A4(G107), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT25), .ZN(new_n460));
  OR2_X1    g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n252), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n207), .A2(G33), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n249), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  AOI22_X1  g0265(.A1(new_n465), .A2(G107), .B1(new_n460), .B2(new_n459), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n439), .A2(new_n458), .A3(new_n461), .A4(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n274), .A2(new_n208), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT19), .ZN(new_n469));
  INV_X1    g0269(.A(G87), .ZN(new_n470));
  INV_X1    g0270(.A(G97), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n470), .A2(new_n471), .A3(new_n420), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n383), .A2(new_n208), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n469), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NOR3_X1   g0274(.A1(new_n383), .A2(KEYINPUT19), .A3(G20), .ZN(new_n475));
  OAI22_X1  g0275(.A1(new_n218), .A2(new_n468), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT79), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  OAI221_X1 g0278(.A(KEYINPUT79), .B1(new_n474), .B2(new_n475), .C1(new_n218), .C2(new_n468), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n478), .A2(new_n479), .A3(new_n252), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n298), .A2(new_n248), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n480), .B(new_n481), .C1(new_n298), .C2(new_n464), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n219), .A2(new_n267), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n274), .B(new_n483), .C1(G244), .C2(new_n267), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n272), .B1(new_n484), .B2(new_n422), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT78), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n277), .B1(new_n486), .B2(new_n440), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(new_n449), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n486), .B(G250), .C1(new_n448), .C2(G1), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n273), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n288), .B1(new_n485), .B2(new_n490), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n485), .A2(new_n490), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(new_n410), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n482), .A2(new_n491), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n492), .A2(G190), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n495), .B1(new_n415), .B2(new_n492), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n465), .A2(G87), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n480), .A2(new_n481), .A3(new_n497), .ZN(new_n498));
  OR2_X1    g0298(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  AND3_X1   g0299(.A1(new_n467), .A2(new_n494), .A3(new_n499), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n249), .A2(G97), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n464), .A2(new_n471), .ZN(new_n502));
  OAI21_X1  g0302(.A(G107), .B1(new_n341), .B2(new_n342), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT6), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n471), .A2(new_n420), .ZN(new_n505));
  NOR2_X1   g0305(.A1(G97), .A2(G107), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n420), .A2(KEYINPUT6), .A3(G97), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(G20), .ZN(new_n510));
  OAI211_X1 g0310(.A(new_n503), .B(new_n510), .C1(new_n300), .C2(new_n259), .ZN(new_n511));
  AOI211_X1 g0311(.A(new_n501), .B(new_n502), .C1(new_n511), .C2(new_n252), .ZN(new_n512));
  INV_X1    g0312(.A(G257), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n455), .B1(new_n513), .B2(new_n452), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n266), .A2(new_n440), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT4), .ZN(new_n516));
  OAI21_X1  g0316(.A(G1698), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n274), .A2(G244), .ZN(new_n518));
  AOI22_X1  g0318(.A1(new_n518), .A2(new_n516), .B1(G33), .B2(G283), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n274), .A2(KEYINPUT4), .A3(G244), .A4(new_n267), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n517), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n514), .B1(new_n521), .B2(new_n273), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(G190), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n521), .A2(new_n273), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT76), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n518), .A2(new_n516), .ZN(new_n527));
  NAND2_X1  g0327(.A1(G33), .A2(G283), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n527), .A2(new_n528), .A3(new_n520), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n274), .A2(G250), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n267), .B1(new_n530), .B2(KEYINPUT4), .ZN(new_n531));
  OAI211_X1 g0331(.A(KEYINPUT76), .B(new_n273), .C1(new_n529), .C2(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n514), .B1(new_n526), .B2(new_n532), .ZN(new_n533));
  OAI211_X1 g0333(.A(new_n512), .B(new_n523), .C1(new_n533), .C2(new_n415), .ZN(new_n534));
  INV_X1    g0334(.A(new_n514), .ZN(new_n535));
  INV_X1    g0335(.A(new_n532), .ZN(new_n536));
  AOI21_X1  g0336(.A(KEYINPUT76), .B1(new_n521), .B2(new_n273), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n410), .B(new_n535), .C1(new_n536), .C2(new_n537), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n501), .B1(new_n511), .B2(new_n252), .ZN(new_n539));
  INV_X1    g0339(.A(new_n502), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  OR2_X1    g0341(.A1(new_n522), .A2(G169), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n538), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n534), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(G264), .A2(G1698), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n274), .B(new_n545), .C1(new_n513), .C2(G1698), .ZN(new_n546));
  INV_X1    g0346(.A(G303), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n266), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n546), .A2(new_n273), .A3(new_n548), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n549), .B(new_n455), .C1(new_n214), .C2(new_n452), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n249), .A2(G116), .A3(new_n462), .A4(new_n463), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n248), .A2(new_n213), .ZN(new_n552));
  AOI22_X1  g0352(.A1(new_n251), .A2(new_n224), .B1(G20), .B2(new_n213), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n528), .B(new_n208), .C1(G33), .C2(new_n471), .ZN(new_n554));
  AND3_X1   g0354(.A1(new_n553), .A2(KEYINPUT20), .A3(new_n554), .ZN(new_n555));
  AOI21_X1  g0355(.A(KEYINPUT20), .B1(new_n553), .B2(new_n554), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n551), .B(new_n552), .C1(new_n555), .C2(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n550), .A2(G169), .A3(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT21), .ZN(new_n559));
  AND3_X1   g0359(.A1(new_n558), .A2(KEYINPUT80), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g0360(.A(KEYINPUT80), .B1(new_n558), .B2(new_n559), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AND3_X1   g0362(.A1(new_n550), .A2(KEYINPUT21), .A3(G169), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n550), .A2(new_n410), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n557), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n550), .A2(G200), .ZN(new_n566));
  INV_X1    g0366(.A(new_n557), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n566), .B(new_n567), .C1(new_n282), .C2(new_n550), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n562), .A2(new_n565), .A3(new_n568), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n544), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n439), .A2(new_n461), .A3(new_n466), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n456), .A2(G179), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n572), .B1(new_n288), .B2(new_n456), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n500), .A2(new_n570), .A3(new_n574), .ZN(new_n575));
  NOR4_X1   g0375(.A1(new_n293), .A2(new_n323), .A3(new_n417), .A4(new_n575), .ZN(G372));
  NOR3_X1   g0376(.A1(new_n293), .A2(new_n323), .A3(new_n417), .ZN(new_n577));
  XNOR2_X1  g0377(.A(new_n491), .B(KEYINPUT84), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n578), .A2(new_n493), .A3(new_n482), .ZN(new_n579));
  INV_X1    g0379(.A(new_n579), .ZN(new_n580));
  AND2_X1   g0380(.A1(new_n534), .A2(new_n543), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n498), .A2(KEYINPUT85), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT85), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n480), .A2(new_n583), .A3(new_n481), .A4(new_n497), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n496), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  AND3_X1   g0386(.A1(new_n581), .A2(new_n467), .A3(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT86), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n562), .A2(new_n588), .A3(new_n565), .ZN(new_n589));
  INV_X1    g0389(.A(new_n589), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n588), .B1(new_n562), .B2(new_n565), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n574), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n580), .B1(new_n587), .B2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT87), .ZN(new_n594));
  NOR3_X1   g0394(.A1(new_n580), .A2(new_n585), .A3(new_n543), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n594), .B1(new_n595), .B2(KEYINPUT26), .ZN(new_n596));
  INV_X1    g0396(.A(new_n543), .ZN(new_n597));
  AND3_X1   g0397(.A1(new_n597), .A2(new_n494), .A3(new_n499), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(KEYINPUT26), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n586), .A2(new_n597), .A3(new_n579), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT26), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n600), .A2(KEYINPUT87), .A3(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n596), .A2(new_n599), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n593), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n577), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n362), .A2(new_n363), .ZN(new_n606));
  INV_X1    g0406(.A(new_n407), .ZN(new_n607));
  INV_X1    g0407(.A(new_n413), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n607), .B1(new_n608), .B2(new_n416), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n371), .A2(new_n374), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n606), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n291), .B1(new_n287), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n605), .A2(new_n612), .ZN(G369));
  NOR2_X1   g0413(.A1(new_n247), .A2(G20), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(new_n207), .ZN(new_n615));
  OR2_X1    g0415(.A1(new_n615), .A2(KEYINPUT27), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(KEYINPUT27), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n616), .A2(G213), .A3(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(G343), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n571), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(new_n467), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(new_n574), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n623), .B1(new_n574), .B2(new_n620), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n562), .A2(new_n565), .ZN(new_n625));
  INV_X1    g0425(.A(new_n620), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n574), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n628), .B1(new_n629), .B2(new_n626), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n625), .A2(KEYINPUT86), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n626), .A2(new_n567), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n631), .A2(new_n589), .A3(new_n632), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n633), .B1(new_n569), .B2(new_n632), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(G330), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n635), .A2(new_n624), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n630), .A2(new_n637), .ZN(G399));
  INV_X1    g0438(.A(new_n209), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n639), .A2(G41), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n472), .A2(G116), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n641), .A2(G1), .A3(new_n642), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n643), .B1(new_n227), .B2(new_n641), .ZN(new_n644));
  XNOR2_X1  g0444(.A(new_n644), .B(KEYINPUT28), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n604), .A2(new_n626), .ZN(new_n646));
  OR2_X1    g0446(.A1(new_n646), .A2(KEYINPUT29), .ZN(new_n647));
  OAI21_X1  g0447(.A(KEYINPUT31), .B1(new_n575), .B2(new_n620), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n564), .A2(new_n522), .A3(new_n454), .A4(new_n492), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT30), .ZN(new_n650));
  OR2_X1    g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n649), .A2(new_n650), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n535), .B1(new_n536), .B2(new_n537), .ZN(new_n653));
  INV_X1    g0453(.A(new_n492), .ZN(new_n654));
  AND2_X1   g0454(.A1(new_n550), .A2(new_n410), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n653), .A2(new_n456), .A3(new_n654), .A4(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n651), .A2(new_n652), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(new_n620), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n648), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n656), .A2(new_n652), .ZN(new_n660));
  XOR2_X1   g0460(.A(new_n660), .B(KEYINPUT88), .Z(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(new_n651), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n662), .A2(KEYINPUT31), .A3(new_n620), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n659), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(G330), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n587), .B1(new_n625), .B2(new_n629), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n595), .A2(KEYINPUT26), .ZN(new_n667));
  OAI211_X1 g0467(.A(new_n667), .B(KEYINPUT89), .C1(KEYINPUT26), .C2(new_n598), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n579), .B1(new_n667), .B2(KEYINPUT89), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n626), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(KEYINPUT29), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n647), .A2(new_n665), .A3(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n645), .B1(new_n674), .B2(G1), .ZN(G364));
  NOR2_X1   g0475(.A1(new_n208), .A2(new_n282), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n410), .A2(G200), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(G322), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n266), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n410), .A2(new_n415), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n208), .A2(G190), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(G317), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(KEYINPUT33), .ZN(new_n686));
  OR2_X1    g0486(.A1(new_n685), .A2(KEYINPUT33), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n684), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n415), .A2(G179), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n676), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(G311), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n682), .A2(new_n677), .ZN(new_n692));
  OAI221_X1 g0492(.A(new_n688), .B1(new_n547), .B2(new_n690), .C1(new_n691), .C2(new_n692), .ZN(new_n693));
  NOR2_X1   g0493(.A1(G179), .A2(G200), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n682), .A2(new_n694), .ZN(new_n695));
  OR2_X1    g0495(.A1(new_n695), .A2(KEYINPUT92), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n695), .A2(KEYINPUT92), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  AOI211_X1 g0499(.A(new_n680), .B(new_n693), .C1(G329), .C2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n676), .A2(new_n681), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(G326), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n208), .B1(new_n694), .B2(G190), .ZN(new_n704));
  AND2_X1   g0504(.A1(new_n704), .A2(KEYINPUT93), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n704), .A2(KEYINPUT93), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(G294), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n703), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(KEYINPUT94), .ZN(new_n710));
  AND2_X1   g0510(.A1(new_n700), .A2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(G283), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n682), .A2(new_n689), .ZN(new_n713));
  OAI221_X1 g0513(.A(new_n711), .B1(KEYINPUT94), .B2(new_n709), .C1(new_n712), .C2(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n713), .A2(new_n420), .ZN(new_n715));
  INV_X1    g0515(.A(new_n690), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n266), .B1(new_n716), .B2(G87), .ZN(new_n717));
  OAI221_X1 g0517(.A(new_n717), .B1(new_n202), .B2(new_n701), .C1(new_n218), .C2(new_n683), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT32), .ZN(new_n719));
  INV_X1    g0519(.A(G159), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n698), .A2(new_n720), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n718), .B1(new_n719), .B2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n721), .ZN(new_n723));
  INV_X1    g0523(.A(new_n707), .ZN(new_n724));
  AOI22_X1  g0524(.A1(new_n723), .A2(KEYINPUT32), .B1(G97), .B2(new_n724), .ZN(new_n725));
  XNOR2_X1  g0525(.A(new_n678), .B(KEYINPUT90), .ZN(new_n726));
  INV_X1    g0526(.A(new_n692), .ZN(new_n727));
  AOI22_X1  g0527(.A1(new_n726), .A2(G58), .B1(G77), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(KEYINPUT91), .ZN(new_n729));
  OR2_X1    g0529(.A1(new_n728), .A2(KEYINPUT91), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n722), .A2(new_n725), .A3(new_n729), .A4(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n714), .B1(new_n715), .B2(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n224), .B1(G20), .B2(new_n288), .ZN(new_n733));
  NOR2_X1   g0533(.A1(G13), .A2(G33), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(G20), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(new_n733), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n639), .A2(new_n274), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n228), .A2(new_n448), .ZN(new_n739));
  OAI211_X1 g0539(.A(new_n738), .B(new_n739), .C1(new_n245), .C2(new_n448), .ZN(new_n740));
  INV_X1    g0540(.A(G355), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n274), .A2(new_n209), .ZN(new_n742));
  OAI221_X1 g0542(.A(new_n740), .B1(G116), .B2(new_n209), .C1(new_n741), .C2(new_n742), .ZN(new_n743));
  AOI22_X1  g0543(.A1(new_n732), .A2(new_n733), .B1(new_n737), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n614), .A2(G45), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n641), .A2(G1), .A3(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n736), .ZN(new_n748));
  OAI211_X1 g0548(.A(new_n744), .B(new_n747), .C1(new_n634), .C2(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n634), .A2(G330), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n635), .A2(new_n746), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n749), .B1(new_n750), .B2(new_n751), .ZN(G396));
  NAND2_X1  g0552(.A1(new_n304), .A2(new_n620), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n322), .A2(new_n413), .A3(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(KEYINPUT97), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  OR2_X1    g0556(.A1(new_n413), .A2(new_n753), .ZN(new_n757));
  NAND4_X1  g0557(.A1(new_n322), .A2(new_n413), .A3(KEYINPUT97), .A4(new_n753), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n756), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  AND3_X1   g0559(.A1(new_n596), .A2(new_n599), .A3(new_n602), .ZN(new_n760));
  AOI22_X1  g0560(.A1(new_n631), .A2(new_n589), .B1(new_n571), .B2(new_n573), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n581), .A2(new_n467), .A3(new_n586), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n579), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  OAI211_X1 g0563(.A(new_n626), .B(new_n759), .C1(new_n760), .C2(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(KEYINPUT98), .ZN(new_n765));
  XNOR2_X1  g0565(.A(new_n665), .B(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n759), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n646), .A2(new_n767), .ZN(new_n768));
  XOR2_X1   g0568(.A(new_n766), .B(new_n768), .Z(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(new_n746), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n726), .A2(G143), .ZN(new_n771));
  AOI22_X1  g0571(.A1(new_n702), .A2(G137), .B1(new_n684), .B2(G150), .ZN(new_n772));
  OAI211_X1 g0572(.A(new_n771), .B(new_n772), .C1(new_n720), .C2(new_n692), .ZN(new_n773));
  INV_X1    g0573(.A(KEYINPUT34), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(G58), .ZN(new_n776));
  OAI221_X1 g0576(.A(new_n274), .B1(new_n202), .B2(new_n690), .C1(new_n707), .C2(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n773), .A2(new_n774), .ZN(new_n779));
  INV_X1    g0579(.A(new_n713), .ZN(new_n780));
  AOI22_X1  g0580(.A1(new_n699), .A2(G132), .B1(G68), .B2(new_n780), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n778), .A2(new_n779), .A3(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n692), .A2(new_n213), .ZN(new_n783));
  OAI22_X1  g0583(.A1(new_n701), .A2(new_n547), .B1(new_n678), .B2(new_n708), .ZN(new_n784));
  OAI22_X1  g0584(.A1(new_n683), .A2(new_n712), .B1(new_n713), .B2(new_n470), .ZN(new_n785));
  AOI211_X1 g0585(.A(new_n784), .B(new_n785), .C1(new_n724), .C2(G97), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n266), .B1(new_n690), .B2(new_n420), .ZN(new_n787));
  XNOR2_X1  g0587(.A(new_n787), .B(KEYINPUT95), .ZN(new_n788));
  OAI211_X1 g0588(.A(new_n786), .B(new_n788), .C1(new_n691), .C2(new_n698), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n782), .B1(new_n783), .B2(new_n789), .ZN(new_n790));
  XOR2_X1   g0590(.A(new_n790), .B(KEYINPUT96), .Z(new_n791));
  AOI21_X1  g0591(.A(new_n746), .B1(new_n791), .B2(new_n733), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n733), .A2(new_n734), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(new_n300), .ZN(new_n794));
  OAI211_X1 g0594(.A(new_n792), .B(new_n794), .C1(new_n735), .C2(new_n759), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n770), .A2(new_n795), .ZN(G384));
  INV_X1    g0596(.A(KEYINPUT102), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n406), .A2(new_n620), .ZN(new_n798));
  INV_X1    g0598(.A(KEYINPUT101), .ZN(new_n799));
  AND3_X1   g0599(.A1(new_n396), .A2(new_n799), .A3(new_n406), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n799), .B1(new_n396), .B2(new_n406), .ZN(new_n801));
  OAI211_X1 g0601(.A(new_n416), .B(new_n798), .C1(new_n800), .C2(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n607), .A2(new_n620), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n797), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n802), .A2(new_n797), .A3(new_n803), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n657), .A2(KEYINPUT31), .A3(new_n620), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n659), .A2(new_n808), .ZN(new_n809));
  AND3_X1   g0609(.A1(new_n807), .A2(new_n809), .A3(new_n759), .ZN(new_n810));
  INV_X1    g0610(.A(KEYINPUT107), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n373), .A2(new_n347), .A3(new_n345), .ZN(new_n812));
  INV_X1    g0612(.A(new_n618), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n348), .A2(new_n813), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n812), .A2(new_n360), .A3(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n815), .A2(KEYINPUT37), .ZN(new_n816));
  AND3_X1   g0616(.A1(new_n345), .A2(KEYINPUT103), .A3(new_n347), .ZN(new_n817));
  AOI21_X1  g0617(.A(KEYINPUT103), .B1(new_n345), .B2(new_n347), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n359), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n813), .B1(new_n817), .B2(new_n818), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n819), .A2(new_n820), .A3(new_n812), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n816), .B1(new_n821), .B2(KEYINPUT37), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  AOI211_X1 g0623(.A(KEYINPUT75), .B(KEYINPUT18), .C1(new_n348), .C2(new_n359), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n610), .A2(new_n824), .ZN(new_n825));
  AOI211_X1 g0625(.A(KEYINPUT104), .B(new_n820), .C1(new_n825), .C2(new_n364), .ZN(new_n826));
  INV_X1    g0626(.A(KEYINPUT104), .ZN(new_n827));
  INV_X1    g0627(.A(new_n820), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n827), .B1(new_n378), .B2(new_n828), .ZN(new_n829));
  OAI211_X1 g0629(.A(KEYINPUT38), .B(new_n823), .C1(new_n826), .C2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(KEYINPUT38), .ZN(new_n831));
  XOR2_X1   g0631(.A(new_n815), .B(KEYINPUT37), .Z(new_n832));
  AOI21_X1  g0632(.A(new_n814), .B1(new_n375), .B2(new_n606), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n831), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n830), .A2(new_n834), .ZN(new_n835));
  NAND4_X1  g0635(.A1(new_n810), .A2(new_n811), .A3(KEYINPUT40), .A4(new_n835), .ZN(new_n836));
  NAND4_X1  g0636(.A1(new_n807), .A2(new_n809), .A3(KEYINPUT40), .A4(new_n759), .ZN(new_n837));
  INV_X1    g0637(.A(new_n835), .ZN(new_n838));
  OAI21_X1  g0638(.A(KEYINPUT107), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT40), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n807), .A2(new_n809), .A3(new_n759), .ZN(new_n841));
  AND3_X1   g0641(.A1(new_n362), .A2(KEYINPUT75), .A3(new_n363), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n377), .A2(new_n371), .A3(new_n374), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n828), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(KEYINPUT104), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n378), .A2(new_n827), .A3(new_n828), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(KEYINPUT38), .B1(new_n847), .B2(new_n823), .ZN(new_n848));
  AOI211_X1 g0648(.A(new_n831), .B(new_n822), .C1(new_n845), .C2(new_n846), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n840), .B1(new_n841), .B2(new_n850), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n836), .A2(new_n839), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n577), .A2(new_n809), .ZN(new_n853));
  XOR2_X1   g0653(.A(new_n852), .B(new_n853), .Z(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(G330), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT106), .ZN(new_n856));
  OAI21_X1  g0656(.A(KEYINPUT39), .B1(new_n848), .B2(new_n849), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT39), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n830), .A2(new_n858), .A3(new_n834), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n859), .A2(KEYINPUT105), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT105), .ZN(new_n861));
  NAND4_X1  g0661(.A1(new_n830), .A2(new_n861), .A3(new_n858), .A4(new_n834), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n857), .A2(new_n860), .A3(new_n862), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n800), .A2(new_n801), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(new_n626), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n863), .A2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n850), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n413), .A2(new_n620), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  AND3_X1   g0670(.A1(new_n764), .A2(KEYINPUT100), .A3(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(KEYINPUT100), .B1(new_n764), .B2(new_n870), .ZN(new_n872));
  OAI211_X1 g0672(.A(new_n868), .B(new_n807), .C1(new_n871), .C2(new_n872), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n606), .A2(new_n813), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  AND4_X1   g0675(.A1(new_n856), .A2(new_n867), .A3(new_n873), .A4(new_n875), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n874), .B1(new_n863), .B2(new_n866), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n856), .B1(new_n877), .B2(new_n873), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  XNOR2_X1  g0679(.A(new_n855), .B(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n647), .A2(new_n672), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(new_n577), .ZN(new_n882));
  AND2_X1   g0682(.A1(new_n882), .A2(new_n612), .ZN(new_n883));
  XNOR2_X1  g0683(.A(new_n880), .B(new_n883), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n884), .B1(new_n207), .B2(new_n614), .ZN(new_n885));
  XNOR2_X1  g0685(.A(new_n509), .B(KEYINPUT99), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n213), .B1(new_n886), .B2(KEYINPUT35), .ZN(new_n887));
  OAI211_X1 g0687(.A(new_n887), .B(new_n225), .C1(KEYINPUT35), .C2(new_n886), .ZN(new_n888));
  XNOR2_X1  g0688(.A(new_n888), .B(KEYINPUT36), .ZN(new_n889));
  OAI21_X1  g0689(.A(G77), .B1(new_n776), .B2(new_n218), .ZN(new_n890));
  OAI22_X1  g0690(.A1(new_n227), .A2(new_n890), .B1(G50), .B2(new_n218), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n891), .A2(G1), .A3(new_n247), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n885), .A2(new_n889), .A3(new_n892), .ZN(G367));
  AOI21_X1  g0693(.A(new_n544), .B1(new_n541), .B2(new_n620), .ZN(new_n894));
  XNOR2_X1  g0694(.A(new_n894), .B(KEYINPUT109), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(new_n629), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n620), .B1(new_n896), .B2(new_n543), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n543), .A2(new_n626), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n895), .A2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(new_n628), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n897), .B1(new_n901), .B2(KEYINPUT42), .ZN(new_n902));
  OR2_X1    g0702(.A1(new_n902), .A2(KEYINPUT110), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(KEYINPUT110), .ZN(new_n904));
  OAI211_X1 g0704(.A(new_n903), .B(new_n904), .C1(KEYINPUT42), .C2(new_n901), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n582), .A2(new_n584), .A3(new_n620), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n586), .A2(new_n579), .A3(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n907), .B1(new_n579), .B2(new_n906), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(KEYINPUT43), .ZN(new_n909));
  XNOR2_X1  g0709(.A(new_n908), .B(KEYINPUT108), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT43), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n905), .A2(new_n909), .A3(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n913), .B1(new_n905), .B2(new_n912), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n637), .A2(new_n899), .ZN(new_n915));
  INV_X1    g0715(.A(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  OAI211_X1 g0717(.A(new_n913), .B(new_n915), .C1(new_n905), .C2(new_n912), .ZN(new_n918));
  XNOR2_X1  g0718(.A(new_n640), .B(KEYINPUT41), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n630), .A2(new_n900), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n921), .B(KEYINPUT44), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n630), .A2(new_n900), .ZN(new_n923));
  XOR2_X1   g0723(.A(KEYINPUT111), .B(KEYINPUT45), .Z(new_n924));
  XNOR2_X1  g0724(.A(new_n923), .B(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n922), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(new_n636), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n922), .A2(new_n637), .A3(new_n925), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n624), .B(new_n627), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n929), .B(new_n635), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n930), .A2(new_n673), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n927), .A2(new_n928), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n920), .B1(new_n932), .B2(new_n674), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n745), .A2(G1), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n917), .B(new_n918), .C1(new_n933), .C2(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(new_n726), .ZN(new_n936));
  OAI22_X1  g0736(.A1(new_n936), .A2(new_n547), .B1(new_n420), .B2(new_n707), .ZN(new_n937));
  AOI21_X1  g0737(.A(KEYINPUT46), .B1(new_n716), .B2(G116), .ZN(new_n938));
  AND3_X1   g0738(.A1(new_n716), .A2(KEYINPUT46), .A3(G116), .ZN(new_n939));
  XNOR2_X1  g0739(.A(KEYINPUT112), .B(G311), .ZN(new_n940));
  AOI211_X1 g0740(.A(new_n938), .B(new_n939), .C1(new_n702), .C2(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n266), .B1(new_n713), .B2(new_n471), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n942), .B1(G283), .B2(new_n727), .ZN(new_n943));
  OAI211_X1 g0743(.A(new_n941), .B(new_n943), .C1(new_n685), .C2(new_n698), .ZN(new_n944));
  AOI211_X1 g0744(.A(new_n937), .B(new_n944), .C1(G294), .C2(new_n684), .ZN(new_n945));
  AOI22_X1  g0745(.A1(G159), .A2(new_n684), .B1(new_n727), .B2(G50), .ZN(new_n946));
  OR2_X1    g0746(.A1(new_n946), .A2(KEYINPUT113), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n699), .A2(G137), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n946), .A2(KEYINPUT113), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n947), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(new_n678), .ZN(new_n951));
  AOI22_X1  g0751(.A1(G143), .A2(new_n702), .B1(new_n951), .B2(G150), .ZN(new_n952));
  OAI221_X1 g0752(.A(new_n952), .B1(new_n776), .B2(new_n690), .C1(new_n300), .C2(new_n713), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n707), .A2(new_n218), .ZN(new_n954));
  NOR4_X1   g0754(.A1(new_n950), .A2(new_n953), .A3(new_n266), .A4(new_n954), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n945), .A2(new_n955), .ZN(new_n956));
  XOR2_X1   g0756(.A(new_n956), .B(KEYINPUT47), .Z(new_n957));
  AOI21_X1  g0757(.A(new_n746), .B1(new_n957), .B2(new_n733), .ZN(new_n958));
  INV_X1    g0758(.A(new_n738), .ZN(new_n959));
  OAI221_X1 g0759(.A(new_n737), .B1(new_n209), .B2(new_n298), .C1(new_n237), .C2(new_n959), .ZN(new_n960));
  OAI211_X1 g0760(.A(new_n958), .B(new_n960), .C1(new_n908), .C2(new_n748), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n935), .A2(new_n961), .ZN(G387));
  NOR2_X1   g0762(.A1(new_n707), .A2(new_n298), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n699), .A2(G150), .ZN(new_n965));
  OAI22_X1  g0765(.A1(new_n701), .A2(new_n720), .B1(new_n713), .B2(new_n471), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n274), .B1(new_n678), .B2(new_n202), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n690), .A2(new_n300), .ZN(new_n968));
  NOR3_X1   g0768(.A1(new_n966), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(new_n261), .ZN(new_n970));
  AOI22_X1  g0770(.A1(new_n970), .A2(new_n684), .B1(new_n727), .B2(G68), .ZN(new_n971));
  NAND4_X1  g0771(.A1(new_n964), .A2(new_n965), .A3(new_n969), .A4(new_n971), .ZN(new_n972));
  AOI22_X1  g0772(.A1(new_n702), .A2(G322), .B1(new_n727), .B2(G303), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n973), .B1(new_n936), .B2(new_n685), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n974), .B1(new_n684), .B2(new_n940), .ZN(new_n975));
  XOR2_X1   g0775(.A(new_n975), .B(KEYINPUT48), .Z(new_n976));
  OAI221_X1 g0776(.A(new_n976), .B1(new_n712), .B2(new_n707), .C1(new_n708), .C2(new_n690), .ZN(new_n977));
  XNOR2_X1  g0777(.A(KEYINPUT114), .B(KEYINPUT49), .ZN(new_n978));
  OR2_X1    g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n977), .A2(new_n978), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n274), .B1(new_n699), .B2(G326), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n979), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n713), .A2(new_n213), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n972), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n738), .B1(new_n233), .B2(new_n448), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n985), .B1(new_n642), .B2(new_n742), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n218), .A2(new_n300), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n970), .A2(new_n202), .ZN(new_n988));
  AOI211_X1 g0788(.A(G116), .B(new_n472), .C1(new_n988), .C2(KEYINPUT50), .ZN(new_n989));
  OAI211_X1 g0789(.A(new_n989), .B(new_n448), .C1(KEYINPUT50), .C2(new_n988), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n986), .B1(new_n987), .B2(new_n990), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n991), .B1(G107), .B2(new_n209), .ZN(new_n992));
  AOI22_X1  g0792(.A1(new_n984), .A2(new_n733), .B1(new_n737), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n624), .A2(new_n736), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n993), .A2(new_n747), .A3(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(new_n934), .ZN(new_n996));
  INV_X1    g0796(.A(new_n930), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n640), .B1(new_n997), .B2(new_n674), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n995), .B1(new_n996), .B2(new_n930), .C1(new_n998), .C2(new_n931), .ZN(G393));
  AOI22_X1  g0799(.A1(new_n241), .A2(new_n738), .B1(G97), .B2(new_n639), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n1000), .A2(new_n737), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n698), .A2(new_n679), .ZN(new_n1002));
  OAI22_X1  g0802(.A1(new_n683), .A2(new_n547), .B1(new_n692), .B2(new_n708), .ZN(new_n1003));
  NOR4_X1   g0803(.A1(new_n1002), .A2(new_n274), .A3(new_n715), .A4(new_n1003), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n1004), .B1(new_n213), .B2(new_n707), .C1(new_n712), .C2(new_n690), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n701), .A2(new_n685), .B1(new_n678), .B2(new_n691), .ZN(new_n1006));
  XOR2_X1   g0806(.A(new_n1006), .B(KEYINPUT52), .Z(new_n1007));
  OAI22_X1  g0807(.A1(new_n202), .A2(new_n683), .B1(new_n690), .B2(new_n218), .ZN(new_n1008));
  AOI211_X1 g0808(.A(new_n266), .B(new_n1008), .C1(G87), .C2(new_n780), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n724), .A2(G77), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n727), .A2(new_n970), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n699), .A2(G143), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n1009), .A2(new_n1010), .A3(new_n1011), .A4(new_n1012), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n701), .A2(new_n257), .B1(new_n678), .B2(new_n720), .ZN(new_n1014));
  XOR2_X1   g0814(.A(new_n1014), .B(KEYINPUT51), .Z(new_n1015));
  OAI22_X1  g0815(.A1(new_n1005), .A2(new_n1007), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n746), .B1(new_n1016), .B2(new_n733), .ZN(new_n1017));
  OAI211_X1 g0817(.A(new_n1001), .B(new_n1017), .C1(new_n900), .C2(new_n748), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n927), .A2(new_n928), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1018), .B1(new_n1019), .B2(new_n996), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n931), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n641), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1020), .B1(new_n932), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n1023), .ZN(G390));
  OAI21_X1  g0824(.A(new_n807), .B1(new_n871), .B2(new_n872), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1025), .A2(new_n865), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n863), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  AND2_X1   g0828(.A1(new_n759), .A2(G330), .ZN(new_n1029));
  AND2_X1   g0829(.A1(new_n664), .A2(new_n1029), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n671), .A2(new_n767), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n1031), .A2(new_n869), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n806), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n1033), .A2(new_n804), .ZN(new_n1034));
  OAI211_X1 g0834(.A(new_n865), .B(new_n835), .C1(new_n1032), .C2(new_n1034), .ZN(new_n1035));
  NAND4_X1  g0835(.A1(new_n1028), .A2(new_n807), .A3(new_n1030), .A4(new_n1035), .ZN(new_n1036));
  AND2_X1   g0836(.A1(new_n1028), .A2(new_n1035), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n809), .A2(new_n1029), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n1038), .A2(new_n1034), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1036), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n577), .A2(G330), .A3(new_n809), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n882), .A2(new_n612), .A3(new_n1041), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n1030), .A2(new_n807), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n1043), .A2(new_n1039), .B1(new_n872), .B2(new_n871), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1030), .A2(new_n807), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1038), .A2(new_n1034), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1045), .A2(new_n1032), .A3(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1042), .B1(new_n1044), .B2(new_n1047), .ZN(new_n1048));
  OR2_X1    g0848(.A1(new_n1040), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1040), .A2(new_n1048), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1049), .A2(new_n640), .A3(new_n1050), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n724), .A2(G159), .B1(G137), .B2(new_n684), .ZN(new_n1052));
  XOR2_X1   g0852(.A(KEYINPUT54), .B(G143), .Z(new_n1053));
  INV_X1    g0853(.A(new_n1053), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1052), .B1(new_n692), .B2(new_n1054), .ZN(new_n1055));
  XOR2_X1   g0855(.A(new_n1055), .B(KEYINPUT115), .Z(new_n1056));
  NOR2_X1   g0856(.A1(new_n690), .A2(new_n257), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1057), .B(KEYINPUT53), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n266), .B1(new_n951), .B2(G132), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n702), .A2(G128), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n1059), .B(new_n1060), .C1(new_n202), .C2(new_n713), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1061), .B1(G125), .B2(new_n699), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1056), .A2(new_n1058), .A3(new_n1062), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1063), .B(KEYINPUT116), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n683), .A2(new_n420), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n701), .A2(new_n712), .B1(new_n690), .B2(new_n470), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n274), .B(new_n1066), .C1(G116), .C2(new_n951), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n218), .A2(new_n713), .B1(new_n692), .B2(new_n471), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1068), .B1(new_n699), .B2(G294), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1067), .A2(new_n1069), .A3(new_n1010), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1064), .B1(new_n1065), .B2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n746), .B1(new_n1071), .B2(new_n733), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1072), .B1(new_n863), .B2(new_n735), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1073), .B1(new_n261), .B2(new_n793), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1074), .B1(new_n1040), .B2(new_n934), .ZN(new_n1075));
  AND2_X1   g0875(.A1(new_n1075), .A2(KEYINPUT117), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n1075), .A2(KEYINPUT117), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1051), .B1(new_n1076), .B2(new_n1077), .ZN(G378));
  INV_X1    g0878(.A(KEYINPUT120), .ZN(new_n1079));
  NAND4_X1  g0879(.A1(new_n836), .A2(new_n839), .A3(G330), .A4(new_n851), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1080), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1081), .B1(new_n876), .B2(new_n878), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n293), .B(KEYINPUT55), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n263), .A2(new_n618), .ZN(new_n1084));
  XNOR2_X1  g0884(.A(new_n1084), .B(KEYINPUT56), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1083), .B(new_n1085), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n867), .A2(new_n873), .A3(new_n875), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1087), .A2(KEYINPUT106), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n877), .A2(new_n856), .A3(new_n873), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1088), .A2(new_n1089), .A3(new_n1080), .ZN(new_n1090));
  AND3_X1   g0890(.A1(new_n1082), .A2(new_n1086), .A3(new_n1090), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1086), .B1(new_n1082), .B2(new_n1090), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1079), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1086), .ZN(new_n1094));
  AND3_X1   g0894(.A1(new_n1088), .A2(new_n1089), .A3(new_n1080), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1080), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1094), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1082), .A2(new_n1090), .A3(new_n1086), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1097), .A2(KEYINPUT120), .A3(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1093), .A2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1044), .A2(new_n1047), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1042), .B1(new_n1040), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(KEYINPUT57), .B1(new_n1100), .B2(new_n1103), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1103), .A2(new_n1105), .A3(KEYINPUT57), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1106), .A2(new_n640), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n1104), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1086), .A2(new_n734), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n793), .A2(new_n202), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n701), .A2(new_n213), .B1(new_n678), .B2(new_n420), .ZN(new_n1111));
  NOR4_X1   g0911(.A1(new_n954), .A2(G41), .A3(new_n968), .A4(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n274), .B1(new_n780), .B2(G58), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n699), .A2(G283), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n298), .A2(new_n692), .B1(new_n471), .B2(new_n683), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(new_n1115), .B(KEYINPUT118), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n1112), .A2(new_n1113), .A3(new_n1114), .A4(new_n1116), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n1117), .B(KEYINPUT58), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n202), .B1(new_n264), .B2(G41), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n724), .A2(G150), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n727), .A2(G137), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(G125), .A2(new_n702), .B1(new_n951), .B2(G128), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(G132), .A2(new_n684), .B1(new_n716), .B2(new_n1053), .ZN(new_n1123));
  NAND4_X1  g0923(.A1(new_n1120), .A2(new_n1121), .A3(new_n1122), .A4(new_n1123), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n1125));
  OR2_X1    g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1127));
  AOI21_X1  g0927(.A(G33), .B1(new_n780), .B2(G159), .ZN(new_n1128));
  AOI21_X1  g0928(.A(G41), .B1(new_n699), .B2(G124), .ZN(new_n1129));
  NAND4_X1  g0929(.A1(new_n1126), .A2(new_n1127), .A3(new_n1128), .A4(new_n1129), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1118), .A2(new_n1119), .A3(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n746), .B1(new_n1131), .B2(new_n733), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1109), .A2(new_n1110), .A3(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1134), .B1(new_n1100), .B2(new_n934), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n1108), .A2(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(G375));
  AOI21_X1  g0938(.A(new_n996), .B1(new_n1044), .B2(new_n1047), .ZN(new_n1139));
  OR2_X1    g0939(.A1(new_n1139), .A2(KEYINPUT121), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n684), .A2(new_n1053), .B1(new_n727), .B2(G150), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n702), .A2(G132), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n1141), .B(new_n1142), .C1(new_n720), .C2(new_n690), .ZN(new_n1143));
  AOI211_X1 g0943(.A(new_n266), .B(new_n1143), .C1(G128), .C2(new_n699), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n724), .A2(G50), .B1(G137), .B2(new_n726), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n1144), .B(new_n1145), .C1(new_n776), .C2(new_n713), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n963), .B1(G283), .B2(new_n951), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1147), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n1148), .A2(KEYINPUT124), .ZN(new_n1149));
  AOI211_X1 g0949(.A(new_n274), .B(new_n1149), .C1(G97), .C2(new_n716), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(new_n699), .A2(G303), .B1(G77), .B2(new_n780), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1148), .A2(KEYINPUT124), .ZN(new_n1152));
  OAI22_X1  g0952(.A1(new_n683), .A2(new_n213), .B1(new_n692), .B2(new_n420), .ZN(new_n1153));
  OR2_X1    g0953(.A1(new_n1153), .A2(KEYINPUT122), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1153), .A2(KEYINPUT122), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n1154), .B(new_n1155), .C1(new_n708), .C2(new_n701), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT123), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  NAND4_X1  g0958(.A1(new_n1150), .A2(new_n1151), .A3(new_n1152), .A4(new_n1158), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1146), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n1161), .A2(new_n733), .B1(new_n218), .B2(new_n793), .ZN(new_n1162));
  OAI211_X1 g0962(.A(new_n747), .B(new_n1162), .C1(new_n807), .C2(new_n735), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1139), .A2(KEYINPUT121), .ZN(new_n1164));
  AND3_X1   g0964(.A1(new_n1140), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1042), .A2(new_n1044), .A3(new_n1047), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1166), .A2(new_n919), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1165), .B1(new_n1048), .B2(new_n1167), .ZN(G381));
  AND2_X1   g0968(.A1(new_n1051), .A2(new_n1075), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(G381), .A2(G384), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1137), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n935), .A2(new_n961), .A3(new_n1023), .ZN(new_n1172));
  OR4_X1    g0972(.A1(G396), .A2(new_n1171), .A3(G393), .A4(new_n1172), .ZN(G407));
  NAND3_X1  g0973(.A1(new_n1137), .A2(new_n619), .A3(new_n1169), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(G407), .A2(G213), .A3(new_n1174), .ZN(G409));
  XNOR2_X1  g0975(.A(G393), .B(G396), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT126), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1172), .A2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1023), .B1(new_n935), .B2(new_n961), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1177), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1180), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1182), .A2(new_n1178), .A3(new_n1172), .A4(new_n1176), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1181), .A2(new_n1183), .ZN(new_n1184));
  OAI211_X1 g0984(.A(G378), .B(new_n1135), .C1(new_n1104), .C2(new_n1107), .ZN(new_n1185));
  AOI211_X1 g0985(.A(new_n920), .B(new_n1102), .C1(new_n1093), .C2(new_n1099), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1105), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1133), .B1(new_n1187), .B2(new_n996), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1169), .B1(new_n1186), .B2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1185), .A2(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(G213), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n1191), .A2(G343), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1190), .A2(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT60), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1166), .B1(new_n1048), .B2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT125), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  OR2_X1    g0998(.A1(new_n1166), .A2(new_n1195), .ZN(new_n1199));
  OAI211_X1 g0999(.A(KEYINPUT125), .B(new_n1166), .C1(new_n1048), .C2(new_n1195), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n1198), .A2(new_n640), .A3(new_n1199), .A4(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1201), .A2(new_n1165), .ZN(new_n1202));
  INV_X1    g1002(.A(G384), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1201), .A2(G384), .A3(new_n1165), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1206), .A2(G2897), .A3(new_n1192), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1192), .A2(G2897), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1204), .A2(new_n1205), .A3(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1207), .A2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1194), .A2(new_n1211), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1190), .A2(new_n1204), .A3(new_n1205), .A4(new_n1193), .ZN(new_n1213));
  AOI21_X1  g1013(.A(KEYINPUT62), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT61), .ZN(new_n1215));
  AOI211_X1 g1015(.A(new_n1192), .B(new_n1206), .C1(new_n1185), .C2(new_n1189), .ZN(new_n1216));
  INV_X1    g1016(.A(KEYINPUT62), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1215), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1184), .B1(new_n1214), .B2(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1210), .B1(new_n1193), .B2(new_n1190), .ZN(new_n1220));
  OAI21_X1  g1020(.A(KEYINPUT63), .B1(new_n1220), .B2(new_n1216), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT63), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1184), .B1(new_n1213), .B2(new_n1222), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1221), .A2(new_n1223), .A3(new_n1215), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1219), .A2(new_n1224), .ZN(G405));
  NAND2_X1  g1025(.A1(G375), .A2(new_n1169), .ZN(new_n1226));
  OAI211_X1 g1026(.A(new_n1226), .B(new_n1185), .C1(KEYINPUT127), .C2(new_n1206), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1206), .A2(KEYINPUT127), .ZN(new_n1228));
  XNOR2_X1  g1028(.A(new_n1184), .B(new_n1228), .ZN(new_n1229));
  XNOR2_X1  g1029(.A(new_n1227), .B(new_n1229), .ZN(G402));
endmodule


