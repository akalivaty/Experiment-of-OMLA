//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 1 0 1 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 0 0 1 1 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 0 0 1 1 0 0 1 1 1 0 0 0 0 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:49 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n579, new_n580, new_n581, new_n582,
    new_n583, new_n584, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n603, new_n604, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n615, new_n616, new_n617, new_n619, new_n620, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n631,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n648, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n798, new_n799, new_n800,
    new_n801, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n837, new_n838,
    new_n839, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT31), .ZN(new_n189));
  INV_X1    g003(.A(G119), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G116), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT68), .B(G116), .ZN(new_n192));
  OAI21_X1  g006(.A(new_n191), .B1(new_n192), .B2(new_n190), .ZN(new_n193));
  XNOR2_X1  g007(.A(KEYINPUT2), .B(G113), .ZN(new_n194));
  XOR2_X1   g008(.A(new_n193), .B(new_n194), .Z(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G143), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n197), .A2(G146), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(KEYINPUT65), .ZN(new_n199));
  INV_X1    g013(.A(G146), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G143), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT65), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  AOI22_X1  g017(.A1(new_n199), .A2(new_n203), .B1(new_n197), .B2(G146), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT1), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n204), .A2(new_n205), .A3(G128), .ZN(new_n206));
  INV_X1    g020(.A(G128), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n207), .B1(new_n201), .B2(KEYINPUT1), .ZN(new_n208));
  INV_X1    g022(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n197), .A2(G146), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n201), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n206), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G134), .ZN(new_n214));
  OAI21_X1  g028(.A(KEYINPUT66), .B1(new_n214), .B2(G137), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(KEYINPUT11), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n214), .A2(G137), .ZN(new_n217));
  INV_X1    g031(.A(G137), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G134), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT11), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n219), .A2(KEYINPUT66), .A3(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n216), .A2(new_n217), .A3(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(G131), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  AND3_X1   g038(.A1(new_n217), .A2(new_n219), .A3(G131), .ZN(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  AOI21_X1  g040(.A(KEYINPUT69), .B1(new_n224), .B2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT69), .ZN(new_n228));
  AOI211_X1 g042(.A(new_n228), .B(new_n225), .C1(new_n222), .C2(new_n223), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n213), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT70), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n204), .A2(KEYINPUT0), .A3(G128), .ZN(new_n233));
  NAND2_X1  g047(.A1(KEYINPUT0), .A2(G128), .ZN(new_n234));
  OR2_X1    g048(.A1(KEYINPUT0), .A2(G128), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n211), .A2(KEYINPUT64), .A3(new_n234), .A4(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n211), .A2(new_n234), .A3(new_n235), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT64), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  AND3_X1   g053(.A1(new_n233), .A2(new_n236), .A3(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(KEYINPUT67), .A2(G131), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  XNOR2_X1  g056(.A(new_n222), .B(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n240), .A2(new_n243), .ZN(new_n244));
  OAI211_X1 g058(.A(KEYINPUT70), .B(new_n213), .C1(new_n227), .C2(new_n229), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n232), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(KEYINPUT30), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT30), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n224), .A2(new_n226), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n213), .A2(new_n249), .ZN(new_n250));
  AND3_X1   g064(.A1(new_n244), .A2(new_n248), .A3(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n247), .A2(new_n252), .ZN(new_n253));
  AND2_X1   g067(.A1(new_n232), .A2(new_n245), .ZN(new_n254));
  NAND4_X1  g068(.A1(new_n254), .A2(KEYINPUT71), .A3(new_n195), .A4(new_n244), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n232), .A2(new_n195), .A3(new_n244), .A4(new_n245), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT71), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  AOI22_X1  g072(.A1(new_n196), .A2(new_n253), .B1(new_n255), .B2(new_n258), .ZN(new_n259));
  XNOR2_X1  g073(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n260));
  XNOR2_X1  g074(.A(new_n260), .B(G101), .ZN(new_n261));
  INV_X1    g075(.A(G237), .ZN(new_n262));
  INV_X1    g076(.A(G953), .ZN(new_n263));
  AND3_X1   g077(.A1(new_n262), .A2(new_n263), .A3(G210), .ZN(new_n264));
  XOR2_X1   g078(.A(new_n261), .B(new_n264), .Z(new_n265));
  AOI21_X1  g079(.A(new_n189), .B1(new_n259), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n253), .A2(new_n196), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n255), .A2(new_n258), .ZN(new_n268));
  NAND4_X1  g082(.A1(new_n267), .A2(new_n268), .A3(new_n189), .A4(new_n265), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  OAI21_X1  g084(.A(KEYINPUT72), .B1(new_n266), .B2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT72), .ZN(new_n272));
  AND2_X1   g086(.A1(new_n256), .A2(new_n257), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n256), .A2(new_n257), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n251), .B1(new_n246), .B2(KEYINPUT30), .ZN(new_n275));
  OAI22_X1  g089(.A1(new_n273), .A2(new_n274), .B1(new_n275), .B2(new_n195), .ZN(new_n276));
  INV_X1    g090(.A(new_n265), .ZN(new_n277));
  OAI21_X1  g091(.A(KEYINPUT31), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n244), .A2(new_n230), .A3(new_n195), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT28), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n195), .B1(new_n244), .B2(new_n250), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n282), .B1(new_n255), .B2(new_n258), .ZN(new_n283));
  XOR2_X1   g097(.A(KEYINPUT73), .B(KEYINPUT28), .Z(new_n284));
  OAI21_X1  g098(.A(new_n281), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  AOI22_X1  g099(.A1(new_n272), .A2(new_n278), .B1(new_n285), .B2(new_n277), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n188), .B1(new_n271), .B2(new_n286), .ZN(new_n287));
  XOR2_X1   g101(.A(KEYINPUT74), .B(KEYINPUT32), .Z(new_n288));
  OAI21_X1  g102(.A(KEYINPUT75), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n287), .A2(KEYINPUT32), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n278), .A2(new_n272), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n285), .A2(new_n277), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n272), .B1(new_n278), .B2(new_n269), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n187), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT75), .ZN(new_n296));
  INV_X1    g110(.A(new_n288), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n295), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n281), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n246), .A2(new_n196), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT76), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n246), .A2(KEYINPUT76), .A3(new_n196), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n268), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n299), .B1(new_n304), .B2(KEYINPUT28), .ZN(new_n305));
  NAND4_X1  g119(.A1(new_n305), .A2(KEYINPUT77), .A3(KEYINPUT29), .A4(new_n265), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n302), .A2(new_n303), .ZN(new_n307));
  XNOR2_X1  g121(.A(new_n256), .B(KEYINPUT71), .ZN(new_n308));
  OAI21_X1  g122(.A(KEYINPUT28), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND4_X1  g123(.A1(new_n309), .A2(KEYINPUT29), .A3(new_n265), .A4(new_n281), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT77), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  OAI211_X1 g126(.A(new_n265), .B(new_n281), .C1(new_n283), .C2(new_n284), .ZN(new_n313));
  AOI21_X1  g127(.A(KEYINPUT29), .B1(new_n276), .B2(new_n277), .ZN(new_n314));
  AOI21_X1  g128(.A(G902), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n306), .A2(new_n312), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(G472), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n289), .A2(new_n290), .A3(new_n298), .A4(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(G125), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n319), .A2(G140), .ZN(new_n320));
  XNOR2_X1  g134(.A(G125), .B(G140), .ZN(new_n321));
  MUX2_X1   g135(.A(new_n320), .B(new_n321), .S(KEYINPUT16), .Z(new_n322));
  XNOR2_X1  g136(.A(new_n322), .B(G146), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n190), .A2(G128), .ZN(new_n325));
  XNOR2_X1  g139(.A(new_n325), .B(KEYINPUT78), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n326), .B1(G119), .B2(new_n207), .ZN(new_n327));
  XOR2_X1   g141(.A(KEYINPUT24), .B(G110), .Z(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n207), .A2(G119), .ZN(new_n330));
  XNOR2_X1  g144(.A(new_n330), .B(KEYINPUT23), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(new_n325), .ZN(new_n332));
  XOR2_X1   g146(.A(new_n332), .B(KEYINPUT79), .Z(new_n333));
  INV_X1    g147(.A(G110), .ZN(new_n334));
  OAI211_X1 g148(.A(new_n324), .B(new_n329), .C1(new_n333), .C2(new_n334), .ZN(new_n335));
  OR2_X1    g149(.A1(new_n322), .A2(new_n200), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n321), .A2(new_n200), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n327), .A2(new_n328), .ZN(new_n338));
  NOR2_X1   g152(.A1(KEYINPUT80), .A2(G110), .ZN(new_n339));
  AND2_X1   g153(.A1(KEYINPUT80), .A2(G110), .ZN(new_n340));
  NOR3_X1   g154(.A1(new_n332), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  OAI211_X1 g155(.A(new_n336), .B(new_n337), .C1(new_n338), .C2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n335), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n263), .A2(G221), .A3(G234), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n344), .B(KEYINPUT22), .ZN(new_n345));
  XNOR2_X1  g159(.A(new_n345), .B(new_n218), .ZN(new_n346));
  OR2_X1    g160(.A1(new_n343), .A2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(G902), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n343), .A2(new_n346), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n347), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(G217), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n351), .B1(G234), .B2(new_n348), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT25), .ZN(new_n354));
  XNOR2_X1  g168(.A(new_n350), .B(new_n354), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n353), .B1(new_n355), .B2(new_n352), .ZN(new_n356));
  OAI21_X1  g170(.A(G214), .B1(G237), .B2(G902), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(G104), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n359), .A2(G107), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT84), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT3), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n360), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(G107), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n361), .A2(new_n364), .A3(G104), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(KEYINPUT3), .ZN(new_n366));
  OAI211_X1 g180(.A(new_n363), .B(new_n366), .C1(G104), .C2(new_n364), .ZN(new_n367));
  AND2_X1   g181(.A1(KEYINPUT85), .A2(G101), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT4), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  OR2_X1    g185(.A1(new_n367), .A2(G101), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n367), .A2(KEYINPUT4), .A3(new_n368), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n196), .A2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT87), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n364), .A2(G104), .ZN(new_n378));
  OAI21_X1  g192(.A(G101), .B1(new_n378), .B2(new_n360), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n372), .A2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT5), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n381), .A2(new_n190), .A3(G116), .ZN(new_n382));
  OAI211_X1 g196(.A(G113), .B(new_n382), .C1(new_n193), .C2(new_n381), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n383), .B1(new_n194), .B2(new_n193), .ZN(new_n384));
  OR2_X1    g198(.A1(new_n380), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n196), .A2(new_n374), .A3(KEYINPUT87), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n377), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  XOR2_X1   g201(.A(G110), .B(G122), .Z(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(new_n388), .ZN(new_n390));
  NAND4_X1  g204(.A1(new_n377), .A2(new_n390), .A3(new_n385), .A4(new_n386), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n389), .A2(KEYINPUT6), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n240), .A2(G125), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n213), .A2(new_n319), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(G224), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n396), .A2(G953), .ZN(new_n397));
  OR2_X1    g211(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n395), .A2(new_n397), .ZN(new_n399));
  AND2_X1   g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT6), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n387), .A2(new_n401), .A3(new_n388), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n392), .A2(new_n400), .A3(new_n402), .ZN(new_n403));
  OAI211_X1 g217(.A(new_n398), .B(new_n399), .C1(KEYINPUT7), .C2(new_n397), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n380), .B(new_n384), .ZN(new_n405));
  XOR2_X1   g219(.A(new_n388), .B(KEYINPUT8), .Z(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  OR3_X1    g221(.A1(new_n395), .A2(KEYINPUT7), .A3(new_n397), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n404), .A2(new_n391), .A3(new_n407), .A4(new_n408), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n403), .A2(new_n348), .A3(new_n409), .ZN(new_n410));
  OAI21_X1  g224(.A(G210), .B1(G237), .B2(G902), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  NAND4_X1  g227(.A1(new_n403), .A2(new_n348), .A3(new_n411), .A4(new_n409), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n358), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  XNOR2_X1  g229(.A(KEYINPUT9), .B(G234), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n416), .B(KEYINPUT81), .ZN(new_n417));
  OAI21_X1  g231(.A(G221), .B1(new_n417), .B2(G902), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n418), .B(KEYINPUT82), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  AND2_X1   g234(.A1(new_n372), .A2(new_n379), .ZN(new_n421));
  OR3_X1    g235(.A1(new_n204), .A2(KEYINPUT86), .A3(new_n208), .ZN(new_n422));
  OAI21_X1  g236(.A(KEYINPUT86), .B1(new_n204), .B2(new_n208), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n422), .A2(new_n206), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n421), .A2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT10), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n243), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n374), .A2(new_n240), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n421), .A2(KEYINPUT10), .A3(new_n213), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n427), .A2(new_n428), .A3(new_n429), .A4(new_n430), .ZN(new_n431));
  XNOR2_X1  g245(.A(G110), .B(G140), .ZN(new_n432));
  AND2_X1   g246(.A1(new_n263), .A2(G227), .ZN(new_n433));
  XOR2_X1   g247(.A(new_n432), .B(new_n433), .Z(new_n434));
  AND2_X1   g248(.A1(new_n431), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n380), .A2(new_n212), .A3(new_n206), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n425), .A2(new_n436), .ZN(new_n437));
  AND3_X1   g251(.A1(new_n437), .A2(KEYINPUT12), .A3(new_n243), .ZN(new_n438));
  AOI21_X1  g252(.A(KEYINPUT12), .B1(new_n437), .B2(new_n243), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n435), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n427), .A2(new_n429), .A3(new_n430), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(new_n243), .ZN(new_n442));
  AND2_X1   g256(.A1(new_n442), .A2(new_n431), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n440), .B1(new_n443), .B2(new_n434), .ZN(new_n444));
  INV_X1    g258(.A(G469), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n444), .A2(new_n445), .A3(new_n348), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n431), .B1(new_n438), .B2(new_n439), .ZN(new_n447));
  XOR2_X1   g261(.A(new_n434), .B(KEYINPUT83), .Z(new_n448));
  AOI22_X1  g262(.A1(new_n447), .A2(new_n448), .B1(new_n435), .B2(new_n442), .ZN(new_n449));
  OAI21_X1  g263(.A(G469), .B1(new_n449), .B2(G902), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n420), .B1(new_n446), .B2(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n262), .A2(new_n263), .A3(G214), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n452), .B(new_n197), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n453), .A2(KEYINPUT17), .A3(G131), .ZN(new_n454));
  OAI21_X1  g268(.A(KEYINPUT88), .B1(new_n453), .B2(G131), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n453), .A2(G131), .ZN(new_n456));
  XNOR2_X1  g270(.A(new_n452), .B(G143), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT88), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n457), .A2(new_n458), .A3(new_n223), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n455), .A2(new_n456), .A3(new_n459), .ZN(new_n460));
  OAI211_X1 g274(.A(new_n323), .B(new_n454), .C1(new_n460), .C2(KEYINPUT17), .ZN(new_n461));
  XNOR2_X1  g275(.A(G113), .B(G122), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n462), .B(new_n359), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT18), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n457), .B1(new_n464), .B2(new_n223), .ZN(new_n465));
  XNOR2_X1  g279(.A(new_n321), .B(new_n200), .ZN(new_n466));
  OAI211_X1 g280(.A(new_n465), .B(new_n466), .C1(new_n464), .C2(new_n456), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n461), .A2(new_n463), .A3(new_n467), .ZN(new_n468));
  XOR2_X1   g282(.A(new_n321), .B(KEYINPUT19), .Z(new_n469));
  OAI211_X1 g283(.A(new_n460), .B(new_n336), .C1(G146), .C2(new_n469), .ZN(new_n470));
  AND2_X1   g284(.A1(new_n470), .A2(new_n467), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n468), .B1(new_n471), .B2(new_n463), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT20), .ZN(new_n473));
  INV_X1    g287(.A(G475), .ZN(new_n474));
  NAND4_X1  g288(.A1(new_n472), .A2(new_n473), .A3(new_n474), .A4(new_n348), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT89), .ZN(new_n476));
  OR2_X1    g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(new_n468), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n463), .B1(new_n470), .B2(new_n467), .ZN(new_n479));
  OAI211_X1 g293(.A(new_n474), .B(new_n348), .C1(new_n478), .C2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(KEYINPUT20), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n481), .A2(new_n475), .A3(new_n476), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n463), .B1(new_n461), .B2(new_n467), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n348), .B1(new_n478), .B2(new_n483), .ZN(new_n484));
  XNOR2_X1  g298(.A(KEYINPUT90), .B(G475), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n477), .A2(new_n482), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(G234), .A2(G237), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n488), .A2(G952), .A3(new_n263), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  XOR2_X1   g304(.A(KEYINPUT21), .B(G898), .Z(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n488), .A2(G902), .A3(G953), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n490), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n197), .A2(G128), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT13), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n197), .A2(G128), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  OAI211_X1 g313(.A(new_n499), .B(KEYINPUT91), .C1(new_n497), .C2(new_n498), .ZN(new_n500));
  OAI211_X1 g314(.A(new_n500), .B(G134), .C1(KEYINPUT91), .C2(new_n499), .ZN(new_n501));
  INV_X1    g315(.A(new_n498), .ZN(new_n502));
  OR3_X1    g316(.A1(new_n502), .A2(G134), .A3(new_n496), .ZN(new_n503));
  INV_X1    g317(.A(G116), .ZN(new_n504));
  MUX2_X1   g318(.A(new_n504), .B(new_n192), .S(G122), .Z(new_n505));
  AND2_X1   g319(.A1(new_n505), .A2(new_n364), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n505), .A2(new_n364), .ZN(new_n507));
  OAI211_X1 g321(.A(new_n501), .B(new_n503), .C1(new_n506), .C2(new_n507), .ZN(new_n508));
  OAI21_X1  g322(.A(G134), .B1(new_n502), .B2(new_n496), .ZN(new_n509));
  AOI22_X1  g323(.A1(new_n505), .A2(new_n364), .B1(new_n503), .B2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT92), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT14), .ZN(new_n512));
  INV_X1    g326(.A(G122), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(G116), .ZN(new_n514));
  OAI211_X1 g328(.A(new_n512), .B(new_n514), .C1(new_n192), .C2(new_n513), .ZN(new_n515));
  OR2_X1    g329(.A1(new_n192), .A2(new_n513), .ZN(new_n516));
  OAI211_X1 g330(.A(G107), .B(new_n515), .C1(new_n516), .C2(new_n512), .ZN(new_n517));
  AND3_X1   g331(.A1(new_n510), .A2(new_n511), .A3(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n511), .B1(new_n510), .B2(new_n517), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n508), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NOR3_X1   g334(.A1(new_n417), .A2(new_n351), .A3(G953), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n508), .B(new_n521), .C1(new_n518), .C2(new_n519), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(new_n348), .ZN(new_n526));
  INV_X1    g340(.A(G478), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n527), .A2(KEYINPUT15), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n526), .B(new_n528), .ZN(new_n529));
  NOR3_X1   g343(.A1(new_n487), .A2(new_n495), .A3(new_n529), .ZN(new_n530));
  AND3_X1   g344(.A1(new_n415), .A2(new_n451), .A3(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n318), .A2(new_n356), .A3(new_n531), .ZN(new_n532));
  XNOR2_X1  g346(.A(KEYINPUT93), .B(G101), .ZN(new_n533));
  XNOR2_X1  g347(.A(new_n532), .B(new_n533), .ZN(G3));
  OAI21_X1  g348(.A(new_n348), .B1(new_n293), .B2(new_n294), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(G472), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT94), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n287), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n446), .A2(new_n450), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(new_n419), .ZN(new_n540));
  INV_X1    g354(.A(new_n356), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n535), .A2(KEYINPUT94), .A3(G472), .ZN(new_n543));
  INV_X1    g357(.A(new_n495), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n415), .A2(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(KEYINPUT95), .B1(new_n523), .B2(new_n524), .ZN(new_n546));
  XNOR2_X1  g360(.A(new_n546), .B(KEYINPUT33), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n547), .A2(G478), .A3(new_n348), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n526), .A2(new_n527), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(new_n487), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n545), .A2(new_n551), .ZN(new_n552));
  NAND4_X1  g366(.A1(new_n538), .A2(new_n542), .A3(new_n543), .A4(new_n552), .ZN(new_n553));
  XOR2_X1   g367(.A(KEYINPUT34), .B(G104), .Z(new_n554));
  XNOR2_X1  g368(.A(new_n553), .B(new_n554), .ZN(G6));
  AOI21_X1  g369(.A(G902), .B1(new_n271), .B2(new_n286), .ZN(new_n556));
  INV_X1    g370(.A(G472), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n537), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND4_X1  g372(.A1(new_n558), .A2(new_n542), .A3(new_n543), .A4(new_n295), .ZN(new_n559));
  AOI22_X1  g373(.A1(new_n481), .A2(new_n475), .B1(new_n484), .B2(new_n485), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(new_n529), .ZN(new_n561));
  NOR3_X1   g375(.A1(new_n559), .A2(new_n545), .A3(new_n561), .ZN(new_n562));
  XNOR2_X1  g376(.A(KEYINPUT35), .B(G107), .ZN(new_n563));
  XNOR2_X1  g377(.A(new_n563), .B(KEYINPUT96), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n562), .B(new_n564), .ZN(G9));
  NAND4_X1  g379(.A1(new_n558), .A2(new_n531), .A3(new_n543), .A4(new_n295), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n355), .A2(new_n352), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n346), .A2(KEYINPUT36), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n343), .B(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  NOR3_X1   g384(.A1(new_n570), .A2(G902), .A3(new_n352), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n567), .A2(new_n572), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n573), .B(KEYINPUT97), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  OR2_X1    g389(.A1(new_n566), .A2(new_n575), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n576), .B(KEYINPUT37), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n577), .B(new_n334), .ZN(G12));
  INV_X1    g392(.A(new_n415), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n579), .A2(new_n540), .ZN(new_n580));
  INV_X1    g394(.A(G900), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n490), .B1(new_n494), .B2(new_n581), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n561), .A2(new_n582), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n318), .A2(new_n580), .A3(new_n574), .A4(new_n583), .ZN(new_n584));
  XNOR2_X1  g398(.A(new_n584), .B(G128), .ZN(G30));
  OAI21_X1  g399(.A(new_n348), .B1(new_n304), .B2(new_n265), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n259), .A2(new_n277), .ZN(new_n587));
  OAI21_X1  g401(.A(G472), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n289), .A2(new_n290), .A3(new_n298), .A4(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n573), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n487), .A2(new_n529), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n591), .A2(new_n358), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n413), .A2(new_n414), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n593), .B(KEYINPUT38), .ZN(new_n594));
  NAND4_X1  g408(.A1(new_n589), .A2(new_n590), .A3(new_n592), .A4(new_n594), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n595), .B(KEYINPUT98), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n582), .B(KEYINPUT39), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n540), .A2(new_n597), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n598), .B(KEYINPUT99), .ZN(new_n599));
  XOR2_X1   g413(.A(new_n599), .B(KEYINPUT40), .Z(new_n600));
  NAND2_X1  g414(.A1(new_n596), .A2(new_n600), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n601), .B(G143), .ZN(G45));
  NOR2_X1   g416(.A1(new_n551), .A2(new_n582), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n318), .A2(new_n580), .A3(new_n574), .A4(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n604), .B(G146), .ZN(G48));
  NAND2_X1  g419(.A1(new_n444), .A2(new_n348), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n606), .A2(G469), .ZN(new_n607));
  AND2_X1   g421(.A1(new_n607), .A2(new_n446), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(new_n418), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n318), .A2(new_n552), .A3(new_n356), .A4(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(KEYINPUT41), .B(G113), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n612), .B(KEYINPUT100), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n611), .B(new_n613), .ZN(G15));
  AND2_X1   g428(.A1(new_n318), .A2(new_n356), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n545), .A2(new_n561), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n615), .A2(new_n616), .A3(new_n610), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n617), .B(G116), .ZN(G18));
  NOR2_X1   g432(.A1(new_n609), .A2(new_n579), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n318), .A2(new_n530), .A3(new_n574), .A4(new_n619), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n620), .B(G119), .ZN(G21));
  INV_X1    g435(.A(KEYINPUT101), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n591), .B(new_n622), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n623), .A2(new_n545), .ZN(new_n624));
  OR2_X1    g438(.A1(new_n305), .A2(new_n265), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n266), .A2(new_n270), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n188), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n627), .B1(G472), .B2(new_n535), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n624), .A2(new_n628), .A3(new_n356), .A4(new_n610), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(G122), .ZN(G24));
  NAND4_X1  g444(.A1(new_n619), .A2(new_n628), .A3(new_n573), .A4(new_n603), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n631), .B(G125), .ZN(G27));
  INV_X1    g446(.A(KEYINPUT32), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n295), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n290), .A2(new_n317), .A3(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(new_n356), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n539), .A2(new_n418), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n593), .A2(new_n358), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n638), .A2(new_n603), .A3(new_n639), .ZN(new_n640));
  OAI21_X1  g454(.A(KEYINPUT42), .B1(new_n636), .B2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n603), .ZN(new_n642));
  INV_X1    g456(.A(new_n639), .ZN(new_n643));
  NOR3_X1   g457(.A1(new_n642), .A2(new_n643), .A3(KEYINPUT42), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n644), .A2(new_n318), .A3(new_n356), .A4(new_n638), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n641), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(new_n223), .ZN(G33));
  NAND4_X1  g461(.A1(new_n615), .A2(new_n583), .A3(new_n638), .A4(new_n639), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(G134), .ZN(G36));
  AOI21_X1  g463(.A(new_n487), .B1(new_n549), .B2(new_n548), .ZN(new_n650));
  XOR2_X1   g464(.A(new_n650), .B(KEYINPUT43), .Z(new_n651));
  AOI21_X1  g465(.A(new_n651), .B1(new_n538), .B2(new_n543), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(new_n573), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(KEYINPUT44), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(new_n639), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(KEYINPUT103), .ZN(new_n656));
  XOR2_X1   g470(.A(new_n449), .B(KEYINPUT45), .Z(new_n657));
  OAI21_X1  g471(.A(G469), .B1(new_n657), .B2(G902), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(KEYINPUT46), .ZN(new_n659));
  XOR2_X1   g473(.A(new_n659), .B(KEYINPUT102), .Z(new_n660));
  OAI211_X1 g474(.A(new_n660), .B(new_n446), .C1(KEYINPUT46), .C2(new_n658), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(new_n418), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n662), .A2(new_n597), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n656), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(G137), .ZN(G39));
  XOR2_X1   g479(.A(KEYINPUT104), .B(KEYINPUT47), .Z(new_n666));
  NAND3_X1  g480(.A1(new_n661), .A2(new_n418), .A3(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT104), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n669), .A2(KEYINPUT47), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n670), .B1(new_n661), .B2(new_n418), .ZN(new_n671));
  OR2_X1    g485(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  NOR4_X1   g486(.A1(new_n318), .A2(new_n356), .A3(new_n642), .A4(new_n643), .ZN(new_n673));
  XOR2_X1   g487(.A(new_n673), .B(KEYINPUT105), .Z(new_n674));
  NOR2_X1   g488(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  XOR2_X1   g489(.A(new_n675), .B(G140), .Z(G42));
  INV_X1    g490(.A(KEYINPUT115), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n589), .A2(new_n541), .ZN(new_n678));
  INV_X1    g492(.A(new_n608), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n419), .B1(new_n679), .B2(KEYINPUT49), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n680), .B1(KEYINPUT49), .B2(new_n679), .ZN(new_n681));
  INV_X1    g495(.A(new_n594), .ZN(new_n682));
  AND2_X1   g496(.A1(new_n682), .A2(new_n650), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n678), .A2(new_n681), .A3(new_n357), .A4(new_n683), .ZN(new_n684));
  XOR2_X1   g498(.A(new_n684), .B(KEYINPUT106), .Z(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(new_n487), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(new_n529), .ZN(new_n688));
  OR2_X1    g502(.A1(new_n545), .A2(new_n688), .ZN(new_n689));
  OAI22_X1  g503(.A1(new_n575), .A2(new_n566), .B1(new_n559), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(KEYINPUT107), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n617), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n611), .B1(new_n690), .B2(KEYINPUT107), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n620), .A2(new_n532), .A3(new_n553), .A4(new_n629), .ZN(new_n694));
  NOR3_X1   g508(.A1(new_n692), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  AND2_X1   g509(.A1(new_n584), .A2(new_n631), .ZN(new_n696));
  NOR3_X1   g510(.A1(new_n623), .A2(new_n579), .A3(new_n582), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n589), .A2(new_n697), .A3(new_n590), .A4(new_n638), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n696), .A2(KEYINPUT52), .A3(new_n604), .A4(new_n698), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n584), .A2(new_n604), .A3(new_n698), .A4(new_n631), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT52), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(new_n646), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n695), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  NOR3_X1   g519(.A1(new_n540), .A2(new_n529), .A3(new_n582), .ZN(new_n706));
  AND4_X1   g520(.A1(new_n318), .A2(new_n560), .A3(new_n574), .A4(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n628), .A2(new_n573), .ZN(new_n708));
  NOR3_X1   g522(.A1(new_n708), .A2(new_n642), .A3(new_n637), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n639), .B1(new_n707), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(new_n648), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT108), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n710), .A2(KEYINPUT108), .A3(new_n648), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  OAI21_X1  g529(.A(KEYINPUT53), .B1(new_n705), .B2(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(new_n714), .ZN(new_n717));
  AOI21_X1  g531(.A(KEYINPUT108), .B1(new_n710), .B2(new_n648), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NOR4_X1   g533(.A1(new_n692), .A2(new_n693), .A3(new_n646), .A4(new_n694), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT53), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n719), .A2(new_n720), .A3(new_n721), .A4(new_n703), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n703), .A2(KEYINPUT109), .A3(new_n721), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n716), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n719), .A2(new_n703), .A3(new_n720), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n724), .B1(new_n725), .B2(new_n723), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(KEYINPUT54), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n716), .A2(new_n722), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT54), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n727), .A2(new_n730), .ZN(new_n731));
  AND4_X1   g545(.A1(new_n490), .A2(new_n678), .A3(new_n610), .A4(new_n639), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n732), .A2(new_n487), .A3(new_n550), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n628), .A2(new_n356), .ZN(new_n734));
  NOR3_X1   g548(.A1(new_n734), .A2(new_n651), .A3(new_n489), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(new_n619), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n733), .A2(G952), .A3(new_n263), .A4(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(KEYINPUT113), .ZN(new_n738));
  NOR4_X1   g552(.A1(new_n651), .A2(new_n489), .A3(new_n609), .A4(new_n643), .ZN(new_n739));
  INV_X1    g553(.A(new_n636), .ZN(new_n740));
  AND2_X1   g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  OR2_X1    g555(.A1(new_n741), .A2(KEYINPUT48), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(KEYINPUT48), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n738), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(KEYINPUT114), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n682), .A2(new_n358), .A3(new_n610), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(KEYINPUT111), .ZN(new_n747));
  INV_X1    g561(.A(new_n735), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  XOR2_X1   g563(.A(new_n749), .B(KEYINPUT50), .Z(new_n750));
  NAND4_X1  g564(.A1(new_n732), .A2(new_n687), .A3(new_n549), .A4(new_n548), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(KEYINPUT112), .ZN(new_n752));
  INV_X1    g566(.A(new_n708), .ZN(new_n753));
  AOI211_X1 g567(.A(new_n750), .B(new_n752), .C1(new_n753), .C2(new_n739), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n748), .A2(new_n643), .ZN(new_n755));
  INV_X1    g569(.A(new_n672), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n679), .A2(new_n419), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(KEYINPUT110), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n755), .B1(new_n756), .B2(new_n758), .ZN(new_n759));
  AOI21_X1  g573(.A(KEYINPUT51), .B1(new_n754), .B2(new_n759), .ZN(new_n760));
  NOR3_X1   g574(.A1(new_n731), .A2(new_n745), .A3(new_n760), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n672), .B1(new_n419), .B2(new_n679), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(new_n755), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n754), .A2(KEYINPUT51), .A3(new_n763), .ZN(new_n764));
  AND2_X1   g578(.A1(new_n761), .A2(new_n764), .ZN(new_n765));
  NOR2_X1   g579(.A1(G952), .A2(G953), .ZN(new_n766));
  OAI211_X1 g580(.A(new_n677), .B(new_n686), .C1(new_n765), .C2(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(G952), .ZN(new_n768));
  AOI22_X1  g582(.A1(new_n761), .A2(new_n764), .B1(new_n768), .B2(new_n263), .ZN(new_n769));
  OAI21_X1  g583(.A(KEYINPUT115), .B1(new_n769), .B2(new_n685), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n767), .A2(new_n770), .ZN(G75));
  NOR2_X1   g585(.A1(new_n263), .A2(G952), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n392), .A2(new_n402), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(new_n400), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(KEYINPUT116), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(KEYINPUT55), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n716), .A2(new_n722), .A3(G902), .ZN(new_n777));
  INV_X1    g591(.A(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(G210), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT56), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n776), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  OR2_X1    g595(.A1(new_n778), .A2(KEYINPUT117), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n778), .A2(KEYINPUT117), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n782), .A2(new_n412), .A3(new_n783), .ZN(new_n784));
  AND2_X1   g598(.A1(new_n776), .A2(new_n780), .ZN(new_n785));
  AOI211_X1 g599(.A(new_n772), .B(new_n781), .C1(new_n784), .C2(new_n785), .ZN(G51));
  INV_X1    g600(.A(KEYINPUT118), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n716), .A2(new_n722), .A3(KEYINPUT54), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n730), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n728), .A2(KEYINPUT118), .A3(new_n729), .ZN(new_n790));
  NAND2_X1  g604(.A1(G469), .A2(G902), .ZN(new_n791));
  XOR2_X1   g605(.A(new_n791), .B(KEYINPUT57), .Z(new_n792));
  NAND3_X1  g606(.A1(new_n789), .A2(new_n790), .A3(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(new_n444), .ZN(new_n794));
  XOR2_X1   g608(.A(new_n794), .B(KEYINPUT119), .Z(new_n795));
  NAND4_X1  g609(.A1(new_n782), .A2(G469), .A3(new_n657), .A4(new_n783), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n772), .B1(new_n795), .B2(new_n796), .ZN(G54));
  NAND4_X1  g611(.A1(new_n782), .A2(KEYINPUT58), .A3(G475), .A4(new_n783), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n478), .A2(new_n479), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n798), .A2(new_n799), .ZN(new_n801));
  NOR3_X1   g615(.A1(new_n800), .A2(new_n801), .A3(new_n772), .ZN(G60));
  NAND2_X1  g616(.A1(G478), .A2(G902), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(KEYINPUT59), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n789), .A2(new_n547), .A3(new_n790), .A4(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(new_n772), .ZN(new_n806));
  AND3_X1   g620(.A1(new_n805), .A2(KEYINPUT120), .A3(new_n806), .ZN(new_n807));
  AOI21_X1  g621(.A(KEYINPUT120), .B1(new_n805), .B2(new_n806), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n547), .B1(new_n731), .B2(new_n804), .ZN(new_n809));
  NOR3_X1   g623(.A1(new_n807), .A2(new_n808), .A3(new_n809), .ZN(G63));
  NAND2_X1  g624(.A1(G217), .A2(G902), .ZN(new_n811));
  XOR2_X1   g625(.A(new_n811), .B(KEYINPUT60), .Z(new_n812));
  NAND3_X1  g626(.A1(new_n716), .A2(new_n722), .A3(new_n812), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n813), .A2(new_n570), .ZN(new_n814));
  INV_X1    g628(.A(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n347), .A2(new_n349), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n813), .A2(new_n816), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n815), .A2(KEYINPUT61), .A3(new_n806), .A4(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT122), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n819), .B1(new_n817), .B2(new_n806), .ZN(new_n820));
  AOI211_X1 g634(.A(KEYINPUT122), .B(new_n772), .C1(new_n813), .C2(new_n816), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n820), .A2(new_n821), .A3(new_n814), .ZN(new_n822));
  XNOR2_X1  g636(.A(KEYINPUT121), .B(KEYINPUT61), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n822), .A2(KEYINPUT123), .A3(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT123), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n817), .A2(new_n806), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(KEYINPUT122), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n817), .A2(new_n819), .A3(new_n806), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n827), .A2(new_n815), .A3(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(new_n823), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n825), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n818), .B1(new_n824), .B2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT124), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  OAI211_X1 g648(.A(KEYINPUT124), .B(new_n818), .C1(new_n824), .C2(new_n831), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(G66));
  OAI21_X1  g650(.A(G953), .B1(new_n492), .B2(new_n396), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n837), .B1(new_n695), .B2(G953), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n773), .B1(G898), .B2(new_n263), .ZN(new_n839));
  XNOR2_X1  g653(.A(new_n838), .B(new_n839), .ZN(G69));
  INV_X1    g654(.A(new_n648), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n696), .A2(new_n604), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n675), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n636), .A2(new_n579), .A3(new_n623), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n663), .B1(new_n656), .B2(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n843), .A2(new_n704), .A3(new_n845), .ZN(new_n846));
  OR2_X1    g660(.A1(new_n846), .A2(KEYINPUT127), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(KEYINPUT127), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n847), .A2(new_n263), .A3(new_n848), .ZN(new_n849));
  XNOR2_X1  g663(.A(new_n275), .B(KEYINPUT125), .ZN(new_n850));
  XNOR2_X1  g664(.A(new_n850), .B(new_n469), .ZN(new_n851));
  INV_X1    g665(.A(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(G900), .A2(G953), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n849), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(new_n842), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n601), .A2(KEYINPUT62), .A3(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n601), .A2(new_n855), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT62), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n675), .B1(new_n856), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n688), .A2(new_n551), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n615), .A2(new_n598), .A3(new_n639), .A4(new_n861), .ZN(new_n862));
  AND3_X1   g676(.A1(new_n860), .A2(new_n664), .A3(new_n862), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n851), .B1(new_n863), .B2(G953), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n864), .A2(KEYINPUT126), .ZN(new_n865));
  OR2_X1    g679(.A1(new_n864), .A2(KEYINPUT126), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n854), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n263), .B1(G227), .B2(G900), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(new_n868), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n854), .A2(new_n870), .A3(new_n865), .A4(new_n866), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n869), .A2(new_n871), .ZN(G72));
  NAND2_X1  g686(.A1(G472), .A2(G902), .ZN(new_n873));
  XOR2_X1   g687(.A(new_n873), .B(KEYINPUT63), .Z(new_n874));
  INV_X1    g688(.A(new_n874), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n875), .B1(new_n863), .B2(new_n695), .ZN(new_n876));
  INV_X1    g690(.A(new_n587), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n806), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(new_n726), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n259), .A2(new_n265), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n276), .A2(new_n277), .ZN(new_n881));
  AOI211_X1 g695(.A(new_n875), .B(new_n879), .C1(new_n880), .C2(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n847), .A2(new_n695), .A3(new_n848), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n265), .B1(new_n883), .B2(new_n874), .ZN(new_n884));
  AOI211_X1 g698(.A(new_n878), .B(new_n882), .C1(new_n884), .C2(new_n259), .ZN(G57));
endmodule


