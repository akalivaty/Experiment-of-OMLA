//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 1 1 1 0 1 1 0 0 1 1 0 1 0 1 0 0 0 1 1 1 0 1 1 1 1 0 0 1 1 1 0 1 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:57 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n450, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n576, new_n577, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n592, new_n594, new_n595, new_n596,
    new_n597, new_n598, new_n599, new_n600, new_n602, new_n603, new_n604,
    new_n605, new_n607, new_n608, new_n609, new_n610, new_n611, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n636, new_n639,
    new_n641, new_n642, new_n643, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1223, new_n1224;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT65), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT66), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(KEYINPUT67), .B(KEYINPUT2), .Z(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  INV_X1    g034(.A(G567), .ZN(new_n460));
  OAI21_X1  g035(.A(new_n459), .B1(new_n460), .B2(new_n455), .ZN(new_n461));
  XOR2_X1   g036(.A(new_n461), .B(KEYINPUT68), .Z(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(KEYINPUT69), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n464), .B1(new_n465), .B2(G2105), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n467), .A2(KEYINPUT69), .A3(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G101), .ZN(new_n470));
  OR2_X1    g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n473), .A2(G137), .A3(new_n467), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n470), .A2(new_n474), .ZN(new_n475));
  AND2_X1   g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  NOR2_X1   g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  OAI21_X1  g052(.A(G125), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(G113), .A2(G2104), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n467), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n475), .A2(new_n480), .ZN(G160));
  NAND2_X1  g056(.A1(new_n473), .A2(G2105), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  AOI21_X1  g059(.A(G2105), .B1(new_n471), .B2(new_n472), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G136), .ZN(new_n486));
  OR2_X1    g061(.A1(G100), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G112), .C2(new_n467), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n484), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G162));
  NAND2_X1  g065(.A1(G126), .A2(G2105), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT71), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(KEYINPUT4), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n467), .A2(G138), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n491), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(new_n473), .ZN(new_n496));
  OAI211_X1 g071(.A(G138), .B(new_n467), .C1(new_n476), .C2(new_n477), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(new_n493), .ZN(new_n498));
  OAI21_X1  g073(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(G114), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n501), .A2(KEYINPUT70), .A3(G2105), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT70), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n503), .B1(new_n467), .B2(G114), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n500), .A2(new_n502), .A3(new_n504), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n496), .A2(new_n498), .A3(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(G164));
  AND3_X1   g082(.A1(KEYINPUT73), .A2(KEYINPUT5), .A3(G543), .ZN(new_n508));
  AOI21_X1  g083(.A(KEYINPUT5), .B1(KEYINPUT73), .B2(G543), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G62), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AND2_X1   g087(.A1(new_n512), .A2(KEYINPUT76), .ZN(new_n513));
  NAND2_X1  g088(.A1(G75), .A2(G543), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n514), .B1(new_n512), .B2(KEYINPUT76), .ZN(new_n515));
  OAI21_X1  g090(.A(G651), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT72), .ZN(new_n517));
  XNOR2_X1  g092(.A(KEYINPUT6), .B(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G543), .ZN(new_n519));
  INV_X1    g094(.A(G50), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n517), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(G543), .ZN(new_n522));
  OR2_X1    g097(.A1(KEYINPUT6), .A2(G651), .ZN(new_n523));
  NAND2_X1  g098(.A1(KEYINPUT6), .A2(G651), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n525), .A2(KEYINPUT72), .A3(G50), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n521), .A2(new_n526), .ZN(new_n527));
  AND2_X1   g102(.A1(KEYINPUT6), .A2(G651), .ZN(new_n528));
  NOR2_X1   g103(.A1(KEYINPUT6), .A2(G651), .ZN(new_n529));
  OAI22_X1  g104(.A1(new_n508), .A2(new_n509), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT74), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(KEYINPUT73), .A2(G543), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT5), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g110(.A1(KEYINPUT73), .A2(KEYINPUT5), .A3(G543), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n537), .A2(KEYINPUT74), .A3(new_n518), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n532), .A2(G88), .A3(new_n538), .ZN(new_n539));
  AND3_X1   g114(.A1(new_n527), .A2(KEYINPUT75), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g115(.A(KEYINPUT75), .B1(new_n527), .B2(new_n539), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n516), .B1(new_n540), .B2(new_n541), .ZN(G303));
  INV_X1    g117(.A(G303), .ZN(G166));
  AND2_X1   g118(.A1(G63), .A2(G651), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n525), .A2(G51), .B1(new_n537), .B2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(new_n545), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n532), .A2(G89), .A3(new_n538), .ZN(new_n547));
  NAND3_X1  g122(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT7), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT77), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n547), .A2(KEYINPUT77), .A3(new_n549), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n546), .B1(new_n552), .B2(new_n553), .ZN(G168));
  AOI22_X1  g129(.A1(new_n537), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n555));
  INV_X1    g130(.A(G651), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n525), .A2(G52), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n532), .A2(new_n538), .ZN(new_n559));
  INV_X1    g134(.A(G90), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NOR2_X1   g136(.A1(new_n561), .A2(KEYINPUT78), .ZN(new_n562));
  INV_X1    g137(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n561), .A2(KEYINPUT78), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n557), .B1(new_n563), .B2(new_n564), .ZN(G171));
  INV_X1    g140(.A(new_n559), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G81), .ZN(new_n567));
  NAND2_X1  g142(.A1(G68), .A2(G543), .ZN(new_n568));
  INV_X1    g143(.A(G56), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n568), .B1(new_n510), .B2(new_n569), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n570), .A2(G651), .B1(G43), .B2(new_n525), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n567), .A2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n573), .A2(G860), .ZN(G153));
  NAND4_X1  g149(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g150(.A1(G1), .A2(G3), .ZN(new_n576));
  XNOR2_X1  g151(.A(new_n576), .B(KEYINPUT8), .ZN(new_n577));
  NAND4_X1  g152(.A1(G319), .A2(G483), .A3(G661), .A4(new_n577), .ZN(G188));
  NAND3_X1  g153(.A1(new_n532), .A2(G91), .A3(new_n538), .ZN(new_n579));
  OAI211_X1 g154(.A(G53), .B(G543), .C1(new_n528), .C2(new_n529), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n580), .A2(KEYINPUT79), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT79), .ZN(new_n582));
  NAND4_X1  g157(.A1(new_n518), .A2(new_n582), .A3(G53), .A4(G543), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n581), .A2(new_n583), .A3(KEYINPUT9), .ZN(new_n584));
  INV_X1    g159(.A(G65), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n585), .B1(new_n535), .B2(new_n536), .ZN(new_n586));
  AND2_X1   g161(.A1(G78), .A2(G543), .ZN(new_n587));
  OAI21_X1  g162(.A(G651), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT9), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n580), .A2(KEYINPUT79), .A3(new_n589), .ZN(new_n590));
  NAND4_X1  g165(.A1(new_n579), .A2(new_n584), .A3(new_n588), .A4(new_n590), .ZN(G299));
  INV_X1    g166(.A(new_n564), .ZN(new_n592));
  OAI22_X1  g167(.A1(new_n592), .A2(new_n562), .B1(new_n556), .B2(new_n555), .ZN(G301));
  INV_X1    g168(.A(new_n553), .ZN(new_n594));
  AOI21_X1  g169(.A(KEYINPUT77), .B1(new_n547), .B2(new_n549), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n545), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n596), .A2(KEYINPUT80), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT80), .ZN(new_n598));
  NAND2_X1  g173(.A1(G168), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(G286));
  INV_X1    g176(.A(G74), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n510), .A2(new_n602), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n603), .A2(G651), .B1(G49), .B2(new_n525), .ZN(new_n604));
  INV_X1    g179(.A(G87), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n559), .B2(new_n605), .ZN(G288));
  NAND2_X1  g181(.A1(G73), .A2(G543), .ZN(new_n607));
  INV_X1    g182(.A(G61), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n510), .B2(new_n608), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n609), .A2(G651), .B1(G48), .B2(new_n525), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n532), .A2(G86), .A3(new_n538), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(G305));
  AOI22_X1  g187(.A1(new_n537), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n613));
  NOR2_X1   g188(.A1(new_n613), .A2(new_n556), .ZN(new_n614));
  INV_X1    g189(.A(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n525), .A2(G47), .ZN(new_n616));
  INV_X1    g191(.A(G85), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n559), .B2(new_n617), .ZN(new_n618));
  AND2_X1   g193(.A1(new_n618), .A2(KEYINPUT81), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n618), .A2(KEYINPUT81), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n615), .B1(new_n619), .B2(new_n620), .ZN(G290));
  NAND2_X1  g196(.A1(G301), .A2(G868), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n566), .A2(KEYINPUT10), .A3(G92), .ZN(new_n623));
  INV_X1    g198(.A(KEYINPUT10), .ZN(new_n624));
  INV_X1    g199(.A(G92), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n624), .B1(new_n559), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n623), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(G79), .A2(G543), .ZN(new_n628));
  XNOR2_X1  g203(.A(KEYINPUT82), .B(G66), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n628), .B1(new_n510), .B2(new_n629), .ZN(new_n630));
  AOI22_X1  g205(.A1(new_n630), .A2(G651), .B1(G54), .B2(new_n525), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n627), .A2(new_n631), .ZN(new_n632));
  INV_X1    g207(.A(new_n632), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n622), .B1(G868), .B2(new_n633), .ZN(G284));
  OAI21_X1  g209(.A(new_n622), .B1(G868), .B2(new_n633), .ZN(G321));
  NOR2_X1   g210(.A1(G299), .A2(G868), .ZN(new_n636));
  AOI21_X1  g211(.A(new_n636), .B1(new_n600), .B2(G868), .ZN(G297));
  AOI21_X1  g212(.A(new_n636), .B1(new_n600), .B2(G868), .ZN(G280));
  INV_X1    g213(.A(G559), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n633), .B1(new_n639), .B2(G860), .ZN(G148));
  NOR2_X1   g215(.A1(new_n572), .A2(G868), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n633), .A2(new_n639), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT83), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n641), .B1(new_n643), .B2(G868), .ZN(G323));
  XNOR2_X1  g219(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g220(.A1(new_n483), .A2(G123), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT84), .ZN(new_n647));
  OAI21_X1  g222(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n648));
  INV_X1    g223(.A(G111), .ZN(new_n649));
  AOI21_X1  g224(.A(new_n648), .B1(new_n649), .B2(G2105), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n650), .B1(G135), .B2(new_n485), .ZN(new_n651));
  AND2_X1   g226(.A1(new_n647), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(G2096), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n469), .A2(new_n473), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT12), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT13), .ZN(new_n656));
  INV_X1    g231(.A(G2100), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n656), .A2(new_n657), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n653), .A2(new_n658), .A3(new_n659), .ZN(G156));
  XOR2_X1   g235(.A(KEYINPUT15), .B(G2435), .Z(new_n661));
  XNOR2_X1  g236(.A(KEYINPUT86), .B(G2438), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2427), .B(G2430), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  OR2_X1    g240(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(KEYINPUT85), .B(KEYINPUT14), .Z(new_n667));
  NAND2_X1  g242(.A1(new_n663), .A2(new_n665), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n666), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G2451), .B(G2454), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT16), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1341), .B(G1348), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n669), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G2443), .B(G2446), .ZN(new_n675));
  OR2_X1    g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n674), .A2(new_n675), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n676), .A2(new_n677), .A3(G14), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT87), .ZN(G401));
  INV_X1    g254(.A(KEYINPUT18), .ZN(new_n680));
  XOR2_X1   g255(.A(G2084), .B(G2090), .Z(new_n681));
  XNOR2_X1  g256(.A(G2067), .B(G2678), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n683), .A2(KEYINPUT17), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n681), .A2(new_n682), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n680), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(new_n657), .ZN(new_n687));
  XOR2_X1   g262(.A(G2072), .B(G2078), .Z(new_n688));
  AOI21_X1  g263(.A(new_n688), .B1(new_n683), .B2(KEYINPUT18), .ZN(new_n689));
  XOR2_X1   g264(.A(new_n689), .B(G2096), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n687), .B(new_n690), .ZN(G227));
  XNOR2_X1  g266(.A(G1956), .B(G2474), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1961), .B(G1966), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  OR2_X1    g270(.A1(new_n695), .A2(KEYINPUT89), .ZN(new_n696));
  XNOR2_X1  g271(.A(G1971), .B(G1976), .ZN(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT88), .B(KEYINPUT19), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n695), .A2(KEYINPUT89), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n696), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  XOR2_X1   g276(.A(KEYINPUT90), .B(KEYINPUT20), .Z(new_n702));
  OR2_X1    g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n701), .A2(new_n702), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n699), .A2(new_n692), .A3(new_n693), .ZN(new_n705));
  INV_X1    g280(.A(new_n699), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n692), .A2(new_n693), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n706), .A2(new_n695), .A3(new_n707), .ZN(new_n708));
  NAND4_X1  g283(.A1(new_n703), .A2(new_n704), .A3(new_n705), .A4(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT91), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n709), .B(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(G1991), .B(G1996), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(G1981), .B(G1986), .ZN(new_n715));
  OR2_X1    g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n714), .A2(new_n715), .ZN(new_n717));
  AND2_X1   g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(G229));
  INV_X1    g294(.A(G290), .ZN(new_n720));
  XOR2_X1   g295(.A(KEYINPUT93), .B(G16), .Z(new_n721));
  INV_X1    g296(.A(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  OR2_X1    g298(.A1(new_n722), .A2(G24), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n725), .A2(KEYINPUT94), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT94), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n723), .A2(new_n727), .A3(new_n724), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(G1986), .ZN(new_n730));
  INV_X1    g305(.A(G29), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n731), .A2(G25), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n485), .A2(G131), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n467), .A2(G107), .ZN(new_n734));
  OAI21_X1  g309(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n735));
  INV_X1    g310(.A(G119), .ZN(new_n736));
  OAI221_X1 g311(.A(new_n733), .B1(new_n734), .B2(new_n735), .C1(new_n736), .C2(new_n482), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT92), .Z(new_n738));
  INV_X1    g313(.A(new_n738), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n732), .B1(new_n739), .B2(new_n731), .ZN(new_n740));
  XOR2_X1   g315(.A(KEYINPUT35), .B(G1991), .Z(new_n741));
  XOR2_X1   g316(.A(new_n740), .B(new_n741), .Z(new_n742));
  NAND2_X1  g317(.A1(new_n721), .A2(G22), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(G166), .B2(new_n721), .ZN(new_n744));
  OR2_X1    g319(.A1(new_n744), .A2(G1971), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n744), .A2(G1971), .ZN(new_n746));
  MUX2_X1   g321(.A(G6), .B(G305), .S(G16), .Z(new_n747));
  XOR2_X1   g322(.A(KEYINPUT32), .B(G1981), .Z(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(G16), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n750), .A2(G23), .ZN(new_n751));
  INV_X1    g326(.A(G288), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n751), .B1(new_n752), .B2(new_n750), .ZN(new_n753));
  XNOR2_X1  g328(.A(KEYINPUT33), .B(G1976), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT95), .Z(new_n755));
  XNOR2_X1  g330(.A(new_n753), .B(new_n755), .ZN(new_n756));
  NAND4_X1  g331(.A1(new_n745), .A2(new_n746), .A3(new_n749), .A4(new_n756), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n742), .B1(new_n757), .B2(KEYINPUT34), .ZN(new_n758));
  OR2_X1    g333(.A1(new_n757), .A2(KEYINPUT34), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n730), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT36), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n750), .A2(G21), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G168), .B2(new_n750), .ZN(new_n763));
  OR2_X1    g338(.A1(new_n763), .A2(G1966), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n731), .A2(G32), .ZN(new_n765));
  NAND3_X1  g340(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT26), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(new_n483), .B2(G129), .ZN(new_n768));
  AOI22_X1  g343(.A1(G141), .A2(new_n485), .B1(new_n469), .B2(G105), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(new_n770), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n765), .B1(new_n771), .B2(new_n731), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT27), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(G1996), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n763), .A2(G1966), .ZN(new_n775));
  INV_X1    g350(.A(G11), .ZN(new_n776));
  OR2_X1    g351(.A1(new_n776), .A2(KEYINPUT31), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n776), .A2(KEYINPUT31), .ZN(new_n778));
  INV_X1    g353(.A(KEYINPUT30), .ZN(new_n779));
  AND2_X1   g354(.A1(new_n779), .A2(G28), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n731), .B1(new_n779), .B2(G28), .ZN(new_n781));
  OAI211_X1 g356(.A(new_n777), .B(new_n778), .C1(new_n780), .C2(new_n781), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(new_n652), .B2(G29), .ZN(new_n783));
  INV_X1    g358(.A(G2084), .ZN(new_n784));
  INV_X1    g359(.A(KEYINPUT24), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n731), .B1(new_n785), .B2(G34), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(new_n785), .B2(G34), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(G160), .B2(G29), .ZN(new_n788));
  INV_X1    g363(.A(new_n788), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n783), .B1(new_n784), .B2(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(G2078), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n731), .A2(G27), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(G164), .B2(new_n731), .ZN(new_n793));
  INV_X1    g368(.A(new_n793), .ZN(new_n794));
  AOI22_X1  g369(.A1(new_n791), .A2(new_n794), .B1(new_n789), .B2(new_n784), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(new_n791), .B2(new_n794), .ZN(new_n796));
  INV_X1    g371(.A(KEYINPUT97), .ZN(new_n797));
  OR3_X1    g372(.A1(new_n797), .A2(G29), .A3(G33), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n797), .B1(G29), .B2(G33), .ZN(new_n799));
  INV_X1    g374(.A(KEYINPUT25), .ZN(new_n800));
  NAND2_X1  g375(.A1(G103), .A2(G2104), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n800), .B1(new_n801), .B2(G2105), .ZN(new_n802));
  NAND4_X1  g377(.A1(new_n467), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n803));
  AOI22_X1  g378(.A1(new_n485), .A2(G139), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  AOI22_X1  g379(.A1(new_n473), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n804), .B1(new_n467), .B2(new_n805), .ZN(new_n806));
  OAI211_X1 g381(.A(new_n798), .B(new_n799), .C1(new_n806), .C2(new_n731), .ZN(new_n807));
  XOR2_X1   g382(.A(new_n807), .B(G2072), .Z(new_n808));
  NOR3_X1   g383(.A1(new_n790), .A2(new_n796), .A3(new_n808), .ZN(new_n809));
  AND4_X1   g384(.A1(new_n764), .A2(new_n774), .A3(new_n775), .A4(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n750), .A2(G5), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(G171), .B2(new_n750), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT98), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n813), .A2(G1961), .ZN(new_n814));
  INV_X1    g389(.A(KEYINPUT99), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  AOI21_X1  g391(.A(KEYINPUT99), .B1(new_n813), .B2(G1961), .ZN(new_n817));
  OAI221_X1 g392(.A(new_n810), .B1(G1961), .B2(new_n813), .C1(new_n816), .C2(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n818), .A2(KEYINPUT100), .ZN(new_n819));
  NOR2_X1   g394(.A1(G29), .A2(G35), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n820), .B1(G162), .B2(G29), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT29), .ZN(new_n822));
  INV_X1    g397(.A(G2090), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n721), .A2(G20), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT23), .ZN(new_n826));
  INV_X1    g401(.A(G299), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n826), .B1(new_n827), .B2(new_n750), .ZN(new_n828));
  INV_X1    g403(.A(G1956), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n828), .B(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n485), .A2(G140), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n467), .A2(G116), .ZN(new_n832));
  OAI21_X1  g407(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n833));
  INV_X1    g408(.A(G128), .ZN(new_n834));
  OAI221_X1 g409(.A(new_n831), .B1(new_n832), .B2(new_n833), .C1(new_n834), .C2(new_n482), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n835), .A2(G29), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n731), .A2(G26), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT28), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(G2067), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n722), .A2(G19), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n841), .B1(new_n573), .B2(new_n722), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(G1341), .ZN(new_n843));
  INV_X1    g418(.A(G1348), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n633), .A2(G16), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n845), .B1(G4), .B2(G16), .ZN(new_n846));
  AOI211_X1 g421(.A(new_n840), .B(new_n843), .C1(new_n844), .C2(new_n846), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n847), .B1(new_n844), .B2(new_n846), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT96), .ZN(new_n849));
  OAI211_X1 g424(.A(new_n824), .B(new_n830), .C1(new_n848), .C2(new_n849), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n850), .B1(new_n849), .B2(new_n848), .ZN(new_n851));
  OR2_X1    g426(.A1(new_n818), .A2(KEYINPUT100), .ZN(new_n852));
  NAND4_X1  g427(.A1(new_n761), .A2(new_n819), .A3(new_n851), .A4(new_n852), .ZN(G150));
  INV_X1    g428(.A(G150), .ZN(G311));
  NAND3_X1  g429(.A1(new_n532), .A2(G93), .A3(new_n538), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n525), .A2(G55), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n857), .A2(KEYINPUT101), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT101), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n855), .A2(new_n859), .A3(new_n856), .ZN(new_n860));
  NAND2_X1  g435(.A1(G80), .A2(G543), .ZN(new_n861));
  INV_X1    g436(.A(G67), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n861), .B1(new_n510), .B2(new_n862), .ZN(new_n863));
  AOI22_X1  g438(.A1(new_n858), .A2(new_n860), .B1(G651), .B2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT102), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n572), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n863), .A2(G651), .ZN(new_n867));
  INV_X1    g442(.A(new_n860), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n859), .B1(new_n855), .B2(new_n856), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n867), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n870), .A2(KEYINPUT102), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n866), .A2(new_n871), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n573), .B1(new_n870), .B2(KEYINPUT102), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n864), .A2(new_n865), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(KEYINPUT38), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n633), .A2(G559), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n877), .B(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT39), .ZN(new_n880));
  AOI21_X1  g455(.A(G860), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n881), .B1(new_n880), .B2(new_n879), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n870), .A2(G860), .ZN(new_n883));
  XOR2_X1   g458(.A(new_n883), .B(KEYINPUT37), .Z(new_n884));
  NAND2_X1  g459(.A1(new_n882), .A2(new_n884), .ZN(G145));
  INV_X1    g460(.A(G130), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n467), .A2(G118), .ZN(new_n887));
  OAI21_X1  g462(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n888));
  OAI22_X1  g463(.A1(new_n482), .A2(new_n886), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n889), .B1(G142), .B2(new_n485), .ZN(new_n890));
  XOR2_X1   g465(.A(new_n890), .B(new_n655), .Z(new_n891));
  XOR2_X1   g466(.A(new_n770), .B(new_n806), .Z(new_n892));
  XNOR2_X1  g467(.A(new_n891), .B(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n835), .B(G164), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n738), .B(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n893), .B(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n489), .B(G160), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n652), .B(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(G37), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n899), .B1(new_n898), .B2(new_n896), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g476(.A(new_n643), .B(new_n876), .Z(new_n902));
  INV_X1    g477(.A(KEYINPUT103), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n632), .A2(new_n827), .ZN(new_n904));
  AOI21_X1  g479(.A(G299), .B1(new_n627), .B2(new_n631), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n903), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  OAI21_X1  g481(.A(KEYINPUT103), .B1(new_n632), .B2(new_n827), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n906), .A2(KEYINPUT41), .A3(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT104), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n904), .A2(new_n905), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n909), .B1(new_n910), .B2(KEYINPUT41), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n908), .A2(new_n911), .ZN(new_n912));
  NAND4_X1  g487(.A1(new_n906), .A2(new_n909), .A3(new_n907), .A4(KEYINPUT41), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  OR2_X1    g490(.A1(new_n902), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(G290), .A2(G288), .ZN(new_n917));
  OAI211_X1 g492(.A(new_n752), .B(new_n615), .C1(new_n619), .C2(new_n620), .ZN(new_n918));
  AOI21_X1  g493(.A(KEYINPUT105), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  XNOR2_X1  g494(.A(G303), .B(G305), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n917), .A2(new_n918), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT105), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n917), .A2(KEYINPUT105), .A3(new_n918), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n921), .B1(new_n926), .B2(new_n920), .ZN(new_n927));
  XOR2_X1   g502(.A(new_n927), .B(KEYINPUT42), .Z(new_n928));
  AND2_X1   g503(.A1(new_n906), .A2(new_n907), .ZN(new_n929));
  INV_X1    g504(.A(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n902), .A2(new_n930), .ZN(new_n931));
  AND3_X1   g506(.A1(new_n916), .A2(new_n928), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n928), .B1(new_n916), .B2(new_n931), .ZN(new_n933));
  OAI21_X1  g508(.A(G868), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n934), .B1(G868), .B2(new_n864), .ZN(G295));
  OAI21_X1  g510(.A(new_n934), .B1(G868), .B2(new_n864), .ZN(G331));
  NAND2_X1  g511(.A1(new_n600), .A2(G171), .ZN(new_n937));
  NAND2_X1  g512(.A1(G301), .A2(new_n596), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n866), .A2(new_n871), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n873), .A2(new_n874), .ZN(new_n940));
  OAI211_X1 g515(.A(new_n937), .B(new_n938), .C1(new_n939), .C2(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(G301), .B1(new_n597), .B2(new_n599), .ZN(new_n942));
  NOR2_X1   g517(.A1(G171), .A2(G168), .ZN(new_n943));
  OAI211_X1 g518(.A(new_n872), .B(new_n875), .C1(new_n942), .C2(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n929), .B1(new_n941), .B2(new_n944), .ZN(new_n945));
  AND2_X1   g520(.A1(new_n941), .A2(new_n944), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n945), .B1(new_n914), .B2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(new_n927), .ZN(new_n948));
  AOI21_X1  g523(.A(G37), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  XOR2_X1   g524(.A(KEYINPUT107), .B(KEYINPUT43), .Z(new_n950));
  INV_X1    g525(.A(KEYINPUT108), .ZN(new_n951));
  INV_X1    g526(.A(new_n910), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n941), .A2(new_n944), .A3(KEYINPUT41), .A4(new_n952), .ZN(new_n953));
  AND2_X1   g528(.A1(new_n927), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n941), .A2(new_n944), .A3(KEYINPUT41), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(new_n929), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n951), .B1(new_n954), .B2(new_n956), .ZN(new_n957));
  AND4_X1   g532(.A1(new_n951), .A2(new_n956), .A3(new_n927), .A4(new_n953), .ZN(new_n958));
  OAI211_X1 g533(.A(new_n949), .B(new_n950), .C1(new_n957), .C2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(new_n950), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n946), .A2(new_n914), .ZN(new_n961));
  INV_X1    g536(.A(new_n945), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n961), .A2(new_n948), .A3(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(G37), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n947), .A2(new_n948), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n960), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n959), .A2(new_n967), .ZN(new_n968));
  XOR2_X1   g543(.A(KEYINPUT106), .B(KEYINPUT44), .Z(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  OAI211_X1 g545(.A(new_n949), .B(new_n950), .C1(new_n948), .C2(new_n947), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n954), .A2(new_n956), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(KEYINPUT108), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n954), .A2(new_n951), .A3(new_n956), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n965), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT43), .ZN(new_n976));
  OAI211_X1 g551(.A(KEYINPUT44), .B(new_n971), .C1(new_n975), .C2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n970), .A2(new_n977), .ZN(G397));
  INV_X1    g553(.A(KEYINPUT125), .ZN(new_n979));
  INV_X1    g554(.A(G8), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT115), .ZN(new_n981));
  AND2_X1   g556(.A1(new_n470), .A2(new_n474), .ZN(new_n982));
  INV_X1    g557(.A(G125), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n983), .B1(new_n471), .B2(new_n472), .ZN(new_n984));
  INV_X1    g559(.A(new_n479), .ZN(new_n985));
  OAI21_X1  g560(.A(G2105), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n982), .A2(G40), .A3(new_n784), .A4(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(G1384), .ZN(new_n988));
  INV_X1    g563(.A(new_n491), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT4), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n990), .A2(KEYINPUT71), .ZN(new_n991));
  INV_X1    g566(.A(G138), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n992), .A2(G2105), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n989), .B1(new_n991), .B2(new_n993), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n476), .A2(new_n477), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n505), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n991), .B1(new_n485), .B2(G138), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n988), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT50), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  XNOR2_X1  g575(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n1001));
  OAI211_X1 g576(.A(new_n988), .B(new_n1001), .C1(new_n996), .C2(new_n997), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n987), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT45), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n998), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(G40), .ZN(new_n1006));
  NOR3_X1   g581(.A1(new_n475), .A2(new_n1006), .A3(new_n480), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n506), .A2(KEYINPUT45), .A3(new_n988), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1005), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(G1966), .ZN(new_n1010));
  AOI22_X1  g585(.A1(new_n981), .A2(new_n1003), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1012));
  INV_X1    g587(.A(new_n987), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(KEYINPUT115), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n980), .B1(new_n1011), .B2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g591(.A(KEYINPUT124), .B1(G168), .B2(new_n980), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT124), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n596), .A2(new_n1018), .A3(G8), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n979), .B1(new_n1016), .B2(new_n1020), .ZN(new_n1021));
  AND2_X1   g596(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1002), .ZN(new_n1024));
  AOI21_X1  g599(.A(KEYINPUT50), .B1(new_n506), .B2(new_n988), .ZN(new_n1025));
  OAI211_X1 g600(.A(new_n1013), .B(new_n981), .C1(new_n1024), .C2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1023), .A2(new_n1026), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1003), .A2(new_n981), .ZN(new_n1028));
  OAI21_X1  g603(.A(G8), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1022), .A2(new_n1029), .A3(KEYINPUT125), .ZN(new_n1030));
  AND3_X1   g605(.A1(new_n1021), .A2(new_n1030), .A3(KEYINPUT51), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT51), .ZN(new_n1032));
  OAI211_X1 g607(.A(new_n979), .B(new_n1032), .C1(new_n1016), .C2(new_n1020), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1020), .B1(new_n1028), .B2(new_n1027), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  OAI21_X1  g610(.A(KEYINPUT62), .B1(new_n1031), .B2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1021), .A2(new_n1030), .A3(KEYINPUT51), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT62), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1037), .A2(new_n1038), .A3(new_n1033), .A4(new_n1034), .ZN(new_n1039));
  INV_X1    g614(.A(G1981), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n610), .A2(new_n1040), .A3(new_n611), .ZN(new_n1041));
  XNOR2_X1  g616(.A(KEYINPUT113), .B(G86), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n532), .A2(new_n538), .A3(new_n1042), .ZN(new_n1043));
  AND2_X1   g618(.A1(new_n610), .A2(new_n1043), .ZN(new_n1044));
  OAI211_X1 g619(.A(KEYINPUT49), .B(new_n1041), .C1(new_n1044), .C2(new_n1040), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT49), .ZN(new_n1046));
  AND3_X1   g621(.A1(new_n610), .A2(new_n1040), .A3(new_n611), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1040), .B1(new_n610), .B2(new_n1043), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1046), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n986), .A2(G40), .A3(new_n470), .A4(new_n474), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n998), .A2(new_n1050), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1051), .A2(new_n980), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1045), .A2(new_n1049), .A3(new_n1052), .ZN(new_n1053));
  OAI211_X1 g628(.A(new_n604), .B(G1976), .C1(new_n559), .C2(new_n605), .ZN(new_n1054));
  INV_X1    g629(.A(G1976), .ZN(new_n1055));
  AOI21_X1  g630(.A(KEYINPUT52), .B1(G288), .B2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1052), .A2(new_n1054), .A3(new_n1056), .ZN(new_n1057));
  OAI211_X1 g632(.A(new_n1054), .B(G8), .C1(new_n1050), .C2(new_n998), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT112), .ZN(new_n1059));
  AND3_X1   g634(.A1(new_n1058), .A2(new_n1059), .A3(KEYINPUT52), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1059), .B1(new_n1058), .B2(KEYINPUT52), .ZN(new_n1061));
  OAI211_X1 g636(.A(new_n1053), .B(new_n1057), .C1(new_n1060), .C2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1062), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1050), .B1(new_n998), .B2(new_n1004), .ZN(new_n1064));
  AOI21_X1  g639(.A(G1971), .B1(new_n1064), .B2(new_n1008), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1012), .A2(new_n823), .A3(new_n1007), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n980), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1068), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1071), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n506), .A2(new_n999), .A3(new_n988), .ZN(new_n1074));
  AOI21_X1  g649(.A(KEYINPUT70), .B1(new_n501), .B2(G2105), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1075), .A2(new_n499), .ZN(new_n1076));
  AOI22_X1  g651(.A1(new_n473), .A2(new_n495), .B1(new_n1076), .B2(new_n502), .ZN(new_n1077));
  AOI21_X1  g652(.A(G1384), .B1(new_n1077), .B2(new_n498), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1001), .ZN(new_n1079));
  OAI211_X1 g654(.A(new_n1074), .B(new_n1007), .C1(new_n1078), .C2(new_n1079), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1080), .A2(G2090), .ZN(new_n1081));
  OAI21_X1  g656(.A(G8), .B1(new_n1081), .B2(new_n1065), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1073), .A2(new_n1082), .A3(new_n1069), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1063), .A2(new_n1072), .A3(new_n1083), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1007), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT118), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(G1961), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1012), .A2(KEYINPUT118), .A3(new_n1007), .ZN(new_n1089));
  AND3_X1   g664(.A1(new_n1087), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1005), .A2(new_n791), .A3(new_n1007), .A4(new_n1008), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT53), .ZN(new_n1092));
  XNOR2_X1  g667(.A(new_n1091), .B(new_n1092), .ZN(new_n1093));
  OAI21_X1  g668(.A(G171), .B1(new_n1090), .B2(new_n1093), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1084), .A2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1036), .A2(new_n1039), .A3(new_n1095), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1029), .A2(G286), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1097), .A2(new_n1063), .A3(new_n1072), .A4(new_n1083), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT63), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT116), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1098), .A2(KEYINPUT116), .A3(new_n1099), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1072), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1104), .A2(new_n1099), .ZN(new_n1105));
  OR3_X1    g680(.A1(new_n1068), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1105), .A2(new_n1063), .A3(new_n1106), .A4(new_n1097), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1102), .A2(new_n1103), .A3(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1053), .A2(new_n1055), .A3(new_n752), .ZN(new_n1109));
  XNOR2_X1  g684(.A(new_n1047), .B(KEYINPUT114), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  AOI22_X1  g686(.A1(new_n1104), .A2(new_n1063), .B1(new_n1052), .B2(new_n1111), .ZN(new_n1112));
  AND3_X1   g687(.A1(new_n1096), .A2(new_n1108), .A3(new_n1112), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1031), .A2(new_n1035), .ZN(new_n1114));
  AND3_X1   g689(.A1(new_n1063), .A2(new_n1072), .A3(new_n1083), .ZN(new_n1115));
  XNOR2_X1  g690(.A(new_n1091), .B(KEYINPUT53), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1087), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1117));
  AND3_X1   g692(.A1(new_n1116), .A2(G301), .A3(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(G301), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1119));
  NOR3_X1   g694(.A1(new_n1118), .A2(new_n1119), .A3(KEYINPUT54), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT54), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1116), .A2(G301), .A3(new_n1117), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1121), .B1(new_n1094), .B2(new_n1122), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1115), .B1(new_n1120), .B2(new_n1123), .ZN(new_n1124));
  OAI21_X1  g699(.A(KEYINPUT126), .B1(new_n1114), .B2(new_n1124), .ZN(new_n1125));
  OAI21_X1  g700(.A(KEYINPUT54), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1094), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1084), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT126), .ZN(new_n1129));
  OAI211_X1 g704(.A(new_n1128), .B(new_n1129), .C1(new_n1031), .C2(new_n1035), .ZN(new_n1130));
  AND2_X1   g705(.A1(new_n584), .A2(new_n590), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT57), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1131), .A2(new_n1132), .A3(new_n579), .A4(new_n588), .ZN(new_n1133));
  NAND2_X1  g708(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  XNOR2_X1  g710(.A(KEYINPUT56), .B(G2072), .ZN(new_n1136));
  AND4_X1   g711(.A1(new_n1007), .A2(new_n1005), .A3(new_n1008), .A4(new_n1136), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1050), .B1(new_n998), .B2(new_n1001), .ZN(new_n1138));
  AOI21_X1  g713(.A(G1956), .B1(new_n1138), .B2(new_n1074), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1135), .B1(new_n1137), .B2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1087), .A2(new_n844), .A3(new_n1089), .ZN(new_n1141));
  INV_X1    g716(.A(G2067), .ZN(new_n1142));
  AND3_X1   g717(.A1(new_n1051), .A2(KEYINPUT117), .A3(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(KEYINPUT117), .B1(new_n1051), .B2(new_n1142), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  AND2_X1   g720(.A1(new_n1141), .A2(new_n1145), .ZN(new_n1146));
  XNOR2_X1  g721(.A(G299), .B(new_n1132), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1080), .A2(new_n829), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1064), .A2(new_n1008), .A3(new_n1136), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1147), .A2(new_n1148), .A3(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(new_n633), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1140), .B1(new_n1146), .B2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1141), .A2(KEYINPUT60), .A3(new_n1145), .ZN(new_n1153));
  OR2_X1    g728(.A1(new_n1153), .A2(KEYINPUT122), .ZN(new_n1154));
  AND3_X1   g729(.A1(new_n1153), .A2(KEYINPUT122), .A3(new_n632), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n632), .B1(new_n1153), .B2(KEYINPUT122), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1154), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  OR2_X1    g732(.A1(new_n1146), .A2(KEYINPUT60), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT61), .ZN(new_n1160));
  AND3_X1   g735(.A1(new_n1147), .A2(new_n1148), .A3(new_n1149), .ZN(new_n1161));
  AOI22_X1  g736(.A1(new_n1148), .A2(new_n1149), .B1(new_n1134), .B2(new_n1133), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1160), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1163), .A2(KEYINPUT120), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT120), .ZN(new_n1165));
  OAI211_X1 g740(.A(new_n1165), .B(new_n1160), .C1(new_n1161), .C2(new_n1162), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1164), .A2(new_n1166), .ZN(new_n1167));
  XOR2_X1   g742(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n1168));
  INV_X1    g743(.A(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(G1996), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1064), .A2(new_n1170), .A3(new_n1008), .ZN(new_n1171));
  XOR2_X1   g746(.A(KEYINPUT58), .B(G1341), .Z(new_n1172));
  OAI21_X1  g747(.A(new_n1172), .B1(new_n998), .B2(new_n1050), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1171), .A2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1169), .B1(new_n1174), .B2(new_n573), .ZN(new_n1175));
  AOI211_X1 g750(.A(new_n572), .B(new_n1168), .C1(new_n1171), .C2(new_n1173), .ZN(new_n1176));
  NOR2_X1   g751(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1140), .A2(new_n1150), .A3(KEYINPUT61), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT121), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  NAND4_X1  g755(.A1(new_n1140), .A2(new_n1150), .A3(KEYINPUT121), .A4(KEYINPUT61), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n1177), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  AND2_X1   g757(.A1(new_n1167), .A2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1152), .B1(new_n1159), .B2(new_n1183), .ZN(new_n1184));
  OAI211_X1 g759(.A(new_n1125), .B(new_n1130), .C1(new_n1184), .C2(KEYINPUT123), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT123), .ZN(new_n1186));
  AOI211_X1 g761(.A(new_n1186), .B(new_n1152), .C1(new_n1159), .C2(new_n1183), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1113), .B1(new_n1185), .B2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1007), .A2(new_n1004), .A3(new_n998), .ZN(new_n1189));
  XOR2_X1   g764(.A(new_n1189), .B(KEYINPUT110), .Z(new_n1190));
  XNOR2_X1  g765(.A(new_n835), .B(new_n1142), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1191), .B1(new_n1170), .B2(new_n771), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1190), .A2(new_n1192), .ZN(new_n1193));
  NOR2_X1   g768(.A1(new_n1189), .A2(G1996), .ZN(new_n1194));
  INV_X1    g769(.A(new_n1194), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n1193), .B1(new_n770), .B2(new_n1195), .ZN(new_n1196));
  XOR2_X1   g771(.A(new_n738), .B(new_n741), .Z(new_n1197));
  AOI21_X1  g772(.A(new_n1196), .B1(new_n1197), .B2(new_n1190), .ZN(new_n1198));
  INV_X1    g773(.A(new_n1198), .ZN(new_n1199));
  INV_X1    g774(.A(G1986), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n720), .A2(new_n1200), .ZN(new_n1201));
  XNOR2_X1  g776(.A(new_n1201), .B(KEYINPUT109), .ZN(new_n1202));
  INV_X1    g777(.A(new_n1202), .ZN(new_n1203));
  OAI21_X1  g778(.A(new_n1203), .B1(new_n1200), .B2(new_n720), .ZN(new_n1204));
  INV_X1    g779(.A(new_n1189), .ZN(new_n1205));
  AOI21_X1  g780(.A(new_n1199), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1188), .A2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1194), .A2(KEYINPUT46), .ZN(new_n1208));
  XNOR2_X1  g783(.A(new_n1208), .B(KEYINPUT127), .ZN(new_n1209));
  INV_X1    g784(.A(new_n1191), .ZN(new_n1210));
  OAI21_X1  g785(.A(new_n1190), .B1(new_n770), .B2(new_n1210), .ZN(new_n1211));
  OAI211_X1 g786(.A(new_n1209), .B(new_n1211), .C1(KEYINPUT46), .C2(new_n1194), .ZN(new_n1212));
  XOR2_X1   g787(.A(new_n1212), .B(KEYINPUT47), .Z(new_n1213));
  INV_X1    g788(.A(KEYINPUT48), .ZN(new_n1214));
  NOR3_X1   g789(.A1(new_n1203), .A2(new_n1214), .A3(new_n1189), .ZN(new_n1215));
  AOI21_X1  g790(.A(KEYINPUT48), .B1(new_n1202), .B2(new_n1205), .ZN(new_n1216));
  NOR3_X1   g791(.A1(new_n1215), .A2(new_n1199), .A3(new_n1216), .ZN(new_n1217));
  NAND2_X1  g792(.A1(new_n739), .A2(new_n741), .ZN(new_n1218));
  OAI22_X1  g793(.A1(new_n1196), .A2(new_n1218), .B1(G2067), .B2(new_n835), .ZN(new_n1219));
  AOI211_X1 g794(.A(new_n1213), .B(new_n1217), .C1(new_n1190), .C2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g795(.A1(new_n1207), .A2(new_n1220), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g796(.A1(G401), .A2(new_n462), .A3(G227), .ZN(new_n1223));
  AND3_X1   g797(.A1(new_n718), .A2(new_n900), .A3(new_n1223), .ZN(new_n1224));
  NAND2_X1  g798(.A1(new_n968), .A2(new_n1224), .ZN(G225));
  INV_X1    g799(.A(G225), .ZN(G308));
endmodule


