//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 1 0 0 0 1 0 1 0 1 1 1 0 1 0 1 1 1 1 0 1 1 0 1 0 1 0 0 0 1 1 1 1 1 1 1 0 0 1 0 0 1 0 0 0 0 1 0 1 0 0 1 1 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:22 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1247, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  INV_X1    g0003(.A(G97), .ZN(new_n204));
  INV_X1    g0004(.A(G107), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT64), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G68), .A2(G238), .B1(G107), .B2(G264), .ZN(new_n210));
  INV_X1    g0010(.A(G50), .ZN(new_n211));
  INV_X1    g0011(.A(G226), .ZN(new_n212));
  INV_X1    g0012(.A(G87), .ZN(new_n213));
  INV_X1    g0013(.A(G250), .ZN(new_n214));
  OAI221_X1 g0014(.A(new_n210), .B1(new_n211), .B2(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n216));
  INV_X1    g0016(.A(G58), .ZN(new_n217));
  INV_X1    g0017(.A(G232), .ZN(new_n218));
  INV_X1    g0018(.A(G257), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n204), .C2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n209), .B1(new_n215), .B2(new_n220), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(KEYINPUT1), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n209), .A2(G13), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n223), .B(G250), .C1(G257), .C2(G264), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT0), .Z(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  INV_X1    g0026(.A(G20), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(G50), .B1(G58), .B2(G68), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  AOI211_X1 g0030(.A(new_n222), .B(new_n225), .C1(new_n228), .C2(new_n230), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(new_n218), .ZN(new_n233));
  XOR2_X1   g0033(.A(KEYINPUT2), .B(G226), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n235), .B(new_n238), .Z(G358));
  XNOR2_X1  g0039(.A(G50), .B(G68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G58), .B(G77), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n240), .B(new_n241), .Z(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  INV_X1    g0046(.A(KEYINPUT21), .ZN(new_n247));
  INV_X1    g0047(.A(G1), .ZN(new_n248));
  NAND3_X1  g0048(.A1(new_n248), .A2(G13), .A3(G20), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n248), .A2(G33), .ZN(new_n250));
  NAND3_X1  g0050(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n251));
  NAND4_X1  g0051(.A1(new_n249), .A2(new_n250), .A3(new_n226), .A4(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(new_n249), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT79), .ZN(new_n255));
  INV_X1    g0055(.A(G116), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n254), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  OAI21_X1  g0057(.A(KEYINPUT79), .B1(new_n249), .B2(G116), .ZN(new_n258));
  AOI22_X1  g0058(.A1(new_n253), .A2(G116), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  AOI22_X1  g0059(.A1(new_n251), .A2(new_n226), .B1(G20), .B2(new_n256), .ZN(new_n260));
  NAND2_X1  g0060(.A1(G33), .A2(G283), .ZN(new_n261));
  OAI211_X1 g0061(.A(new_n261), .B(new_n227), .C1(G33), .C2(new_n204), .ZN(new_n262));
  AOI21_X1  g0062(.A(KEYINPUT20), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  AND3_X1   g0063(.A1(new_n260), .A2(KEYINPUT20), .A3(new_n262), .ZN(new_n264));
  OAI211_X1 g0064(.A(new_n259), .B(KEYINPUT80), .C1(new_n263), .C2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT80), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n264), .A2(new_n263), .ZN(new_n267));
  INV_X1    g0067(.A(new_n258), .ZN(new_n268));
  NOR3_X1   g0068(.A1(new_n249), .A2(KEYINPUT79), .A3(G116), .ZN(new_n269));
  OAI22_X1  g0069(.A1(new_n268), .A2(new_n269), .B1(new_n256), .B2(new_n252), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n266), .B1(new_n267), .B2(new_n270), .ZN(new_n271));
  AND2_X1   g0071(.A1(new_n265), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G41), .ZN(new_n273));
  OAI211_X1 g0073(.A(new_n248), .B(G45), .C1(new_n273), .C2(KEYINPUT5), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT74), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G45), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n277), .A2(G1), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT5), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(G41), .ZN(new_n280));
  AOI21_X1  g0080(.A(KEYINPUT74), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  OAI21_X1  g0081(.A(KEYINPUT75), .B1(new_n276), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n274), .A2(new_n275), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT75), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n278), .A2(KEYINPUT74), .A3(new_n280), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n283), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(G33), .A2(G41), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n287), .A2(G1), .A3(G13), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n273), .A2(KEYINPUT5), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n288), .A2(G274), .A3(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n282), .A2(new_n286), .A3(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n283), .A2(new_n285), .A3(new_n289), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n293), .A2(G270), .A3(new_n288), .ZN(new_n294));
  XNOR2_X1  g0094(.A(KEYINPUT3), .B(G33), .ZN(new_n295));
  NOR2_X1   g0095(.A1(G257), .A2(G1698), .ZN(new_n296));
  INV_X1    g0096(.A(G1698), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n297), .A2(G264), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n295), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n226), .B1(G33), .B2(G41), .ZN(new_n300));
  OAI211_X1 g0100(.A(new_n299), .B(new_n300), .C1(G303), .C2(new_n295), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n292), .A2(new_n294), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(G169), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n247), .B1(new_n272), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n302), .A2(G200), .ZN(new_n305));
  INV_X1    g0105(.A(G190), .ZN(new_n306));
  OAI211_X1 g0106(.A(new_n272), .B(new_n305), .C1(new_n306), .C2(new_n302), .ZN(new_n307));
  INV_X1    g0107(.A(G179), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n302), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n265), .A2(new_n271), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n310), .A2(KEYINPUT21), .A3(G169), .A4(new_n302), .ZN(new_n312));
  AND4_X1   g0112(.A1(new_n304), .A2(new_n307), .A3(new_n311), .A4(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n251), .A2(new_n226), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT65), .ZN(new_n315));
  INV_X1    g0115(.A(G33), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n315), .A2(new_n227), .A3(new_n316), .ZN(new_n317));
  OAI21_X1  g0117(.A(KEYINPUT65), .B1(G20), .B2(G33), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(G150), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  XNOR2_X1  g0122(.A(KEYINPUT8), .B(G58), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n227), .A2(G33), .ZN(new_n324));
  OAI22_X1  g0124(.A1(new_n323), .A2(new_n324), .B1(new_n227), .B2(new_n201), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n314), .B1(new_n322), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n248), .A2(G20), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(G50), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(new_n249), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n254), .A2(new_n314), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n329), .B1(new_n330), .B2(new_n211), .ZN(new_n331));
  AND2_X1   g0131(.A1(new_n331), .A2(KEYINPUT66), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n331), .A2(KEYINPUT66), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n326), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT9), .ZN(new_n335));
  AND2_X1   g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  OAI211_X1 g0136(.A(KEYINPUT9), .B(new_n326), .C1(new_n332), .C2(new_n333), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n295), .A2(G223), .A3(G1698), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n295), .A2(new_n297), .ZN(new_n339));
  INV_X1    g0139(.A(G222), .ZN(new_n340));
  OAI221_X1 g0140(.A(new_n338), .B1(new_n202), .B2(new_n295), .C1(new_n339), .C2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(new_n300), .ZN(new_n342));
  AOI21_X1  g0142(.A(G1), .B1(new_n273), .B2(new_n277), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n343), .A2(new_n288), .A3(G274), .ZN(new_n344));
  INV_X1    g0144(.A(new_n344), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n248), .B1(G41), .B2(G45), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n288), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n345), .B1(G226), .B2(new_n348), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n342), .A2(G190), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n337), .A2(new_n350), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n336), .A2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT10), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n342), .A2(new_n349), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(G200), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n352), .A2(new_n353), .A3(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT68), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n357), .B1(new_n336), .B2(new_n351), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n334), .A2(new_n335), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n359), .A2(KEYINPUT68), .A3(new_n337), .A4(new_n350), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n358), .A2(new_n360), .A3(new_n355), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT69), .ZN(new_n362));
  AND3_X1   g0162(.A1(new_n361), .A2(new_n362), .A3(KEYINPUT10), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n362), .B1(new_n361), .B2(KEYINPUT10), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n356), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n354), .A2(G179), .ZN(new_n366));
  XNOR2_X1  g0166(.A(new_n366), .B(KEYINPUT67), .ZN(new_n367));
  INV_X1    g0167(.A(new_n354), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n334), .B1(new_n368), .B2(G169), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n365), .A2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n318), .ZN(new_n373));
  NOR3_X1   g0173(.A1(KEYINPUT65), .A2(G20), .A3(G33), .ZN(new_n374));
  OAI21_X1  g0174(.A(G159), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT71), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n319), .A2(KEYINPUT71), .A3(G159), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  AND2_X1   g0179(.A1(KEYINPUT3), .A2(G33), .ZN(new_n380));
  NOR2_X1   g0180(.A1(KEYINPUT3), .A2(G33), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(KEYINPUT7), .B1(new_n382), .B2(new_n227), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT7), .ZN(new_n384));
  NOR4_X1   g0184(.A1(new_n380), .A2(new_n381), .A3(new_n384), .A4(G20), .ZN(new_n385));
  OAI21_X1  g0185(.A(G68), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(G68), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n217), .A2(new_n387), .ZN(new_n388));
  NOR2_X1   g0188(.A1(G58), .A2(G68), .ZN(new_n389));
  OAI21_X1  g0189(.A(G20), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n379), .A2(new_n386), .A3(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT16), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n379), .A2(new_n386), .A3(KEYINPUT16), .A4(new_n390), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n393), .A2(new_n314), .A3(new_n394), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n344), .B1(new_n347), .B2(new_n218), .ZN(new_n396));
  OAI211_X1 g0196(.A(G223), .B(new_n297), .C1(new_n380), .C2(new_n381), .ZN(new_n397));
  OAI211_X1 g0197(.A(G226), .B(G1698), .C1(new_n380), .C2(new_n381), .ZN(new_n398));
  OAI211_X1 g0198(.A(new_n397), .B(new_n398), .C1(new_n316), .C2(new_n213), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n396), .B1(new_n300), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(new_n306), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n401), .B1(G200), .B2(new_n400), .ZN(new_n402));
  INV_X1    g0202(.A(new_n323), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(new_n327), .ZN(new_n404));
  INV_X1    g0204(.A(new_n314), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(new_n249), .ZN(new_n406));
  OAI22_X1  g0206(.A1(new_n404), .A2(new_n406), .B1(new_n249), .B2(new_n403), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n395), .A2(new_n402), .A3(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT17), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n405), .B1(new_n391), .B2(new_n392), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n407), .B1(new_n412), .B2(new_n394), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n413), .A2(KEYINPUT17), .A3(new_n402), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n411), .A2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT18), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n399), .A2(new_n300), .ZN(new_n417));
  INV_X1    g0217(.A(new_n396), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n417), .A2(new_n418), .A3(new_n308), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n419), .B1(new_n400), .B2(G169), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n416), .B1(new_n413), .B2(new_n420), .ZN(new_n421));
  AOI211_X1 g0221(.A(new_n416), .B(new_n420), .C1(new_n395), .C2(new_n408), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n421), .B1(new_n422), .B2(KEYINPUT72), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n420), .B1(new_n395), .B2(new_n408), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT72), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n425), .A2(new_n426), .A3(new_n416), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n415), .B1(new_n423), .B2(new_n427), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n320), .A2(new_n211), .ZN(new_n429));
  OAI22_X1  g0229(.A1(new_n324), .A2(new_n202), .B1(new_n227), .B2(G68), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n314), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT11), .ZN(new_n432));
  AND2_X1   g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(KEYINPUT12), .B1(new_n249), .B2(G68), .ZN(new_n434));
  OR3_X1    g0234(.A1(new_n249), .A2(KEYINPUT12), .A3(G68), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n387), .B1(new_n248), .B2(G20), .ZN(new_n436));
  AOI22_X1  g0236(.A1(new_n434), .A2(new_n435), .B1(new_n330), .B2(new_n436), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n437), .B1(new_n431), .B2(new_n432), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n433), .A2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n295), .A2(G232), .A3(G1698), .ZN(new_n441));
  NAND2_X1  g0241(.A1(G33), .A2(G97), .ZN(new_n442));
  OAI211_X1 g0242(.A(new_n441), .B(new_n442), .C1(new_n339), .C2(new_n212), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(new_n300), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT13), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n345), .B1(G238), .B2(new_n348), .ZN(new_n446));
  AND3_X1   g0246(.A1(new_n444), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n445), .B1(new_n444), .B2(new_n446), .ZN(new_n448));
  OAI21_X1  g0248(.A(G169), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n444), .A2(new_n446), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(KEYINPUT13), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n444), .A2(new_n445), .A3(new_n446), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  OAI22_X1  g0253(.A1(new_n449), .A2(KEYINPUT14), .B1(new_n453), .B2(new_n308), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT14), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n455), .B1(new_n453), .B2(G169), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n440), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n451), .A2(G190), .A3(new_n452), .ZN(new_n458));
  AOI21_X1  g0258(.A(KEYINPUT70), .B1(new_n453), .B2(G200), .ZN(new_n459));
  OAI211_X1 g0259(.A(KEYINPUT70), .B(G200), .C1(new_n447), .C2(new_n448), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n439), .B(new_n458), .C1(new_n459), .C2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n327), .A2(G77), .ZN(new_n463));
  OAI22_X1  g0263(.A1(new_n406), .A2(new_n463), .B1(G77), .B2(new_n249), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n320), .A2(new_n323), .ZN(new_n465));
  XNOR2_X1  g0265(.A(KEYINPUT15), .B(G87), .ZN(new_n466));
  OAI22_X1  g0266(.A1(new_n466), .A2(new_n324), .B1(new_n227), .B2(new_n202), .ZN(new_n467));
  OR2_X1    g0267(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n464), .B1(new_n468), .B2(new_n314), .ZN(new_n469));
  INV_X1    g0269(.A(G169), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n295), .A2(G232), .A3(new_n297), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n295), .A2(G238), .A3(G1698), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n471), .B(new_n472), .C1(new_n205), .C2(new_n295), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(new_n300), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n345), .B1(G244), .B2(new_n348), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n469), .B1(new_n470), .B2(new_n476), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n477), .B1(G179), .B2(new_n476), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n476), .A2(G200), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n479), .B(new_n469), .C1(new_n306), .C2(new_n476), .ZN(new_n480));
  AND2_X1   g0280(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n428), .A2(new_n457), .A3(new_n462), .A4(new_n481), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n372), .A2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT82), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n214), .A2(new_n297), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n219), .A2(G1698), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n485), .B(new_n486), .C1(new_n380), .C2(new_n381), .ZN(new_n487));
  NAND2_X1  g0287(.A1(G33), .A2(G294), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT81), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n487), .A2(KEYINPUT81), .A3(new_n488), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n491), .A2(new_n300), .A3(new_n492), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n293), .A2(G264), .A3(new_n288), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n493), .A2(new_n292), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(G169), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n493), .A2(G179), .A3(new_n292), .A4(new_n494), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n484), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT25), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n499), .B1(new_n249), .B2(G107), .ZN(new_n500));
  NOR3_X1   g0300(.A1(new_n249), .A2(new_n499), .A3(G107), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  AOI22_X1  g0302(.A1(new_n500), .A2(new_n502), .B1(new_n253), .B2(G107), .ZN(new_n503));
  INV_X1    g0303(.A(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(G33), .A2(G116), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n505), .A2(G20), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT23), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n507), .B1(new_n227), .B2(G107), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n205), .A2(KEYINPUT23), .A3(G20), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n506), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT22), .ZN(new_n511));
  OR2_X1    g0311(.A1(KEYINPUT3), .A2(G33), .ZN(new_n512));
  NAND2_X1  g0312(.A1(KEYINPUT3), .A2(G33), .ZN(new_n513));
  AOI21_X1  g0313(.A(G20), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n511), .B1(new_n514), .B2(G87), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n227), .B(G87), .C1(new_n380), .C2(new_n381), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n516), .A2(KEYINPUT22), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n510), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(KEYINPUT24), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT24), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n520), .B(new_n510), .C1(new_n515), .C2(new_n517), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n504), .B1(new_n522), .B2(new_n314), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n498), .A2(new_n523), .ZN(new_n524));
  AND3_X1   g0324(.A1(new_n496), .A2(new_n484), .A3(new_n497), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(G200), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n495), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n493), .A2(new_n306), .A3(new_n292), .A4(new_n494), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  AOI22_X1  g0330(.A1(new_n524), .A2(new_n526), .B1(new_n523), .B2(new_n530), .ZN(new_n531));
  OAI211_X1 g0331(.A(G244), .B(new_n297), .C1(new_n380), .C2(new_n381), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT4), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(new_n261), .ZN(new_n535));
  NAND2_X1  g0335(.A1(G250), .A2(G1698), .ZN(new_n536));
  NAND2_X1  g0336(.A1(KEYINPUT4), .A2(G244), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n536), .B1(new_n537), .B2(G1698), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n535), .B1(new_n295), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n534), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n300), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n293), .A2(G257), .A3(new_n288), .ZN(new_n542));
  AND3_X1   g0342(.A1(new_n292), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  OAI21_X1  g0343(.A(KEYINPUT76), .B1(new_n543), .B2(new_n527), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n204), .A2(G107), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT6), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(KEYINPUT73), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT73), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(KEYINPUT6), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n545), .A2(new_n547), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(G97), .A2(G107), .ZN(new_n551));
  AND2_X1   g0351(.A1(new_n206), .A2(new_n551), .ZN(new_n552));
  XNOR2_X1  g0352(.A(KEYINPUT73), .B(KEYINPUT6), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n550), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  AOI22_X1  g0354(.A1(new_n554), .A2(G20), .B1(G77), .B2(new_n319), .ZN(new_n555));
  OAI21_X1  g0355(.A(G107), .B1(new_n383), .B2(new_n385), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n405), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n249), .A2(G97), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n558), .B1(new_n253), .B2(G97), .ZN(new_n559));
  INV_X1    g0359(.A(new_n559), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n292), .A2(new_n541), .A3(new_n542), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT76), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n562), .A2(new_n563), .A3(G200), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n543), .A2(G190), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n544), .A2(new_n561), .A3(new_n564), .A4(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(G274), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n278), .A2(new_n567), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n214), .B1(new_n277), .B2(G1), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n568), .A2(new_n288), .A3(new_n569), .ZN(new_n570));
  NOR2_X1   g0370(.A1(G238), .A2(G1698), .ZN(new_n571));
  INV_X1    g0371(.A(G244), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n571), .B1(new_n572), .B2(G1698), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n573), .A2(new_n295), .B1(G33), .B2(G116), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n308), .B(new_n570), .C1(new_n574), .C2(new_n288), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT77), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  OR2_X1    g0377(.A1(G238), .A2(G1698), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n572), .A2(G1698), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n578), .B(new_n579), .C1(new_n380), .C2(new_n381), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n288), .B1(new_n580), .B2(new_n505), .ZN(new_n581));
  AND3_X1   g0381(.A1(new_n568), .A2(new_n288), .A3(new_n569), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n583), .A2(KEYINPUT77), .A3(new_n308), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT19), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n227), .B1(new_n442), .B2(new_n585), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n586), .B1(G87), .B2(new_n206), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n227), .B(G68), .C1(new_n380), .C2(new_n381), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n585), .B1(new_n324), .B2(new_n204), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n314), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n466), .A2(new_n254), .ZN(new_n592));
  OR2_X1    g0392(.A1(new_n466), .A2(KEYINPUT78), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n466), .A2(KEYINPUT78), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n593), .A2(new_n253), .A3(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n591), .A2(new_n592), .A3(new_n595), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n570), .B1(new_n574), .B2(new_n288), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n470), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n577), .A2(new_n584), .A3(new_n596), .A4(new_n598), .ZN(new_n599));
  AOI22_X1  g0399(.A1(new_n590), .A2(new_n314), .B1(new_n254), .B2(new_n466), .ZN(new_n600));
  OAI21_X1  g0400(.A(G200), .B1(new_n581), .B2(new_n582), .ZN(new_n601));
  OAI211_X1 g0401(.A(G190), .B(new_n570), .C1(new_n574), .C2(new_n288), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n253), .A2(G87), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n600), .A2(new_n601), .A3(new_n602), .A4(new_n603), .ZN(new_n604));
  AND2_X1   g0404(.A1(new_n599), .A2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(new_n550), .ZN(new_n606));
  AOI22_X1  g0406(.A1(new_n547), .A2(new_n549), .B1(new_n206), .B2(new_n551), .ZN(new_n607));
  OAI21_X1  g0407(.A(G20), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n319), .A2(G77), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(new_n556), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n314), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n559), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n562), .A2(new_n470), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n292), .A2(new_n541), .A3(new_n308), .A4(new_n542), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n613), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  AND3_X1   g0416(.A1(new_n566), .A2(new_n605), .A3(new_n616), .ZN(new_n617));
  AND4_X1   g0417(.A1(new_n313), .A2(new_n483), .A3(new_n531), .A4(new_n617), .ZN(G372));
  INV_X1    g0418(.A(new_n422), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(new_n421), .ZN(new_n620));
  INV_X1    g0420(.A(new_n478), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n449), .A2(KEYINPUT14), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n453), .A2(new_n455), .A3(G169), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n447), .A2(new_n448), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(G179), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n622), .A2(new_n623), .A3(new_n625), .ZN(new_n626));
  AOI22_X1  g0426(.A1(new_n462), .A2(new_n621), .B1(new_n440), .B2(new_n626), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n620), .B1(new_n627), .B2(new_n415), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n370), .B1(new_n365), .B2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n483), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n596), .A2(new_n598), .A3(new_n575), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(new_n604), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n633), .B1(new_n530), .B2(new_n523), .ZN(new_n634));
  AND3_X1   g0434(.A1(new_n634), .A2(new_n616), .A3(new_n566), .ZN(new_n635));
  INV_X1    g0435(.A(new_n523), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n496), .A2(new_n497), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n638), .A2(new_n304), .A3(new_n311), .A4(new_n312), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n632), .B1(new_n635), .B2(new_n639), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n615), .B1(new_n557), .B2(new_n560), .ZN(new_n641));
  AND2_X1   g0441(.A1(new_n562), .A2(new_n470), .ZN(new_n642));
  OAI21_X1  g0442(.A(KEYINPUT83), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT83), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n613), .A2(new_n614), .A3(new_n644), .A4(new_n615), .ZN(new_n645));
  INV_X1    g0445(.A(new_n633), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n643), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT26), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n641), .A2(new_n642), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n650), .A2(new_n605), .A3(KEYINPUT26), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT84), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n599), .A2(new_n604), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n616), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n655), .A2(KEYINPUT84), .A3(KEYINPUT26), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n649), .A2(new_n653), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n640), .A2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n629), .B1(new_n630), .B2(new_n659), .ZN(G369));
  INV_X1    g0460(.A(G13), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n661), .A2(G1), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(new_n227), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(KEYINPUT85), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT27), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT85), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n662), .A2(new_n666), .A3(new_n227), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n664), .A2(new_n665), .A3(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(G213), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n665), .B1(new_n664), .B2(new_n667), .ZN(new_n670));
  OAI21_X1  g0470(.A(KEYINPUT86), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n670), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT86), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n672), .A2(new_n673), .A3(G213), .A4(new_n668), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(G343), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n313), .B1(new_n272), .B2(new_n677), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n304), .A2(new_n311), .A3(new_n312), .ZN(new_n679));
  INV_X1    g0479(.A(new_n677), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n679), .A2(new_n310), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  XOR2_X1   g0482(.A(new_n682), .B(KEYINPUT87), .Z(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(G330), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n531), .B1(new_n523), .B2(new_n677), .ZN(new_n686));
  NOR3_X1   g0486(.A1(new_n525), .A2(new_n498), .A3(new_n523), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(new_n680), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g0489(.A(new_n689), .B(KEYINPUT88), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n685), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n638), .A2(new_n680), .ZN(new_n692));
  AND2_X1   g0492(.A1(new_n679), .A2(new_n677), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n692), .B1(new_n690), .B2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n691), .A2(new_n694), .ZN(G399));
  INV_X1    g0495(.A(new_n223), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n696), .A2(G41), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NOR3_X1   g0498(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n698), .A2(G1), .A3(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n700), .B1(new_n229), .B2(new_n698), .ZN(new_n701));
  XNOR2_X1  g0501(.A(new_n701), .B(KEYINPUT89), .ZN(new_n702));
  XNOR2_X1  g0502(.A(new_n702), .B(KEYINPUT28), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT91), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n647), .A2(KEYINPUT26), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n632), .B1(new_n655), .B2(new_n648), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n687), .A2(new_n679), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n634), .A2(new_n566), .A3(new_n616), .ZN(new_n708));
  OAI211_X1 g0508(.A(new_n705), .B(new_n706), .C1(new_n707), .C2(new_n708), .ZN(new_n709));
  AND4_X1   g0509(.A1(new_n704), .A2(new_n709), .A3(KEYINPUT29), .A4(new_n677), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT29), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n711), .B1(new_n659), .B2(new_n680), .ZN(new_n712));
  AND2_X1   g0512(.A1(new_n705), .A2(new_n706), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n635), .B1(new_n679), .B2(new_n687), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n680), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n704), .B1(new_n715), .B2(KEYINPUT29), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n710), .B1(new_n712), .B2(new_n716), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n531), .A2(new_n313), .A3(new_n617), .A4(new_n677), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n302), .A2(new_n308), .A3(new_n597), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT90), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n302), .A2(KEYINPUT90), .A3(new_n308), .A4(new_n597), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n721), .A2(new_n495), .A3(new_n562), .A4(new_n722), .ZN(new_n723));
  AND3_X1   g0523(.A1(new_n493), .A2(new_n494), .A3(new_n583), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n309), .A2(new_n543), .A3(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT30), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n309), .A2(KEYINPUT30), .A3(new_n543), .A4(new_n724), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n723), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(new_n680), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT31), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n729), .A2(KEYINPUT31), .A3(new_n680), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n718), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(G330), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n717), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n703), .B1(new_n737), .B2(G1), .ZN(G364));
  NOR2_X1   g0538(.A1(new_n661), .A2(G20), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n248), .B1(new_n739), .B2(G45), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n697), .A2(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n685), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n683), .A2(G330), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(G13), .A2(G33), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(G20), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n678), .A2(new_n681), .A3(new_n748), .ZN(new_n749));
  XOR2_X1   g0549(.A(new_n742), .B(KEYINPUT92), .Z(new_n750));
  NOR2_X1   g0550(.A1(new_n696), .A2(new_n382), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(G355), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n752), .B1(G116), .B2(new_n223), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n696), .A2(new_n295), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n755), .B1(new_n277), .B2(new_n230), .ZN(new_n756));
  OR2_X1    g0556(.A1(new_n242), .A2(new_n277), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n753), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n226), .B1(G20), .B2(new_n470), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n748), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n750), .B1(new_n758), .B2(new_n761), .ZN(new_n762));
  XNOR2_X1  g0562(.A(new_n762), .B(KEYINPUT93), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n227), .A2(G179), .ZN(new_n764));
  NOR2_X1   g0564(.A1(G190), .A2(G200), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(G159), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g0568(.A(new_n768), .B(KEYINPUT32), .ZN(new_n769));
  NOR3_X1   g0569(.A1(new_n227), .A2(new_n308), .A3(KEYINPUT94), .ZN(new_n770));
  INV_X1    g0570(.A(KEYINPUT94), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n771), .B1(G20), .B2(G179), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n306), .A2(new_n527), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n769), .B1(new_n211), .B2(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n306), .A2(G200), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n774), .A2(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n527), .A2(G190), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n774), .A2(new_n780), .ZN(new_n781));
  OAI22_X1  g0581(.A1(new_n217), .A2(new_n779), .B1(new_n781), .B2(new_n387), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n775), .A2(new_n764), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n382), .B1(new_n784), .B2(G87), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n764), .A2(new_n780), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n778), .A2(new_n308), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(G20), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  OAI221_X1 g0589(.A(new_n785), .B1(new_n205), .B2(new_n786), .C1(new_n204), .C2(new_n789), .ZN(new_n790));
  NOR3_X1   g0590(.A1(new_n777), .A2(new_n782), .A3(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(KEYINPUT95), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n792), .B1(new_n774), .B2(new_n765), .ZN(new_n793));
  NOR4_X1   g0593(.A1(new_n773), .A2(KEYINPUT95), .A3(G190), .A4(G200), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n791), .B1(new_n202), .B2(new_n795), .ZN(new_n796));
  XOR2_X1   g0596(.A(new_n796), .B(KEYINPUT96), .Z(new_n797));
  INV_X1    g0597(.A(G311), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n795), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(G303), .ZN(new_n800));
  INV_X1    g0600(.A(G294), .ZN(new_n801));
  OAI221_X1 g0601(.A(new_n382), .B1(new_n783), .B2(new_n800), .C1(new_n789), .C2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n781), .ZN(new_n803));
  XNOR2_X1  g0603(.A(KEYINPUT33), .B(G317), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n802), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n779), .ZN(new_n806));
  INV_X1    g0606(.A(new_n776), .ZN(new_n807));
  AOI22_X1  g0607(.A1(G322), .A2(new_n806), .B1(new_n807), .B2(G326), .ZN(new_n808));
  INV_X1    g0608(.A(new_n786), .ZN(new_n809));
  INV_X1    g0609(.A(new_n766), .ZN(new_n810));
  AOI22_X1  g0610(.A1(new_n809), .A2(G283), .B1(new_n810), .B2(G329), .ZN(new_n811));
  XNOR2_X1  g0611(.A(new_n811), .B(KEYINPUT97), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n805), .A2(new_n808), .A3(new_n812), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n797), .B1(new_n799), .B2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(KEYINPUT98), .ZN(new_n815));
  OR2_X1    g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n759), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n817), .B1(new_n814), .B2(new_n815), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n763), .B1(new_n816), .B2(new_n818), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n743), .A2(new_n745), .B1(new_n749), .B2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(G396));
  NAND2_X1  g0621(.A1(new_n621), .A2(new_n677), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n480), .B1(new_n677), .B2(new_n469), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(new_n478), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n825), .B1(new_n659), .B2(new_n680), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n481), .A2(new_n677), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  AND3_X1   g0628(.A1(new_n649), .A2(new_n653), .A3(new_n656), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n523), .B1(new_n496), .B2(new_n497), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n679), .A2(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n631), .B1(new_n831), .B2(new_n708), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n828), .B1(new_n829), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n826), .A2(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n742), .B1(new_n834), .B2(new_n735), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n835), .B1(new_n735), .B2(new_n834), .ZN(new_n836));
  INV_X1    g0636(.A(new_n750), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n759), .A2(new_n746), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n837), .B1(new_n202), .B2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n825), .ZN(new_n840));
  AOI22_X1  g0640(.A1(G137), .A2(new_n807), .B1(new_n803), .B2(G150), .ZN(new_n841));
  XNOR2_X1  g0641(.A(new_n841), .B(KEYINPUT101), .ZN(new_n842));
  XOR2_X1   g0642(.A(KEYINPUT102), .B(G143), .Z(new_n843));
  OAI221_X1 g0643(.A(new_n842), .B1(new_n767), .B2(new_n795), .C1(new_n779), .C2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT34), .ZN(new_n845));
  OR2_X1    g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  AOI22_X1  g0646(.A1(G50), .A2(new_n784), .B1(new_n809), .B2(G68), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n382), .B1(new_n810), .B2(G132), .ZN(new_n848));
  OAI211_X1 g0648(.A(new_n847), .B(new_n848), .C1(new_n217), .C2(new_n789), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n849), .B1(new_n844), .B2(new_n845), .ZN(new_n850));
  AOI22_X1  g0650(.A1(G283), .A2(new_n803), .B1(new_n807), .B2(G303), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n851), .B1(new_n795), .B2(new_n256), .ZN(new_n852));
  XOR2_X1   g0652(.A(new_n852), .B(KEYINPUT99), .Z(new_n853));
  OAI22_X1  g0653(.A1(new_n779), .A2(new_n801), .B1(new_n204), .B2(new_n789), .ZN(new_n854));
  XNOR2_X1  g0654(.A(new_n854), .B(KEYINPUT100), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n382), .B1(new_n786), .B2(new_n213), .ZN(new_n856));
  OAI22_X1  g0656(.A1(new_n783), .A2(new_n205), .B1(new_n766), .B2(new_n798), .ZN(new_n857));
  NOR3_X1   g0657(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  AOI22_X1  g0658(.A1(new_n846), .A2(new_n850), .B1(new_n853), .B2(new_n858), .ZN(new_n859));
  OAI221_X1 g0659(.A(new_n839), .B1(new_n840), .B2(new_n747), .C1(new_n859), .C2(new_n817), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n836), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g0661(.A(new_n861), .B(KEYINPUT103), .ZN(G384));
  INV_X1    g0662(.A(KEYINPUT109), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT37), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n864), .A2(KEYINPUT106), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n865), .B1(new_n413), .B2(new_n402), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n395), .A2(new_n408), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n676), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n864), .A2(KEYINPUT106), .ZN(new_n869));
  NAND4_X1  g0669(.A1(new_n425), .A2(new_n866), .A3(new_n868), .A4(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n409), .ZN(new_n871));
  AOI22_X1  g0671(.A1(new_n395), .A2(new_n408), .B1(new_n675), .B2(new_n420), .ZN(new_n872));
  OAI211_X1 g0672(.A(KEYINPUT106), .B(new_n864), .C1(new_n871), .C2(new_n872), .ZN(new_n873));
  AND2_X1   g0673(.A1(new_n870), .A2(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n874), .B1(new_n428), .B2(new_n868), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT38), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  OAI211_X1 g0677(.A(new_n874), .B(KEYINPUT38), .C1(new_n428), .C2(new_n868), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n458), .A2(new_n439), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT70), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n881), .B1(new_n624), .B2(new_n527), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n880), .B1(new_n882), .B2(new_n460), .ZN(new_n883));
  OAI211_X1 g0683(.A(new_n440), .B(new_n680), .C1(new_n883), .C2(new_n626), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n680), .A2(new_n440), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n457), .A2(new_n462), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(KEYINPUT105), .B1(new_n833), .B2(new_n822), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n827), .B1(new_n640), .B2(new_n657), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT105), .ZN(new_n890));
  INV_X1    g0690(.A(new_n822), .ZN(new_n891));
  NOR3_X1   g0691(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n879), .B(new_n887), .C1(new_n888), .C2(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n619), .A2(new_n421), .A3(new_n675), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n626), .A2(new_n440), .A3(new_n677), .ZN(new_n896));
  INV_X1    g0696(.A(new_n415), .ZN(new_n897));
  AOI21_X1  g0697(.A(KEYINPUT72), .B1(new_n424), .B2(KEYINPUT18), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n424), .A2(KEYINPUT18), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NOR3_X1   g0700(.A1(new_n424), .A2(KEYINPUT72), .A3(KEYINPUT18), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n897), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n868), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(KEYINPUT38), .B1(new_n904), .B2(new_n874), .ZN(new_n905));
  INV_X1    g0705(.A(new_n878), .ZN(new_n906));
  OAI21_X1  g0706(.A(KEYINPUT39), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  XNOR2_X1  g0707(.A(KEYINPUT108), .B(KEYINPUT39), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n870), .A2(new_n873), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT107), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n415), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n411), .A2(KEYINPUT107), .A3(new_n414), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n911), .A2(new_n620), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n909), .B1(new_n913), .B2(new_n903), .ZN(new_n914));
  OAI211_X1 g0714(.A(new_n878), .B(new_n908), .C1(new_n914), .C2(KEYINPUT38), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n896), .B1(new_n907), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n863), .B1(new_n895), .B2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(new_n896), .ZN(new_n918));
  INV_X1    g0718(.A(new_n915), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT39), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n920), .B1(new_n877), .B2(new_n878), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n918), .B1(new_n919), .B2(new_n921), .ZN(new_n922));
  NAND4_X1  g0722(.A1(new_n922), .A2(KEYINPUT109), .A3(new_n893), .A4(new_n894), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n917), .A2(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n629), .B1(new_n717), .B2(new_n630), .ZN(new_n925));
  XOR2_X1   g0725(.A(new_n924), .B(new_n925), .Z(new_n926));
  INV_X1    g0726(.A(KEYINPUT40), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n905), .A2(new_n906), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n825), .B1(new_n884), .B2(new_n886), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n734), .A2(new_n929), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n927), .B1(new_n928), .B2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT110), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n878), .B1(new_n914), .B2(KEYINPUT38), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n734), .A2(new_n929), .A3(KEYINPUT110), .ZN(new_n935));
  NAND4_X1  g0735(.A1(new_n933), .A2(new_n934), .A3(KEYINPUT40), .A4(new_n935), .ZN(new_n936));
  AND2_X1   g0736(.A1(new_n931), .A2(new_n936), .ZN(new_n937));
  AND2_X1   g0737(.A1(new_n483), .A2(new_n734), .ZN(new_n938));
  OR2_X1    g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n937), .A2(new_n938), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n939), .A2(G330), .A3(new_n940), .ZN(new_n941));
  OAI22_X1  g0741(.A1(new_n926), .A2(new_n941), .B1(new_n248), .B2(new_n739), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT111), .ZN(new_n943));
  OR2_X1    g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n942), .A2(new_n943), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n926), .A2(new_n941), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  XOR2_X1   g0747(.A(new_n554), .B(KEYINPUT104), .Z(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT35), .ZN(new_n950));
  OAI211_X1 g0750(.A(G116), .B(new_n228), .C1(new_n949), .C2(new_n950), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n951), .B1(new_n950), .B2(new_n949), .ZN(new_n952));
  XOR2_X1   g0752(.A(new_n952), .B(KEYINPUT36), .Z(new_n953));
  NOR3_X1   g0753(.A1(new_n388), .A2(new_n229), .A3(new_n202), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n387), .A2(G50), .ZN(new_n955));
  OAI211_X1 g0755(.A(G1), .B(new_n661), .C1(new_n954), .C2(new_n955), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n947), .A2(new_n953), .A3(new_n956), .ZN(new_n957));
  XOR2_X1   g0757(.A(new_n957), .B(KEYINPUT112), .Z(G367));
  OAI211_X1 g0758(.A(new_n566), .B(new_n616), .C1(new_n561), .C2(new_n677), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n680), .A2(new_n650), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n690), .A2(new_n693), .A3(new_n961), .ZN(new_n962));
  OR2_X1    g0762(.A1(new_n962), .A2(KEYINPUT42), .ZN(new_n963));
  INV_X1    g0763(.A(new_n687), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n616), .B1(new_n964), .B2(new_n959), .ZN(new_n965));
  AOI22_X1  g0765(.A1(new_n962), .A2(KEYINPUT42), .B1(new_n677), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n963), .A2(new_n966), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n677), .B1(new_n600), .B2(new_n603), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n968), .A2(new_n633), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n969), .B1(new_n632), .B2(new_n968), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT43), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  OR2_X1    g0772(.A1(new_n970), .A2(new_n971), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n967), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  NAND4_X1  g0774(.A1(new_n963), .A2(new_n966), .A3(new_n971), .A4(new_n970), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(new_n961), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n691), .A2(new_n977), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n976), .B(new_n978), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n697), .B(KEYINPUT41), .Z(new_n980));
  INV_X1    g0780(.A(KEYINPUT45), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n690), .A2(new_n693), .ZN(new_n982));
  INV_X1    g0782(.A(new_n692), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n981), .B1(new_n984), .B2(new_n977), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n694), .A2(KEYINPUT45), .A3(new_n961), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n984), .A2(KEYINPUT44), .A3(new_n977), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT44), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n989), .B1(new_n694), .B2(new_n961), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n987), .A2(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(new_n691), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  OR2_X1    g0794(.A1(new_n690), .A2(new_n693), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n995), .A2(new_n982), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n996), .A2(new_n684), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n685), .A2(new_n995), .A3(new_n982), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n999), .A2(new_n736), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n987), .A2(new_n691), .A3(new_n991), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n994), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n980), .B1(new_n1002), .B2(new_n737), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n979), .B1(new_n1003), .B2(new_n741), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n970), .A2(new_n748), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n760), .B1(new_n223), .B2(new_n466), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1006), .B1(new_n754), .B2(new_n238), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n837), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(G283), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n795), .A2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n295), .B1(new_n809), .B2(G97), .ZN(new_n1011));
  INV_X1    g0811(.A(G317), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n1011), .B1(new_n1012), .B2(new_n766), .C1(new_n776), .C2(new_n798), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n784), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT46), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1015), .B1(new_n783), .B2(new_n256), .ZN(new_n1016));
  OAI211_X1 g0816(.A(new_n1014), .B(new_n1016), .C1(new_n205), .C2(new_n789), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n801), .A2(new_n781), .B1(new_n779), .B2(new_n800), .ZN(new_n1018));
  NOR4_X1   g0818(.A1(new_n1010), .A2(new_n1013), .A3(new_n1017), .A4(new_n1018), .ZN(new_n1019));
  XOR2_X1   g0819(.A(new_n1019), .B(KEYINPUT113), .Z(new_n1020));
  AOI22_X1  g0820(.A1(G58), .A2(new_n784), .B1(new_n810), .B2(G137), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n788), .A2(G68), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n809), .A2(G77), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n1021), .A2(new_n295), .A3(new_n1022), .A4(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n806), .A2(G150), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n1025), .B1(new_n767), .B2(new_n781), .C1(new_n776), .C2(new_n843), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n795), .ZN(new_n1027));
  AOI211_X1 g0827(.A(new_n1024), .B(new_n1026), .C1(G50), .C2(new_n1027), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n1020), .A2(new_n1028), .ZN(new_n1029));
  AND2_X1   g0829(.A1(new_n1029), .A2(KEYINPUT47), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n759), .B1(new_n1029), .B2(KEYINPUT47), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n1005), .B(new_n1008), .C1(new_n1030), .C2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1004), .A2(new_n1032), .ZN(G387));
  NOR2_X1   g0833(.A1(new_n999), .A2(new_n740), .ZN(new_n1034));
  XOR2_X1   g0834(.A(new_n1034), .B(KEYINPUT114), .Z(new_n1035));
  INV_X1    g0835(.A(new_n1000), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n999), .A2(new_n736), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1036), .A2(new_n697), .A3(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n403), .A2(new_n211), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1039), .B(KEYINPUT50), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n1040), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n699), .ZN(new_n1042));
  AOI211_X1 g0842(.A(G45), .B(new_n1042), .C1(G68), .C2(G77), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n755), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1044));
  OR2_X1    g0844(.A1(new_n1044), .A2(KEYINPUT115), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1044), .A2(KEYINPUT115), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n1045), .B(new_n1046), .C1(new_n277), .C2(new_n235), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n751), .A2(new_n1042), .B1(new_n205), .B2(new_n696), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1047), .A2(KEYINPUT116), .A3(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1049), .A2(new_n760), .ZN(new_n1050));
  AOI21_X1  g0850(.A(KEYINPUT116), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n750), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n767), .A2(new_n776), .B1(new_n781), .B2(new_n323), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1053), .B1(G50), .B2(new_n806), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n295), .B1(new_n786), .B2(new_n204), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n783), .A2(new_n202), .B1(new_n766), .B2(new_n321), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n593), .A2(new_n594), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n1057), .ZN(new_n1058));
  AOI211_X1 g0858(.A(new_n1055), .B(new_n1056), .C1(new_n1058), .C2(new_n788), .ZN(new_n1059));
  OAI211_X1 g0859(.A(new_n1054), .B(new_n1059), .C1(new_n387), .C2(new_n795), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n789), .A2(new_n1009), .B1(new_n783), .B2(new_n801), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n781), .A2(new_n798), .ZN(new_n1062));
  XOR2_X1   g0862(.A(KEYINPUT117), .B(G322), .Z(new_n1063));
  AOI21_X1  g0863(.A(new_n1062), .B1(new_n807), .B2(new_n1063), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n1064), .B1(new_n800), .B2(new_n795), .C1(new_n1012), .C2(new_n779), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT48), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1061), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1067), .B1(new_n1066), .B2(new_n1065), .ZN(new_n1068));
  XOR2_X1   g0868(.A(new_n1068), .B(KEYINPUT49), .Z(new_n1069));
  OAI21_X1  g0869(.A(new_n382), .B1(new_n786), .B2(new_n256), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(G326), .B2(new_n810), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT118), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1060), .B1(new_n1069), .B2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1052), .B1(new_n1073), .B2(new_n759), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n748), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1074), .B1(new_n690), .B2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1035), .A2(new_n1038), .A3(new_n1076), .ZN(G393));
  INV_X1    g0877(.A(new_n1001), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n691), .B1(new_n987), .B2(new_n991), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n977), .A2(new_n748), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n755), .A2(new_n245), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n760), .B1(new_n223), .B2(new_n204), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n750), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n798), .A2(new_n779), .B1(new_n776), .B2(new_n1012), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1085), .B(KEYINPUT52), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(G283), .A2(new_n784), .B1(new_n810), .B2(new_n1063), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n295), .B1(new_n809), .B2(G107), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n1087), .B(new_n1088), .C1(new_n256), .C2(new_n789), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1089), .B1(G303), .B2(new_n803), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n1086), .B(new_n1090), .C1(new_n801), .C2(new_n795), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n789), .A2(new_n202), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n382), .B1(new_n809), .B2(G87), .ZN(new_n1093));
  OAI221_X1 g0893(.A(new_n1093), .B1(new_n387), .B2(new_n783), .C1(new_n766), .C2(new_n843), .ZN(new_n1094));
  AOI211_X1 g0894(.A(new_n1092), .B(new_n1094), .C1(G50), .C2(new_n803), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1095), .B1(new_n323), .B2(new_n795), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n321), .A2(new_n776), .B1(new_n779), .B2(new_n767), .ZN(new_n1097));
  XOR2_X1   g0897(.A(new_n1097), .B(KEYINPUT51), .Z(new_n1098));
  OAI21_X1  g0898(.A(new_n1091), .B1(new_n1096), .B2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1084), .B1(new_n1099), .B2(new_n759), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(new_n1080), .A2(new_n741), .B1(new_n1081), .B2(new_n1100), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1036), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1102), .A2(new_n1002), .A3(new_n697), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1101), .A2(new_n1103), .ZN(G390));
  AOI21_X1  g0904(.A(new_n837), .B1(new_n323), .B2(new_n838), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n382), .B1(new_n810), .B2(G125), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1106), .B1(new_n211), .B2(new_n786), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(G128), .A2(new_n807), .B1(new_n806), .B2(G132), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT53), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1109), .B1(new_n783), .B2(new_n321), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n784), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n803), .A2(G137), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1108), .A2(new_n1112), .ZN(new_n1113));
  AOI211_X1 g0913(.A(new_n1107), .B(new_n1113), .C1(G159), .C2(new_n788), .ZN(new_n1114));
  XOR2_X1   g0914(.A(KEYINPUT54), .B(G143), .Z(new_n1115));
  NAND2_X1  g0915(.A1(new_n1027), .A2(new_n1115), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(G107), .A2(new_n803), .B1(new_n806), .B2(G116), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1117), .B1(new_n1009), .B2(new_n776), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n382), .B1(new_n783), .B2(new_n213), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n786), .A2(new_n387), .B1(new_n766), .B2(new_n801), .ZN(new_n1120));
  NOR4_X1   g0920(.A1(new_n1118), .A2(new_n1092), .A3(new_n1119), .A4(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1027), .A2(G97), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n1114), .A2(new_n1116), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n907), .A2(new_n915), .ZN(new_n1124));
  OAI221_X1 g0924(.A(new_n1105), .B1(new_n817), .B2(new_n1123), .C1(new_n1124), .C2(new_n747), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(new_n887), .B(KEYINPUT119), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n891), .B1(new_n715), .B2(new_n824), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n896), .B(new_n934), .C1(new_n1127), .C2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n833), .A2(KEYINPUT105), .A3(new_n822), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n890), .B1(new_n889), .B2(new_n891), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n918), .B1(new_n1132), .B2(new_n887), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1129), .B1(new_n1133), .B2(new_n1124), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n734), .A2(G330), .A3(new_n840), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1134), .A2(new_n887), .A3(new_n1136), .ZN(new_n1137));
  AND2_X1   g0937(.A1(new_n734), .A2(G330), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1138), .A2(new_n840), .A3(new_n887), .ZN(new_n1139));
  OAI211_X1 g0939(.A(new_n1129), .B(new_n1139), .C1(new_n1133), .C2(new_n1124), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1137), .A2(new_n1140), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1125), .B1(new_n1141), .B2(new_n740), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n887), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1135), .A2(KEYINPUT120), .A3(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1139), .A2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(KEYINPUT120), .B1(new_n1135), .B2(new_n1143), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1132), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n1139), .B(new_n1128), .C1(new_n1126), .C2(new_n1136), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n483), .A2(new_n1138), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n629), .B(new_n1150), .C1(new_n717), .C2(new_n630), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1149), .A2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n698), .B1(new_n1141), .B2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1151), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1137), .A2(new_n1155), .A3(new_n1140), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1142), .B1(new_n1154), .B2(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(G378));
  NAND2_X1  g0958(.A1(new_n1156), .A2(new_n1152), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n930), .B1(new_n877), .B2(new_n878), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n936), .B(G330), .C1(KEYINPUT40), .C2(new_n1160), .ZN(new_n1161));
  AND2_X1   g0961(.A1(new_n676), .A2(new_n334), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(new_n1162), .B(KEYINPUT121), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1163), .ZN(new_n1164));
  XOR2_X1   g0964(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  AND3_X1   g0966(.A1(new_n365), .A2(new_n371), .A3(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1166), .B1(new_n365), .B2(new_n371), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1164), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n372), .A2(new_n1165), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n365), .A2(new_n371), .A3(new_n1166), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1170), .A2(new_n1163), .A3(new_n1171), .ZN(new_n1172));
  AND2_X1   g0972(.A1(new_n1169), .A2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1161), .A2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1169), .A2(new_n1172), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n1175), .A2(new_n931), .A3(G330), .A4(new_n936), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n917), .A2(new_n1174), .A3(new_n923), .A4(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1174), .A2(new_n1176), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n924), .A2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1159), .A2(new_n1177), .A3(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT57), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n698), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1179), .A2(new_n1177), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1184), .A2(KEYINPUT57), .A3(new_n1159), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1182), .A2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1173), .A2(new_n746), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n838), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n742), .B1(G50), .B2(new_n1188), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(G33), .A2(G41), .ZN(new_n1190));
  AOI211_X1 g0990(.A(G50), .B(new_n1190), .C1(new_n382), .C2(new_n273), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n205), .A2(new_n779), .B1(new_n776), .B2(new_n256), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1192), .B1(G97), .B2(new_n803), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n786), .A2(new_n217), .B1(new_n766), .B2(new_n1009), .ZN(new_n1194));
  OAI211_X1 g0994(.A(new_n273), .B(new_n382), .C1(new_n783), .C2(new_n202), .ZN(new_n1195));
  AOI211_X1 g0995(.A(new_n1194), .B(new_n1195), .C1(G68), .C2(new_n788), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n1193), .B(new_n1196), .C1(new_n1057), .C2(new_n795), .ZN(new_n1197));
  INV_X1    g0997(.A(KEYINPUT58), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1191), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(G125), .A2(new_n807), .B1(new_n806), .B2(G128), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n803), .A2(G132), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(G150), .A2(new_n788), .B1(new_n784), .B2(new_n1115), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1200), .A2(new_n1201), .A3(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(G137), .B2(new_n1027), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1204), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n1205), .A2(KEYINPUT59), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1190), .B1(new_n786), .B2(new_n767), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1207), .B1(G124), .B2(new_n810), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT59), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1208), .B1(new_n1204), .B2(new_n1209), .ZN(new_n1210));
  OAI221_X1 g1010(.A(new_n1199), .B1(new_n1198), .B2(new_n1197), .C1(new_n1206), .C2(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1189), .B1(new_n1211), .B2(new_n759), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1187), .A2(new_n1212), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1213), .B1(new_n1183), .B2(new_n740), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1186), .A2(new_n1215), .ZN(G375));
  NAND2_X1  g1016(.A1(new_n1058), .A2(new_n788), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(G97), .A2(new_n784), .B1(new_n810), .B2(G303), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1217), .A2(new_n382), .A3(new_n1023), .A4(new_n1218), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(G116), .A2(new_n803), .B1(new_n807), .B2(G294), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1220), .B1(new_n1009), .B2(new_n779), .ZN(new_n1221));
  AOI211_X1 g1021(.A(new_n1219), .B(new_n1221), .C1(G107), .C2(new_n1027), .ZN(new_n1222));
  OAI221_X1 g1022(.A(new_n295), .B1(new_n786), .B2(new_n217), .C1(new_n789), .C2(new_n211), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1223), .B1(G132), .B2(new_n807), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(G159), .A2(new_n784), .B1(new_n810), .B2(G128), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1225), .A2(KEYINPUT122), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1226), .B1(G137), .B2(new_n806), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n803), .A2(new_n1115), .B1(new_n1225), .B2(KEYINPUT122), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1224), .A2(new_n1227), .A3(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1229), .B1(G150), .B2(new_n1027), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n759), .B1(new_n1222), .B2(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n837), .B1(new_n387), .B2(new_n838), .ZN(new_n1232));
  OAI211_X1 g1032(.A(new_n1231), .B(new_n1232), .C1(new_n1126), .C2(new_n747), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1149), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1233), .B1(new_n1234), .B2(new_n740), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1235), .ZN(new_n1236));
  OR2_X1    g1036(.A1(new_n1155), .A2(new_n980), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1234), .A2(new_n1151), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1236), .B1(new_n1237), .B2(new_n1239), .ZN(G381));
  NAND4_X1  g1040(.A1(new_n1035), .A2(new_n820), .A3(new_n1038), .A4(new_n1076), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1241), .A2(G384), .ZN(new_n1242));
  XOR2_X1   g1042(.A(new_n1242), .B(KEYINPUT123), .Z(new_n1243));
  NOR3_X1   g1043(.A1(G390), .A2(G378), .A3(G381), .ZN(new_n1244));
  NAND4_X1  g1044(.A1(new_n1243), .A2(new_n1004), .A3(new_n1032), .A4(new_n1244), .ZN(new_n1245));
  OR2_X1    g1045(.A1(new_n1245), .A2(G375), .ZN(G407));
  OR3_X1    g1046(.A1(G375), .A2(G343), .A3(G378), .ZN(new_n1247));
  OAI211_X1 g1047(.A(G213), .B(new_n1247), .C1(new_n1245), .C2(G375), .ZN(G409));
  INV_X1    g1048(.A(G213), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1249), .A2(G343), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1234), .A2(KEYINPUT60), .A3(new_n1151), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(new_n697), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1153), .A2(KEYINPUT60), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1253), .B1(new_n1238), .B2(new_n1254), .ZN(new_n1255));
  OR3_X1    g1055(.A1(new_n1255), .A2(G384), .A3(new_n1235), .ZN(new_n1256));
  OAI21_X1  g1056(.A(G384), .B1(new_n1255), .B2(new_n1235), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1180), .A2(new_n980), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1213), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n740), .B1(new_n1183), .B2(KEYINPUT124), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT124), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1179), .A2(new_n1262), .A3(new_n1177), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1260), .B1(new_n1261), .B2(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1259), .B1(new_n1264), .B2(KEYINPUT125), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1177), .ZN(new_n1266));
  AOI22_X1  g1066(.A1(new_n917), .A2(new_n923), .B1(new_n1174), .B2(new_n1176), .ZN(new_n1267));
  OAI21_X1  g1067(.A(KEYINPUT124), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1268), .A2(new_n741), .A3(new_n1263), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(new_n1213), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT125), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  AOI21_X1  g1072(.A(G378), .B1(new_n1265), .B2(new_n1272), .ZN(new_n1273));
  AOI211_X1 g1073(.A(new_n1157), .B(new_n1214), .C1(new_n1182), .C2(new_n1185), .ZN(new_n1274));
  OAI211_X1 g1074(.A(new_n1251), .B(new_n1258), .C1(new_n1273), .C2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1275), .A2(KEYINPUT62), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT61), .ZN(new_n1277));
  AND2_X1   g1077(.A1(new_n1250), .A2(G2897), .ZN(new_n1278));
  AND3_X1   g1078(.A1(new_n1256), .A2(new_n1257), .A3(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1278), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  OR2_X1    g1081(.A1(new_n1180), .A2(new_n980), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1269), .A2(KEYINPUT125), .A3(new_n1213), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1272), .A2(new_n1282), .A3(new_n1283), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1274), .B1(new_n1284), .B2(new_n1157), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1281), .B1(new_n1285), .B2(new_n1250), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1283), .A2(new_n1282), .ZN(new_n1287));
  AOI21_X1  g1087(.A(KEYINPUT125), .B1(new_n1269), .B2(new_n1213), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1157), .B1(new_n1287), .B2(new_n1288), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1186), .A2(G378), .A3(new_n1215), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT62), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1291), .A2(new_n1292), .A3(new_n1251), .A4(new_n1258), .ZN(new_n1293));
  NAND4_X1  g1093(.A1(new_n1276), .A2(new_n1277), .A3(new_n1286), .A4(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(G390), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(G387), .A2(new_n1295), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1004), .A2(new_n1032), .A3(G390), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(G393), .A2(G396), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1299), .A2(new_n1241), .ZN(new_n1300));
  AOI21_X1  g1100(.A(G390), .B1(new_n1004), .B2(new_n1032), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT127), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1300), .B1(new_n1301), .B2(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1298), .A2(new_n1303), .ZN(new_n1304));
  NAND4_X1  g1104(.A1(new_n1296), .A2(new_n1300), .A3(new_n1302), .A4(new_n1297), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1294), .A2(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1291), .A2(new_n1251), .ZN(new_n1309));
  AOI21_X1  g1109(.A(KEYINPUT61), .B1(new_n1309), .B2(new_n1281), .ZN(new_n1310));
  XOR2_X1   g1110(.A(KEYINPUT126), .B(KEYINPUT63), .Z(new_n1311));
  NAND2_X1  g1111(.A1(new_n1275), .A2(new_n1311), .ZN(new_n1312));
  NAND4_X1  g1112(.A1(new_n1291), .A2(KEYINPUT63), .A3(new_n1251), .A4(new_n1258), .ZN(new_n1313));
  NAND4_X1  g1113(.A1(new_n1310), .A2(new_n1306), .A3(new_n1312), .A4(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1308), .A2(new_n1314), .ZN(G405));
  NAND2_X1  g1115(.A1(G375), .A2(new_n1157), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1316), .A2(new_n1290), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1304), .A2(new_n1258), .A3(new_n1305), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1318), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1258), .B1(new_n1304), .B2(new_n1305), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n1317), .B1(new_n1319), .B2(new_n1320), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1258), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1306), .A2(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1317), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1323), .A2(new_n1324), .A3(new_n1318), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1321), .A2(new_n1325), .ZN(G402));
endmodule


