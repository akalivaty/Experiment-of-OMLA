//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 1 1 0 0 0 1 0 1 0 0 1 0 0 0 0 1 0 0 1 1 0 0 0 0 0 0 0 1 0 0 1 0 0 1 0 1 0 1 0 0 1 1 1 1 1 0 0 0 1 0 0 0 0 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:54 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1264, new_n1265, new_n1266, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(new_n201), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G50), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT66), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G1), .A2(G13), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  XOR2_X1   g0011(.A(new_n211), .B(KEYINPUT65), .Z(new_n212));
  NAND2_X1  g0012(.A1(new_n208), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(KEYINPUT0), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G20), .ZN(new_n215));
  OR3_X1    g0015(.A1(new_n215), .A2(KEYINPUT64), .A3(G13), .ZN(new_n216));
  OAI21_X1  g0016(.A(KEYINPUT64), .B1(new_n215), .B2(G13), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  OAI211_X1 g0018(.A(new_n218), .B(G250), .C1(G257), .C2(G264), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n213), .B1(new_n214), .B2(new_n219), .ZN(new_n220));
  AOI21_X1  g0020(.A(new_n220), .B1(new_n214), .B2(new_n219), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(KEYINPUT67), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n223));
  INV_X1    g0023(.A(G68), .ZN(new_n224));
  INV_X1    g0024(.A(G238), .ZN(new_n225));
  INV_X1    g0025(.A(G87), .ZN(new_n226));
  INV_X1    g0026(.A(G250), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n223), .B1(new_n224), .B2(new_n225), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n229));
  INV_X1    g0029(.A(G77), .ZN(new_n230));
  INV_X1    g0030(.A(G244), .ZN(new_n231));
  INV_X1    g0031(.A(G107), .ZN(new_n232));
  INV_X1    g0032(.A(G264), .ZN(new_n233));
  OAI221_X1 g0033(.A(new_n229), .B1(new_n230), .B2(new_n231), .C1(new_n232), .C2(new_n233), .ZN(new_n234));
  OAI21_X1  g0034(.A(new_n215), .B1(new_n228), .B2(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT1), .ZN(new_n236));
  NOR2_X1   g0036(.A1(new_n222), .A2(new_n236), .ZN(G361));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT2), .B(G226), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G264), .B(G270), .Z(new_n242));
  XNOR2_X1  g0042(.A(G250), .B(G257), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G358));
  XNOR2_X1  g0045(.A(G50), .B(G68), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G58), .B(G77), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n246), .B(new_n247), .Z(new_n248));
  XOR2_X1   g0048(.A(G87), .B(G97), .Z(new_n249));
  XNOR2_X1  g0049(.A(G107), .B(G116), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G351));
  NAND3_X1  g0052(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT69), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n253), .A2(new_n254), .A3(new_n209), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n254), .B1(new_n253), .B2(new_n209), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT71), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT8), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n259), .A2(new_n260), .A3(G58), .ZN(new_n261));
  INV_X1    g0061(.A(G58), .ZN(new_n262));
  NOR3_X1   g0062(.A1(new_n262), .A2(KEYINPUT70), .A3(KEYINPUT71), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT70), .ZN(new_n264));
  OAI21_X1  g0064(.A(KEYINPUT8), .B1(new_n264), .B2(G58), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n261), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT72), .ZN(new_n267));
  INV_X1    g0067(.A(G33), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n267), .B1(new_n268), .B2(G20), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n210), .A2(KEYINPUT72), .A3(G33), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n266), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  NOR2_X1   g0071(.A1(G20), .A2(G33), .ZN(new_n272));
  AOI22_X1  g0072(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n258), .B1(new_n271), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n253), .A2(new_n209), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(KEYINPUT69), .ZN(new_n276));
  INV_X1    g0076(.A(G13), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n277), .A2(G1), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G20), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n276), .A2(new_n255), .A3(new_n279), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n210), .A2(G1), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G50), .ZN(new_n283));
  AOI22_X1  g0083(.A1(new_n280), .A2(G50), .B1(new_n279), .B2(new_n283), .ZN(new_n284));
  OAI21_X1  g0084(.A(KEYINPUT9), .B1(new_n274), .B2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(new_n258), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n269), .A2(new_n270), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n264), .A2(new_n259), .A3(G58), .ZN(new_n288));
  OAI211_X1 g0088(.A(new_n288), .B(KEYINPUT8), .C1(new_n264), .C2(G58), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n287), .B1(new_n289), .B2(new_n261), .ZN(new_n290));
  INV_X1    g0090(.A(new_n273), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n286), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n283), .A2(new_n279), .ZN(new_n293));
  NOR3_X1   g0093(.A1(new_n277), .A2(new_n210), .A3(G1), .ZN(new_n294));
  NOR3_X1   g0094(.A1(new_n256), .A2(new_n257), .A3(new_n294), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n293), .B1(new_n295), .B2(new_n202), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT9), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n292), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n285), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT68), .ZN(new_n300));
  AND2_X1   g0100(.A1(G33), .A2(G41), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n300), .B1(new_n301), .B2(new_n209), .ZN(new_n302));
  NAND2_X1  g0102(.A1(G33), .A2(G41), .ZN(new_n303));
  NAND4_X1  g0103(.A1(new_n303), .A2(KEYINPUT68), .A3(G1), .A4(G13), .ZN(new_n304));
  AND3_X1   g0104(.A1(new_n302), .A2(G274), .A3(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(G41), .ZN(new_n306));
  INV_X1    g0106(.A(G45), .ZN(new_n307));
  AOI21_X1  g0107(.A(G1), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  XNOR2_X1  g0108(.A(KEYINPUT3), .B(G33), .ZN(new_n309));
  NOR2_X1   g0109(.A1(G222), .A2(G1698), .ZN(new_n310));
  INV_X1    g0110(.A(G1698), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n311), .A2(G223), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n309), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n303), .A2(G1), .A3(G13), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT3), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(G33), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n268), .A2(KEYINPUT3), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n314), .B1(new_n318), .B2(new_n230), .ZN(new_n319));
  AOI22_X1  g0119(.A1(new_n305), .A2(new_n308), .B1(new_n313), .B2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n308), .ZN(new_n321));
  NAND4_X1  g0121(.A1(new_n321), .A2(new_n302), .A3(G226), .A4(new_n304), .ZN(new_n322));
  NAND4_X1  g0122(.A1(new_n320), .A2(KEYINPUT74), .A3(G190), .A4(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n319), .A2(new_n313), .ZN(new_n324));
  NAND4_X1  g0124(.A1(new_n302), .A2(G274), .A3(new_n308), .A4(new_n304), .ZN(new_n325));
  NAND4_X1  g0125(.A1(new_n324), .A2(G190), .A3(new_n322), .A4(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT74), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n323), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n299), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n320), .A2(new_n322), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(G200), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  NOR3_X1   g0133(.A1(new_n330), .A2(KEYINPUT10), .A3(new_n333), .ZN(new_n334));
  AOI22_X1  g0134(.A1(new_n285), .A2(new_n298), .B1(new_n323), .B2(new_n328), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT75), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n332), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  AND3_X1   g0137(.A1(new_n299), .A2(new_n336), .A3(new_n329), .ZN(new_n338));
  OAI21_X1  g0138(.A(KEYINPUT10), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT76), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n330), .A2(KEYINPUT75), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n335), .A2(new_n336), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n342), .A2(new_n343), .A3(new_n332), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n344), .A2(KEYINPUT76), .A3(KEYINPUT10), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n334), .B1(new_n341), .B2(new_n345), .ZN(new_n346));
  XNOR2_X1  g0146(.A(KEYINPUT15), .B(G87), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n287), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(KEYINPUT73), .ZN(new_n349));
  XOR2_X1   g0149(.A(KEYINPUT8), .B(G58), .Z(new_n350));
  AOI22_X1  g0150(.A1(new_n350), .A2(new_n272), .B1(G20), .B2(G77), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n348), .A2(KEYINPUT73), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n275), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n294), .A2(new_n275), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n281), .A2(new_n230), .ZN(new_n356));
  AOI22_X1  g0156(.A1(new_n355), .A2(new_n356), .B1(new_n230), .B2(new_n294), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n354), .A2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  AND2_X1   g0159(.A1(new_n302), .A2(new_n304), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n360), .A2(G244), .A3(new_n321), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n314), .B1(new_n318), .B2(new_n232), .ZN(new_n362));
  NOR2_X1   g0162(.A1(G232), .A2(G1698), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n363), .B1(new_n225), .B2(G1698), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n362), .B1(new_n318), .B2(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n361), .A2(new_n325), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(G200), .ZN(new_n367));
  INV_X1    g0167(.A(G190), .ZN(new_n368));
  OAI211_X1 g0168(.A(new_n359), .B(new_n367), .C1(new_n368), .C2(new_n366), .ZN(new_n369));
  INV_X1    g0169(.A(G169), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n331), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n292), .A2(new_n296), .ZN(new_n372));
  OAI211_X1 g0172(.A(new_n371), .B(new_n372), .C1(G179), .C2(new_n331), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n366), .A2(new_n370), .ZN(new_n374));
  OAI211_X1 g0174(.A(new_n358), .B(new_n374), .C1(G179), .C2(new_n366), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n369), .A2(new_n373), .A3(new_n375), .ZN(new_n376));
  OAI21_X1  g0176(.A(KEYINPUT77), .B1(new_n346), .B2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n334), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT10), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n333), .B1(new_n330), .B2(KEYINPUT75), .ZN(new_n380));
  AOI211_X1 g0180(.A(new_n340), .B(new_n379), .C1(new_n380), .C2(new_n343), .ZN(new_n381));
  AOI21_X1  g0181(.A(KEYINPUT76), .B1(new_n344), .B2(KEYINPUT10), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n378), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT77), .ZN(new_n384));
  INV_X1    g0184(.A(new_n376), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n383), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n377), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n309), .A2(G226), .A3(new_n311), .ZN(new_n388));
  NAND2_X1  g0188(.A1(G33), .A2(G97), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n309), .A2(G1698), .ZN(new_n390));
  INV_X1    g0190(.A(G232), .ZN(new_n391));
  OAI211_X1 g0191(.A(new_n388), .B(new_n389), .C1(new_n390), .C2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n314), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n392), .A2(KEYINPUT78), .A3(new_n393), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n321), .A2(new_n302), .A3(G238), .A4(new_n304), .ZN(new_n395));
  AND2_X1   g0195(.A1(new_n395), .A2(new_n325), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(KEYINPUT78), .B1(new_n392), .B2(new_n393), .ZN(new_n398));
  OAI21_X1  g0198(.A(KEYINPUT13), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n392), .A2(new_n393), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT78), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT13), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n402), .A2(new_n403), .A3(new_n394), .A4(new_n396), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n399), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(G169), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(KEYINPUT14), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n399), .A2(G179), .A3(new_n404), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT14), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n405), .A2(new_n409), .A3(G169), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n407), .A2(new_n408), .A3(new_n410), .ZN(new_n411));
  OR3_X1    g0211(.A1(new_n279), .A2(KEYINPUT12), .A3(G68), .ZN(new_n412));
  OAI21_X1  g0212(.A(KEYINPUT12), .B1(new_n279), .B2(G68), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n281), .A2(new_n224), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n412), .A2(new_n413), .B1(new_n355), .B2(new_n414), .ZN(new_n415));
  AOI22_X1  g0215(.A1(new_n272), .A2(G50), .B1(G20), .B2(new_n224), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n416), .B1(new_n287), .B2(new_n230), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n286), .A2(KEYINPUT11), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n415), .A2(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(KEYINPUT11), .B1(new_n286), .B2(new_n417), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n411), .A2(new_n422), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n421), .B1(new_n405), .B2(new_n368), .ZN(new_n424));
  INV_X1    g0224(.A(G200), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n425), .B1(new_n399), .B2(new_n404), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n423), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n266), .A2(new_n282), .ZN(new_n430));
  OAI22_X1  g0230(.A1(new_n430), .A2(new_n280), .B1(new_n266), .B2(new_n279), .ZN(new_n431));
  XNOR2_X1  g0231(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n432));
  XNOR2_X1  g0232(.A(KEYINPUT70), .B(G58), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n206), .B1(new_n433), .B2(new_n224), .ZN(new_n434));
  AOI22_X1  g0234(.A1(new_n434), .A2(G20), .B1(G159), .B2(new_n272), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT82), .ZN(new_n436));
  AOI21_X1  g0236(.A(G20), .B1(new_n316), .B2(new_n317), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n436), .B1(new_n437), .B2(KEYINPUT7), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT7), .ZN(new_n439));
  OAI211_X1 g0239(.A(KEYINPUT82), .B(new_n439), .C1(new_n309), .C2(G20), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  XNOR2_X1  g0241(.A(KEYINPUT79), .B(G33), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n317), .B1(new_n442), .B2(KEYINPUT3), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n439), .A2(G20), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n224), .B1(new_n441), .B2(new_n445), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n435), .B1(new_n446), .B2(KEYINPUT83), .ZN(new_n447));
  AOI22_X1  g0247(.A1(new_n438), .A2(new_n440), .B1(new_n443), .B2(new_n444), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT83), .ZN(new_n449));
  NOR3_X1   g0249(.A1(new_n448), .A2(new_n449), .A3(new_n224), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n432), .B1(new_n447), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n268), .A2(KEYINPUT79), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT79), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(G33), .ZN(new_n454));
  AND3_X1   g0254(.A1(new_n452), .A2(new_n454), .A3(KEYINPUT3), .ZN(new_n455));
  OAI21_X1  g0255(.A(KEYINPUT80), .B1(new_n268), .B2(KEYINPUT3), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT80), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n457), .A2(new_n315), .A3(G33), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n439), .B(new_n210), .C1(new_n455), .C2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(G68), .ZN(new_n461));
  AND2_X1   g0261(.A1(new_n456), .A2(new_n458), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n452), .A2(new_n454), .A3(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n439), .B1(new_n464), .B2(new_n210), .ZN(new_n465));
  OAI211_X1 g0265(.A(KEYINPUT16), .B(new_n435), .C1(new_n461), .C2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(new_n275), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n431), .B1(new_n451), .B2(new_n468), .ZN(new_n469));
  MUX2_X1   g0269(.A(G223), .B(G226), .S(G1698), .Z(new_n470));
  NAND3_X1  g0270(.A1(new_n462), .A2(new_n463), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(G33), .A2(G87), .ZN(new_n472));
  XOR2_X1   g0272(.A(new_n472), .B(KEYINPUT84), .Z(new_n473));
  NAND2_X1  g0273(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(new_n393), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n321), .A2(new_n302), .A3(G232), .A4(new_n304), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(new_n325), .ZN(new_n477));
  INV_X1    g0277(.A(new_n477), .ZN(new_n478));
  AOI21_X1  g0278(.A(G169), .B1(new_n475), .B2(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n314), .B1(new_n471), .B2(new_n473), .ZN(new_n480));
  NOR3_X1   g0280(.A1(new_n480), .A2(G179), .A3(new_n477), .ZN(new_n481));
  OAI21_X1  g0281(.A(KEYINPUT85), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT85), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n370), .B1(new_n480), .B2(new_n477), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n475), .A2(new_n478), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n483), .B(new_n484), .C1(new_n485), .C2(G179), .ZN(new_n486));
  AND2_X1   g0286(.A1(new_n482), .A2(new_n486), .ZN(new_n487));
  OAI21_X1  g0287(.A(KEYINPUT18), .B1(new_n469), .B2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT18), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n482), .A2(new_n486), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n446), .A2(KEYINPUT83), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n449), .B1(new_n448), .B2(new_n224), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n491), .A2(new_n492), .A3(new_n435), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n467), .B1(new_n493), .B2(new_n432), .ZN(new_n494));
  OAI211_X1 g0294(.A(new_n489), .B(new_n490), .C1(new_n494), .C2(new_n431), .ZN(new_n495));
  AND2_X1   g0295(.A1(new_n488), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n451), .A2(new_n468), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n485), .A2(new_n425), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n498), .B1(G190), .B2(new_n485), .ZN(new_n499));
  INV_X1    g0299(.A(new_n431), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n497), .A2(KEYINPUT86), .A3(new_n499), .A4(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT17), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n469), .A2(KEYINPUT86), .A3(KEYINPUT17), .A4(new_n499), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n496), .A2(KEYINPUT87), .A3(new_n503), .A4(new_n504), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n503), .A2(new_n504), .A3(new_n488), .A4(new_n495), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT87), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n429), .B1(new_n505), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n387), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(KEYINPUT88), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT88), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n387), .A2(new_n509), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n302), .A2(G274), .A3(new_n304), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n307), .A2(G1), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT5), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(G41), .ZN(new_n518));
  AND3_X1   g0318(.A1(new_n306), .A2(KEYINPUT90), .A3(KEYINPUT5), .ZN(new_n519));
  AOI21_X1  g0319(.A(KEYINPUT90), .B1(new_n306), .B2(KEYINPUT5), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n516), .B(new_n518), .C1(new_n519), .C2(new_n520), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n515), .A2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n306), .A2(KEYINPUT5), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n516), .A2(new_n518), .A3(new_n524), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n360), .A2(G257), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n523), .A2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT4), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n311), .A2(G244), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n528), .B1(new_n464), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n528), .A2(new_n231), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n309), .A2(new_n311), .A3(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT89), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n309), .A2(KEYINPUT89), .A3(new_n311), .A4(new_n531), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(G33), .A2(G283), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n537), .B1(new_n390), .B2(new_n227), .ZN(new_n538));
  INV_X1    g0338(.A(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n530), .A2(new_n536), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n527), .B1(new_n540), .B2(new_n393), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(G190), .ZN(new_n542));
  INV_X1    g0342(.A(G97), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n294), .A2(new_n543), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n295), .B1(G1), .B2(new_n268), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n544), .B1(new_n545), .B2(new_n543), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n232), .A2(KEYINPUT6), .A3(G97), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n543), .A2(new_n232), .ZN(new_n548));
  NOR2_X1   g0348(.A1(G97), .A2(G107), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n547), .B1(new_n550), .B2(KEYINPUT6), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n551), .A2(G20), .B1(G77), .B2(new_n272), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n552), .B1(new_n448), .B2(new_n232), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n546), .B1(new_n553), .B2(new_n275), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n542), .B(new_n554), .C1(new_n425), .C2(new_n541), .ZN(new_n555));
  INV_X1    g0355(.A(new_n554), .ZN(new_n556));
  INV_X1    g0356(.A(G179), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n541), .A2(new_n557), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n538), .B1(new_n534), .B2(new_n535), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n314), .B1(new_n559), .B2(new_n530), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n370), .B1(new_n560), .B2(new_n527), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n556), .A2(new_n558), .A3(new_n561), .ZN(new_n562));
  AND2_X1   g0362(.A1(new_n555), .A2(new_n562), .ZN(new_n563));
  XOR2_X1   g0363(.A(new_n347), .B(KEYINPUT92), .Z(new_n564));
  OR2_X1    g0364(.A1(new_n545), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n347), .A2(new_n294), .ZN(new_n566));
  XNOR2_X1  g0366(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n210), .B1(new_n567), .B2(new_n389), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n549), .A2(new_n226), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n567), .B1(new_n287), .B2(new_n543), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n462), .A2(new_n210), .A3(new_n463), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n570), .B(new_n571), .C1(new_n572), .C2(new_n224), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(new_n275), .ZN(new_n574));
  AND3_X1   g0374(.A1(new_n565), .A2(new_n566), .A3(new_n574), .ZN(new_n575));
  NOR2_X1   g0375(.A1(G238), .A2(G1698), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n576), .B1(new_n231), .B2(G1698), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n462), .A2(new_n463), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n452), .A2(new_n454), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(G116), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n314), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n302), .A2(new_n304), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n516), .A2(G250), .ZN(new_n583));
  NOR3_X1   g0383(.A1(new_n307), .A2(G1), .A3(G274), .ZN(new_n584));
  NOR3_X1   g0384(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n581), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(new_n557), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n587), .B1(G169), .B2(new_n586), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n586), .A2(G190), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n589), .B1(new_n425), .B2(new_n586), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n574), .B(new_n566), .C1(new_n226), .C2(new_n545), .ZN(new_n591));
  OAI22_X1  g0391(.A1(new_n575), .A2(new_n588), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n227), .A2(new_n311), .ZN(new_n593));
  OR2_X1    g0393(.A1(new_n311), .A2(G257), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n462), .A2(new_n463), .A3(new_n593), .A4(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n579), .A2(G294), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n393), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT95), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n360), .A2(G264), .A3(new_n525), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n314), .B1(new_n595), .B2(new_n596), .ZN(new_n602));
  INV_X1    g0402(.A(new_n600), .ZN(new_n603));
  OAI21_X1  g0403(.A(KEYINPUT95), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n601), .A2(new_n604), .A3(new_n523), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(new_n425), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n598), .A2(new_n368), .A3(new_n523), .A4(new_n600), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n279), .A2(G107), .ZN(new_n609));
  XNOR2_X1  g0409(.A(new_n609), .B(KEYINPUT25), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n610), .B1(new_n545), .B2(new_n232), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(KEYINPUT94), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT94), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n610), .B(new_n613), .C1(new_n545), .C2(new_n232), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n309), .A2(new_n210), .A3(G87), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT22), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT23), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n618), .B1(new_n210), .B2(G107), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n232), .A2(KEYINPUT23), .A3(G20), .ZN(new_n620));
  AOI22_X1  g0420(.A1(new_n616), .A2(new_n617), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  OAI21_X1  g0421(.A(KEYINPUT93), .B1(new_n580), .B2(G20), .ZN(new_n622));
  AND2_X1   g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(KEYINPUT22), .A2(G87), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n572), .A2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(G116), .ZN(new_n627));
  OR4_X1    g0427(.A1(KEYINPUT93), .A2(new_n442), .A3(G20), .A4(new_n627), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n623), .A2(new_n626), .A3(KEYINPUT24), .A4(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT24), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n628), .A2(new_n622), .A3(new_n621), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n630), .B1(new_n631), .B2(new_n625), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n629), .A2(new_n632), .A3(new_n275), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n615), .A2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n592), .B1(new_n608), .B2(new_n635), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n601), .A2(new_n604), .A3(G179), .A4(new_n523), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n598), .A2(new_n523), .A3(new_n600), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(G169), .ZN(new_n639));
  AOI22_X1  g0439(.A1(new_n615), .A2(new_n633), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  NOR2_X1   g0440(.A1(G257), .A2(G1698), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n641), .B1(new_n233), .B2(G1698), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n462), .A2(new_n463), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n318), .A2(G303), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n314), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n525), .A2(new_n302), .A3(G270), .A4(new_n304), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n646), .B1(new_n521), .B2(new_n515), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(G190), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n210), .A2(G116), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n278), .A2(new_n650), .ZN(new_n651));
  OAI211_X1 g0451(.A(new_n355), .B(G116), .C1(G1), .C2(new_n268), .ZN(new_n652));
  OAI211_X1 g0452(.A(new_n537), .B(new_n210), .C1(G33), .C2(new_n543), .ZN(new_n653));
  INV_X1    g0453(.A(new_n650), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n653), .A2(new_n654), .A3(new_n275), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT20), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n655), .A2(new_n656), .ZN(new_n658));
  OAI211_X1 g0458(.A(new_n651), .B(new_n652), .C1(new_n657), .C2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  OAI211_X1 g0460(.A(new_n649), .B(new_n660), .C1(new_n425), .C2(new_n648), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT21), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n659), .A2(G169), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n662), .B1(new_n663), .B2(new_n648), .ZN(new_n664));
  INV_X1    g0464(.A(new_n648), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n665), .A2(KEYINPUT21), .A3(G169), .A4(new_n659), .ZN(new_n666));
  NOR3_X1   g0466(.A1(new_n645), .A2(new_n647), .A3(new_n557), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(new_n659), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n661), .A2(new_n664), .A3(new_n666), .A4(new_n668), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n640), .A2(new_n669), .ZN(new_n670));
  AND4_X1   g0470(.A1(new_n514), .A2(new_n563), .A3(new_n636), .A4(new_n670), .ZN(G372));
  NOR2_X1   g0471(.A1(new_n588), .A2(new_n575), .ZN(new_n672));
  INV_X1    g0472(.A(new_n592), .ZN(new_n673));
  INV_X1    g0473(.A(new_n562), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n673), .A2(KEYINPUT26), .A3(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT26), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n676), .B1(new_n592), .B2(new_n562), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n672), .B1(new_n675), .B2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n640), .ZN(new_n679));
  AND3_X1   g0479(.A1(new_n666), .A2(new_n664), .A3(new_n668), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n681), .A2(new_n636), .A3(new_n563), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n678), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n514), .A2(new_n683), .ZN(new_n684));
  AND3_X1   g0484(.A1(new_n488), .A2(KEYINPUT96), .A3(new_n495), .ZN(new_n685));
  AOI21_X1  g0485(.A(KEYINPUT96), .B1(new_n488), .B2(new_n495), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  AND2_X1   g0487(.A1(new_n503), .A2(new_n504), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(new_n428), .ZN(new_n689));
  AND2_X1   g0489(.A1(new_n423), .A2(new_n375), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n687), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n383), .A2(KEYINPUT97), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT97), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n346), .A2(new_n693), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n691), .A2(new_n692), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(new_n373), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n684), .A2(new_n697), .ZN(G369));
  INV_X1    g0498(.A(new_n278), .ZN(new_n699));
  OR3_X1    g0499(.A1(new_n699), .A2(KEYINPUT27), .A3(G20), .ZN(new_n700));
  OAI21_X1  g0500(.A(KEYINPUT27), .B1(new_n699), .B2(G20), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n700), .A2(G213), .A3(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(G343), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  OR3_X1    g0505(.A1(new_n680), .A2(new_n660), .A3(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n660), .A2(new_n705), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n706), .B1(new_n669), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(G330), .ZN(new_n709));
  XNOR2_X1  g0509(.A(new_n709), .B(KEYINPUT98), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n635), .A2(new_n608), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n711), .B1(new_n635), .B2(new_n705), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(new_n679), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n640), .A2(new_n705), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  OR2_X1    g0515(.A1(new_n710), .A2(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n680), .A2(new_n704), .ZN(new_n717));
  AOI22_X1  g0517(.A1(new_n713), .A2(new_n717), .B1(new_n640), .B2(new_n705), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n716), .A2(new_n718), .ZN(G399));
  INV_X1    g0519(.A(new_n218), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n720), .A2(G41), .ZN(new_n721));
  INV_X1    g0521(.A(G1), .ZN(new_n722));
  NOR4_X1   g0522(.A1(new_n721), .A2(new_n722), .A3(G116), .A4(new_n569), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n723), .B1(new_n208), .B2(new_n721), .ZN(new_n724));
  XOR2_X1   g0524(.A(new_n724), .B(KEYINPUT28), .Z(new_n725));
  XOR2_X1   g0525(.A(KEYINPUT100), .B(KEYINPUT29), .Z(new_n726));
  NOR2_X1   g0526(.A1(KEYINPUT100), .A2(KEYINPUT29), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n704), .B1(new_n678), .B2(new_n682), .ZN(new_n728));
  MUX2_X1   g0528(.A(new_n726), .B(new_n727), .S(new_n728), .Z(new_n729));
  NAND4_X1  g0529(.A1(new_n636), .A2(new_n670), .A3(new_n563), .A4(new_n705), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT30), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n601), .A2(new_n604), .A3(new_n667), .A4(new_n586), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n540), .A2(new_n393), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n733), .A2(new_n523), .A3(new_n526), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n731), .B1(new_n732), .B2(new_n734), .ZN(new_n735));
  AND2_X1   g0535(.A1(new_n601), .A2(new_n604), .ZN(new_n736));
  AND2_X1   g0536(.A1(new_n667), .A2(new_n586), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n736), .A2(KEYINPUT30), .A3(new_n737), .A4(new_n541), .ZN(new_n738));
  NOR3_X1   g0538(.A1(new_n648), .A2(new_n586), .A3(G179), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n734), .A2(new_n605), .A3(new_n739), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n735), .A2(new_n738), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(new_n704), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT31), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g0544(.A(KEYINPUT99), .B(KEYINPUT31), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n741), .A2(new_n704), .A3(new_n746), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n730), .A2(new_n744), .A3(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n729), .B1(G330), .B2(new_n748), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n725), .B1(new_n749), .B2(G1), .ZN(G364));
  NOR2_X1   g0550(.A1(new_n277), .A2(G20), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n722), .B1(new_n751), .B2(G45), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  OAI221_X1 g0553(.A(new_n710), .B1(G330), .B2(new_n708), .C1(new_n721), .C2(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n721), .A2(new_n753), .ZN(new_n755));
  XNOR2_X1  g0555(.A(new_n755), .B(KEYINPUT101), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n218), .A2(new_n309), .ZN(new_n757));
  INV_X1    g0557(.A(G355), .ZN(new_n758));
  OAI22_X1  g0558(.A1(new_n757), .A2(new_n758), .B1(G116), .B2(new_n218), .ZN(new_n759));
  OR2_X1    g0559(.A1(new_n248), .A2(new_n307), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n464), .A2(new_n218), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n761), .B1(new_n307), .B2(new_n208), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n759), .B1(new_n760), .B2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(G13), .A2(G33), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(G20), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n209), .B1(G20), .B2(new_n370), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n756), .B1(new_n763), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(G20), .A2(G179), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(G200), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(G190), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  XNOR2_X1  g0575(.A(KEYINPUT33), .B(G317), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n775), .B1(new_n776), .B2(KEYINPUT104), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n777), .B1(KEYINPUT104), .B2(new_n776), .ZN(new_n778));
  NOR2_X1   g0578(.A1(G190), .A2(G200), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n772), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n309), .B1(new_n781), .B2(G311), .ZN(new_n782));
  NOR2_X1   g0582(.A1(G179), .A2(G200), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NOR3_X1   g0584(.A1(new_n784), .A2(new_n210), .A3(G190), .ZN(new_n785));
  NOR3_X1   g0585(.A1(new_n771), .A2(new_n368), .A3(G200), .ZN(new_n786));
  AOI22_X1  g0586(.A1(new_n785), .A2(G329), .B1(new_n786), .B2(G322), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n773), .A2(new_n368), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n210), .A2(G179), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n789), .A2(new_n368), .A3(G200), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  AOI22_X1  g0591(.A1(G326), .A2(new_n788), .B1(new_n791), .B2(G283), .ZN(new_n792));
  AND4_X1   g0592(.A1(new_n778), .A2(new_n782), .A3(new_n787), .A4(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(G294), .ZN(new_n794));
  OAI21_X1  g0594(.A(G20), .B1(new_n784), .B2(new_n368), .ZN(new_n795));
  INV_X1    g0595(.A(KEYINPUT103), .ZN(new_n796));
  OR2_X1    g0596(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n795), .A2(new_n796), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(G303), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n789), .A2(G190), .A3(G200), .ZN(new_n801));
  INV_X1    g0601(.A(KEYINPUT102), .ZN(new_n802));
  OR2_X1    g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n801), .A2(new_n802), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  OAI221_X1 g0605(.A(new_n793), .B1(new_n794), .B2(new_n799), .C1(new_n800), .C2(new_n805), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n309), .B1(new_n780), .B2(new_n230), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n785), .A2(G159), .ZN(new_n808));
  XNOR2_X1  g0608(.A(new_n808), .B(KEYINPUT32), .ZN(new_n809));
  INV_X1    g0609(.A(new_n433), .ZN(new_n810));
  AOI211_X1 g0610(.A(new_n807), .B(new_n809), .C1(new_n810), .C2(new_n786), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n790), .A2(new_n232), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n775), .A2(new_n224), .ZN(new_n813));
  AOI211_X1 g0613(.A(new_n812), .B(new_n813), .C1(G50), .C2(new_n788), .ZN(new_n814));
  INV_X1    g0614(.A(new_n799), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n815), .A2(G97), .ZN(new_n816));
  INV_X1    g0616(.A(new_n805), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(G87), .ZN(new_n818));
  NAND4_X1  g0618(.A1(new_n811), .A2(new_n814), .A3(new_n816), .A4(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n806), .A2(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n770), .B1(new_n820), .B2(new_n767), .ZN(new_n821));
  INV_X1    g0621(.A(new_n766), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n821), .B1(new_n708), .B2(new_n822), .ZN(new_n823));
  AND2_X1   g0623(.A1(new_n754), .A2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(G396));
  NOR2_X1   g0625(.A1(new_n375), .A2(new_n704), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n369), .B1(new_n359), .B2(new_n705), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n826), .B1(new_n827), .B2(new_n375), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n728), .B(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n748), .A2(G330), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n755), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n831), .B1(new_n830), .B2(new_n829), .ZN(new_n832));
  INV_X1    g0632(.A(new_n767), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(new_n765), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n756), .B1(G77), .B2(new_n834), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n781), .A2(G159), .B1(G143), .B2(new_n786), .ZN(new_n836));
  INV_X1    g0636(.A(G150), .ZN(new_n837));
  INV_X1    g0637(.A(G137), .ZN(new_n838));
  INV_X1    g0638(.A(new_n788), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n836), .B1(new_n775), .B2(new_n837), .C1(new_n838), .C2(new_n839), .ZN(new_n840));
  XOR2_X1   g0640(.A(new_n840), .B(KEYINPUT34), .Z(new_n841));
  AOI21_X1  g0641(.A(new_n464), .B1(G132), .B2(new_n785), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n791), .A2(G68), .ZN(new_n843));
  AND2_X1   g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  OAI221_X1 g0644(.A(new_n844), .B1(new_n202), .B2(new_n805), .C1(new_n433), .C2(new_n799), .ZN(new_n845));
  AOI22_X1  g0645(.A1(G283), .A2(new_n774), .B1(new_n788), .B2(G303), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n309), .B1(new_n781), .B2(G116), .ZN(new_n847));
  AOI22_X1  g0647(.A1(new_n785), .A2(G311), .B1(new_n786), .B2(G294), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n791), .A2(G87), .ZN(new_n849));
  NAND4_X1  g0649(.A1(new_n846), .A2(new_n847), .A3(new_n848), .A4(new_n849), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n816), .B1(new_n232), .B2(new_n805), .ZN(new_n851));
  OAI22_X1  g0651(.A1(new_n841), .A2(new_n845), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n835), .B1(new_n852), .B2(new_n767), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n853), .B1(new_n828), .B2(new_n765), .ZN(new_n854));
  AND2_X1   g0654(.A1(new_n832), .A2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(G384));
  OR2_X1    g0656(.A1(new_n551), .A2(KEYINPUT35), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n551), .A2(KEYINPUT35), .ZN(new_n858));
  NAND4_X1  g0658(.A1(new_n857), .A2(G116), .A3(new_n212), .A4(new_n858), .ZN(new_n859));
  XOR2_X1   g0659(.A(new_n859), .B(KEYINPUT36), .Z(new_n860));
  OAI211_X1 g0660(.A(new_n208), .B(G77), .C1(new_n224), .C2(new_n433), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n202), .A2(G68), .ZN(new_n862));
  AOI211_X1 g0662(.A(new_n722), .B(G13), .C1(new_n861), .C2(new_n862), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n860), .A2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT38), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n435), .B1(new_n461), .B2(new_n465), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n258), .B1(new_n866), .B2(new_n432), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT105), .ZN(new_n868));
  AND2_X1   g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n466), .B1(new_n867), .B2(new_n868), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n500), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n702), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n873), .B1(new_n688), .B2(new_n496), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n871), .A2(new_n490), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n469), .A2(new_n499), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n873), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n872), .B1(new_n494), .B2(new_n431), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n469), .A2(new_n487), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n881), .A2(KEYINPUT37), .ZN(new_n882));
  AOI22_X1  g0682(.A1(new_n877), .A2(KEYINPUT37), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n865), .B1(new_n874), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n877), .A2(KEYINPUT37), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n880), .A2(new_n882), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n506), .A2(new_n872), .A3(new_n871), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n887), .A2(KEYINPUT38), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n884), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n422), .A2(new_n704), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n423), .A2(new_n428), .A3(new_n891), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n422), .B(new_n704), .C1(new_n411), .C2(new_n427), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n728), .A2(new_n828), .ZN(new_n895));
  INV_X1    g0695(.A(new_n826), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n890), .A2(new_n894), .A3(new_n897), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n898), .B1(new_n687), .B2(new_n872), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n878), .B1(new_n687), .B2(new_n688), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n876), .A2(KEYINPUT96), .A3(new_n878), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(KEYINPUT37), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n902), .B1(new_n881), .B2(new_n879), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT96), .ZN(new_n904));
  INV_X1    g0704(.A(new_n881), .ZN(new_n905));
  NAND4_X1  g0705(.A1(new_n880), .A2(new_n904), .A3(KEYINPUT37), .A4(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n903), .A2(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n865), .B1(new_n900), .B2(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(KEYINPUT39), .B1(new_n908), .B2(new_n889), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n884), .A2(new_n889), .A3(KEYINPUT39), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n411), .A2(new_n422), .A3(new_n705), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n899), .B1(new_n912), .B2(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n696), .B1(new_n514), .B2(new_n729), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n915), .B(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT40), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n884), .A2(new_n889), .A3(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(new_n828), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n920), .B1(new_n892), .B2(new_n893), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n742), .A2(new_n745), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n741), .A2(KEYINPUT31), .A3(new_n704), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n730), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n921), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n918), .A2(KEYINPUT106), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n919), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(KEYINPUT106), .B1(new_n921), .B2(new_n924), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n929), .B1(new_n908), .B2(new_n889), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n928), .B1(new_n930), .B2(new_n918), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n931), .A2(new_n514), .A3(new_n924), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT106), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n925), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n488), .A2(new_n495), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(new_n904), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n488), .A2(KEYINPUT96), .A3(new_n495), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n688), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(new_n878), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  AOI22_X1  g0740(.A1(new_n880), .A2(new_n905), .B1(new_n901), .B2(KEYINPUT37), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT37), .ZN(new_n942));
  NOR4_X1   g0742(.A1(new_n879), .A2(new_n881), .A3(KEYINPUT96), .A4(new_n942), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  AOI21_X1  g0744(.A(KEYINPUT38), .B1(new_n940), .B2(new_n944), .ZN(new_n945));
  NOR3_X1   g0745(.A1(new_n874), .A2(new_n883), .A3(new_n865), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n934), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  AOI22_X1  g0747(.A1(new_n947), .A2(KEYINPUT40), .B1(new_n919), .B2(new_n927), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n514), .A2(new_n924), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n932), .A2(G330), .A3(new_n950), .ZN(new_n951));
  OAI22_X1  g0751(.A1(new_n917), .A2(new_n951), .B1(new_n722), .B2(new_n751), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT107), .ZN(new_n953));
  AND2_X1   g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n917), .A2(new_n951), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(new_n952), .B2(new_n953), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n864), .B1(new_n954), .B2(new_n956), .ZN(G367));
  OAI21_X1  g0757(.A(new_n563), .B1(new_n554), .B2(new_n705), .ZN(new_n958));
  OR2_X1    g0758(.A1(new_n958), .A2(new_n679), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n704), .B1(new_n959), .B2(new_n562), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n674), .A2(new_n704), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n958), .A2(new_n961), .ZN(new_n962));
  NAND4_X1  g0762(.A1(new_n962), .A2(new_n714), .A3(new_n713), .A4(new_n717), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n960), .B1(new_n963), .B2(KEYINPUT42), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n964), .B1(KEYINPUT42), .B2(new_n963), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n591), .A2(new_n704), .ZN(new_n966));
  MUX2_X1   g0766(.A(new_n672), .B(new_n673), .S(new_n966), .Z(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(KEYINPUT43), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n968), .B(KEYINPUT108), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n965), .A2(new_n969), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n967), .A2(KEYINPUT43), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n970), .B(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(new_n716), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(new_n962), .ZN(new_n974));
  XOR2_X1   g0774(.A(new_n972), .B(new_n974), .Z(new_n975));
  XOR2_X1   g0775(.A(new_n721), .B(KEYINPUT41), .Z(new_n976));
  XNOR2_X1  g0776(.A(new_n710), .B(new_n715), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(new_n717), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n978), .A2(new_n749), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n718), .A2(new_n962), .ZN(new_n980));
  AND2_X1   g0780(.A1(new_n980), .A2(KEYINPUT44), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n980), .A2(KEYINPUT44), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT109), .ZN(new_n983));
  OR3_X1    g0783(.A1(new_n981), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n982), .A2(new_n983), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n718), .A2(new_n962), .ZN(new_n986));
  XOR2_X1   g0786(.A(new_n986), .B(KEYINPUT45), .Z(new_n987));
  NAND3_X1  g0787(.A1(new_n984), .A2(new_n985), .A3(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n988), .A2(new_n973), .ZN(new_n989));
  INV_X1    g0789(.A(new_n989), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n988), .A2(new_n973), .ZN(new_n991));
  OR3_X1    g0791(.A1(new_n979), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n976), .B1(new_n992), .B2(new_n749), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n975), .B1(new_n993), .B2(new_n753), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n817), .A2(new_n810), .B1(G137), .B2(new_n785), .ZN(new_n995));
  OR2_X1    g0795(.A1(new_n995), .A2(KEYINPUT114), .ZN(new_n996));
  AOI22_X1  g0796(.A1(new_n781), .A2(G50), .B1(G150), .B2(new_n786), .ZN(new_n997));
  INV_X1    g0797(.A(G159), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n997), .B1(new_n998), .B2(new_n775), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n999), .B1(G143), .B2(new_n788), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n815), .A2(G68), .ZN(new_n1001));
  AND2_X1   g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n995), .A2(KEYINPUT114), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n309), .B1(new_n790), .B2(new_n230), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT113), .ZN(new_n1005));
  NAND4_X1  g0805(.A1(new_n996), .A2(new_n1002), .A3(new_n1003), .A4(new_n1005), .ZN(new_n1006));
  AOI21_X1  g0806(.A(KEYINPUT46), .B1(new_n817), .B2(G116), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(KEYINPUT112), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n464), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n775), .A2(new_n794), .B1(new_n543), .B2(new_n790), .ZN(new_n1010));
  AOI211_X1 g0810(.A(new_n1009), .B(new_n1010), .C1(G311), .C2(new_n788), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n817), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n815), .A2(G107), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n786), .ZN(new_n1014));
  INV_X1    g0814(.A(G283), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n1014), .A2(new_n800), .B1(new_n780), .B2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1016), .B1(G317), .B2(new_n785), .ZN(new_n1017));
  NAND4_X1  g0817(.A1(new_n1011), .A2(new_n1012), .A3(new_n1013), .A4(new_n1017), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1006), .B1(new_n1008), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT47), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n833), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1021), .B1(new_n1020), .B2(new_n1019), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n768), .B1(new_n218), .B2(new_n347), .C1(new_n244), .C2(new_n761), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT110), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1024), .A2(new_n756), .ZN(new_n1025));
  XOR2_X1   g0825(.A(new_n1025), .B(KEYINPUT111), .Z(new_n1026));
  OAI211_X1 g0826(.A(new_n1022), .B(new_n1026), .C1(new_n967), .C2(new_n822), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n994), .A2(new_n1027), .ZN(G387));
  INV_X1    g0828(.A(new_n721), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1029), .B1(new_n978), .B2(new_n749), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1030), .B1(new_n749), .B2(new_n978), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n241), .A2(new_n307), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n569), .A2(G116), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n1032), .A2(new_n761), .B1(new_n1033), .B2(new_n757), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n350), .ZN(new_n1035));
  OR3_X1    g0835(.A1(new_n1035), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1036));
  OAI21_X1  g0836(.A(KEYINPUT50), .B1(new_n1035), .B2(G50), .ZN(new_n1037));
  AOI21_X1  g0837(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1038));
  NAND4_X1  g0838(.A1(new_n1036), .A2(new_n1033), .A3(new_n1037), .A4(new_n1038), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n1034), .A2(new_n1039), .B1(new_n232), .B2(new_n720), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n756), .B1(new_n1040), .B2(new_n769), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1041), .B(KEYINPUT115), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n564), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n815), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n817), .A2(G77), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1009), .B1(new_n543), .B2(new_n790), .C1(new_n839), .C2(new_n998), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n785), .A2(G150), .B1(new_n786), .B2(G50), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n774), .A2(new_n266), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n1048), .B(new_n1049), .C1(new_n224), .C2(new_n780), .ZN(new_n1050));
  NOR3_X1   g0850(.A1(new_n1046), .A2(new_n1047), .A3(new_n1050), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n781), .A2(G303), .B1(G317), .B2(new_n786), .ZN(new_n1052));
  INV_X1    g0852(.A(G322), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1052), .B1(new_n1053), .B2(new_n839), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(G311), .B2(new_n774), .ZN(new_n1055));
  XOR2_X1   g0855(.A(new_n1055), .B(KEYINPUT116), .Z(new_n1056));
  INV_X1    g0856(.A(new_n1056), .ZN(new_n1057));
  AND2_X1   g0857(.A1(new_n1057), .A2(KEYINPUT48), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n1057), .A2(KEYINPUT48), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n799), .A2(new_n1015), .B1(new_n805), .B2(new_n794), .ZN(new_n1060));
  NOR3_X1   g0860(.A1(new_n1058), .A2(new_n1059), .A3(new_n1060), .ZN(new_n1061));
  OR2_X1    g0861(.A1(new_n1061), .A2(KEYINPUT49), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1009), .B1(G326), .B2(new_n785), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1063), .B1(new_n627), .B2(new_n790), .ZN(new_n1064));
  XOR2_X1   g0864(.A(new_n1064), .B(KEYINPUT117), .Z(new_n1065));
  AOI21_X1  g0865(.A(new_n1065), .B1(new_n1061), .B2(KEYINPUT49), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1051), .B1(new_n1062), .B2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1042), .B1(new_n1067), .B2(new_n833), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1068), .B1(new_n715), .B2(new_n766), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1069), .B1(new_n978), .B2(new_n753), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1031), .A2(new_n1070), .ZN(G393));
  OAI21_X1  g0871(.A(new_n979), .B1(new_n990), .B2(new_n991), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n992), .A2(new_n721), .A3(new_n1072), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n991), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1074), .A2(new_n753), .A3(new_n989), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n962), .A2(new_n822), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n464), .B1(G143), .B2(new_n785), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n1077), .B(new_n849), .C1(new_n224), .C2(new_n805), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(new_n1078), .B(KEYINPUT118), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n788), .A2(G150), .B1(G159), .B2(new_n786), .ZN(new_n1080));
  XOR2_X1   g0880(.A(new_n1080), .B(KEYINPUT51), .Z(new_n1081));
  NAND2_X1  g0881(.A1(new_n815), .A2(G77), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n774), .A2(G50), .B1(new_n781), .B2(new_n350), .ZN(new_n1083));
  NAND4_X1  g0883(.A1(new_n1079), .A2(new_n1081), .A3(new_n1082), .A4(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n785), .ZN(new_n1085));
  OAI221_X1 g0885(.A(new_n318), .B1(new_n794), .B2(new_n780), .C1(new_n1085), .C2(new_n1053), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n812), .B(new_n1086), .C1(G303), .C2(new_n774), .ZN(new_n1087));
  OAI221_X1 g0887(.A(new_n1087), .B1(new_n627), .B2(new_n799), .C1(new_n1015), .C2(new_n805), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n788), .A2(G317), .B1(G311), .B2(new_n786), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n1089), .B(KEYINPUT52), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1084), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1091), .A2(new_n767), .ZN(new_n1092));
  OAI221_X1 g0892(.A(new_n768), .B1(new_n543), .B2(new_n218), .C1(new_n251), .C2(new_n761), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1092), .A2(new_n756), .A3(new_n1093), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n1073), .B(new_n1075), .C1(new_n1076), .C2(new_n1094), .ZN(G390));
  OAI21_X1  g0895(.A(new_n756), .B1(new_n266), .B2(new_n834), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n1085), .A2(new_n794), .B1(new_n627), .B2(new_n1014), .ZN(new_n1097));
  AOI211_X1 g0897(.A(new_n309), .B(new_n1097), .C1(G97), .C2(new_n781), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n843), .B1(new_n839), .B2(new_n1015), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1099), .B1(G107), .B2(new_n774), .ZN(new_n1100));
  NAND4_X1  g0900(.A1(new_n1098), .A2(new_n818), .A3(new_n1082), .A4(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(G132), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n309), .B1(new_n1014), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(G128), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n839), .A2(new_n1104), .B1(new_n202), .B2(new_n790), .ZN(new_n1105));
  AOI211_X1 g0905(.A(new_n1103), .B(new_n1105), .C1(G125), .C2(new_n785), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(KEYINPUT54), .B(G143), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n775), .A2(new_n838), .B1(new_n780), .B2(new_n1107), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n815), .A2(G159), .B1(new_n1108), .B2(KEYINPUT121), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n1106), .B(new_n1109), .C1(KEYINPUT121), .C2(new_n1108), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n817), .A2(G150), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(new_n1111), .B(KEYINPUT53), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1101), .B1(new_n1110), .B2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1096), .B1(new_n1113), .B2(new_n767), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(new_n1114), .B(KEYINPUT122), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1115), .B1(new_n912), .B2(new_n765), .ZN(new_n1116));
  AND2_X1   g0916(.A1(new_n924), .A2(G330), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1117), .A2(new_n921), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n914), .B1(new_n897), .B2(new_n894), .ZN(new_n1120));
  INV_X1    g0920(.A(KEYINPUT39), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1121), .B1(new_n945), .B2(new_n946), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1120), .B1(new_n1122), .B2(new_n910), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n826), .B1(new_n728), .B2(new_n828), .ZN(new_n1124));
  AND2_X1   g0924(.A1(new_n892), .A2(new_n893), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n913), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1126), .B1(new_n889), .B2(new_n908), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1119), .B1(new_n1123), .B2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1126), .B1(new_n909), .B2(new_n911), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1120), .B1(new_n946), .B2(new_n945), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n894), .A2(G330), .A3(new_n748), .A4(new_n828), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1129), .A2(new_n1130), .A3(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1128), .A2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1116), .B1(new_n1133), .B2(new_n752), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT123), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(new_n1134), .B(new_n1135), .ZN(new_n1136));
  AND3_X1   g0936(.A1(new_n387), .A2(new_n509), .A3(new_n512), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n512), .B1(new_n387), .B2(new_n509), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n729), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1117), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n924), .A2(G330), .A3(new_n828), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(new_n1125), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1142), .A2(new_n1131), .A3(new_n1124), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n748), .A2(G330), .A3(new_n828), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n1117), .A2(new_n921), .B1(new_n1144), .B2(new_n1125), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1143), .B1(new_n1145), .B2(new_n1124), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n1139), .A2(new_n1140), .A3(new_n1146), .A4(new_n697), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1147), .A2(KEYINPUT119), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT119), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n916), .A2(new_n1149), .A3(new_n1140), .A4(new_n1146), .ZN(new_n1150));
  AND2_X1   g0950(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1029), .B1(new_n1151), .B2(new_n1133), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1133), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(KEYINPUT120), .B1(new_n1152), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1131), .ZN(new_n1157));
  NOR3_X1   g0957(.A1(new_n1123), .A2(new_n1127), .A3(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1118), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n1150), .B(new_n1148), .C1(new_n1158), .C2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1160), .A2(new_n721), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1133), .B1(new_n1150), .B2(new_n1148), .ZN(new_n1162));
  INV_X1    g0962(.A(KEYINPUT120), .ZN(new_n1163));
  NOR3_X1   g0963(.A1(new_n1161), .A2(new_n1162), .A3(new_n1163), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1136), .B1(new_n1156), .B2(new_n1164), .ZN(G378));
  INV_X1    g0965(.A(KEYINPUT57), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n692), .A2(new_n694), .A3(new_n373), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n372), .A2(new_n872), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1167), .A2(new_n1169), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n692), .A2(new_n694), .A3(new_n373), .A4(new_n1168), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1172));
  AND3_X1   g0972(.A1(new_n1170), .A2(new_n1171), .A3(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1172), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(G330), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1175), .B1(new_n948), .B2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1172), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1170), .A2(new_n1171), .A3(new_n1172), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n931), .A2(G330), .A3(new_n1182), .ZN(new_n1183));
  AND3_X1   g0983(.A1(new_n1177), .A2(new_n915), .A3(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n915), .B1(new_n1177), .B2(new_n1183), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1139), .A2(new_n1140), .A3(new_n697), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1187), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1166), .B1(new_n1186), .B2(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1187), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1190), .B1(new_n1151), .B2(new_n1133), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1122), .A2(new_n910), .ZN(new_n1192));
  OAI221_X1 g0992(.A(new_n898), .B1(new_n687), .B2(new_n872), .C1(new_n1192), .C2(new_n913), .ZN(new_n1193));
  NOR3_X1   g0993(.A1(new_n948), .A2(new_n1175), .A3(new_n1176), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1182), .B1(new_n931), .B2(G330), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1193), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1177), .A2(new_n915), .A3(new_n1183), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1166), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1029), .B1(new_n1191), .B2(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT125), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1189), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  OAI21_X1  g1001(.A(KEYINPUT57), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n1200), .B(new_n721), .C1(new_n1202), .C2(new_n1188), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1203), .ZN(new_n1204));
  OR2_X1    g1004(.A1(new_n1201), .A2(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1186), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1175), .A2(new_n764), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n755), .B1(G50), .B2(new_n834), .ZN(new_n1208));
  XOR2_X1   g1008(.A(new_n1208), .B(KEYINPUT124), .Z(new_n1209));
  NOR2_X1   g1009(.A1(new_n790), .A2(new_n433), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n464), .B1(new_n775), .B2(new_n543), .ZN(new_n1211));
  AOI211_X1 g1011(.A(new_n1210), .B(new_n1211), .C1(G116), .C2(new_n788), .ZN(new_n1212));
  OAI221_X1 g1012(.A(new_n306), .B1(new_n232), .B2(new_n1014), .C1(new_n1085), .C2(new_n1015), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(new_n1043), .B2(new_n781), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n1212), .A2(new_n1001), .A3(new_n1045), .A4(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1216), .A2(KEYINPUT58), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n306), .B1(new_n464), .B2(new_n268), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1218), .A2(new_n202), .ZN(new_n1219));
  AND2_X1   g1019(.A1(new_n1217), .A2(new_n1219), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n1014), .A2(new_n1104), .B1(new_n780), .B2(new_n838), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n775), .A2(new_n1102), .ZN(new_n1222));
  AOI211_X1 g1022(.A(new_n1221), .B(new_n1222), .C1(G125), .C2(new_n788), .ZN(new_n1223));
  OAI221_X1 g1023(.A(new_n1223), .B1(new_n837), .B2(new_n799), .C1(new_n805), .C2(new_n1107), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n1224), .A2(KEYINPUT59), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1224), .A2(KEYINPUT59), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n791), .A2(G159), .ZN(new_n1227));
  AOI211_X1 g1027(.A(G33), .B(G41), .C1(new_n785), .C2(G124), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1226), .A2(new_n1227), .A3(new_n1228), .ZN(new_n1229));
  OAI221_X1 g1029(.A(new_n1220), .B1(KEYINPUT58), .B2(new_n1216), .C1(new_n1225), .C2(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1209), .B1(new_n1230), .B2(new_n767), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(new_n1206), .A2(new_n753), .B1(new_n1207), .B2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1205), .A2(new_n1232), .ZN(G375));
  NAND2_X1  g1033(.A1(new_n1146), .A2(new_n753), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n756), .B1(G68), .B2(new_n834), .ZN(new_n1235));
  OAI22_X1  g1035(.A1(new_n1085), .A2(new_n800), .B1(new_n1015), .B2(new_n1014), .ZN(new_n1236));
  AOI211_X1 g1036(.A(new_n309), .B(new_n1236), .C1(G107), .C2(new_n781), .ZN(new_n1237));
  OAI22_X1  g1037(.A1(new_n775), .A2(new_n627), .B1(new_n230), .B2(new_n790), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1238), .B1(G294), .B2(new_n788), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n817), .A2(G97), .ZN(new_n1240));
  NAND4_X1  g1040(.A1(new_n1237), .A2(new_n1044), .A3(new_n1239), .A4(new_n1240), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n1014), .A2(new_n838), .B1(new_n780), .B2(new_n837), .ZN(new_n1242));
  OAI22_X1  g1042(.A1(new_n1102), .A2(new_n839), .B1(new_n775), .B2(new_n1107), .ZN(new_n1243));
  AOI211_X1 g1043(.A(new_n1242), .B(new_n1243), .C1(G128), .C2(new_n785), .ZN(new_n1244));
  OAI221_X1 g1044(.A(new_n1244), .B1(new_n202), .B2(new_n799), .C1(new_n998), .C2(new_n805), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n464), .A2(new_n1210), .ZN(new_n1246));
  XOR2_X1   g1046(.A(new_n1246), .B(KEYINPUT126), .Z(new_n1247));
  OAI21_X1  g1047(.A(new_n1241), .B1(new_n1245), .B2(new_n1247), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1235), .B1(new_n1248), .B2(new_n767), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1249), .B1(new_n894), .B2(new_n765), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1234), .A2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1146), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1187), .A2(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  OR2_X1    g1055(.A1(new_n1255), .A2(new_n976), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1252), .B1(new_n1256), .B2(new_n1154), .ZN(G381));
  NOR2_X1   g1057(.A1(G393), .A2(G396), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1258), .A2(new_n855), .ZN(new_n1259));
  NOR4_X1   g1059(.A1(G387), .A2(G390), .A3(G381), .A4(new_n1259), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1261), .A2(new_n1134), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1260), .A2(new_n1232), .A3(new_n1205), .A4(new_n1262), .ZN(G407));
  NAND2_X1  g1063(.A1(new_n703), .A2(G213), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1262), .A2(new_n1265), .ZN(new_n1266));
  OAI211_X1 g1066(.A(G407), .B(G213), .C1(G375), .C2(new_n1266), .ZN(G409));
  XNOR2_X1  g1067(.A(G393), .B(new_n824), .ZN(new_n1268));
  OR2_X1    g1068(.A1(new_n1268), .A2(G390), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1268), .A2(G390), .ZN(new_n1270));
  AND4_X1   g1070(.A1(new_n994), .A2(new_n1269), .A3(new_n1027), .A4(new_n1270), .ZN(new_n1271));
  AOI22_X1  g1071(.A1(new_n1269), .A2(new_n1270), .B1(new_n994), .B2(new_n1027), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT63), .ZN(new_n1274));
  OAI211_X1 g1074(.A(G378), .B(new_n1232), .C1(new_n1201), .C2(new_n1204), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1206), .A2(new_n1191), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1232), .B1(new_n1276), .B2(new_n976), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1277), .A2(new_n1262), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1275), .A2(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1279), .A2(new_n1264), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1148), .A2(new_n1150), .A3(KEYINPUT60), .ZN(new_n1281));
  AND2_X1   g1081(.A1(new_n1281), .A2(new_n1254), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT60), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n721), .B1(new_n1254), .B2(new_n1283), .ZN(new_n1284));
  OAI211_X1 g1084(.A(G384), .B(new_n1252), .C1(new_n1282), .C2(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1284), .B1(new_n1281), .B2(new_n1254), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n855), .B1(new_n1286), .B2(new_n1251), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1285), .A2(new_n1287), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1274), .B1(new_n1280), .B2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(G2897), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1264), .A2(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT127), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1292), .B1(new_n1288), .B2(new_n1293), .ZN(new_n1294));
  AOI211_X1 g1094(.A(KEYINPUT127), .B(new_n1291), .C1(new_n1285), .C2(new_n1287), .ZN(new_n1295));
  OAI22_X1  g1095(.A1(new_n1294), .A2(new_n1295), .B1(new_n1293), .B2(new_n1288), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1296), .ZN(new_n1297));
  AOI21_X1  g1097(.A(KEYINPUT61), .B1(new_n1280), .B2(new_n1297), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1265), .B1(new_n1275), .B2(new_n1278), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1288), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1299), .A2(KEYINPUT63), .A3(new_n1300), .ZN(new_n1301));
  NAND4_X1  g1101(.A1(new_n1273), .A2(new_n1289), .A3(new_n1298), .A4(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT62), .ZN(new_n1303));
  AND3_X1   g1103(.A1(new_n1299), .A2(new_n1303), .A3(new_n1300), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT61), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1305), .B1(new_n1299), .B2(new_n1296), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1303), .B1(new_n1299), .B2(new_n1300), .ZN(new_n1307));
  NOR3_X1   g1107(.A1(new_n1304), .A2(new_n1306), .A3(new_n1307), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1302), .B1(new_n1308), .B2(new_n1273), .ZN(G405));
  INV_X1    g1109(.A(new_n1273), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1262), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1311), .B1(new_n1205), .B2(new_n1232), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1312), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1313), .A2(new_n1288), .A3(new_n1275), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1275), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1300), .B1(new_n1312), .B2(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1314), .A2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1310), .A2(new_n1317), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1273), .A2(new_n1316), .A3(new_n1314), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1318), .A2(new_n1319), .ZN(G402));
endmodule


