//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 0 0 1 1 1 0 0 0 1 1 1 1 1 1 0 1 0 0 1 1 1 0 1 1 1 0 0 1 0 0 0 1 1 1 0 1 0 1 0 0 1 1 1 0 0 1 0 1 1 0 0 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:19 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n764, new_n766, new_n767, new_n768, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n780, new_n781, new_n782, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n796, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008;
  INV_X1    g000(.A(G472), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  XNOR2_X1  g002(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT71), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n189), .B(new_n190), .ZN(new_n191));
  NOR2_X1   g005(.A1(G237), .A2(G953), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G210), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n191), .A2(new_n194), .ZN(new_n195));
  XNOR2_X1  g009(.A(new_n189), .B(KEYINPUT71), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(new_n193), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  XNOR2_X1  g012(.A(KEYINPUT26), .B(G101), .ZN(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n198), .A2(new_n200), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n195), .A2(new_n197), .A3(new_n199), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT28), .ZN(new_n204));
  INV_X1    g018(.A(G146), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G143), .ZN(new_n206));
  INV_X1    g020(.A(G143), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G146), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  OAI211_X1 g023(.A(KEYINPUT67), .B(KEYINPUT1), .C1(new_n207), .C2(G146), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G128), .ZN(new_n211));
  AOI21_X1  g025(.A(KEYINPUT67), .B1(new_n206), .B2(KEYINPUT1), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n209), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT1), .ZN(new_n214));
  AND4_X1   g028(.A1(new_n214), .A2(new_n206), .A3(new_n208), .A4(G128), .ZN(new_n215));
  INV_X1    g029(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n213), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(G131), .ZN(new_n218));
  INV_X1    g032(.A(G137), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G134), .ZN(new_n220));
  INV_X1    g034(.A(G134), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G137), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n218), .B1(new_n220), .B2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT11), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n224), .B1(new_n221), .B2(G137), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n219), .A2(KEYINPUT11), .A3(G134), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n225), .A2(new_n226), .A3(new_n222), .ZN(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n223), .B1(new_n228), .B2(new_n218), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n217), .A2(new_n229), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n218), .A2(KEYINPUT66), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n227), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(new_n231), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n233), .A2(new_n225), .A3(new_n226), .A4(new_n222), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  AND2_X1   g049(.A1(KEYINPUT0), .A2(G128), .ZN(new_n236));
  AND3_X1   g050(.A1(new_n206), .A2(new_n208), .A3(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n236), .B1(new_n206), .B2(new_n208), .ZN(new_n238));
  OAI21_X1  g052(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  NOR3_X1   g054(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n237), .B1(new_n238), .B2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT65), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n235), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n242), .A2(new_n238), .ZN(new_n246));
  INV_X1    g060(.A(new_n237), .ZN(new_n247));
  AND3_X1   g061(.A1(new_n246), .A2(new_n244), .A3(new_n247), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n230), .B1(new_n245), .B2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(G116), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n250), .A2(G119), .ZN(new_n251));
  INV_X1    g065(.A(G119), .ZN(new_n252));
  OAI21_X1  g066(.A(KEYINPUT68), .B1(new_n252), .B2(G116), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT68), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n254), .A2(new_n250), .A3(G119), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n251), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  XOR2_X1   g070(.A(KEYINPUT2), .B(G113), .Z(new_n257));
  XNOR2_X1  g071(.A(new_n256), .B(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n249), .A2(new_n258), .ZN(new_n259));
  AOI22_X1  g073(.A1(new_n217), .A2(new_n229), .B1(new_n235), .B2(new_n243), .ZN(new_n260));
  INV_X1    g074(.A(new_n258), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n204), .B1(new_n259), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n235), .A2(new_n243), .ZN(new_n264));
  OAI21_X1  g078(.A(KEYINPUT1), .B1(new_n207), .B2(G146), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT67), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n267), .A2(G128), .A3(new_n210), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n215), .B1(new_n268), .B2(new_n209), .ZN(new_n269));
  INV_X1    g083(.A(new_n223), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n270), .B1(new_n227), .B2(G131), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n264), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n258), .B1(new_n272), .B2(KEYINPUT73), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT73), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n260), .A2(new_n274), .ZN(new_n275));
  AOI21_X1  g089(.A(KEYINPUT28), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n203), .B1(new_n263), .B2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT30), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n249), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n230), .A2(KEYINPUT30), .A3(new_n264), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT69), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n260), .A2(KEYINPUT69), .A3(KEYINPUT30), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n279), .A2(new_n282), .A3(new_n258), .A4(new_n283), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n272), .A2(new_n258), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n203), .A2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT31), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n284), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n287), .B1(new_n284), .B2(new_n286), .ZN(new_n289));
  OAI211_X1 g103(.A(new_n277), .B(new_n288), .C1(new_n289), .C2(KEYINPUT72), .ZN(new_n290));
  AND2_X1   g104(.A1(new_n289), .A2(KEYINPUT72), .ZN(new_n291));
  OAI211_X1 g105(.A(new_n187), .B(new_n188), .C1(new_n290), .C2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT32), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  AND2_X1   g108(.A1(new_n284), .A2(new_n286), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n246), .A2(new_n247), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(KEYINPUT65), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n243), .A2(new_n244), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n297), .A2(new_n235), .A3(new_n298), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n261), .B1(new_n299), .B2(new_n230), .ZN(new_n300));
  OAI21_X1  g114(.A(KEYINPUT28), .B1(new_n300), .B2(new_n285), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n261), .B1(new_n260), .B2(new_n274), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n272), .A2(KEYINPUT73), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n204), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  AOI22_X1  g119(.A1(new_n295), .A2(new_n287), .B1(new_n305), .B2(new_n203), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n284), .A2(new_n286), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(KEYINPUT31), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT72), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n289), .A2(KEYINPUT72), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n306), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  NAND4_X1  g126(.A1(new_n312), .A2(KEYINPUT32), .A3(new_n187), .A4(new_n188), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n272), .A2(new_n258), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(new_n262), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(KEYINPUT28), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(new_n304), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT29), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n203), .A2(new_n319), .ZN(new_n320));
  AOI21_X1  g134(.A(G902), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  AND2_X1   g135(.A1(new_n284), .A2(new_n262), .ZN(new_n322));
  INV_X1    g136(.A(new_n203), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n319), .B1(new_n305), .B2(new_n203), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n321), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(G472), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n294), .A2(new_n313), .A3(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT74), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT82), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT81), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n332), .A2(KEYINPUT25), .ZN(new_n333));
  INV_X1    g147(.A(G953), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n334), .A2(G221), .A3(G234), .ZN(new_n335));
  XNOR2_X1  g149(.A(new_n335), .B(KEYINPUT80), .ZN(new_n336));
  XNOR2_X1  g150(.A(KEYINPUT22), .B(G137), .ZN(new_n337));
  XNOR2_X1  g151(.A(new_n336), .B(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT23), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n340), .B1(new_n252), .B2(G128), .ZN(new_n341));
  INV_X1    g155(.A(G128), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n342), .A2(KEYINPUT23), .A3(G119), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n252), .A2(G128), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n341), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  XNOR2_X1  g159(.A(G119), .B(G128), .ZN(new_n346));
  INV_X1    g160(.A(G110), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(KEYINPUT24), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT24), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(G110), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  AOI22_X1  g165(.A1(new_n345), .A2(G110), .B1(new_n346), .B2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(G140), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(G125), .ZN(new_n354));
  INV_X1    g168(.A(G125), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(G140), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n354), .A2(new_n356), .A3(KEYINPUT16), .ZN(new_n357));
  OR3_X1    g171(.A1(new_n355), .A2(KEYINPUT16), .A3(G140), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n357), .A2(new_n358), .A3(G146), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(G146), .B1(new_n357), .B2(new_n358), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n352), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT76), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  OAI211_X1 g178(.A(new_n352), .B(KEYINPUT76), .C1(new_n360), .C2(new_n361), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n342), .A2(G119), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(new_n344), .ZN(new_n367));
  XNOR2_X1  g181(.A(KEYINPUT24), .B(G110), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND4_X1  g183(.A1(new_n341), .A2(new_n343), .A3(new_n347), .A4(new_n344), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(KEYINPUT77), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT77), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n369), .A2(new_n370), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n354), .A2(new_n356), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(KEYINPUT78), .ZN(new_n376));
  XNOR2_X1  g190(.A(G125), .B(G140), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT78), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n376), .A2(new_n379), .A3(new_n205), .ZN(new_n380));
  NAND4_X1  g194(.A1(new_n372), .A2(new_n374), .A3(new_n380), .A4(new_n359), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(KEYINPUT79), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n205), .B1(new_n377), .B2(new_n378), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n375), .A2(KEYINPUT78), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n359), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT79), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n386), .A2(new_n387), .A3(new_n374), .A4(new_n372), .ZN(new_n388));
  AOI221_X4 g202(.A(new_n339), .B1(new_n364), .B2(new_n365), .C1(new_n382), .C2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n382), .A2(new_n388), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n364), .A2(new_n365), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n338), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n389), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n333), .B1(new_n393), .B2(new_n188), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n373), .B1(new_n369), .B2(new_n370), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n385), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n387), .B1(new_n396), .B2(new_n374), .ZN(new_n397));
  AND3_X1   g211(.A1(new_n369), .A2(new_n373), .A3(new_n370), .ZN(new_n398));
  NOR4_X1   g212(.A1(new_n385), .A2(new_n398), .A3(new_n395), .A4(KEYINPUT79), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n391), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(new_n339), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n390), .A2(new_n391), .A3(new_n338), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n401), .A2(new_n188), .A3(new_n402), .A4(new_n333), .ZN(new_n403));
  INV_X1    g217(.A(G217), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n404), .B1(G234), .B2(new_n188), .ZN(new_n405));
  XOR2_X1   g219(.A(new_n405), .B(KEYINPUT75), .Z(new_n406));
  NAND2_X1  g220(.A1(new_n403), .A2(new_n406), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n331), .B1(new_n394), .B2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n333), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n401), .A2(new_n402), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n409), .B1(new_n410), .B2(G902), .ZN(new_n411));
  NAND4_X1  g225(.A1(new_n411), .A2(KEYINPUT82), .A3(new_n403), .A4(new_n406), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n405), .A2(G902), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n393), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n408), .A2(new_n412), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(KEYINPUT83), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT83), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n408), .A2(new_n412), .A3(new_n417), .A4(new_n414), .ZN(new_n418));
  AND2_X1   g232(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n192), .A2(G143), .A3(G214), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  AOI21_X1  g235(.A(G143), .B1(new_n192), .B2(G214), .ZN(new_n422));
  OAI21_X1  g236(.A(G131), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT17), .ZN(new_n424));
  INV_X1    g238(.A(G237), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n425), .A2(new_n334), .A3(G214), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(new_n207), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n427), .A2(new_n218), .A3(new_n420), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n423), .A2(new_n424), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(KEYINPUT95), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n360), .A2(new_n361), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT95), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n423), .A2(new_n432), .A3(new_n424), .A4(new_n428), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n427), .A2(new_n420), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n434), .A2(KEYINPUT17), .A3(G131), .ZN(new_n435));
  NAND4_X1  g249(.A1(new_n430), .A2(new_n431), .A3(new_n433), .A4(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT92), .ZN(new_n437));
  NAND2_X1  g251(.A1(KEYINPUT18), .A2(G131), .ZN(new_n438));
  OR3_X1    g252(.A1(new_n434), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n438), .B1(new_n434), .B2(new_n437), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n375), .A2(G146), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n380), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  XOR2_X1   g258(.A(G113), .B(G122), .Z(new_n445));
  XOR2_X1   g259(.A(KEYINPUT94), .B(G104), .Z(new_n446));
  XOR2_X1   g260(.A(new_n445), .B(new_n446), .Z(new_n447));
  AND3_X1   g261(.A1(new_n436), .A2(new_n444), .A3(new_n447), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n447), .B1(new_n436), .B2(new_n444), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n188), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(G475), .ZN(new_n451));
  INV_X1    g265(.A(G478), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n452), .A2(KEYINPUT15), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT97), .ZN(new_n455));
  XNOR2_X1  g269(.A(G116), .B(G122), .ZN(new_n456));
  INV_X1    g270(.A(G107), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n207), .A2(G128), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n342), .A2(G143), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n459), .A2(new_n460), .A3(new_n221), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n221), .B1(new_n459), .B2(new_n460), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n458), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n250), .A2(G122), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT14), .ZN(new_n466));
  OAI21_X1  g280(.A(G107), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n467), .B1(new_n466), .B2(new_n456), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n455), .B1(new_n464), .B2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(G122), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(G116), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n465), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(G107), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n462), .B1(new_n473), .B2(new_n458), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT96), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT13), .ZN(new_n476));
  OAI211_X1 g290(.A(new_n475), .B(new_n476), .C1(new_n342), .C2(G143), .ZN(new_n477));
  OAI211_X1 g291(.A(new_n477), .B(new_n460), .C1(new_n476), .C2(new_n459), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n475), .B1(new_n459), .B2(new_n476), .ZN(new_n479));
  OAI21_X1  g293(.A(G134), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n474), .A2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(new_n463), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(new_n461), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n470), .A2(G116), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n457), .B1(new_n484), .B2(KEYINPUT14), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n485), .B1(new_n472), .B2(KEYINPUT14), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n483), .A2(new_n486), .A3(KEYINPUT97), .A4(new_n458), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n469), .A2(new_n481), .A3(new_n487), .ZN(new_n488));
  XNOR2_X1  g302(.A(KEYINPUT9), .B(G234), .ZN(new_n489));
  NOR3_X1   g303(.A1(new_n489), .A2(new_n404), .A3(G953), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n469), .A2(new_n481), .A3(new_n487), .A4(new_n490), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n454), .B1(new_n494), .B2(new_n188), .ZN(new_n495));
  AOI211_X1 g309(.A(G902), .B(new_n453), .C1(new_n492), .C2(new_n493), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n436), .A2(new_n444), .A3(new_n447), .ZN(new_n498));
  INV_X1    g312(.A(new_n447), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT19), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n377), .A2(new_n378), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT93), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  OAI21_X1  g317(.A(KEYINPUT78), .B1(new_n502), .B2(new_n500), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n377), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(G146), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n423), .A2(new_n428), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(new_n359), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  AOI22_X1  g323(.A1(new_n439), .A2(new_n440), .B1(new_n380), .B2(new_n442), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n499), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n498), .A2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT20), .ZN(new_n513));
  NOR2_X1   g327(.A1(G475), .A2(G902), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n512), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n513), .B1(new_n512), .B2(new_n514), .ZN(new_n517));
  OAI211_X1 g331(.A(new_n451), .B(new_n497), .C1(new_n516), .C2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(G234), .A2(G237), .ZN(new_n519));
  AND3_X1   g333(.A1(new_n519), .A2(G952), .A3(new_n334), .ZN(new_n520));
  AND3_X1   g334(.A1(new_n519), .A2(G902), .A3(G953), .ZN(new_n521));
  XNOR2_X1  g335(.A(KEYINPUT21), .B(G898), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  OAI21_X1  g337(.A(KEYINPUT98), .B1(new_n518), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n512), .A2(new_n514), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(KEYINPUT20), .ZN(new_n526));
  AOI22_X1  g340(.A1(new_n526), .A2(new_n515), .B1(G475), .B2(new_n450), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT98), .ZN(new_n528));
  INV_X1    g342(.A(new_n523), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n527), .A2(new_n528), .A3(new_n529), .A4(new_n497), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n524), .A2(new_n530), .ZN(new_n531));
  OAI21_X1  g345(.A(G221), .B1(new_n489), .B2(G902), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n457), .A2(G104), .ZN(new_n534));
  OR2_X1    g348(.A1(KEYINPUT86), .A2(KEYINPUT3), .ZN(new_n535));
  NAND2_X1  g349(.A1(KEYINPUT86), .A2(KEYINPUT3), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(G104), .ZN(new_n538));
  OAI22_X1  g352(.A1(new_n538), .A2(G107), .B1(KEYINPUT86), .B2(KEYINPUT3), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(G107), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  OAI21_X1  g355(.A(G101), .B1(new_n537), .B2(new_n541), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n538), .A2(G107), .ZN(new_n543));
  INV_X1    g357(.A(new_n536), .ZN(new_n544));
  NOR2_X1   g358(.A1(KEYINPUT86), .A2(KEYINPUT3), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(G101), .ZN(new_n547));
  NAND4_X1  g361(.A1(new_n546), .A2(new_n547), .A3(new_n539), .A4(new_n540), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n542), .A2(KEYINPUT4), .A3(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT4), .ZN(new_n550));
  OAI211_X1 g364(.A(new_n550), .B(G101), .C1(new_n537), .C2(new_n541), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n549), .A2(new_n243), .A3(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT10), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n265), .A2(KEYINPUT87), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT87), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n206), .A2(new_n555), .A3(KEYINPUT1), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n554), .A2(G128), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n215), .B1(new_n557), .B2(new_n209), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n547), .B1(new_n534), .B2(new_n540), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n548), .A2(new_n560), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n553), .B1(new_n558), .B2(new_n561), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n537), .A2(new_n541), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n559), .B1(new_n563), .B2(new_n547), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n564), .A2(KEYINPUT10), .A3(new_n217), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n552), .A2(new_n562), .A3(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n235), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT88), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n269), .A2(new_n561), .A3(new_n569), .ZN(new_n570));
  OAI21_X1  g384(.A(KEYINPUT88), .B1(new_n558), .B2(new_n561), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n564), .A2(new_n217), .ZN(new_n572));
  OAI211_X1 g386(.A(new_n235), .B(new_n570), .C1(new_n571), .C2(new_n572), .ZN(new_n573));
  AOI22_X1  g387(.A1(new_n567), .A2(new_n568), .B1(new_n573), .B2(KEYINPUT12), .ZN(new_n574));
  XNOR2_X1  g388(.A(G110), .B(G140), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n334), .A2(G227), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n575), .B(new_n576), .ZN(new_n577));
  XNOR2_X1  g391(.A(KEYINPUT84), .B(KEYINPUT85), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n577), .B(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n209), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n214), .B1(G143), .B2(new_n205), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n342), .B1(new_n582), .B2(new_n555), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n581), .B1(new_n583), .B2(new_n554), .ZN(new_n584));
  OAI211_X1 g398(.A(new_n548), .B(new_n560), .C1(new_n584), .C2(new_n215), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n269), .A2(new_n561), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n585), .A2(KEYINPUT88), .A3(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT12), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n587), .A2(new_n588), .A3(new_n235), .A4(new_n570), .ZN(new_n589));
  NAND4_X1  g403(.A1(new_n574), .A2(KEYINPUT90), .A3(new_n580), .A4(new_n589), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n571), .A2(new_n572), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n570), .A2(new_n235), .ZN(new_n592));
  OAI21_X1  g406(.A(KEYINPUT12), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n552), .A2(new_n562), .A3(new_n565), .A4(new_n568), .ZN(new_n594));
  NAND4_X1  g408(.A1(new_n593), .A2(new_n594), .A3(new_n580), .A4(new_n589), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT90), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n566), .A2(new_n235), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n580), .B1(new_n598), .B2(new_n594), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n590), .A2(new_n597), .A3(new_n600), .ZN(new_n601));
  XNOR2_X1  g415(.A(KEYINPUT89), .B(G469), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n601), .A2(new_n188), .A3(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n574), .A2(new_n579), .A3(new_n589), .ZN(new_n605));
  INV_X1    g419(.A(new_n598), .ZN(new_n606));
  INV_X1    g420(.A(new_n594), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n580), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g423(.A(G469), .B1(new_n609), .B2(G902), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n533), .B1(new_n604), .B2(new_n610), .ZN(new_n611));
  OAI21_X1  g425(.A(G214), .B1(G237), .B2(G902), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n258), .A2(new_n549), .A3(new_n551), .ZN(new_n614));
  XNOR2_X1  g428(.A(KEYINPUT91), .B(KEYINPUT5), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n256), .A2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(G113), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n618), .B1(new_n615), .B2(new_n251), .ZN(new_n619));
  AOI22_X1  g433(.A1(new_n617), .A2(new_n619), .B1(new_n256), .B2(new_n257), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n564), .ZN(new_n621));
  XNOR2_X1  g435(.A(G110), .B(G122), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n614), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n243), .A2(G125), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n624), .B1(G125), .B2(new_n269), .ZN(new_n625));
  INV_X1    g439(.A(G224), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n626), .A2(G953), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n625), .A2(KEYINPUT7), .A3(new_n628), .ZN(new_n629));
  XOR2_X1   g443(.A(new_n622), .B(KEYINPUT8), .Z(new_n630));
  AOI21_X1  g444(.A(new_n630), .B1(new_n620), .B2(new_n561), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n256), .A2(new_n257), .ZN(new_n632));
  AND2_X1   g446(.A1(new_n256), .A2(KEYINPUT5), .ZN(new_n633));
  INV_X1    g447(.A(new_n619), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n632), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(new_n564), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n631), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n628), .A2(KEYINPUT7), .ZN(new_n638));
  OAI211_X1 g452(.A(new_n624), .B(new_n638), .C1(G125), .C2(new_n269), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n623), .A2(new_n629), .A3(new_n637), .A4(new_n639), .ZN(new_n640));
  AND2_X1   g454(.A1(new_n640), .A2(new_n188), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n614), .A2(new_n621), .ZN(new_n642));
  INV_X1    g456(.A(new_n622), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n644), .A2(KEYINPUT6), .A3(new_n623), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT6), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n642), .A2(new_n646), .A3(new_n643), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n625), .B(new_n628), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n645), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n641), .A2(new_n649), .ZN(new_n650));
  OAI21_X1  g464(.A(G210), .B1(G237), .B2(G902), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n641), .A2(new_n649), .A3(new_n651), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n613), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  AND3_X1   g469(.A1(new_n531), .A2(new_n611), .A3(new_n655), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n294), .A2(new_n313), .A3(KEYINPUT74), .A4(new_n327), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n330), .A2(new_n419), .A3(new_n656), .A4(new_n657), .ZN(new_n658));
  XOR2_X1   g472(.A(KEYINPUT99), .B(G101), .Z(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G3));
  AOI21_X1  g474(.A(G478), .B1(new_n494), .B2(new_n188), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT103), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n494), .A2(KEYINPUT102), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(KEYINPUT33), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n188), .A2(G478), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n663), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(new_n527), .ZN(new_n668));
  AND2_X1   g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(KEYINPUT104), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT101), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n671), .B1(new_n650), .B2(new_n652), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n613), .B1(new_n672), .B2(new_n654), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n641), .A2(new_n649), .A3(new_n671), .A4(new_n651), .ZN(new_n674));
  AND2_X1   g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(new_n529), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n670), .A2(new_n676), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n188), .B1(new_n290), .B2(new_n291), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT100), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n678), .A2(new_n679), .A3(G472), .ZN(new_n680));
  OAI211_X1 g494(.A(new_n312), .B(new_n188), .C1(KEYINPUT100), .C2(new_n187), .ZN(new_n681));
  AND3_X1   g495(.A1(new_n611), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  AND2_X1   g496(.A1(new_n419), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n677), .A2(new_n683), .ZN(new_n684));
  XOR2_X1   g498(.A(KEYINPUT34), .B(G104), .Z(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(G6));
  INV_X1    g500(.A(new_n497), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n527), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n676), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n683), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(KEYINPUT105), .ZN(new_n691));
  XOR2_X1   g505(.A(KEYINPUT35), .B(G107), .Z(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(G9));
  OR2_X1    g507(.A1(new_n339), .A2(KEYINPUT36), .ZN(new_n694));
  XOR2_X1   g508(.A(new_n400), .B(new_n694), .Z(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(new_n413), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n408), .A2(new_n412), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(KEYINPUT106), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT106), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n408), .A2(new_n412), .A3(new_n699), .A4(new_n696), .ZN(new_n700));
  AND3_X1   g514(.A1(new_n698), .A2(new_n531), .A3(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n680), .A2(new_n681), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n611), .A2(new_n655), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  XOR2_X1   g519(.A(KEYINPUT37), .B(G110), .Z(new_n706));
  XNOR2_X1  g520(.A(new_n705), .B(new_n706), .ZN(G12));
  NAND3_X1  g521(.A1(new_n330), .A2(new_n657), .A3(new_n675), .ZN(new_n708));
  INV_X1    g522(.A(G900), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n520), .B1(new_n521), .B2(new_n709), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n688), .A2(new_n710), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n698), .A2(new_n611), .A3(new_n700), .A4(new_n711), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n708), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(new_n342), .ZN(G30));
  AND2_X1   g528(.A1(new_n653), .A2(new_n654), .ZN(new_n715));
  XOR2_X1   g529(.A(KEYINPUT107), .B(KEYINPUT38), .Z(new_n716));
  XNOR2_X1  g530(.A(new_n715), .B(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n527), .A2(new_n497), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(new_n612), .ZN(new_n720));
  NOR3_X1   g534(.A1(new_n718), .A2(new_n697), .A3(new_n720), .ZN(new_n721));
  XOR2_X1   g535(.A(new_n710), .B(KEYINPUT39), .Z(new_n722));
  NAND2_X1  g536(.A1(new_n611), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(KEYINPUT40), .ZN(new_n724));
  OR2_X1    g538(.A1(new_n723), .A2(KEYINPUT40), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n322), .A2(new_n203), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n188), .B1(new_n323), .B2(new_n315), .ZN(new_n727));
  OAI21_X1  g541(.A(G472), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n294), .A2(new_n313), .A3(new_n728), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n721), .A2(new_n724), .A3(new_n725), .A4(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G143), .ZN(G45));
  AND3_X1   g545(.A1(new_n330), .A2(new_n657), .A3(new_n675), .ZN(new_n732));
  INV_X1    g546(.A(new_n710), .ZN(new_n733));
  AND3_X1   g547(.A1(new_n667), .A2(new_n668), .A3(new_n733), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n698), .A2(new_n734), .A3(new_n611), .A4(new_n700), .ZN(new_n735));
  INV_X1    g549(.A(new_n735), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n732), .A2(KEYINPUT108), .A3(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT108), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n738), .B1(new_n708), .B2(new_n735), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G146), .ZN(G48));
  AND3_X1   g555(.A1(new_n330), .A2(new_n419), .A3(new_n657), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT109), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n601), .A2(new_n743), .A3(new_n188), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(G469), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n599), .B1(new_n595), .B2(new_n596), .ZN(new_n746));
  AOI21_X1  g560(.A(G902), .B1(new_n746), .B2(new_n590), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n747), .A2(new_n743), .ZN(new_n748));
  OAI211_X1 g562(.A(new_n532), .B(new_n604), .C1(new_n745), .C2(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(KEYINPUT110), .ZN(new_n750));
  AOI211_X1 g564(.A(G902), .B(new_n602), .C1(new_n746), .C2(new_n590), .ZN(new_n751));
  INV_X1    g565(.A(G469), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n752), .B1(new_n747), .B2(new_n743), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n601), .A2(new_n188), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(KEYINPUT109), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n751), .B1(new_n753), .B2(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT110), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n756), .A2(new_n757), .A3(new_n532), .ZN(new_n758));
  AND2_X1   g572(.A1(new_n750), .A2(new_n758), .ZN(new_n759));
  AND2_X1   g573(.A1(new_n742), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(new_n677), .ZN(new_n761));
  XNOR2_X1  g575(.A(KEYINPUT41), .B(G113), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n761), .B(new_n762), .ZN(G15));
  NAND2_X1  g577(.A1(new_n760), .A2(new_n689), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G116), .ZN(G18));
  INV_X1    g579(.A(new_n749), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n701), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n708), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(new_n252), .ZN(G21));
  NAND2_X1  g583(.A1(new_n187), .A2(new_n188), .ZN(new_n770));
  AOI22_X1  g584(.A1(new_n317), .A2(new_n203), .B1(new_n307), .B2(KEYINPUT31), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n770), .B1(new_n771), .B2(new_n288), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n772), .B1(new_n678), .B2(G472), .ZN(new_n773));
  AND3_X1   g587(.A1(new_n408), .A2(new_n412), .A3(new_n414), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n673), .A2(new_n529), .A3(new_n674), .A4(new_n719), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n777), .A2(new_n750), .A3(new_n758), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G122), .ZN(G24));
  NAND3_X1  g593(.A1(new_n756), .A2(new_n675), .A3(new_n532), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n734), .A2(new_n773), .A3(new_n697), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(new_n355), .ZN(G27));
  AND2_X1   g597(.A1(new_n715), .A2(new_n612), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(new_n611), .ZN(new_n785));
  INV_X1    g599(.A(new_n734), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  AND3_X1   g601(.A1(new_n328), .A2(KEYINPUT111), .A3(new_n774), .ZN(new_n788));
  AOI21_X1  g602(.A(KEYINPUT111), .B1(new_n328), .B2(new_n774), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n787), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  AND3_X1   g604(.A1(new_n611), .A2(new_n612), .A3(new_n715), .ZN(new_n791));
  AND4_X1   g605(.A1(new_n330), .A2(new_n419), .A3(new_n657), .A4(new_n791), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n786), .A2(KEYINPUT42), .ZN(new_n793));
  AOI22_X1  g607(.A1(KEYINPUT42), .A2(new_n790), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(G131), .ZN(G33));
  NAND2_X1  g609(.A1(new_n792), .A2(new_n711), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(G134), .ZN(G36));
  AND2_X1   g611(.A1(new_n667), .A2(new_n527), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(KEYINPUT43), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n799), .A2(new_n702), .A3(new_n697), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT44), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n784), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  OR2_X1    g616(.A1(new_n802), .A2(KEYINPUT112), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n609), .A2(KEYINPUT45), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n609), .A2(KEYINPUT45), .ZN(new_n805));
  NOR3_X1   g619(.A1(new_n804), .A2(new_n805), .A3(new_n752), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n806), .B1(G469), .B2(G902), .ZN(new_n807));
  AND2_X1   g621(.A1(new_n807), .A2(KEYINPUT46), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n604), .B1(new_n807), .B2(KEYINPUT46), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n532), .B(new_n722), .C1(new_n808), .C2(new_n809), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n810), .B1(new_n800), .B2(new_n801), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n802), .A2(KEYINPUT112), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n803), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(G137), .ZN(G39));
  OAI21_X1  g628(.A(new_n532), .B1(new_n808), .B2(new_n809), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT47), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n815), .B(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n330), .A2(new_n657), .ZN(new_n818));
  INV_X1    g632(.A(new_n419), .ZN(new_n819));
  AND4_X1   g633(.A1(new_n818), .A2(new_n819), .A3(new_n734), .A4(new_n784), .ZN(new_n820));
  AOI21_X1  g634(.A(KEYINPUT113), .B1(new_n817), .B2(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n817), .A2(KEYINPUT113), .A3(new_n820), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n824), .B(G140), .ZN(G42));
  NAND2_X1  g639(.A1(new_n766), .A2(new_n784), .ZN(new_n826));
  XOR2_X1   g640(.A(new_n826), .B(KEYINPUT117), .Z(new_n827));
  INV_X1    g641(.A(new_n520), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n819), .A2(new_n729), .A3(new_n828), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n667), .A2(new_n668), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n832), .B(KEYINPUT118), .ZN(new_n833));
  AND3_X1   g647(.A1(new_n827), .A2(new_n520), .A3(new_n799), .ZN(new_n834));
  AND2_X1   g648(.A1(new_n773), .A2(new_n697), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  AND4_X1   g650(.A1(new_n774), .A2(new_n799), .A3(new_n520), .A4(new_n773), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n837), .A2(new_n613), .A3(new_n718), .A4(new_n766), .ZN(new_n838));
  XOR2_X1   g652(.A(new_n838), .B(KEYINPUT50), .Z(new_n839));
  XOR2_X1   g653(.A(new_n756), .B(KEYINPUT115), .Z(new_n840));
  NOR2_X1   g654(.A1(new_n840), .A2(new_n532), .ZN(new_n841));
  OAI211_X1 g655(.A(new_n784), .B(new_n837), .C1(new_n817), .C2(new_n841), .ZN(new_n842));
  AND4_X1   g656(.A1(new_n833), .A2(new_n836), .A3(new_n839), .A4(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n843), .A2(KEYINPUT51), .ZN(new_n844));
  OR2_X1    g658(.A1(new_n788), .A2(new_n789), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n834), .A2(new_n845), .ZN(new_n846));
  XNOR2_X1  g660(.A(KEYINPUT119), .B(KEYINPUT48), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n846), .A2(new_n847), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n334), .A2(G952), .ZN(new_n850));
  INV_X1    g664(.A(new_n780), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n850), .B1(new_n837), .B2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(new_n830), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n852), .B1(new_n853), .B2(new_n670), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n849), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n844), .A2(new_n848), .A3(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT52), .ZN(new_n857));
  OAI22_X1  g671(.A1(new_n708), .A2(new_n712), .B1(new_n780), .B2(new_n781), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n858), .B1(new_n737), .B2(new_n739), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n675), .A2(new_n719), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n697), .A2(new_n710), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n860), .A2(new_n611), .A3(new_n729), .A4(new_n861), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n857), .B1(new_n859), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n655), .A2(new_n529), .ZN(new_n864));
  AOI22_X1  g678(.A1(KEYINPUT116), .A2(new_n688), .B1(new_n667), .B2(new_n668), .ZN(new_n865));
  OR2_X1    g679(.A1(new_n688), .A2(KEYINPUT116), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n864), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n419), .A2(new_n867), .A3(new_n682), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n658), .A2(new_n778), .A3(new_n705), .A4(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n869), .A2(new_n768), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n835), .A2(new_n669), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n698), .A2(new_n497), .A3(new_n527), .A4(new_n700), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n871), .B1(new_n818), .B2(new_n872), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n785), .A2(new_n710), .ZN(new_n874));
  AOI22_X1  g688(.A1(new_n873), .A2(new_n874), .B1(new_n792), .B2(new_n711), .ZN(new_n875));
  OAI211_X1 g689(.A(new_n742), .B(new_n759), .C1(new_n677), .C2(new_n689), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n870), .A2(new_n794), .A3(new_n875), .A4(new_n876), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n863), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n859), .A2(new_n857), .A3(new_n862), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT53), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n878), .A2(KEYINPUT53), .A3(new_n879), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  XNOR2_X1  g698(.A(new_n884), .B(KEYINPUT54), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n843), .A2(KEYINPUT51), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n856), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  NOR2_X1   g701(.A1(G952), .A2(G953), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n840), .A2(KEYINPUT49), .ZN(new_n889));
  AND4_X1   g703(.A1(new_n774), .A2(new_n798), .A3(new_n532), .A4(new_n612), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n718), .B1(new_n890), .B2(KEYINPUT114), .ZN(new_n891));
  AOI211_X1 g705(.A(new_n729), .B(new_n891), .C1(KEYINPUT114), .C2(new_n890), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n840), .A2(KEYINPUT49), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  OAI22_X1  g708(.A1(new_n887), .A2(new_n888), .B1(new_n889), .B2(new_n894), .ZN(G75));
  NOR2_X1   g709(.A1(new_n334), .A2(G952), .ZN(new_n896));
  INV_X1    g710(.A(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT56), .ZN(new_n898));
  AOI21_X1  g712(.A(KEYINPUT53), .B1(new_n878), .B2(new_n879), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n873), .A2(new_n874), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n790), .A2(KEYINPUT42), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n792), .A2(new_n793), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n900), .A2(new_n901), .A3(new_n902), .A4(new_n796), .ZN(new_n903));
  AND4_X1   g717(.A1(new_n658), .A2(new_n778), .A3(new_n705), .A4(new_n868), .ZN(new_n904));
  INV_X1    g718(.A(new_n768), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n904), .A2(new_n905), .A3(new_n876), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n903), .A2(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(new_n712), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n782), .B1(new_n732), .B2(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(KEYINPUT108), .B1(new_n732), .B2(new_n736), .ZN(new_n910));
  NOR3_X1   g724(.A1(new_n708), .A2(new_n738), .A3(new_n735), .ZN(new_n911));
  OAI211_X1 g725(.A(new_n909), .B(new_n862), .C1(new_n910), .C2(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(KEYINPUT52), .ZN(new_n913));
  AND4_X1   g727(.A1(KEYINPUT53), .A2(new_n907), .A3(new_n879), .A4(new_n913), .ZN(new_n914));
  OAI21_X1  g728(.A(G902), .B1(new_n899), .B2(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(G210), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n898), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n645), .A2(new_n647), .ZN(new_n918));
  XOR2_X1   g732(.A(new_n918), .B(new_n648), .Z(new_n919));
  XNOR2_X1  g733(.A(new_n919), .B(KEYINPUT55), .ZN(new_n920));
  AND3_X1   g734(.A1(new_n917), .A2(KEYINPUT120), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g735(.A(KEYINPUT120), .B1(new_n917), .B2(new_n920), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n897), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT121), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n924), .B1(new_n884), .B2(G902), .ZN(new_n925));
  OAI211_X1 g739(.A(new_n924), .B(G902), .C1(new_n899), .C2(new_n914), .ZN(new_n926));
  INV_X1    g740(.A(new_n926), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(new_n652), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT122), .ZN(new_n930));
  INV_X1    g744(.A(new_n920), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n929), .A2(new_n930), .A3(new_n898), .A4(new_n931), .ZN(new_n932));
  NOR3_X1   g746(.A1(new_n925), .A2(new_n927), .A3(new_n651), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n931), .A2(new_n898), .ZN(new_n934));
  OAI21_X1  g748(.A(KEYINPUT122), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n923), .B1(new_n932), .B2(new_n935), .ZN(G51));
  NAND2_X1  g750(.A1(G469), .A2(G902), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n937), .B(KEYINPUT57), .Z(new_n938));
  NAND2_X1  g752(.A1(new_n885), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n939), .A2(new_n601), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n928), .A2(new_n806), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n896), .B1(new_n940), .B2(new_n941), .ZN(G54));
  NAND2_X1  g756(.A1(new_n915), .A2(KEYINPUT121), .ZN(new_n943));
  AND2_X1   g757(.A1(KEYINPUT58), .A2(G475), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n943), .A2(new_n926), .A3(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT124), .ZN(new_n946));
  INV_X1    g760(.A(new_n512), .ZN(new_n947));
  AND3_X1   g761(.A1(new_n945), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n946), .B1(new_n945), .B2(new_n947), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n897), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n943), .A2(new_n512), .A3(new_n926), .A4(new_n944), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT123), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n951), .B(new_n952), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n950), .A2(new_n953), .ZN(G60));
  NAND2_X1  g768(.A1(G478), .A2(G902), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n955), .B(KEYINPUT59), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n885), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n957), .A2(new_n665), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n958), .A2(new_n897), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n957), .A2(new_n665), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n959), .A2(new_n960), .ZN(G63));
  NAND2_X1  g775(.A1(G217), .A2(G902), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n962), .B(KEYINPUT60), .Z(new_n963));
  NAND3_X1  g777(.A1(new_n884), .A2(new_n695), .A3(new_n963), .ZN(new_n964));
  AND2_X1   g778(.A1(new_n884), .A2(new_n963), .ZN(new_n965));
  OAI211_X1 g779(.A(new_n897), .B(new_n964), .C1(new_n965), .C2(new_n393), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n966), .B(KEYINPUT61), .Z(G66));
  OAI21_X1  g781(.A(G953), .B1(new_n522), .B2(new_n626), .ZN(new_n968));
  INV_X1    g782(.A(new_n906), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n968), .B1(new_n969), .B2(G953), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n918), .B1(G898), .B2(new_n334), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n971), .B(KEYINPUT125), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n970), .B(new_n972), .ZN(G69));
  NAND3_X1  g787(.A1(new_n279), .A2(new_n282), .A3(new_n283), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n503), .A2(new_n505), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n974), .B(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n865), .A2(new_n866), .ZN(new_n977));
  AND2_X1   g791(.A1(new_n977), .A2(new_n784), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n742), .A2(new_n611), .A3(new_n722), .A4(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(new_n823), .ZN(new_n980));
  OAI211_X1 g794(.A(new_n813), .B(new_n979), .C1(new_n980), .C2(new_n821), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n859), .A2(new_n730), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n982), .B(KEYINPUT62), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n976), .B1(new_n984), .B2(G953), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n976), .B1(G900), .B2(G953), .ZN(new_n986));
  INV_X1    g800(.A(new_n810), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n987), .A2(new_n845), .A3(new_n860), .ZN(new_n988));
  AND3_X1   g802(.A1(new_n813), .A2(new_n796), .A3(new_n988), .ZN(new_n989));
  NAND4_X1  g803(.A1(new_n824), .A2(new_n794), .A3(new_n859), .A4(new_n989), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n986), .B1(new_n990), .B2(G953), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n985), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n992), .A2(KEYINPUT126), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n334), .B1(G227), .B2(G900), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT126), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n985), .A2(new_n995), .A3(new_n991), .ZN(new_n996));
  AND3_X1   g810(.A1(new_n993), .A2(new_n994), .A3(new_n996), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n994), .B1(new_n993), .B2(new_n996), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n997), .A2(new_n998), .ZN(G72));
  NAND2_X1  g813(.A1(new_n984), .A2(new_n969), .ZN(new_n1000));
  XNOR2_X1  g814(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n1001));
  NAND2_X1  g815(.A1(G472), .A2(G902), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n1001), .B(new_n1002), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1000), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1004), .A2(new_n726), .ZN(new_n1005));
  OAI211_X1 g819(.A(new_n884), .B(new_n1003), .C1(new_n295), .C2(new_n324), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n1003), .B1(new_n990), .B2(new_n906), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n1007), .A2(new_n203), .A3(new_n322), .ZN(new_n1008));
  AND4_X1   g822(.A1(new_n897), .A2(new_n1005), .A3(new_n1006), .A4(new_n1008), .ZN(G57));
endmodule


