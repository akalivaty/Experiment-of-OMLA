

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590;

  XNOR2_X1 U326 ( .A(n338), .B(n375), .ZN(n339) );
  XOR2_X1 U327 ( .A(G176GAT), .B(G64GAT), .Z(n360) );
  XNOR2_X1 U328 ( .A(n367), .B(n366), .ZN(n368) );
  XNOR2_X1 U329 ( .A(n369), .B(n368), .ZN(n373) );
  XNOR2_X1 U330 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U331 ( .A(n403), .B(n549), .Z(n588) );
  NOR2_X1 U332 ( .A1(n529), .A2(n455), .ZN(n456) );
  INV_X1 U333 ( .A(G190GAT), .ZN(n463) );
  XOR2_X1 U334 ( .A(KEYINPUT80), .B(n566), .Z(n549) );
  XNOR2_X1 U335 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U336 ( .A(n466), .B(n465), .ZN(G1351GAT) );
  XOR2_X1 U337 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n295) );
  XNOR2_X1 U338 ( .A(KEYINPUT86), .B(G183GAT), .ZN(n294) );
  XNOR2_X1 U339 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U340 ( .A(KEYINPUT19), .B(n296), .Z(n324) );
  XOR2_X1 U341 ( .A(G15GAT), .B(G127GAT), .Z(n388) );
  XOR2_X1 U342 ( .A(G113GAT), .B(KEYINPUT0), .Z(n421) );
  XOR2_X1 U343 ( .A(n388), .B(n421), .Z(n298) );
  NAND2_X1 U344 ( .A1(G227GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U345 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U346 ( .A(G120GAT), .B(G71GAT), .Z(n363) );
  XOR2_X1 U347 ( .A(n299), .B(n363), .Z(n307) );
  XOR2_X1 U348 ( .A(G99GAT), .B(G190GAT), .Z(n301) );
  XNOR2_X1 U349 ( .A(G43GAT), .B(G134GAT), .ZN(n300) );
  XNOR2_X1 U350 ( .A(n301), .B(n300), .ZN(n305) );
  XOR2_X1 U351 ( .A(G176GAT), .B(KEYINPUT85), .Z(n303) );
  XNOR2_X1 U352 ( .A(G169GAT), .B(KEYINPUT20), .ZN(n302) );
  XNOR2_X1 U353 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U354 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U355 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U356 ( .A(n324), .B(n308), .Z(n539) );
  INV_X1 U357 ( .A(n539), .ZN(n529) );
  XOR2_X1 U358 ( .A(KEYINPUT96), .B(n360), .Z(n310) );
  XOR2_X1 U359 ( .A(G169GAT), .B(G8GAT), .Z(n347) );
  XNOR2_X1 U360 ( .A(n347), .B(G92GAT), .ZN(n309) );
  XNOR2_X1 U361 ( .A(n310), .B(n309), .ZN(n320) );
  XOR2_X1 U362 ( .A(KEYINPUT97), .B(KEYINPUT95), .Z(n318) );
  XOR2_X1 U363 ( .A(KEYINPUT21), .B(G211GAT), .Z(n312) );
  XNOR2_X1 U364 ( .A(KEYINPUT88), .B(G204GAT), .ZN(n311) );
  XNOR2_X1 U365 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U366 ( .A(G197GAT), .B(n313), .Z(n452) );
  INV_X1 U367 ( .A(n452), .ZN(n316) );
  XOR2_X1 U368 ( .A(KEYINPUT79), .B(G218GAT), .Z(n315) );
  XNOR2_X1 U369 ( .A(G36GAT), .B(G190GAT), .ZN(n314) );
  XNOR2_X1 U370 ( .A(n315), .B(n314), .ZN(n333) );
  XOR2_X1 U371 ( .A(n316), .B(n333), .Z(n317) );
  XNOR2_X1 U372 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U373 ( .A(n320), .B(n319), .Z(n322) );
  NAND2_X1 U374 ( .A1(G226GAT), .A2(G233GAT), .ZN(n321) );
  XNOR2_X1 U375 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U376 ( .A(n324), .B(n323), .Z(n506) );
  INV_X1 U377 ( .A(n506), .ZN(n527) );
  XOR2_X1 U378 ( .A(KEYINPUT9), .B(KEYINPUT10), .Z(n326) );
  XNOR2_X1 U379 ( .A(KEYINPUT76), .B(KEYINPUT65), .ZN(n325) );
  XOR2_X1 U380 ( .A(n326), .B(n325), .Z(n342) );
  XOR2_X1 U381 ( .A(KEYINPUT77), .B(KEYINPUT11), .Z(n328) );
  NAND2_X1 U382 ( .A1(G232GAT), .A2(G233GAT), .ZN(n327) );
  XNOR2_X1 U383 ( .A(n328), .B(n327), .ZN(n330) );
  INV_X1 U384 ( .A(KEYINPUT64), .ZN(n329) );
  XNOR2_X1 U385 ( .A(n330), .B(n329), .ZN(n335) );
  XOR2_X1 U386 ( .A(G29GAT), .B(G43GAT), .Z(n332) );
  XNOR2_X1 U387 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n331) );
  XNOR2_X1 U388 ( .A(n332), .B(n331), .ZN(n355) );
  XNOR2_X1 U389 ( .A(n355), .B(n333), .ZN(n334) );
  XNOR2_X1 U390 ( .A(n335), .B(n334), .ZN(n340) );
  XOR2_X1 U391 ( .A(G50GAT), .B(G162GAT), .Z(n443) );
  XOR2_X1 U392 ( .A(G134GAT), .B(KEYINPUT78), .Z(n420) );
  XOR2_X1 U393 ( .A(n443), .B(n420), .Z(n338) );
  XOR2_X1 U394 ( .A(G92GAT), .B(G85GAT), .Z(n337) );
  XNOR2_X1 U395 ( .A(G99GAT), .B(G106GAT), .ZN(n336) );
  XNOR2_X1 U396 ( .A(n337), .B(n336), .ZN(n375) );
  XNOR2_X1 U397 ( .A(n342), .B(n341), .ZN(n566) );
  XOR2_X1 U398 ( .A(KEYINPUT46), .B(KEYINPUT112), .Z(n379) );
  XOR2_X1 U399 ( .A(G22GAT), .B(G141GAT), .Z(n344) );
  XNOR2_X1 U400 ( .A(G15GAT), .B(G113GAT), .ZN(n343) );
  XNOR2_X1 U401 ( .A(n344), .B(n343), .ZN(n359) );
  XOR2_X1 U402 ( .A(KEYINPUT67), .B(KEYINPUT30), .Z(n346) );
  XNOR2_X1 U403 ( .A(G197GAT), .B(KEYINPUT29), .ZN(n345) );
  XNOR2_X1 U404 ( .A(n346), .B(n345), .ZN(n351) );
  XOR2_X1 U405 ( .A(G36GAT), .B(G50GAT), .Z(n349) );
  XOR2_X1 U406 ( .A(G1GAT), .B(KEYINPUT68), .Z(n383) );
  XNOR2_X1 U407 ( .A(n383), .B(n347), .ZN(n348) );
  XNOR2_X1 U408 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U409 ( .A(n351), .B(n350), .Z(n353) );
  NAND2_X1 U410 ( .A1(G229GAT), .A2(G233GAT), .ZN(n352) );
  XNOR2_X1 U411 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U412 ( .A(n354), .B(KEYINPUT66), .Z(n357) );
  XNOR2_X1 U413 ( .A(n355), .B(KEYINPUT69), .ZN(n356) );
  XNOR2_X1 U414 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U415 ( .A(n359), .B(n358), .ZN(n469) );
  XOR2_X1 U416 ( .A(KEYINPUT74), .B(n360), .Z(n362) );
  XOR2_X1 U417 ( .A(G148GAT), .B(G78GAT), .Z(n440) );
  XNOR2_X1 U418 ( .A(G204GAT), .B(n440), .ZN(n361) );
  XNOR2_X1 U419 ( .A(n362), .B(n361), .ZN(n369) );
  XOR2_X1 U420 ( .A(n363), .B(KEYINPUT71), .Z(n367) );
  XOR2_X1 U421 ( .A(KEYINPUT75), .B(KEYINPUT73), .Z(n365) );
  NAND2_X1 U422 ( .A1(G230GAT), .A2(G233GAT), .ZN(n364) );
  XNOR2_X1 U423 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U424 ( .A(KEYINPUT31), .B(KEYINPUT33), .Z(n371) );
  XNOR2_X1 U425 ( .A(KEYINPUT32), .B(KEYINPUT72), .ZN(n370) );
  XNOR2_X1 U426 ( .A(n371), .B(n370), .ZN(n372) );
  XOR2_X1 U427 ( .A(n373), .B(n372), .Z(n377) );
  XNOR2_X1 U428 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n374) );
  XNOR2_X1 U429 ( .A(n374), .B(KEYINPUT70), .ZN(n386) );
  XNOR2_X1 U430 ( .A(n375), .B(n386), .ZN(n376) );
  XNOR2_X1 U431 ( .A(n377), .B(n376), .ZN(n580) );
  XNOR2_X1 U432 ( .A(n580), .B(KEYINPUT41), .ZN(n513) );
  NOR2_X1 U433 ( .A1(n469), .A2(n513), .ZN(n378) );
  XNOR2_X1 U434 ( .A(n379), .B(n378), .ZN(n400) );
  XOR2_X1 U435 ( .A(G78GAT), .B(G211GAT), .Z(n381) );
  XNOR2_X1 U436 ( .A(G183GAT), .B(G71GAT), .ZN(n380) );
  XNOR2_X1 U437 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U438 ( .A(n382), .B(G64GAT), .Z(n385) );
  XNOR2_X1 U439 ( .A(n383), .B(G8GAT), .ZN(n384) );
  XNOR2_X1 U440 ( .A(n385), .B(n384), .ZN(n387) );
  XOR2_X1 U441 ( .A(n387), .B(n386), .Z(n390) );
  XOR2_X1 U442 ( .A(G22GAT), .B(G155GAT), .Z(n446) );
  XNOR2_X1 U443 ( .A(n388), .B(n446), .ZN(n389) );
  XNOR2_X1 U444 ( .A(n390), .B(n389), .ZN(n394) );
  XOR2_X1 U445 ( .A(KEYINPUT84), .B(KEYINPUT83), .Z(n392) );
  NAND2_X1 U446 ( .A1(G231GAT), .A2(G233GAT), .ZN(n391) );
  XNOR2_X1 U447 ( .A(n392), .B(n391), .ZN(n393) );
  XOR2_X1 U448 ( .A(n394), .B(n393), .Z(n399) );
  XOR2_X1 U449 ( .A(KEYINPUT14), .B(KEYINPUT82), .Z(n396) );
  XNOR2_X1 U450 ( .A(KEYINPUT12), .B(KEYINPUT81), .ZN(n395) );
  XNOR2_X1 U451 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U452 ( .A(n397), .B(KEYINPUT15), .ZN(n398) );
  XOR2_X1 U453 ( .A(n399), .B(n398), .Z(n494) );
  AND2_X1 U454 ( .A1(n400), .A2(n494), .ZN(n401) );
  NAND2_X1 U455 ( .A1(n566), .A2(n401), .ZN(n402) );
  XNOR2_X1 U456 ( .A(n402), .B(KEYINPUT47), .ZN(n408) );
  XNOR2_X1 U457 ( .A(KEYINPUT36), .B(KEYINPUT104), .ZN(n403) );
  NOR2_X1 U458 ( .A1(n588), .A2(n494), .ZN(n404) );
  XNOR2_X1 U459 ( .A(n404), .B(KEYINPUT45), .ZN(n406) );
  INV_X1 U460 ( .A(n469), .ZN(n574) );
  NOR2_X1 U461 ( .A1(n574), .A2(n580), .ZN(n405) );
  AND2_X1 U462 ( .A1(n406), .A2(n405), .ZN(n407) );
  NOR2_X1 U463 ( .A1(n408), .A2(n407), .ZN(n409) );
  XNOR2_X1 U464 ( .A(n409), .B(KEYINPUT48), .ZN(n538) );
  NOR2_X1 U465 ( .A1(n527), .A2(n538), .ZN(n411) );
  XNOR2_X1 U466 ( .A(KEYINPUT120), .B(KEYINPUT54), .ZN(n410) );
  XNOR2_X1 U467 ( .A(n411), .B(n410), .ZN(n435) );
  XOR2_X1 U468 ( .A(KEYINPUT4), .B(KEYINPUT92), .Z(n413) );
  XNOR2_X1 U469 ( .A(G148GAT), .B(KEYINPUT5), .ZN(n412) );
  XNOR2_X1 U470 ( .A(n413), .B(n412), .ZN(n417) );
  XOR2_X1 U471 ( .A(G85GAT), .B(G155GAT), .Z(n415) );
  XNOR2_X1 U472 ( .A(G120GAT), .B(G127GAT), .ZN(n414) );
  XNOR2_X1 U473 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U474 ( .A(n417), .B(n416), .ZN(n434) );
  XOR2_X1 U475 ( .A(KEYINPUT1), .B(KEYINPUT6), .Z(n419) );
  XNOR2_X1 U476 ( .A(G1GAT), .B(G57GAT), .ZN(n418) );
  XNOR2_X1 U477 ( .A(n419), .B(n418), .ZN(n425) );
  XOR2_X1 U478 ( .A(n420), .B(G162GAT), .Z(n423) );
  XNOR2_X1 U479 ( .A(G29GAT), .B(n421), .ZN(n422) );
  XNOR2_X1 U480 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U481 ( .A(n425), .B(n424), .Z(n427) );
  NAND2_X1 U482 ( .A1(G225GAT), .A2(G233GAT), .ZN(n426) );
  XNOR2_X1 U483 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U484 ( .A(n428), .B(KEYINPUT94), .Z(n432) );
  XOR2_X1 U485 ( .A(KEYINPUT89), .B(KEYINPUT3), .Z(n430) );
  XNOR2_X1 U486 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n429) );
  XNOR2_X1 U487 ( .A(n430), .B(n429), .ZN(n442) );
  XNOR2_X1 U488 ( .A(n442), .B(KEYINPUT93), .ZN(n431) );
  XNOR2_X1 U489 ( .A(n432), .B(n431), .ZN(n433) );
  XOR2_X1 U490 ( .A(n434), .B(n433), .Z(n501) );
  INV_X1 U491 ( .A(n501), .ZN(n525) );
  NAND2_X1 U492 ( .A1(n435), .A2(n525), .ZN(n573) );
  XOR2_X1 U493 ( .A(KEYINPUT91), .B(KEYINPUT90), .Z(n437) );
  XNOR2_X1 U494 ( .A(KEYINPUT22), .B(KEYINPUT23), .ZN(n436) );
  XNOR2_X1 U495 ( .A(n437), .B(n436), .ZN(n451) );
  XOR2_X1 U496 ( .A(KEYINPUT87), .B(KEYINPUT24), .Z(n439) );
  XNOR2_X1 U497 ( .A(G218GAT), .B(G106GAT), .ZN(n438) );
  XNOR2_X1 U498 ( .A(n439), .B(n438), .ZN(n441) );
  XOR2_X1 U499 ( .A(n441), .B(n440), .Z(n449) );
  XOR2_X1 U500 ( .A(n443), .B(n442), .Z(n445) );
  NAND2_X1 U501 ( .A1(G228GAT), .A2(G233GAT), .ZN(n444) );
  XNOR2_X1 U502 ( .A(n445), .B(n444), .ZN(n447) );
  XNOR2_X1 U503 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U504 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U505 ( .A(n451), .B(n450), .ZN(n453) );
  XOR2_X1 U506 ( .A(n453), .B(n452), .Z(n478) );
  NOR2_X1 U507 ( .A1(n573), .A2(n478), .ZN(n454) );
  XNOR2_X1 U508 ( .A(n454), .B(KEYINPUT55), .ZN(n455) );
  XOR2_X1 U509 ( .A(KEYINPUT121), .B(n456), .Z(n570) );
  INV_X1 U510 ( .A(n513), .ZN(n557) );
  NAND2_X1 U511 ( .A1(n570), .A2(n557), .ZN(n459) );
  XOR2_X1 U512 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n457) );
  XNOR2_X1 U513 ( .A(n457), .B(G176GAT), .ZN(n458) );
  XNOR2_X1 U514 ( .A(n459), .B(n458), .ZN(G1349GAT) );
  INV_X1 U515 ( .A(n494), .ZN(n584) );
  NAND2_X1 U516 ( .A1(n570), .A2(n584), .ZN(n462) );
  XOR2_X1 U517 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n460) );
  XNOR2_X1 U518 ( .A(n460), .B(G183GAT), .ZN(n461) );
  XNOR2_X1 U519 ( .A(n462), .B(n461), .ZN(G1350GAT) );
  NAND2_X1 U520 ( .A1(n570), .A2(n549), .ZN(n466) );
  XOR2_X1 U521 ( .A(KEYINPUT124), .B(KEYINPUT58), .Z(n464) );
  XOR2_X1 U522 ( .A(KEYINPUT100), .B(KEYINPUT34), .Z(n468) );
  XNOR2_X1 U523 ( .A(G1GAT), .B(KEYINPUT101), .ZN(n467) );
  XNOR2_X1 U524 ( .A(n468), .B(n467), .ZN(n486) );
  NOR2_X1 U525 ( .A1(n580), .A2(n469), .ZN(n498) );
  NOR2_X1 U526 ( .A1(n529), .A2(n527), .ZN(n470) );
  NOR2_X1 U527 ( .A1(n478), .A2(n470), .ZN(n471) );
  XNOR2_X1 U528 ( .A(n471), .B(KEYINPUT25), .ZN(n475) );
  NAND2_X1 U529 ( .A1(n478), .A2(n529), .ZN(n472) );
  XNOR2_X1 U530 ( .A(n472), .B(KEYINPUT26), .ZN(n473) );
  XNOR2_X1 U531 ( .A(KEYINPUT98), .B(n473), .ZN(n572) );
  INV_X1 U532 ( .A(n572), .ZN(n554) );
  XNOR2_X1 U533 ( .A(KEYINPUT27), .B(n506), .ZN(n479) );
  NAND2_X1 U534 ( .A1(n554), .A2(n479), .ZN(n474) );
  NAND2_X1 U535 ( .A1(n475), .A2(n474), .ZN(n476) );
  XOR2_X1 U536 ( .A(KEYINPUT99), .B(n476), .Z(n477) );
  NAND2_X1 U537 ( .A1(n477), .A2(n525), .ZN(n482) );
  XOR2_X1 U538 ( .A(KEYINPUT28), .B(n478), .Z(n533) );
  INV_X1 U539 ( .A(n533), .ZN(n542) );
  NAND2_X1 U540 ( .A1(n501), .A2(n479), .ZN(n537) );
  NOR2_X1 U541 ( .A1(n542), .A2(n537), .ZN(n480) );
  NAND2_X1 U542 ( .A1(n480), .A2(n529), .ZN(n481) );
  NAND2_X1 U543 ( .A1(n482), .A2(n481), .ZN(n493) );
  OR2_X1 U544 ( .A1(n494), .A2(n549), .ZN(n483) );
  XOR2_X1 U545 ( .A(KEYINPUT16), .B(n483), .Z(n484) );
  AND2_X1 U546 ( .A1(n493), .A2(n484), .ZN(n514) );
  NAND2_X1 U547 ( .A1(n498), .A2(n514), .ZN(n491) );
  NOR2_X1 U548 ( .A1(n525), .A2(n491), .ZN(n485) );
  XOR2_X1 U549 ( .A(n486), .B(n485), .Z(G1324GAT) );
  NOR2_X1 U550 ( .A1(n527), .A2(n491), .ZN(n487) );
  XOR2_X1 U551 ( .A(G8GAT), .B(n487), .Z(G1325GAT) );
  NOR2_X1 U552 ( .A1(n529), .A2(n491), .ZN(n489) );
  XNOR2_X1 U553 ( .A(KEYINPUT102), .B(KEYINPUT35), .ZN(n488) );
  XNOR2_X1 U554 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U555 ( .A(G15GAT), .B(n490), .ZN(G1326GAT) );
  NOR2_X1 U556 ( .A1(n533), .A2(n491), .ZN(n492) );
  XOR2_X1 U557 ( .A(G22GAT), .B(n492), .Z(G1327GAT) );
  XOR2_X1 U558 ( .A(KEYINPUT106), .B(KEYINPUT38), .Z(n500) );
  NAND2_X1 U559 ( .A1(n494), .A2(n493), .ZN(n495) );
  NOR2_X1 U560 ( .A1(n588), .A2(n495), .ZN(n497) );
  XNOR2_X1 U561 ( .A(KEYINPUT37), .B(KEYINPUT105), .ZN(n496) );
  XNOR2_X1 U562 ( .A(n497), .B(n496), .ZN(n524) );
  NAND2_X1 U563 ( .A1(n498), .A2(n524), .ZN(n499) );
  XNOR2_X1 U564 ( .A(n500), .B(n499), .ZN(n511) );
  NAND2_X1 U565 ( .A1(n501), .A2(n511), .ZN(n505) );
  XOR2_X1 U566 ( .A(KEYINPUT103), .B(KEYINPUT39), .Z(n503) );
  XNOR2_X1 U567 ( .A(G29GAT), .B(KEYINPUT107), .ZN(n502) );
  XNOR2_X1 U568 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U569 ( .A(n505), .B(n504), .ZN(G1328GAT) );
  XNOR2_X1 U570 ( .A(G36GAT), .B(KEYINPUT108), .ZN(n508) );
  NAND2_X1 U571 ( .A1(n506), .A2(n511), .ZN(n507) );
  XNOR2_X1 U572 ( .A(n508), .B(n507), .ZN(G1329GAT) );
  NAND2_X1 U573 ( .A1(n511), .A2(n539), .ZN(n509) );
  XNOR2_X1 U574 ( .A(n509), .B(KEYINPUT40), .ZN(n510) );
  XNOR2_X1 U575 ( .A(G43GAT), .B(n510), .ZN(G1330GAT) );
  NAND2_X1 U576 ( .A1(n511), .A2(n542), .ZN(n512) );
  XNOR2_X1 U577 ( .A(n512), .B(G50GAT), .ZN(G1331GAT) );
  NOR2_X1 U578 ( .A1(n574), .A2(n513), .ZN(n523) );
  NAND2_X1 U579 ( .A1(n523), .A2(n514), .ZN(n520) );
  NOR2_X1 U580 ( .A1(n525), .A2(n520), .ZN(n516) );
  XNOR2_X1 U581 ( .A(KEYINPUT109), .B(KEYINPUT42), .ZN(n515) );
  XNOR2_X1 U582 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U583 ( .A(G57GAT), .B(n517), .ZN(G1332GAT) );
  NOR2_X1 U584 ( .A1(n527), .A2(n520), .ZN(n518) );
  XOR2_X1 U585 ( .A(G64GAT), .B(n518), .Z(G1333GAT) );
  NOR2_X1 U586 ( .A1(n529), .A2(n520), .ZN(n519) );
  XOR2_X1 U587 ( .A(G71GAT), .B(n519), .Z(G1334GAT) );
  NOR2_X1 U588 ( .A1(n533), .A2(n520), .ZN(n522) );
  XNOR2_X1 U589 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n521) );
  XNOR2_X1 U590 ( .A(n522), .B(n521), .ZN(G1335GAT) );
  NAND2_X1 U591 ( .A1(n524), .A2(n523), .ZN(n532) );
  NOR2_X1 U592 ( .A1(n525), .A2(n532), .ZN(n526) );
  XOR2_X1 U593 ( .A(G85GAT), .B(n526), .Z(G1336GAT) );
  NOR2_X1 U594 ( .A1(n527), .A2(n532), .ZN(n528) );
  XOR2_X1 U595 ( .A(G92GAT), .B(n528), .Z(G1337GAT) );
  NOR2_X1 U596 ( .A1(n529), .A2(n532), .ZN(n530) );
  XOR2_X1 U597 ( .A(KEYINPUT110), .B(n530), .Z(n531) );
  XNOR2_X1 U598 ( .A(G99GAT), .B(n531), .ZN(G1338GAT) );
  NOR2_X1 U599 ( .A1(n533), .A2(n532), .ZN(n535) );
  XNOR2_X1 U600 ( .A(KEYINPUT44), .B(KEYINPUT111), .ZN(n534) );
  XNOR2_X1 U601 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U602 ( .A(G106GAT), .B(n536), .ZN(G1339GAT) );
  NOR2_X1 U603 ( .A1(n538), .A2(n537), .ZN(n553) );
  NAND2_X1 U604 ( .A1(n539), .A2(n553), .ZN(n540) );
  XOR2_X1 U605 ( .A(KEYINPUT113), .B(n540), .Z(n541) );
  NOR2_X1 U606 ( .A1(n542), .A2(n541), .ZN(n550) );
  NAND2_X1 U607 ( .A1(n550), .A2(n574), .ZN(n543) );
  XNOR2_X1 U608 ( .A(n543), .B(KEYINPUT114), .ZN(n544) );
  XNOR2_X1 U609 ( .A(G113GAT), .B(n544), .ZN(G1340GAT) );
  XOR2_X1 U610 ( .A(G120GAT), .B(KEYINPUT49), .Z(n546) );
  NAND2_X1 U611 ( .A1(n550), .A2(n557), .ZN(n545) );
  XNOR2_X1 U612 ( .A(n546), .B(n545), .ZN(G1341GAT) );
  NAND2_X1 U613 ( .A1(n550), .A2(n584), .ZN(n547) );
  XNOR2_X1 U614 ( .A(n547), .B(KEYINPUT50), .ZN(n548) );
  XNOR2_X1 U615 ( .A(G127GAT), .B(n548), .ZN(G1342GAT) );
  XOR2_X1 U616 ( .A(G134GAT), .B(KEYINPUT51), .Z(n552) );
  NAND2_X1 U617 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n552), .B(n551), .ZN(G1343GAT) );
  NAND2_X1 U619 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U620 ( .A(n555), .B(KEYINPUT115), .Z(n565) );
  INV_X1 U621 ( .A(n565), .ZN(n562) );
  NAND2_X1 U622 ( .A1(n574), .A2(n562), .ZN(n556) );
  XNOR2_X1 U623 ( .A(G141GAT), .B(n556), .ZN(G1344GAT) );
  XNOR2_X1 U624 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n561) );
  XOR2_X1 U625 ( .A(KEYINPUT116), .B(KEYINPUT52), .Z(n559) );
  NAND2_X1 U626 ( .A1(n562), .A2(n557), .ZN(n558) );
  XNOR2_X1 U627 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U628 ( .A(n561), .B(n560), .ZN(G1345GAT) );
  XOR2_X1 U629 ( .A(G155GAT), .B(KEYINPUT117), .Z(n564) );
  NAND2_X1 U630 ( .A1(n562), .A2(n584), .ZN(n563) );
  XNOR2_X1 U631 ( .A(n564), .B(n563), .ZN(G1346GAT) );
  NOR2_X1 U632 ( .A1(n566), .A2(n565), .ZN(n568) );
  XNOR2_X1 U633 ( .A(KEYINPUT118), .B(KEYINPUT119), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U635 ( .A(G162GAT), .B(n569), .ZN(G1347GAT) );
  NAND2_X1 U636 ( .A1(n574), .A2(n570), .ZN(n571) );
  XNOR2_X1 U637 ( .A(G169GAT), .B(n571), .ZN(G1348GAT) );
  XOR2_X1 U638 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n576) );
  NOR2_X1 U639 ( .A1(n573), .A2(n572), .ZN(n586) );
  NAND2_X1 U640 ( .A1(n586), .A2(n574), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U642 ( .A(G197GAT), .B(n577), .ZN(G1352GAT) );
  XOR2_X1 U643 ( .A(KEYINPUT61), .B(KEYINPUT127), .Z(n579) );
  XNOR2_X1 U644 ( .A(G204GAT), .B(KEYINPUT126), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n579), .B(n578), .ZN(n583) );
  NAND2_X1 U646 ( .A1(n586), .A2(n580), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n581), .B(KEYINPUT125), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(G1353GAT) );
  NAND2_X1 U649 ( .A1(n586), .A2(n584), .ZN(n585) );
  XNOR2_X1 U650 ( .A(n585), .B(G211GAT), .ZN(G1354GAT) );
  INV_X1 U651 ( .A(n586), .ZN(n587) );
  NOR2_X1 U652 ( .A1(n588), .A2(n587), .ZN(n589) );
  XOR2_X1 U653 ( .A(KEYINPUT62), .B(n589), .Z(n590) );
  XNOR2_X1 U654 ( .A(G218GAT), .B(n590), .ZN(G1355GAT) );
endmodule

