//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 1 1 0 1 0 0 0 1 1 0 1 1 0 1 0 1 0 0 1 1 0 0 1 1 0 1 1 1 0 0 1 1 1 1 1 1 0 0 0 1 0 0 0 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:38 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n691, new_n692, new_n693,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n733, new_n735,
    new_n736, new_n737, new_n738, new_n740, new_n741, new_n742, new_n743,
    new_n745, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n765, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n831, new_n832, new_n834, new_n835,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n900, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n914, new_n915, new_n916, new_n917, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n936, new_n937,
    new_n938, new_n939, new_n941, new_n942, new_n943, new_n944, new_n946,
    new_n947, new_n948;
  INV_X1    g000(.A(KEYINPUT15), .ZN(new_n202));
  NOR2_X1   g001(.A1(G43gat), .A2(G50gat), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(G43gat), .A2(G50gat), .ZN(new_n205));
  AOI21_X1  g004(.A(new_n202), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(G29gat), .ZN(new_n208));
  INV_X1    g007(.A(G36gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NOR3_X1   g009(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n211));
  INV_X1    g010(.A(new_n211), .ZN(new_n212));
  OAI21_X1  g011(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT92), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT93), .ZN(new_n216));
  OAI211_X1 g015(.A(KEYINPUT92), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n217));
  AND3_X1   g016(.A1(new_n215), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  AOI21_X1  g017(.A(new_n216), .B1(new_n215), .B2(new_n217), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n212), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n210), .B1(new_n220), .B2(KEYINPUT94), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT94), .ZN(new_n222));
  OAI211_X1 g021(.A(new_n222), .B(new_n212), .C1(new_n218), .C2(new_n219), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n207), .B1(new_n221), .B2(new_n223), .ZN(new_n224));
  XOR2_X1   g023(.A(KEYINPUT95), .B(G50gat), .Z(new_n225));
  OAI211_X1 g024(.A(new_n202), .B(new_n205), .C1(new_n225), .C2(G43gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n215), .A2(new_n217), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(new_n212), .ZN(new_n228));
  INV_X1    g027(.A(new_n210), .ZN(new_n229));
  NAND4_X1  g028(.A1(new_n226), .A2(new_n207), .A3(new_n228), .A4(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n224), .A2(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(G15gat), .B(G22gat), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n233), .A2(G1gat), .ZN(new_n234));
  INV_X1    g033(.A(G15gat), .ZN(new_n235));
  INV_X1    g034(.A(G22gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(G15gat), .A2(G22gat), .ZN(new_n238));
  INV_X1    g037(.A(G1gat), .ZN(new_n239));
  AOI22_X1  g038(.A1(new_n237), .A2(new_n238), .B1(KEYINPUT16), .B2(new_n239), .ZN(new_n240));
  OAI21_X1  g039(.A(KEYINPUT97), .B1(new_n234), .B2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(G8gat), .ZN(new_n242));
  OR2_X1    g041(.A1(new_n240), .A2(KEYINPUT97), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n241), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT98), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n241), .A2(new_n243), .A3(KEYINPUT98), .A4(new_n242), .ZN(new_n247));
  OR2_X1    g046(.A1(new_n234), .A2(new_n240), .ZN(new_n248));
  AOI22_X1  g047(.A1(new_n246), .A2(new_n247), .B1(G8gat), .B2(new_n248), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n232), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT17), .ZN(new_n251));
  OR2_X1    g050(.A1(new_n251), .A2(KEYINPUT96), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(KEYINPUT96), .ZN(new_n253));
  OAI211_X1 g052(.A(new_n252), .B(new_n253), .C1(new_n224), .C2(new_n231), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n227), .A2(KEYINPUT93), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n215), .A2(new_n216), .A3(new_n217), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n211), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n229), .B1(new_n257), .B2(new_n222), .ZN(new_n258));
  INV_X1    g057(.A(new_n223), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n206), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND4_X1  g059(.A1(new_n260), .A2(KEYINPUT96), .A3(new_n251), .A4(new_n230), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n254), .A2(new_n261), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n250), .B1(new_n262), .B2(new_n249), .ZN(new_n263));
  NAND2_X1  g062(.A1(G229gat), .A2(G233gat), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT99), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n264), .B1(new_n265), .B2(KEYINPUT18), .ZN(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n263), .A2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT18), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n269), .A2(KEYINPUT99), .ZN(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n268), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n249), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n273), .B1(new_n254), .B2(new_n261), .ZN(new_n274));
  NOR4_X1   g073(.A1(new_n274), .A2(new_n250), .A3(new_n271), .A4(new_n266), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n230), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n277), .B(new_n249), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n264), .B(KEYINPUT13), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n272), .A2(new_n276), .A3(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(G113gat), .B(G141gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n283), .B(G197gat), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n284), .B(KEYINPUT11), .ZN(new_n285));
  INV_X1    g084(.A(G169gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n285), .B(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(KEYINPUT91), .B(KEYINPUT12), .ZN(new_n288));
  XOR2_X1   g087(.A(new_n287), .B(new_n288), .Z(new_n289));
  NAND2_X1  g088(.A1(new_n282), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n270), .B1(new_n263), .B2(new_n267), .ZN(new_n291));
  NOR3_X1   g090(.A1(new_n291), .A2(new_n275), .A3(new_n280), .ZN(new_n292));
  INV_X1    g091(.A(new_n289), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n290), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(G71gat), .A2(G78gat), .ZN(new_n297));
  OR2_X1    g096(.A1(G71gat), .A2(G78gat), .ZN(new_n298));
  XNOR2_X1  g097(.A(G57gat), .B(G64gat), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT9), .ZN(new_n300));
  OAI211_X1 g099(.A(new_n297), .B(new_n298), .C1(new_n299), .C2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT101), .ZN(new_n302));
  NAND2_X1  g101(.A1(KEYINPUT100), .A2(G57gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(G64gat), .ZN(new_n304));
  INV_X1    g103(.A(G64gat), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n305), .A2(KEYINPUT100), .A3(G57gat), .ZN(new_n306));
  AOI22_X1  g105(.A1(new_n304), .A2(new_n306), .B1(new_n298), .B2(new_n297), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n297), .A2(new_n300), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n302), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n304), .A2(new_n306), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n298), .A2(new_n297), .ZN(new_n311));
  AND4_X1   g110(.A1(new_n302), .A2(new_n310), .A3(new_n308), .A4(new_n311), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n301), .B1(new_n309), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(G85gat), .A2(G92gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(KEYINPUT7), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT7), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n316), .A2(G85gat), .A3(G92gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  XNOR2_X1  g117(.A(G99gat), .B(G106gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(G99gat), .A2(G106gat), .ZN(new_n320));
  INV_X1    g119(.A(G85gat), .ZN(new_n321));
  INV_X1    g120(.A(G92gat), .ZN(new_n322));
  AOI22_X1  g121(.A1(KEYINPUT8), .A2(new_n320), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  AND3_X1   g122(.A1(new_n318), .A2(new_n319), .A3(new_n323), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n319), .B1(new_n318), .B2(new_n323), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n313), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT10), .ZN(new_n329));
  OAI211_X1 g128(.A(new_n326), .B(new_n301), .C1(new_n309), .C2(new_n312), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n328), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(new_n313), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n332), .A2(KEYINPUT10), .A3(new_n326), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(G230gat), .A2(G233gat), .ZN(new_n335));
  XOR2_X1   g134(.A(new_n335), .B(KEYINPUT105), .Z(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n334), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n328), .A2(new_n330), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(new_n336), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  XNOR2_X1  g140(.A(G120gat), .B(G148gat), .ZN(new_n342));
  XNOR2_X1  g141(.A(new_n342), .B(KEYINPUT106), .ZN(new_n343));
  INV_X1    g142(.A(G176gat), .ZN(new_n344));
  XNOR2_X1  g143(.A(new_n343), .B(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(G204gat), .ZN(new_n346));
  XNOR2_X1  g145(.A(new_n345), .B(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n341), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n338), .A2(new_n340), .A3(new_n347), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n296), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n332), .A2(KEYINPUT21), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n249), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(KEYINPUT104), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT104), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n249), .A2(new_n357), .A3(new_n354), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(G231gat), .ZN(new_n360));
  INV_X1    g159(.A(G233gat), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n359), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND4_X1  g161(.A1(new_n356), .A2(G231gat), .A3(G233gat), .A4(new_n358), .ZN(new_n363));
  XNOR2_X1  g162(.A(KEYINPUT102), .B(KEYINPUT103), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n362), .A2(new_n363), .A3(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n365), .B1(new_n362), .B2(new_n363), .ZN(new_n368));
  XOR2_X1   g167(.A(G127gat), .B(G155gat), .Z(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n332), .A2(KEYINPUT21), .ZN(new_n371));
  XNOR2_X1  g170(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n372));
  XNOR2_X1  g171(.A(new_n371), .B(new_n372), .ZN(new_n373));
  XNOR2_X1  g172(.A(G183gat), .B(G211gat), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(new_n372), .ZN(new_n376));
  XNOR2_X1  g175(.A(new_n371), .B(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(new_n374), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n370), .B1(new_n375), .B2(new_n379), .ZN(new_n380));
  AND3_X1   g179(.A1(new_n375), .A2(new_n379), .A3(new_n370), .ZN(new_n381));
  OAI22_X1  g180(.A1(new_n367), .A2(new_n368), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(new_n368), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n381), .A2(new_n380), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n383), .A2(new_n384), .A3(new_n366), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n382), .A2(new_n385), .ZN(new_n386));
  AOI21_X1  g185(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n387));
  XNOR2_X1  g186(.A(new_n387), .B(G162gat), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  XNOR2_X1  g188(.A(G190gat), .B(G218gat), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n262), .A2(new_n327), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n232), .A2(new_n327), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n392), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(G134gat), .ZN(new_n397));
  INV_X1    g196(.A(new_n395), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n398), .B1(new_n262), .B2(new_n327), .ZN(new_n399));
  INV_X1    g198(.A(G134gat), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n399), .A2(new_n400), .A3(new_n394), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n391), .B1(new_n397), .B2(new_n401), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n400), .B1(new_n399), .B2(new_n394), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n326), .B1(new_n254), .B2(new_n261), .ZN(new_n404));
  NOR4_X1   g203(.A1(new_n404), .A2(G134gat), .A3(new_n393), .A4(new_n398), .ZN(new_n405));
  NOR3_X1   g204(.A1(new_n403), .A2(new_n405), .A3(new_n390), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n389), .B1(new_n402), .B2(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n397), .A2(new_n401), .A3(new_n391), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n390), .B1(new_n403), .B2(new_n405), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n408), .A2(new_n409), .A3(new_n388), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n386), .A2(new_n407), .A3(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT73), .ZN(new_n412));
  INV_X1    g211(.A(G148gat), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n412), .B1(new_n413), .B2(G141gat), .ZN(new_n414));
  INV_X1    g213(.A(G141gat), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n415), .A2(KEYINPUT73), .A3(G148gat), .ZN(new_n416));
  OAI211_X1 g215(.A(new_n414), .B(new_n416), .C1(new_n415), .C2(G148gat), .ZN(new_n417));
  OR3_X1    g216(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n418));
  NAND2_X1  g217(.A1(G155gat), .A2(G162gat), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n417), .A2(new_n420), .ZN(new_n421));
  XNOR2_X1  g220(.A(G141gat), .B(G148gat), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT2), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n423), .A2(KEYINPUT72), .ZN(new_n424));
  OAI22_X1  g223(.A1(new_n422), .A2(new_n424), .B1(G155gat), .B2(G162gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(new_n419), .B(KEYINPUT72), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n421), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  XNOR2_X1  g226(.A(G197gat), .B(G204gat), .ZN(new_n428));
  AND2_X1   g227(.A1(G211gat), .A2(G218gat), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n428), .B1(KEYINPUT22), .B2(new_n429), .ZN(new_n430));
  XNOR2_X1  g229(.A(G211gat), .B(G218gat), .ZN(new_n431));
  XNOR2_X1  g230(.A(new_n430), .B(new_n431), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n432), .A2(KEYINPUT29), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n427), .B1(new_n433), .B2(KEYINPUT3), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT3), .ZN(new_n436));
  OAI211_X1 g235(.A(new_n421), .B(new_n436), .C1(new_n425), .C2(new_n426), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT29), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  AND2_X1   g238(.A1(new_n439), .A2(new_n432), .ZN(new_n440));
  INV_X1    g239(.A(G228gat), .ZN(new_n441));
  OAI22_X1  g240(.A1(new_n435), .A2(new_n440), .B1(new_n441), .B2(new_n361), .ZN(new_n442));
  INV_X1    g241(.A(new_n432), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n439), .A2(KEYINPUT81), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT81), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n437), .A2(new_n445), .A3(new_n438), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n443), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT82), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n441), .A2(new_n361), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n434), .B1(new_n447), .B2(new_n448), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n442), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(G22gat), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT83), .ZN(new_n455));
  OAI211_X1 g254(.A(new_n442), .B(new_n236), .C1(new_n451), .C2(new_n452), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n454), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  XOR2_X1   g256(.A(KEYINPUT80), .B(G50gat), .Z(new_n458));
  XNOR2_X1  g257(.A(G78gat), .B(G106gat), .ZN(new_n459));
  XNOR2_X1  g258(.A(new_n458), .B(new_n459), .ZN(new_n460));
  XOR2_X1   g259(.A(KEYINPUT79), .B(KEYINPUT31), .Z(new_n461));
  XNOR2_X1  g260(.A(new_n460), .B(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n453), .A2(KEYINPUT83), .A3(G22gat), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n457), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT85), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n462), .B1(new_n456), .B2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT84), .ZN(new_n467));
  OAI211_X1 g266(.A(new_n467), .B(G22gat), .C1(new_n453), .C2(new_n465), .ZN(new_n468));
  OR2_X1    g267(.A1(new_n451), .A2(new_n452), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n467), .A2(G22gat), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n469), .A2(KEYINPUT85), .A3(new_n442), .A4(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n466), .A2(new_n468), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n464), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(KEYINPUT86), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT86), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n464), .A2(new_n472), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT68), .ZN(new_n478));
  NAND2_X1  g277(.A1(G183gat), .A2(G190gat), .ZN(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(KEYINPUT24), .ZN(new_n481));
  AND2_X1   g280(.A1(KEYINPUT64), .A2(KEYINPUT24), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n479), .B1(KEYINPUT64), .B2(KEYINPUT24), .ZN(new_n483));
  OAI221_X1 g282(.A(new_n481), .B1(G183gat), .B2(G190gat), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  OR3_X1    g283(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n485));
  OAI21_X1  g284(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n486));
  AOI22_X1  g285(.A1(new_n485), .A2(new_n486), .B1(G169gat), .B2(G176gat), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n484), .A2(KEYINPUT25), .A3(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT65), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n481), .B1(G183gat), .B2(G190gat), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n480), .A2(KEYINPUT24), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n487), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT25), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n484), .A2(KEYINPUT65), .A3(KEYINPUT25), .A4(new_n487), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n490), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  XOR2_X1   g296(.A(KEYINPUT27), .B(G183gat), .Z(new_n498));
  OAI21_X1  g297(.A(KEYINPUT28), .B1(new_n498), .B2(G190gat), .ZN(new_n499));
  INV_X1    g298(.A(G183gat), .ZN(new_n500));
  OR3_X1    g299(.A1(new_n500), .A2(KEYINPUT66), .A3(KEYINPUT27), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT28), .ZN(new_n502));
  INV_X1    g301(.A(G190gat), .ZN(new_n503));
  OAI21_X1  g302(.A(KEYINPUT27), .B1(new_n500), .B2(KEYINPUT66), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n501), .A2(new_n502), .A3(new_n503), .A4(new_n504), .ZN(new_n505));
  OR3_X1    g304(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n506));
  OAI21_X1  g305(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n507));
  OAI211_X1 g306(.A(new_n506), .B(new_n507), .C1(new_n286), .C2(new_n344), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n499), .A2(new_n479), .A3(new_n505), .A4(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n497), .A2(new_n509), .ZN(new_n510));
  XOR2_X1   g309(.A(G113gat), .B(G120gat), .Z(new_n511));
  INV_X1    g310(.A(KEYINPUT1), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT67), .ZN(new_n515));
  INV_X1    g314(.A(G127gat), .ZN(new_n516));
  NOR3_X1   g315(.A1(new_n515), .A2(new_n516), .A3(G134gat), .ZN(new_n517));
  XNOR2_X1  g316(.A(G127gat), .B(G134gat), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n517), .B1(new_n515), .B2(new_n518), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n514), .A2(new_n519), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n513), .A2(new_n518), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n478), .B1(new_n510), .B2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(new_n521), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n525), .B1(new_n514), .B2(new_n519), .ZN(new_n526));
  AOI211_X1 g325(.A(KEYINPUT68), .B(new_n526), .C1(new_n497), .C2(new_n509), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n510), .A2(new_n522), .ZN(new_n529));
  INV_X1    g328(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(G227gat), .A2(G233gat), .ZN(new_n531));
  NAND4_X1  g330(.A1(new_n524), .A2(new_n528), .A3(new_n530), .A4(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT34), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n532), .B(new_n533), .ZN(new_n534));
  XNOR2_X1  g333(.A(G15gat), .B(G43gat), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n535), .B(G71gat), .ZN(new_n536));
  XOR2_X1   g335(.A(new_n536), .B(G99gat), .Z(new_n537));
  OR2_X1    g336(.A1(new_n537), .A2(KEYINPUT69), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(KEYINPUT69), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n538), .A2(new_n539), .A3(KEYINPUT33), .ZN(new_n540));
  NOR3_X1   g339(.A1(new_n523), .A2(new_n527), .A3(new_n529), .ZN(new_n541));
  OAI211_X1 g340(.A(KEYINPUT32), .B(new_n540), .C1(new_n541), .C2(new_n531), .ZN(new_n542));
  INV_X1    g341(.A(new_n537), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n524), .A2(new_n528), .A3(new_n530), .ZN(new_n544));
  INV_X1    g343(.A(new_n531), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT32), .ZN(new_n546));
  AOI22_X1  g345(.A1(new_n544), .A2(new_n545), .B1(new_n546), .B2(KEYINPUT33), .ZN(new_n547));
  OAI211_X1 g346(.A(new_n534), .B(new_n542), .C1(new_n543), .C2(new_n547), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n542), .B1(new_n547), .B2(new_n543), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n532), .B(KEYINPUT34), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n548), .A2(KEYINPUT70), .A3(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT70), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n549), .A2(new_n553), .A3(new_n550), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT35), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n477), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  AND2_X1   g356(.A1(G226gat), .A2(G233gat), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n510), .A2(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(KEYINPUT29), .B1(new_n497), .B2(new_n509), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n559), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(new_n432), .ZN(new_n562));
  OAI211_X1 g361(.A(new_n559), .B(new_n443), .C1(new_n558), .C2(new_n560), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n562), .A2(KEYINPUT71), .A3(new_n563), .ZN(new_n564));
  OR2_X1    g363(.A1(new_n563), .A2(KEYINPUT71), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(G8gat), .B(G36gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(new_n305), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n568), .B(new_n322), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n566), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n564), .A2(new_n565), .A3(new_n569), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n571), .A2(KEYINPUT30), .A3(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT30), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n566), .A2(new_n574), .A3(new_n570), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT74), .ZN(new_n577));
  OAI211_X1 g376(.A(new_n525), .B(new_n577), .C1(new_n514), .C2(new_n519), .ZN(new_n578));
  OAI21_X1  g377(.A(KEYINPUT74), .B1(new_n520), .B2(new_n521), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n427), .A2(KEYINPUT3), .ZN(new_n580));
  NAND4_X1  g379(.A1(new_n578), .A2(new_n579), .A3(new_n580), .A4(new_n437), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(G225gat), .A2(G233gat), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(KEYINPUT76), .B(KEYINPUT5), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n522), .A2(new_n427), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT4), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n427), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n526), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n592), .A2(KEYINPUT4), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT78), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n590), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n594), .B1(new_n590), .B2(new_n593), .ZN(new_n597));
  OAI211_X1 g396(.A(new_n585), .B(new_n587), .C1(new_n596), .C2(new_n597), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n578), .A2(new_n579), .A3(new_n427), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(KEYINPUT75), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT75), .ZN(new_n601));
  NAND4_X1  g400(.A1(new_n578), .A2(new_n579), .A3(new_n601), .A4(new_n427), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n600), .A2(new_n592), .A3(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n587), .B1(new_n603), .B2(new_n584), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT77), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n588), .A2(new_n589), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n592), .A2(KEYINPUT4), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n585), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  AND3_X1   g407(.A1(new_n604), .A2(new_n605), .A3(new_n608), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n605), .B1(new_n604), .B2(new_n608), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n598), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(G1gat), .B(G29gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(KEYINPUT0), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(G57gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(new_n321), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n611), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT6), .ZN(new_n618));
  OAI211_X1 g417(.A(new_n615), .B(new_n598), .C1(new_n609), .C2(new_n610), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n617), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n611), .A2(KEYINPUT6), .A3(new_n616), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n576), .B1(new_n621), .B2(new_n623), .ZN(new_n624));
  OAI21_X1  g423(.A(KEYINPUT90), .B1(new_n557), .B2(new_n624), .ZN(new_n625));
  AND2_X1   g424(.A1(new_n548), .A2(new_n551), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n477), .A2(new_n626), .ZN(new_n627));
  OAI21_X1  g426(.A(KEYINPUT35), .B1(new_n627), .B2(new_n624), .ZN(new_n628));
  INV_X1    g427(.A(new_n576), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n629), .B1(new_n622), .B2(new_n620), .ZN(new_n630));
  AOI22_X1  g429(.A1(new_n474), .A2(new_n476), .B1(new_n552), .B2(new_n554), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT90), .ZN(new_n632));
  NAND4_X1  g431(.A1(new_n630), .A2(new_n631), .A3(new_n632), .A4(new_n556), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n625), .A2(new_n628), .A3(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT89), .ZN(new_n635));
  OR2_X1    g434(.A1(new_n603), .A2(new_n584), .ZN(new_n636));
  OAI21_X1  g435(.A(KEYINPUT78), .B1(new_n606), .B2(new_n607), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n582), .B1(new_n637), .B2(new_n595), .ZN(new_n638));
  OAI211_X1 g437(.A(new_n636), .B(KEYINPUT39), .C1(new_n638), .C2(new_n583), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n581), .B1(new_n596), .B2(new_n597), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT39), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n640), .A2(new_n641), .A3(new_n584), .ZN(new_n642));
  NAND4_X1  g441(.A1(new_n639), .A2(KEYINPUT40), .A3(new_n642), .A4(new_n615), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT87), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n638), .A2(new_n583), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n616), .B1(new_n646), .B2(new_n641), .ZN(new_n647));
  NAND4_X1  g446(.A1(new_n647), .A2(KEYINPUT87), .A3(KEYINPUT40), .A4(new_n639), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n649), .A2(new_n617), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n647), .A2(new_n639), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT40), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n653), .A2(new_n575), .A3(new_n573), .ZN(new_n654));
  INV_X1    g453(.A(new_n476), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n475), .B1(new_n464), .B2(new_n472), .ZN(new_n656));
  OAI22_X1  g455(.A1(new_n650), .A2(new_n654), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  XOR2_X1   g456(.A(KEYINPUT88), .B(KEYINPUT37), .Z(new_n658));
  NAND2_X1  g457(.A1(new_n566), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n562), .A2(new_n563), .ZN(new_n660));
  AOI21_X1  g459(.A(KEYINPUT38), .B1(new_n660), .B2(KEYINPUT37), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n659), .A2(new_n569), .A3(new_n661), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n620), .A2(new_n622), .A3(new_n662), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n564), .A2(new_n565), .A3(KEYINPUT37), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n659), .A2(new_n569), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n665), .A2(KEYINPUT38), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n666), .A2(new_n571), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n663), .A2(new_n667), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n635), .B1(new_n657), .B2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n477), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n626), .A2(KEYINPUT36), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT36), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n552), .A2(new_n672), .A3(new_n554), .ZN(new_n673));
  AOI22_X1  g472(.A1(new_n670), .A2(new_n624), .B1(new_n671), .B2(new_n673), .ZN(new_n674));
  NAND4_X1  g473(.A1(new_n629), .A2(new_n617), .A3(new_n649), .A4(new_n653), .ZN(new_n675));
  AOI22_X1  g474(.A1(new_n665), .A2(KEYINPUT38), .B1(new_n566), .B2(new_n570), .ZN(new_n676));
  NAND4_X1  g475(.A1(new_n676), .A2(new_n622), .A3(new_n620), .A4(new_n662), .ZN(new_n677));
  NAND4_X1  g476(.A1(new_n675), .A2(new_n677), .A3(KEYINPUT89), .A4(new_n477), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n669), .A2(new_n674), .A3(new_n678), .ZN(new_n679));
  AOI211_X1 g478(.A(new_n353), .B(new_n411), .C1(new_n634), .C2(new_n679), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n621), .A2(new_n623), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g482(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n680), .A2(new_n629), .A3(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT16), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n685), .B1(new_n686), .B2(new_n242), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n242), .B1(new_n680), .B2(new_n629), .ZN(new_n688));
  OAI21_X1  g487(.A(KEYINPUT42), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n689), .B1(KEYINPUT42), .B2(new_n687), .ZN(G1325gat));
  AOI21_X1  g489(.A(G15gat), .B1(new_n680), .B2(new_n555), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n671), .A2(new_n673), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n692), .A2(new_n235), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n691), .B1(new_n680), .B2(new_n693), .ZN(G1326gat));
  NAND2_X1  g493(.A1(new_n680), .A2(new_n670), .ZN(new_n695));
  XNOR2_X1  g494(.A(KEYINPUT43), .B(G22gat), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n695), .B(new_n696), .ZN(G1327gat));
  NAND2_X1  g496(.A1(new_n634), .A2(new_n679), .ZN(new_n698));
  INV_X1    g497(.A(new_n386), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n407), .A2(new_n410), .ZN(new_n700));
  AND4_X1   g499(.A1(new_n352), .A2(new_n698), .A3(new_n699), .A4(new_n700), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n701), .A2(new_n208), .A3(new_n681), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(KEYINPUT45), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n386), .B(KEYINPUT107), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n351), .B(KEYINPUT108), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  AND2_X1   g505(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT44), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n708), .B1(new_n698), .B2(new_n700), .ZN(new_n709));
  INV_X1    g508(.A(new_n700), .ZN(new_n710));
  AOI211_X1 g509(.A(KEYINPUT44), .B(new_n710), .C1(new_n634), .C2(new_n679), .ZN(new_n711));
  OAI211_X1 g510(.A(new_n295), .B(new_n707), .C1(new_n709), .C2(new_n711), .ZN(new_n712));
  NOR3_X1   g511(.A1(new_n712), .A2(new_n623), .A3(new_n621), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n703), .B1(new_n208), .B2(new_n713), .ZN(G1328gat));
  NAND3_X1  g513(.A1(new_n701), .A2(new_n209), .A3(new_n629), .ZN(new_n715));
  XOR2_X1   g514(.A(new_n715), .B(KEYINPUT46), .Z(new_n716));
  OAI21_X1  g515(.A(G36gat), .B1(new_n712), .B2(new_n576), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(G1329gat));
  OAI21_X1  g517(.A(G43gat), .B1(new_n712), .B2(new_n692), .ZN(new_n719));
  INV_X1    g518(.A(G43gat), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n701), .A2(new_n720), .A3(new_n555), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT47), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n722), .B(new_n723), .ZN(G1330gat));
  OAI21_X1  g523(.A(new_n225), .B1(new_n712), .B2(new_n477), .ZN(new_n725));
  INV_X1    g524(.A(new_n225), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n701), .A2(new_n726), .A3(new_n670), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT48), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n728), .B(new_n729), .ZN(G1331gat));
  INV_X1    g529(.A(new_n411), .ZN(new_n731));
  AND4_X1   g530(.A1(new_n296), .A2(new_n698), .A3(new_n731), .A4(new_n705), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(new_n681), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g533(.A(new_n576), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(KEYINPUT109), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n732), .A2(new_n736), .ZN(new_n737));
  NOR2_X1   g536(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n738));
  XOR2_X1   g537(.A(new_n737), .B(new_n738), .Z(G1333gat));
  INV_X1    g538(.A(new_n692), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n732), .A2(new_n740), .ZN(new_n741));
  AOI21_X1  g540(.A(G71gat), .B1(new_n552), .B2(new_n554), .ZN(new_n742));
  AOI22_X1  g541(.A1(new_n741), .A2(G71gat), .B1(new_n732), .B2(new_n742), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g543(.A1(new_n732), .A2(new_n670), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(G78gat), .ZN(G1335gat));
  INV_X1    g545(.A(new_n351), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n295), .A2(new_n747), .ZN(new_n748));
  OAI211_X1 g547(.A(new_n699), .B(new_n748), .C1(new_n709), .C2(new_n711), .ZN(new_n749));
  NOR3_X1   g548(.A1(new_n749), .A2(new_n623), .A3(new_n621), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n698), .A2(new_n296), .A3(new_n699), .A4(new_n700), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT51), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n751), .B(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(new_n753), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n681), .A2(new_n321), .A3(new_n351), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(KEYINPUT110), .ZN(new_n756));
  OAI22_X1  g555(.A1(new_n750), .A2(new_n321), .B1(new_n754), .B2(new_n756), .ZN(G1336gat));
  NAND4_X1  g556(.A1(new_n753), .A2(new_n322), .A3(new_n629), .A4(new_n705), .ZN(new_n758));
  OAI21_X1  g557(.A(G92gat), .B1(new_n749), .B2(new_n576), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(KEYINPUT52), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT52), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n758), .A2(new_n762), .A3(new_n759), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n761), .A2(new_n763), .ZN(G1337gat));
  XNOR2_X1  g563(.A(KEYINPUT111), .B(G99gat), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n765), .B1(new_n749), .B2(new_n692), .ZN(new_n766));
  INV_X1    g565(.A(new_n765), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n555), .A2(new_n351), .A3(new_n767), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n766), .B1(new_n754), .B2(new_n768), .ZN(G1338gat));
  INV_X1    g568(.A(new_n709), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n698), .A2(new_n708), .A3(new_n700), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n386), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT114), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n772), .A2(new_n773), .A3(new_n670), .A4(new_n748), .ZN(new_n774));
  OAI21_X1  g573(.A(KEYINPUT114), .B1(new_n749), .B2(new_n477), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n774), .A2(new_n775), .A3(G106gat), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT53), .ZN(new_n777));
  NOR3_X1   g576(.A1(new_n477), .A2(G106gat), .A3(new_n706), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n778), .B(KEYINPUT112), .ZN(new_n779));
  AND2_X1   g578(.A1(new_n751), .A2(new_n752), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n751), .A2(new_n752), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n779), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n776), .A2(new_n777), .A3(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT113), .ZN(new_n784));
  OAI21_X1  g583(.A(G106gat), .B1(new_n749), .B2(new_n477), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(new_n782), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n784), .B1(new_n786), .B2(KEYINPUT53), .ZN(new_n787));
  AOI211_X1 g586(.A(KEYINPUT113), .B(new_n777), .C1(new_n785), .C2(new_n782), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n783), .B1(new_n787), .B2(new_n788), .ZN(G1339gat));
  AOI21_X1  g588(.A(new_n336), .B1(new_n331), .B2(new_n333), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT54), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n347), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(new_n792), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n331), .A2(new_n333), .A3(new_n336), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n338), .A2(KEYINPUT54), .A3(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT115), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n338), .A2(KEYINPUT115), .A3(KEYINPUT54), .A4(new_n794), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n793), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n350), .B1(new_n799), .B2(KEYINPUT55), .ZN(new_n800));
  AND3_X1   g599(.A1(new_n331), .A2(new_n333), .A3(new_n336), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n801), .A2(new_n790), .ZN(new_n802));
  AOI21_X1  g601(.A(KEYINPUT115), .B1(new_n802), .B2(KEYINPUT54), .ZN(new_n803));
  INV_X1    g602(.A(new_n798), .ZN(new_n804));
  OAI211_X1 g603(.A(KEYINPUT55), .B(new_n792), .C1(new_n803), .C2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT116), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n799), .A2(KEYINPUT116), .A3(KEYINPUT55), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n800), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n278), .A2(new_n279), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n810), .B1(new_n264), .B2(new_n263), .ZN(new_n811));
  AOI22_X1  g610(.A1(new_n292), .A2(new_n293), .B1(new_n287), .B2(new_n811), .ZN(new_n812));
  AND3_X1   g611(.A1(new_n408), .A2(new_n409), .A3(new_n388), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n388), .B1(new_n408), .B2(new_n409), .ZN(new_n814));
  OAI211_X1 g613(.A(new_n809), .B(new_n812), .C1(new_n813), .C2(new_n814), .ZN(new_n815));
  AOI22_X1  g614(.A1(new_n295), .A2(new_n809), .B1(new_n812), .B2(new_n351), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n815), .B1(new_n816), .B2(new_n700), .ZN(new_n817));
  AND2_X1   g616(.A1(new_n817), .A2(new_n704), .ZN(new_n818));
  NOR3_X1   g617(.A1(new_n411), .A2(new_n351), .A3(new_n295), .ZN(new_n819));
  OR2_X1    g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(new_n681), .ZN(new_n821));
  INV_X1    g620(.A(new_n631), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n821), .A2(new_n629), .A3(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(G113gat), .B1(new_n824), .B2(new_n296), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n821), .A2(new_n629), .ZN(new_n826));
  INV_X1    g625(.A(new_n627), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  OR2_X1    g627(.A1(new_n296), .A2(G113gat), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n825), .B1(new_n828), .B2(new_n829), .ZN(G1340gat));
  OAI21_X1  g629(.A(G120gat), .B1(new_n824), .B2(new_n706), .ZN(new_n831));
  OR2_X1    g630(.A1(new_n747), .A2(G120gat), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n831), .B1(new_n828), .B2(new_n832), .ZN(G1341gat));
  NAND3_X1  g632(.A1(new_n826), .A2(new_n386), .A3(new_n827), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n704), .A2(new_n516), .ZN(new_n835));
  AOI22_X1  g634(.A1(new_n834), .A2(new_n516), .B1(new_n823), .B2(new_n835), .ZN(G1342gat));
  NAND2_X1  g635(.A1(new_n700), .A2(new_n576), .ZN(new_n837));
  NOR4_X1   g636(.A1(new_n821), .A2(G134gat), .A3(new_n627), .A4(new_n837), .ZN(new_n838));
  XNOR2_X1  g637(.A(new_n838), .B(KEYINPUT56), .ZN(new_n839));
  OAI21_X1  g638(.A(G134gat), .B1(new_n824), .B2(new_n710), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n840), .A2(KEYINPUT117), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n840), .A2(KEYINPUT117), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n839), .B1(new_n841), .B2(new_n842), .ZN(G1343gat));
  INV_X1    g642(.A(KEYINPUT58), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n819), .B1(new_n817), .B2(new_n699), .ZN(new_n845));
  OAI21_X1  g644(.A(KEYINPUT57), .B1(new_n845), .B2(new_n477), .ZN(new_n846));
  AND3_X1   g645(.A1(new_n692), .A2(new_n681), .A3(new_n576), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n820), .A2(new_n670), .ZN(new_n848));
  OAI211_X1 g647(.A(new_n846), .B(new_n847), .C1(new_n848), .C2(KEYINPUT57), .ZN(new_n849));
  OAI21_X1  g648(.A(G141gat), .B1(new_n849), .B2(new_n296), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n844), .B1(new_n850), .B2(KEYINPUT120), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT118), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n821), .A2(new_n852), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n740), .A2(new_n477), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n820), .A2(KEYINPUT118), .A3(new_n681), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n853), .A2(new_n576), .A3(new_n854), .A4(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n295), .A2(new_n415), .ZN(new_n857));
  XOR2_X1   g656(.A(new_n857), .B(KEYINPUT119), .Z(new_n858));
  OAI21_X1  g657(.A(new_n850), .B1(new_n856), .B2(new_n858), .ZN(new_n859));
  XNOR2_X1  g658(.A(new_n851), .B(new_n859), .ZN(G1344gat));
  INV_X1    g659(.A(KEYINPUT59), .ZN(new_n861));
  OAI211_X1 g660(.A(new_n861), .B(G148gat), .C1(new_n849), .C2(new_n747), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT123), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT121), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n812), .A2(new_n351), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n807), .A2(new_n808), .ZN(new_n866));
  INV_X1    g665(.A(new_n800), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n291), .A2(new_n275), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n293), .B1(new_n868), .B2(new_n281), .ZN(new_n869));
  NOR4_X1   g668(.A1(new_n291), .A2(new_n275), .A3(new_n280), .A4(new_n289), .ZN(new_n870));
  OAI211_X1 g669(.A(new_n866), .B(new_n867), .C1(new_n869), .C2(new_n870), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n700), .B1(new_n865), .B2(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(new_n815), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n699), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(new_n819), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n477), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n864), .B1(new_n876), .B2(KEYINPUT57), .ZN(new_n877));
  OAI211_X1 g676(.A(KEYINPUT57), .B(new_n670), .C1(new_n818), .C2(new_n819), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT57), .ZN(new_n879));
  OAI211_X1 g678(.A(KEYINPUT121), .B(new_n879), .C1(new_n845), .C2(new_n477), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n877), .A2(new_n878), .A3(new_n880), .ZN(new_n881));
  AND2_X1   g680(.A1(new_n847), .A2(new_n351), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT122), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n413), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n881), .A2(KEYINPUT122), .A3(new_n882), .ZN(new_n886));
  AOI211_X1 g685(.A(new_n863), .B(new_n861), .C1(new_n885), .C2(new_n886), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n883), .A2(new_n884), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n888), .A2(G148gat), .A3(new_n886), .ZN(new_n889));
  AOI21_X1  g688(.A(KEYINPUT123), .B1(new_n889), .B2(KEYINPUT59), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n862), .B1(new_n887), .B2(new_n890), .ZN(new_n891));
  OR3_X1    g690(.A1(new_n856), .A2(G148gat), .A3(new_n747), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(G1345gat));
  INV_X1    g692(.A(G155gat), .ZN(new_n894));
  NOR3_X1   g693(.A1(new_n849), .A2(new_n894), .A3(new_n704), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n856), .A2(new_n699), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT124), .ZN(new_n897));
  XNOR2_X1  g696(.A(new_n896), .B(new_n897), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n895), .B1(new_n898), .B2(new_n894), .ZN(G1346gat));
  OAI21_X1  g698(.A(G162gat), .B1(new_n849), .B2(new_n710), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n837), .A2(G162gat), .ZN(new_n901));
  NAND4_X1  g700(.A1(new_n853), .A2(new_n854), .A3(new_n855), .A4(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n900), .A2(new_n902), .ZN(G1347gat));
  NOR2_X1   g702(.A1(new_n681), .A2(new_n576), .ZN(new_n904));
  AND3_X1   g703(.A1(new_n820), .A2(new_n631), .A3(new_n904), .ZN(new_n905));
  INV_X1    g704(.A(new_n905), .ZN(new_n906));
  OAI21_X1  g705(.A(G169gat), .B1(new_n906), .B2(new_n296), .ZN(new_n907));
  AND3_X1   g706(.A1(new_n820), .A2(new_n827), .A3(new_n904), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n908), .A2(new_n286), .A3(new_n295), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n907), .A2(new_n909), .ZN(G1348gat));
  AOI21_X1  g709(.A(G176gat), .B1(new_n908), .B2(new_n351), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n706), .A2(new_n344), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n911), .B1(new_n905), .B2(new_n912), .ZN(G1349gat));
  NOR2_X1   g712(.A1(new_n699), .A2(new_n498), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n908), .A2(new_n914), .ZN(new_n915));
  OAI21_X1  g714(.A(G183gat), .B1(new_n906), .B2(new_n704), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  XNOR2_X1  g716(.A(new_n917), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g717(.A1(new_n908), .A2(new_n503), .A3(new_n700), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT61), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n905), .A2(new_n700), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n920), .B1(new_n921), .B2(G190gat), .ZN(new_n922));
  AOI211_X1 g721(.A(KEYINPUT61), .B(new_n503), .C1(new_n905), .C2(new_n700), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n919), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  XNOR2_X1  g723(.A(new_n924), .B(KEYINPUT125), .ZN(G1351gat));
  INV_X1    g724(.A(G197gat), .ZN(new_n926));
  INV_X1    g725(.A(new_n881), .ZN(new_n927));
  AND2_X1   g726(.A1(new_n904), .A2(new_n692), .ZN(new_n928));
  XNOR2_X1  g727(.A(new_n928), .B(KEYINPUT126), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n926), .B1(new_n930), .B2(new_n295), .ZN(new_n931));
  INV_X1    g730(.A(new_n848), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(new_n928), .ZN(new_n933));
  NOR3_X1   g732(.A1(new_n933), .A2(G197gat), .A3(new_n296), .ZN(new_n934));
  OR2_X1    g733(.A1(new_n931), .A2(new_n934), .ZN(G1352gat));
  NOR3_X1   g734(.A1(new_n933), .A2(G204gat), .A3(new_n747), .ZN(new_n936));
  XNOR2_X1  g735(.A(KEYINPUT127), .B(KEYINPUT62), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n936), .B(new_n937), .ZN(new_n938));
  NOR3_X1   g737(.A1(new_n927), .A2(new_n706), .A3(new_n929), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n938), .B1(new_n346), .B2(new_n939), .ZN(G1353gat));
  OR3_X1    g739(.A1(new_n933), .A2(G211gat), .A3(new_n699), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n930), .A2(new_n386), .ZN(new_n942));
  AND3_X1   g741(.A1(new_n942), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n943));
  AOI21_X1  g742(.A(KEYINPUT63), .B1(new_n942), .B2(G211gat), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n941), .B1(new_n943), .B2(new_n944), .ZN(G1354gat));
  INV_X1    g744(.A(G218gat), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n710), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n932), .A2(new_n700), .A3(new_n928), .ZN(new_n948));
  AOI22_X1  g747(.A1(new_n930), .A2(new_n947), .B1(new_n948), .B2(new_n946), .ZN(G1355gat));
endmodule


