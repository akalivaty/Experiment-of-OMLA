//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 0 0 1 0 0 1 0 0 0 1 0 0 0 0 1 1 1 1 1 0 1 0 0 1 1 1 0 1 0 0 0 0 0 1 1 0 1 0 1 1 1 1 1 1 0 1 0 1 1 1 1 0 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:30 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n644, new_n645,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n675,
    new_n676, new_n677, new_n679, new_n680, new_n681, new_n682, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n708, new_n709, new_n710, new_n711, new_n713, new_n714, new_n715,
    new_n717, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n816, new_n817, new_n818, new_n819, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n827, new_n828, new_n829,
    new_n830, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n874,
    new_n875, new_n876, new_n878, new_n879, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n888, new_n889, new_n891, new_n892,
    new_n893, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n924, new_n925;
  XNOR2_X1  g000(.A(G127gat), .B(G155gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G211gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(G15gat), .B(G22gat), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT16), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n204), .B1(new_n205), .B2(G1gat), .ZN(new_n206));
  OAI211_X1 g005(.A(new_n206), .B(KEYINPUT92), .C1(G1gat), .C2(new_n204), .ZN(new_n207));
  INV_X1    g006(.A(G8gat), .ZN(new_n208));
  XNOR2_X1  g007(.A(new_n207), .B(new_n208), .ZN(new_n209));
  NOR2_X1   g008(.A1(G71gat), .A2(G78gat), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT94), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n210), .B(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G57gat), .ZN(new_n213));
  AND2_X1   g012(.A1(new_n213), .A2(G64gat), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n213), .A2(G64gat), .ZN(new_n215));
  OAI21_X1  g014(.A(KEYINPUT9), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(G71gat), .A2(G78gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n212), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT95), .ZN(new_n219));
  XNOR2_X1  g018(.A(new_n218), .B(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n210), .A2(KEYINPUT9), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(new_n217), .ZN(new_n222));
  XNOR2_X1  g021(.A(new_n215), .B(KEYINPUT96), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n222), .B1(new_n223), .B2(new_n214), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n220), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT21), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n209), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(new_n227), .B(G183gat), .ZN(new_n228));
  AOI21_X1  g027(.A(KEYINPUT21), .B1(new_n220), .B2(new_n224), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n228), .B(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(G231gat), .ZN(new_n232));
  INV_X1    g031(.A(G233gat), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n231), .A2(new_n234), .ZN(new_n235));
  NOR3_X1   g034(.A1(new_n230), .A2(new_n232), .A3(new_n233), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n203), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  XNOR2_X1  g036(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n231), .A2(new_n234), .ZN(new_n239));
  INV_X1    g038(.A(new_n203), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n230), .B1(new_n232), .B2(new_n233), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n239), .A2(new_n240), .A3(new_n241), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n237), .A2(new_n238), .A3(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n238), .B1(new_n237), .B2(new_n242), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT14), .ZN(new_n248));
  INV_X1    g047(.A(G29gat), .ZN(new_n249));
  INV_X1    g048(.A(G36gat), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n248), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  OAI21_X1  g050(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n252));
  AOI22_X1  g051(.A1(new_n251), .A2(new_n252), .B1(G29gat), .B2(G36gat), .ZN(new_n253));
  XNOR2_X1  g052(.A(G43gat), .B(G50gat), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(KEYINPUT15), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  AND2_X1   g055(.A1(new_n256), .A2(KEYINPUT90), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n256), .A2(KEYINPUT90), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n251), .B(KEYINPUT91), .ZN(new_n259));
  INV_X1    g058(.A(new_n252), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n255), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  OAI22_X1  g060(.A1(new_n254), .A2(KEYINPUT15), .B1(new_n249), .B2(new_n250), .ZN(new_n262));
  OAI22_X1  g061(.A1(new_n257), .A2(new_n258), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NOR2_X1   g062(.A1(KEYINPUT93), .A2(KEYINPUT17), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(KEYINPUT93), .A2(KEYINPUT17), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n265), .B(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(G85gat), .A2(G92gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n268), .B(KEYINPUT7), .ZN(new_n269));
  INV_X1    g068(.A(G99gat), .ZN(new_n270));
  INV_X1    g069(.A(G106gat), .ZN(new_n271));
  OAI21_X1  g070(.A(KEYINPUT8), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  OAI211_X1 g071(.A(new_n269), .B(new_n272), .C1(G85gat), .C2(G92gat), .ZN(new_n273));
  XNOR2_X1  g072(.A(G99gat), .B(G106gat), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n273), .B(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n267), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g076(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n263), .A2(new_n275), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n277), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  XOR2_X1   g079(.A(G190gat), .B(G218gat), .Z(new_n281));
  XNOR2_X1  g080(.A(new_n280), .B(new_n281), .ZN(new_n282));
  XOR2_X1   g081(.A(G134gat), .B(G162gat), .Z(new_n283));
  AOI21_X1  g082(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n283), .B(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(new_n282), .B(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(G15gat), .B(G43gat), .ZN(new_n288));
  XNOR2_X1  g087(.A(G71gat), .B(G99gat), .ZN(new_n289));
  XOR2_X1   g088(.A(new_n288), .B(new_n289), .Z(new_n290));
  AND2_X1   g089(.A1(G227gat), .A2(G233gat), .ZN(new_n291));
  XNOR2_X1  g090(.A(G127gat), .B(G134gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(KEYINPUT67), .ZN(new_n293));
  INV_X1    g092(.A(G134gat), .ZN(new_n294));
  OR3_X1    g093(.A1(new_n294), .A2(KEYINPUT67), .A3(G127gat), .ZN(new_n295));
  XNOR2_X1  g094(.A(G113gat), .B(G120gat), .ZN(new_n296));
  OAI211_X1 g095(.A(new_n293), .B(new_n295), .C1(KEYINPUT1), .C2(new_n296), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n292), .B1(new_n296), .B2(KEYINPUT68), .ZN(new_n298));
  AOI21_X1  g097(.A(KEYINPUT1), .B1(new_n296), .B2(KEYINPUT68), .ZN(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n297), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT27), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(G183gat), .ZN(new_n304));
  INV_X1    g103(.A(G183gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(KEYINPUT27), .ZN(new_n306));
  INV_X1    g105(.A(G190gat), .ZN(new_n307));
  NAND4_X1  g106(.A1(new_n304), .A2(new_n306), .A3(KEYINPUT28), .A4(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT66), .ZN(new_n309));
  XNOR2_X1  g108(.A(new_n308), .B(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT28), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT64), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n312), .B1(new_n304), .B2(new_n306), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n312), .B1(new_n305), .B2(KEYINPUT27), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(new_n307), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n311), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT65), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  OAI211_X1 g117(.A(KEYINPUT65), .B(new_n311), .C1(new_n313), .C2(new_n315), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n310), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(G169gat), .ZN(new_n321));
  INV_X1    g120(.A(G176gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT26), .ZN(new_n324));
  NAND2_X1  g123(.A1(G169gat), .A2(G176gat), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n323), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(G183gat), .A2(G190gat), .ZN(new_n327));
  OAI211_X1 g126(.A(new_n326), .B(new_n327), .C1(new_n324), .C2(new_n323), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n320), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT23), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n331), .A2(new_n321), .A3(new_n322), .ZN(new_n332));
  OAI21_X1  g131(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n305), .A2(new_n307), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n335), .A2(KEYINPUT24), .A3(new_n327), .ZN(new_n336));
  INV_X1    g135(.A(new_n327), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT24), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND4_X1  g138(.A1(new_n334), .A2(new_n336), .A3(new_n325), .A4(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(KEYINPUT25), .ZN(new_n341));
  AOI22_X1  g140(.A1(new_n332), .A2(new_n333), .B1(new_n337), .B2(new_n338), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT25), .ZN(new_n343));
  NAND4_X1  g142(.A1(new_n342), .A2(new_n343), .A3(new_n325), .A4(new_n336), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n341), .A2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n302), .B1(new_n330), .B2(new_n346), .ZN(new_n347));
  AOI211_X1 g146(.A(new_n301), .B(new_n345), .C1(new_n320), .C2(new_n329), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n291), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT69), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  OAI211_X1 g150(.A(KEYINPUT69), .B(new_n291), .C1(new_n347), .C2(new_n348), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n290), .B1(new_n354), .B2(KEYINPUT33), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  NOR3_X1   g155(.A1(new_n347), .A2(new_n348), .A3(new_n291), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT70), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n359), .A2(KEYINPUT34), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT32), .ZN(new_n361));
  AOI221_X4 g160(.A(new_n361), .B1(new_n357), .B2(new_n358), .C1(new_n351), .C2(new_n352), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n357), .A2(new_n358), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n363), .B1(new_n353), .B2(KEYINPUT32), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n360), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n345), .B1(new_n320), .B2(new_n329), .ZN(new_n366));
  XNOR2_X1  g165(.A(new_n366), .B(new_n302), .ZN(new_n367));
  AOI21_X1  g166(.A(KEYINPUT69), .B1(new_n367), .B2(new_n291), .ZN(new_n368));
  INV_X1    g167(.A(new_n352), .ZN(new_n369));
  OAI21_X1  g168(.A(KEYINPUT32), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(new_n363), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n360), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n353), .A2(KEYINPUT32), .A3(new_n363), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n372), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n356), .B1(new_n365), .B2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n365), .A2(new_n375), .A3(new_n356), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n377), .A2(KEYINPUT87), .A3(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT3), .ZN(new_n380));
  XNOR2_X1  g179(.A(G197gat), .B(G204gat), .ZN(new_n381));
  INV_X1    g180(.A(G211gat), .ZN(new_n382));
  INV_X1    g181(.A(G218gat), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n381), .B1(KEYINPUT22), .B2(new_n384), .ZN(new_n385));
  XNOR2_X1  g184(.A(G211gat), .B(G218gat), .ZN(new_n386));
  XNOR2_X1  g185(.A(new_n385), .B(new_n386), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n380), .B1(new_n387), .B2(KEYINPUT29), .ZN(new_n388));
  INV_X1    g187(.A(G141gat), .ZN(new_n389));
  OAI21_X1  g188(.A(KEYINPUT75), .B1(new_n389), .B2(G148gat), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT75), .ZN(new_n391));
  INV_X1    g190(.A(G148gat), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n391), .A2(new_n392), .A3(G141gat), .ZN(new_n393));
  OAI211_X1 g192(.A(new_n390), .B(new_n393), .C1(G141gat), .C2(new_n392), .ZN(new_n394));
  XNOR2_X1  g193(.A(G155gat), .B(G162gat), .ZN(new_n395));
  INV_X1    g194(.A(G155gat), .ZN(new_n396));
  INV_X1    g195(.A(G162gat), .ZN(new_n397));
  OAI21_X1  g196(.A(KEYINPUT2), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n394), .A2(new_n395), .A3(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n395), .ZN(new_n400));
  XNOR2_X1  g199(.A(G141gat), .B(G148gat), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n400), .B1(KEYINPUT2), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n399), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n388), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(G228gat), .A2(G233gat), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n403), .A2(KEYINPUT3), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n387), .B1(new_n406), .B2(KEYINPUT29), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n404), .A2(new_n405), .A3(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT76), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n403), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n399), .A2(KEYINPUT76), .A3(new_n402), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n388), .A2(new_n412), .ZN(new_n413));
  AND2_X1   g212(.A1(new_n413), .A2(new_n407), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n408), .B1(new_n414), .B2(new_n405), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(G22gat), .ZN(new_n416));
  INV_X1    g215(.A(G22gat), .ZN(new_n417));
  OAI211_X1 g216(.A(new_n408), .B(new_n417), .C1(new_n414), .C2(new_n405), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n416), .A2(KEYINPUT83), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(KEYINPUT84), .ZN(new_n420));
  XOR2_X1   g219(.A(KEYINPUT81), .B(KEYINPUT31), .Z(new_n421));
  XNOR2_X1  g220(.A(G78gat), .B(G106gat), .ZN(new_n422));
  XNOR2_X1  g221(.A(new_n421), .B(new_n422), .ZN(new_n423));
  XOR2_X1   g222(.A(KEYINPUT82), .B(G50gat), .Z(new_n424));
  XNOR2_X1  g223(.A(new_n423), .B(new_n424), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n420), .A2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT84), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n416), .A2(new_n427), .A3(new_n418), .ZN(new_n428));
  AND2_X1   g227(.A1(new_n420), .A2(new_n428), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n426), .B1(new_n429), .B2(new_n425), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT87), .ZN(new_n431));
  AND3_X1   g230(.A1(new_n365), .A2(new_n375), .A3(new_n356), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n431), .B1(new_n432), .B2(new_n376), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n379), .A2(new_n430), .A3(new_n433), .ZN(new_n434));
  XNOR2_X1  g233(.A(G8gat), .B(G36gat), .ZN(new_n435));
  XNOR2_X1  g234(.A(G64gat), .B(G92gat), .ZN(new_n436));
  XNOR2_X1  g235(.A(new_n435), .B(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(G226gat), .A2(G233gat), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n439), .B1(new_n366), .B2(KEYINPUT29), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT72), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  OAI211_X1 g241(.A(KEYINPUT72), .B(new_n439), .C1(new_n366), .C2(KEYINPUT29), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n387), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n330), .A2(new_n346), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(KEYINPUT71), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT71), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n366), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n439), .ZN(new_n450));
  AOI21_X1  g249(.A(KEYINPUT73), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n447), .B1(new_n330), .B2(new_n346), .ZN(new_n452));
  AOI211_X1 g251(.A(KEYINPUT71), .B(new_n345), .C1(new_n320), .C2(new_n329), .ZN(new_n453));
  OAI211_X1 g252(.A(KEYINPUT73), .B(new_n450), .C1(new_n452), .C2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(new_n454), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n444), .B1(new_n451), .B2(new_n455), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n450), .A2(KEYINPUT29), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n457), .B1(new_n452), .B2(new_n453), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n366), .A2(new_n450), .ZN(new_n459));
  AND3_X1   g258(.A1(new_n458), .A2(new_n387), .A3(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n438), .B1(new_n456), .B2(new_n461), .ZN(new_n462));
  AND3_X1   g261(.A1(new_n456), .A2(new_n461), .A3(new_n438), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n462), .B1(new_n463), .B2(KEYINPUT30), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n456), .A2(new_n461), .A3(new_n438), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT30), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT74), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n406), .B1(new_n412), .B2(KEYINPUT3), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n302), .A2(KEYINPUT77), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT77), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n301), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n470), .A2(new_n474), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n299), .B(new_n292), .C1(KEYINPUT68), .C2(new_n296), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n476), .A2(new_n402), .A3(new_n399), .A4(new_n297), .ZN(new_n477));
  XNOR2_X1  g276(.A(new_n477), .B(KEYINPUT4), .ZN(new_n478));
  NAND2_X1  g277(.A1(G225gat), .A2(G233gat), .ZN(new_n479));
  XOR2_X1   g278(.A(new_n479), .B(KEYINPUT78), .Z(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n475), .A2(new_n478), .A3(new_n481), .ZN(new_n482));
  AOI22_X1  g281(.A1(new_n471), .A2(new_n473), .B1(new_n410), .B2(new_n411), .ZN(new_n483));
  INV_X1    g282(.A(new_n477), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n480), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n482), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(KEYINPUT5), .ZN(new_n487));
  XNOR2_X1  g286(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n488));
  XNOR2_X1  g287(.A(G57gat), .B(G85gat), .ZN(new_n489));
  XNOR2_X1  g288(.A(new_n488), .B(new_n489), .ZN(new_n490));
  XNOR2_X1  g289(.A(G1gat), .B(G29gat), .ZN(new_n491));
  XOR2_X1   g290(.A(new_n490), .B(new_n491), .Z(new_n492));
  INV_X1    g291(.A(KEYINPUT5), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n482), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n487), .A2(new_n492), .A3(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(new_n492), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n493), .B1(new_n482), .B2(new_n485), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT4), .ZN(new_n498));
  XNOR2_X1  g297(.A(new_n477), .B(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n499), .B1(new_n474), .B2(new_n470), .ZN(new_n500));
  AOI21_X1  g299(.A(KEYINPUT5), .B1(new_n500), .B2(new_n481), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n496), .B1(new_n497), .B2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT6), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n495), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n487), .A2(KEYINPUT6), .A3(new_n492), .A4(new_n494), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n465), .A2(KEYINPUT74), .A3(new_n466), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n464), .A2(new_n469), .A3(new_n506), .A4(new_n507), .ZN(new_n508));
  OR2_X1    g307(.A1(new_n508), .A2(KEYINPUT35), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n434), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n508), .A2(KEYINPUT80), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n450), .B1(new_n452), .B2(new_n453), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT73), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(new_n454), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n460), .B1(new_n516), .B2(new_n444), .ZN(new_n517));
  AOI211_X1 g316(.A(new_n468), .B(KEYINPUT30), .C1(new_n517), .C2(new_n438), .ZN(new_n518));
  AOI21_X1  g317(.A(KEYINPUT74), .B1(new_n465), .B2(new_n466), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT80), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n520), .A2(new_n521), .A3(new_n506), .A4(new_n464), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n512), .A2(new_n522), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n430), .B1(new_n432), .B2(new_n376), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT88), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  OAI211_X1 g325(.A(KEYINPUT88), .B(new_n430), .C1(new_n432), .C2(new_n376), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n523), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT89), .ZN(new_n529));
  AND3_X1   g328(.A1(new_n528), .A2(new_n529), .A3(KEYINPUT35), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n529), .B1(new_n528), .B2(KEYINPUT35), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n511), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(new_n506), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n442), .A2(new_n443), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n516), .A2(new_n534), .A3(new_n387), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n458), .A2(new_n459), .ZN(new_n536));
  OAI211_X1 g335(.A(new_n535), .B(KEYINPUT37), .C1(new_n387), .C2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT38), .ZN(new_n538));
  XOR2_X1   g337(.A(KEYINPUT85), .B(KEYINPUT37), .Z(new_n539));
  NAND2_X1  g338(.A1(new_n517), .A2(new_n539), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n537), .A2(new_n538), .A3(new_n540), .A4(new_n437), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n437), .ZN(new_n542));
  INV_X1    g341(.A(new_n517), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n542), .B1(new_n543), .B2(KEYINPUT37), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n463), .A2(KEYINPUT38), .ZN(new_n545));
  OAI211_X1 g344(.A(new_n533), .B(new_n541), .C1(new_n544), .C2(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n464), .A2(new_n469), .A3(new_n507), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n500), .A2(new_n481), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT39), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n492), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NOR3_X1   g349(.A1(new_n483), .A2(new_n480), .A3(new_n484), .ZN(new_n551));
  OR2_X1    g350(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n550), .B1(new_n552), .B2(new_n549), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n553), .B(KEYINPUT40), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n547), .A2(new_n495), .A3(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n546), .A2(new_n430), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(KEYINPUT86), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT86), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n546), .A2(new_n555), .A3(new_n558), .A4(new_n430), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n523), .A2(new_n430), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n377), .A2(KEYINPUT36), .A3(new_n378), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT36), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n564), .B1(new_n432), .B2(new_n376), .ZN(new_n565));
  NAND4_X1  g364(.A1(new_n560), .A2(new_n562), .A3(new_n563), .A4(new_n565), .ZN(new_n566));
  AOI211_X1 g365(.A(new_n247), .B(new_n287), .C1(new_n532), .C2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n267), .A2(new_n209), .ZN(new_n568));
  INV_X1    g367(.A(new_n209), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n569), .A2(new_n263), .ZN(new_n570));
  AND2_X1   g369(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(G229gat), .A2(G233gat), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n571), .A2(KEYINPUT18), .A3(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n263), .B(new_n209), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n572), .B(KEYINPUT13), .ZN(new_n575));
  OR2_X1    g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n568), .A2(new_n570), .A3(new_n572), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT18), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n573), .A2(new_n576), .A3(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(G113gat), .B(G141gat), .ZN(new_n581));
  INV_X1    g380(.A(G197gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n581), .B(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(KEYINPUT11), .B(G169gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n583), .B(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(KEYINPUT12), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  OR2_X1    g386(.A1(new_n580), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n580), .A2(new_n587), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n225), .B(new_n275), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT10), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n225), .A2(new_n276), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n595), .A2(KEYINPUT10), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n596), .A2(KEYINPUT97), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT97), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n595), .A2(new_n598), .A3(KEYINPUT10), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n594), .A2(new_n597), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(G230gat), .A2(G233gat), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT102), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n592), .A2(new_n601), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(KEYINPUT98), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n600), .A2(KEYINPUT102), .A3(new_n601), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n604), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(G120gat), .B(G148gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(KEYINPUT101), .ZN(new_n610));
  XOR2_X1   g409(.A(KEYINPUT99), .B(KEYINPUT100), .Z(new_n611));
  XNOR2_X1  g410(.A(new_n610), .B(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(G176gat), .B(G204gat), .ZN(new_n613));
  XOR2_X1   g412(.A(new_n612), .B(new_n613), .Z(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n608), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n606), .A2(new_n602), .A3(new_n614), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n591), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n567), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n620), .A2(new_n506), .ZN(new_n621));
  XOR2_X1   g420(.A(KEYINPUT103), .B(G1gat), .Z(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(G1324gat));
  INV_X1    g422(.A(new_n547), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n620), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n205), .A2(new_n208), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n625), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT42), .ZN(new_n629));
  OR2_X1    g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n628), .A2(new_n629), .ZN(new_n631));
  OAI211_X1 g430(.A(new_n630), .B(new_n631), .C1(new_n208), .C2(new_n625), .ZN(G1325gat));
  INV_X1    g431(.A(G15gat), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n563), .A2(new_n565), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n634), .A2(KEYINPUT104), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT104), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n563), .A2(new_n636), .A3(new_n565), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  NOR3_X1   g437(.A1(new_n620), .A2(new_n633), .A3(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n379), .A2(new_n433), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n567), .A2(new_n619), .A3(new_n641), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n639), .B1(new_n633), .B2(new_n642), .ZN(G1326gat));
  NOR2_X1   g442(.A1(new_n620), .A2(new_n430), .ZN(new_n644));
  XOR2_X1   g443(.A(KEYINPUT43), .B(G22gat), .Z(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(G1327gat));
  AOI21_X1  g445(.A(new_n286), .B1(new_n532), .B2(new_n566), .ZN(new_n647));
  AND3_X1   g446(.A1(new_n647), .A2(new_n619), .A3(new_n247), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n648), .A2(new_n249), .A3(new_n533), .ZN(new_n649));
  OR2_X1    g448(.A1(new_n649), .A2(KEYINPUT105), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(KEYINPUT105), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT45), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT44), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n528), .A2(KEYINPUT35), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n656), .A2(KEYINPUT89), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n528), .A2(new_n529), .A3(KEYINPUT35), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n510), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  AND3_X1   g458(.A1(new_n560), .A2(new_n562), .A3(new_n638), .ZN(new_n660));
  OAI211_X1 g459(.A(new_n655), .B(new_n287), .C1(new_n659), .C2(new_n660), .ZN(new_n661));
  OAI211_X1 g460(.A(new_n661), .B(KEYINPUT108), .C1(new_n655), .C2(new_n647), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n618), .B(KEYINPUT107), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n663), .A2(new_n591), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n560), .A2(new_n562), .A3(new_n638), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n532), .A2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT108), .ZN(new_n667));
  NAND4_X1  g466(.A1(new_n666), .A2(new_n667), .A3(new_n655), .A4(new_n287), .ZN(new_n668));
  XOR2_X1   g467(.A(new_n246), .B(KEYINPUT106), .Z(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NAND4_X1  g469(.A1(new_n662), .A2(new_n664), .A3(new_n668), .A4(new_n670), .ZN(new_n671));
  OAI21_X1  g470(.A(G29gat), .B1(new_n671), .B2(new_n506), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n650), .A2(KEYINPUT45), .A3(new_n651), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n654), .A2(new_n672), .A3(new_n673), .ZN(G1328gat));
  NAND3_X1  g473(.A1(new_n648), .A2(new_n250), .A3(new_n547), .ZN(new_n675));
  XOR2_X1   g474(.A(new_n675), .B(KEYINPUT46), .Z(new_n676));
  OAI21_X1  g475(.A(G36gat), .B1(new_n671), .B2(new_n624), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(G1329gat));
  INV_X1    g477(.A(new_n638), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n679), .A2(G43gat), .ZN(new_n680));
  AND2_X1   g479(.A1(new_n648), .A2(new_n641), .ZN(new_n681));
  OAI22_X1  g480(.A1(new_n671), .A2(new_n680), .B1(new_n681), .B2(G43gat), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g482(.A(G50gat), .B1(new_n671), .B2(new_n430), .ZN(new_n684));
  INV_X1    g483(.A(G50gat), .ZN(new_n685));
  INV_X1    g484(.A(new_n430), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n648), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT109), .ZN(new_n689));
  AOI21_X1  g488(.A(KEYINPUT48), .B1(new_n687), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  OAI211_X1 g490(.A(new_n684), .B(new_n687), .C1(new_n689), .C2(KEYINPUT48), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(G1331gat));
  INV_X1    g492(.A(KEYINPUT111), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n237), .A2(new_n242), .ZN(new_n695));
  INV_X1    g494(.A(new_n238), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND4_X1  g496(.A1(new_n697), .A2(new_n591), .A3(new_n243), .A4(new_n286), .ZN(new_n698));
  INV_X1    g497(.A(new_n663), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(KEYINPUT110), .ZN(new_n701));
  AND3_X1   g500(.A1(new_n666), .A2(new_n694), .A3(new_n701), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n694), .B1(new_n666), .B2(new_n701), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(new_n533), .ZN(new_n705));
  XNOR2_X1  g504(.A(KEYINPUT112), .B(G57gat), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n705), .B(new_n706), .ZN(G1332gat));
  NOR3_X1   g506(.A1(new_n702), .A2(new_n703), .A3(new_n624), .ZN(new_n708));
  NOR2_X1   g507(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n709));
  AND2_X1   g508(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n708), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n711), .B1(new_n708), .B2(new_n709), .ZN(G1333gat));
  NAND3_X1  g511(.A1(new_n704), .A2(G71gat), .A3(new_n679), .ZN(new_n713));
  NOR3_X1   g512(.A1(new_n702), .A2(new_n703), .A3(new_n640), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n713), .B1(G71gat), .B2(new_n714), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g515(.A1(new_n704), .A2(new_n686), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(G78gat), .ZN(G1335gat));
  INV_X1    g517(.A(new_n668), .ZN(new_n719));
  INV_X1    g518(.A(new_n566), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n287), .B1(new_n720), .B2(new_n659), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n667), .B1(new_n721), .B2(KEYINPUT44), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n719), .B1(new_n722), .B2(new_n661), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n246), .A2(new_n590), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(new_n618), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n723), .A2(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(G85gat), .B1(new_n727), .B2(new_n506), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n666), .A2(new_n287), .A3(new_n724), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT51), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND4_X1  g530(.A1(new_n666), .A2(KEYINPUT51), .A3(new_n287), .A4(new_n724), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  OR2_X1    g532(.A1(new_n733), .A2(KEYINPUT113), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(KEYINPUT113), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n734), .A2(new_n618), .A3(new_n735), .ZN(new_n736));
  OR2_X1    g535(.A1(new_n506), .A2(G85gat), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n728), .B1(new_n736), .B2(new_n737), .ZN(G1336gat));
  INV_X1    g537(.A(KEYINPUT115), .ZN(new_n739));
  NAND4_X1  g538(.A1(new_n662), .A2(new_n547), .A3(new_n668), .A4(new_n726), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n739), .B1(new_n740), .B2(G92gat), .ZN(new_n741));
  NOR3_X1   g540(.A1(new_n699), .A2(G92gat), .A3(new_n624), .ZN(new_n742));
  XOR2_X1   g541(.A(new_n742), .B(KEYINPUT114), .Z(new_n743));
  AOI21_X1  g542(.A(new_n743), .B1(new_n731), .B2(new_n732), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n744), .B1(new_n740), .B2(G92gat), .ZN(new_n745));
  NOR3_X1   g544(.A1(new_n741), .A2(new_n745), .A3(KEYINPUT52), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT52), .ZN(new_n747));
  AOI221_X4 g546(.A(new_n744), .B1(new_n739), .B2(new_n747), .C1(G92gat), .C2(new_n740), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n746), .A2(new_n748), .ZN(G1337gat));
  OAI21_X1  g548(.A(G99gat), .B1(new_n727), .B2(new_n638), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n641), .A2(new_n270), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n750), .B1(new_n736), .B2(new_n751), .ZN(G1338gat));
  NAND4_X1  g551(.A1(new_n723), .A2(KEYINPUT117), .A3(new_n686), .A4(new_n726), .ZN(new_n753));
  NAND4_X1  g552(.A1(new_n662), .A2(new_n686), .A3(new_n668), .A4(new_n726), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT117), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n753), .A2(G106gat), .A3(new_n756), .ZN(new_n757));
  NOR3_X1   g556(.A1(new_n699), .A2(G106gat), .A3(new_n430), .ZN(new_n758));
  AOI21_X1  g557(.A(KEYINPUT53), .B1(new_n733), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  AND2_X1   g559(.A1(new_n754), .A2(G106gat), .ZN(new_n761));
  XOR2_X1   g560(.A(new_n758), .B(KEYINPUT116), .Z(new_n762));
  AOI21_X1  g561(.A(new_n762), .B1(new_n731), .B2(new_n732), .ZN(new_n763));
  OAI21_X1  g562(.A(KEYINPUT53), .B1(new_n761), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n760), .A2(new_n764), .ZN(G1339gat));
  NOR3_X1   g564(.A1(new_n244), .A2(new_n245), .A3(new_n287), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT118), .ZN(new_n767));
  INV_X1    g566(.A(new_n618), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n766), .A2(new_n767), .A3(new_n768), .A4(new_n591), .ZN(new_n769));
  OAI21_X1  g568(.A(KEYINPUT118), .B1(new_n698), .B2(new_n618), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  OR3_X1    g570(.A1(new_n571), .A2(KEYINPUT121), .A3(new_n572), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n574), .A2(new_n575), .ZN(new_n773));
  OAI21_X1  g572(.A(KEYINPUT121), .B1(new_n571), .B2(new_n572), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n772), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(new_n585), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(new_n588), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(KEYINPUT122), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT122), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n776), .A2(new_n588), .A3(new_n779), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n286), .B1(new_n778), .B2(new_n780), .ZN(new_n781));
  AOI21_X1  g580(.A(KEYINPUT54), .B1(new_n604), .B2(new_n607), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n782), .A2(new_n614), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT55), .ZN(new_n784));
  INV_X1    g583(.A(new_n601), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n594), .A2(new_n785), .A3(new_n597), .A4(new_n599), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n602), .A2(KEYINPUT54), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(KEYINPUT119), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT119), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n602), .A2(new_n789), .A3(KEYINPUT54), .A4(new_n786), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  AND3_X1   g590(.A1(new_n783), .A2(new_n784), .A3(new_n791), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n784), .B1(new_n783), .B2(new_n791), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n617), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT120), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  OAI211_X1 g595(.A(KEYINPUT120), .B(new_n617), .C1(new_n792), .C2(new_n793), .ZN(new_n797));
  AND3_X1   g596(.A1(new_n781), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n796), .A2(new_n590), .A3(new_n797), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n776), .A2(new_n588), .A3(new_n618), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n798), .B1(new_n801), .B2(new_n286), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n771), .B1(new_n802), .B2(new_n669), .ZN(new_n803));
  AND2_X1   g602(.A1(new_n526), .A2(new_n527), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NOR3_X1   g604(.A1(new_n805), .A2(new_n506), .A3(new_n547), .ZN(new_n806));
  INV_X1    g605(.A(G113gat), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n806), .A2(new_n807), .A3(new_n590), .ZN(new_n808));
  INV_X1    g607(.A(new_n434), .ZN(new_n809));
  AND2_X1   g608(.A1(new_n803), .A2(new_n809), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n547), .A2(new_n506), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n810), .A2(new_n590), .A3(new_n811), .ZN(new_n812));
  AND3_X1   g611(.A1(new_n812), .A2(KEYINPUT123), .A3(G113gat), .ZN(new_n813));
  AOI21_X1  g612(.A(KEYINPUT123), .B1(new_n812), .B2(G113gat), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n808), .B1(new_n813), .B2(new_n814), .ZN(G1340gat));
  NAND2_X1  g614(.A1(new_n810), .A2(new_n811), .ZN(new_n816));
  OAI21_X1  g615(.A(G120gat), .B1(new_n816), .B2(new_n699), .ZN(new_n817));
  INV_X1    g616(.A(G120gat), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n806), .A2(new_n818), .A3(new_n618), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n817), .A2(new_n819), .ZN(G1341gat));
  OAI21_X1  g619(.A(G127gat), .B1(new_n816), .B2(new_n670), .ZN(new_n821));
  INV_X1    g620(.A(G127gat), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n806), .A2(new_n822), .A3(new_n246), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT124), .ZN(new_n825));
  XNOR2_X1  g624(.A(new_n824), .B(new_n825), .ZN(G1342gat));
  NAND3_X1  g625(.A1(new_n806), .A2(new_n294), .A3(new_n287), .ZN(new_n827));
  OR2_X1    g626(.A1(new_n827), .A2(KEYINPUT56), .ZN(new_n828));
  OAI21_X1  g627(.A(G134gat), .B1(new_n816), .B2(new_n286), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n827), .A2(KEYINPUT56), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n828), .A2(new_n829), .A3(new_n830), .ZN(G1343gat));
  NAND2_X1  g630(.A1(new_n638), .A2(new_n811), .ZN(new_n832));
  INV_X1    g631(.A(new_n832), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n800), .B1(new_n794), .B2(new_n591), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(new_n286), .ZN(new_n835));
  INV_X1    g634(.A(new_n835), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n247), .B1(new_n836), .B2(new_n798), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(new_n771), .ZN(new_n838));
  NAND4_X1  g637(.A1(new_n838), .A2(KEYINPUT125), .A3(KEYINPUT57), .A4(new_n686), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n781), .A2(new_n796), .A3(new_n797), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n246), .B1(new_n835), .B2(new_n840), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n769), .A2(new_n770), .ZN(new_n842));
  OAI211_X1 g641(.A(KEYINPUT57), .B(new_n686), .C1(new_n841), .C2(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT125), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n839), .A2(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(KEYINPUT57), .B1(new_n803), .B2(new_n686), .ZN(new_n847));
  OAI211_X1 g646(.A(new_n590), .B(new_n833), .C1(new_n846), .C2(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(G141gat), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n803), .A2(new_n686), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n850), .A2(new_n832), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n851), .A2(new_n389), .A3(new_n590), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n849), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(KEYINPUT58), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT58), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n849), .A2(new_n852), .A3(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n854), .A2(new_n856), .ZN(G1344gat));
  INV_X1    g656(.A(KEYINPUT59), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n833), .B1(new_n846), .B2(new_n847), .ZN(new_n859));
  OAI211_X1 g658(.A(new_n858), .B(G148gat), .C1(new_n859), .C2(new_n768), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n850), .A2(KEYINPUT57), .ZN(new_n861));
  AOI211_X1 g660(.A(new_n286), .B(new_n794), .C1(new_n778), .C2(new_n780), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n247), .B1(new_n836), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n863), .B1(new_n618), .B2(new_n698), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT57), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n864), .A2(new_n865), .A3(new_n686), .ZN(new_n866));
  AND2_X1   g665(.A1(new_n861), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n832), .A2(new_n768), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n392), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n860), .B1(new_n869), .B2(new_n858), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n851), .A2(new_n392), .A3(new_n618), .ZN(new_n871));
  XNOR2_X1  g670(.A(new_n871), .B(KEYINPUT126), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n870), .A2(new_n872), .ZN(G1345gat));
  AOI21_X1  g672(.A(G155gat), .B1(new_n851), .B2(new_n246), .ZN(new_n874));
  INV_X1    g673(.A(new_n859), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n670), .A2(new_n396), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n874), .B1(new_n875), .B2(new_n876), .ZN(G1346gat));
  AOI21_X1  g676(.A(G162gat), .B1(new_n851), .B2(new_n287), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n286), .A2(new_n397), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n878), .B1(new_n875), .B2(new_n879), .ZN(G1347gat));
  NOR2_X1   g679(.A1(new_n624), .A2(new_n533), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n810), .A2(new_n881), .ZN(new_n882));
  OAI21_X1  g681(.A(G169gat), .B1(new_n882), .B2(new_n591), .ZN(new_n883));
  INV_X1    g682(.A(new_n881), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n805), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n885), .A2(new_n321), .A3(new_n590), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n883), .A2(new_n886), .ZN(G1348gat));
  NOR3_X1   g686(.A1(new_n882), .A2(new_n322), .A3(new_n699), .ZN(new_n888));
  AOI21_X1  g687(.A(G176gat), .B1(new_n885), .B2(new_n618), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n888), .A2(new_n889), .ZN(G1349gat));
  OAI21_X1  g689(.A(G183gat), .B1(new_n882), .B2(new_n670), .ZN(new_n891));
  NAND4_X1  g690(.A1(new_n885), .A2(new_n304), .A3(new_n306), .A4(new_n246), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  XNOR2_X1  g692(.A(new_n893), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g693(.A1(new_n810), .A2(new_n287), .A3(new_n881), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n895), .A2(G190gat), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(KEYINPUT127), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT127), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n895), .A2(new_n898), .A3(G190gat), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n897), .A2(KEYINPUT61), .A3(new_n899), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n885), .A2(new_n307), .A3(new_n287), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT61), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n896), .A2(KEYINPUT127), .A3(new_n902), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n900), .A2(new_n901), .A3(new_n903), .ZN(G1351gat));
  NOR2_X1   g703(.A1(new_n679), .A2(new_n884), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n867), .A2(new_n905), .ZN(new_n906));
  OAI21_X1  g705(.A(G197gat), .B1(new_n906), .B2(new_n591), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n803), .A2(new_n686), .A3(new_n905), .ZN(new_n908));
  INV_X1    g707(.A(new_n908), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n909), .A2(new_n582), .A3(new_n590), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n907), .A2(new_n910), .ZN(G1352gat));
  OAI21_X1  g710(.A(G204gat), .B1(new_n906), .B2(new_n699), .ZN(new_n912));
  NOR3_X1   g711(.A1(new_n908), .A2(G204gat), .A3(new_n768), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT62), .ZN(new_n914));
  OR2_X1    g713(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n913), .A2(new_n914), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n912), .A2(new_n915), .A3(new_n916), .ZN(G1353gat));
  NAND3_X1  g716(.A1(new_n909), .A2(new_n382), .A3(new_n246), .ZN(new_n918));
  NAND4_X1  g717(.A1(new_n861), .A2(new_n246), .A3(new_n866), .A4(new_n905), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n919), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n920));
  INV_X1    g719(.A(new_n920), .ZN(new_n921));
  AOI21_X1  g720(.A(KEYINPUT63), .B1(new_n919), .B2(G211gat), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n918), .B1(new_n921), .B2(new_n922), .ZN(G1354gat));
  OAI21_X1  g722(.A(G218gat), .B1(new_n906), .B2(new_n286), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n909), .A2(new_n383), .A3(new_n287), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(G1355gat));
endmodule


