

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762;

  OR2_X1 U373 ( .A1(n612), .A2(n406), .ZN(n643) );
  XNOR2_X1 U374 ( .A(n411), .B(n451), .ZN(n762) );
  NAND2_X1 U375 ( .A1(n591), .A2(n590), .ZN(n422) );
  AND2_X1 U376 ( .A1(n390), .A2(n389), .ZN(n388) );
  AND2_X2 U377 ( .A1(n417), .A2(n413), .ZN(n404) );
  NAND2_X2 U378 ( .A1(n350), .A2(n355), .ZN(n402) );
  NAND2_X1 U379 ( .A1(n605), .A2(n426), .ZN(n350) );
  NAND2_X1 U380 ( .A1(n599), .A2(n598), .ZN(n421) );
  NOR2_X1 U381 ( .A1(n661), .A2(n659), .ZN(n699) );
  XNOR2_X2 U382 ( .A(n421), .B(n600), .ZN(n608) );
  INV_X2 U383 ( .A(n601), .ZN(n351) );
  NAND2_X1 U384 ( .A1(n436), .A2(n439), .ZN(n704) );
  XNOR2_X1 U385 ( .A(n562), .B(KEYINPUT6), .ZN(n609) );
  XNOR2_X1 U386 ( .A(n561), .B(n492), .ZN(n603) );
  XNOR2_X1 U387 ( .A(n511), .B(n510), .ZN(n568) );
  XOR2_X1 U388 ( .A(n531), .B(KEYINPUT59), .Z(n627) );
  XNOR2_X1 U389 ( .A(n396), .B(n541), .ZN(n740) );
  INV_X2 U390 ( .A(G953), .ZN(n754) );
  BUF_X1 U391 ( .A(n761), .Z(n352) );
  XNOR2_X1 U392 ( .A(n444), .B(n443), .ZN(n761) );
  XNOR2_X1 U393 ( .A(n401), .B(n585), .ZN(n384) );
  XNOR2_X2 U394 ( .A(n573), .B(n572), .ZN(n591) );
  XNOR2_X1 U395 ( .A(n403), .B(n471), .ZN(n409) );
  XNOR2_X2 U396 ( .A(n424), .B(G110), .ZN(n508) );
  XNOR2_X2 U397 ( .A(G104), .B(KEYINPUT75), .ZN(n424) );
  NOR2_X1 U398 ( .A1(n717), .A2(n622), .ZN(n480) );
  NAND2_X1 U399 ( .A1(n380), .A2(n378), .ZN(n579) );
  NAND2_X1 U400 ( .A1(n379), .A2(KEYINPUT47), .ZN(n378) );
  AND2_X1 U401 ( .A1(n429), .A2(n428), .ZN(n570) );
  XNOR2_X1 U402 ( .A(n665), .B(n430), .ZN(n429) );
  XNOR2_X1 U403 ( .A(G902), .B(KEYINPUT15), .ZN(n623) );
  NAND2_X1 U404 ( .A1(n704), .A2(n594), .ZN(n368) );
  NOR2_X1 U405 ( .A1(n704), .A2(n594), .ZN(n367) );
  NAND2_X1 U406 ( .A1(n682), .A2(n683), .ZN(n617) );
  XNOR2_X1 U407 ( .A(n561), .B(G472), .ZN(n562) );
  INV_X1 U408 ( .A(n608), .ZN(n398) );
  XNOR2_X1 U409 ( .A(G125), .B(G146), .ZN(n475) );
  XNOR2_X1 U410 ( .A(n534), .B(n486), .ZN(n748) );
  XNOR2_X1 U411 ( .A(n475), .B(KEYINPUT10), .ZN(n514) );
  INV_X1 U412 ( .A(n758), .ZN(n432) );
  NAND2_X1 U413 ( .A1(n404), .A2(n412), .ZN(n401) );
  XNOR2_X1 U414 ( .A(n506), .B(n505), .ZN(n507) );
  INV_X1 U415 ( .A(G107), .ZN(n505) );
  XOR2_X1 U416 ( .A(G137), .B(G140), .Z(n515) );
  XOR2_X1 U417 ( .A(KEYINPUT4), .B(G101), .Z(n504) );
  XOR2_X1 U418 ( .A(KEYINPUT77), .B(KEYINPUT18), .Z(n473) );
  XOR2_X1 U419 ( .A(G143), .B(G128), .Z(n482) );
  XNOR2_X1 U420 ( .A(n435), .B(n434), .ZN(n605) );
  INV_X1 U421 ( .A(KEYINPUT66), .ZN(n434) );
  AND2_X1 U422 ( .A1(n683), .A2(n593), .ZN(n441) );
  OR2_X1 U423 ( .A1(n609), .A2(n593), .ZN(n438) );
  INV_X1 U424 ( .A(n623), .ZN(n622) );
  AND2_X1 U425 ( .A1(n603), .A2(n563), .ZN(n551) );
  XNOR2_X1 U426 ( .A(n748), .B(G146), .ZN(n503) );
  XNOR2_X1 U427 ( .A(n409), .B(n504), .ZN(n377) );
  NOR2_X1 U428 ( .A1(G953), .A2(G237), .ZN(n489) );
  XNOR2_X1 U429 ( .A(G116), .B(G137), .ZN(n487) );
  XOR2_X1 U430 ( .A(KEYINPUT5), .B(KEYINPUT96), .Z(n488) );
  INV_X1 U431 ( .A(KEYINPUT3), .ZN(n468) );
  INV_X1 U432 ( .A(G119), .ZN(n467) );
  XNOR2_X1 U433 ( .A(n508), .B(KEYINPUT16), .ZN(n396) );
  XNOR2_X1 U434 ( .A(n423), .B(G116), .ZN(n541) );
  XNOR2_X1 U435 ( .A(G107), .B(G122), .ZN(n423) );
  XNOR2_X1 U436 ( .A(G143), .B(G113), .ZN(n457) );
  NAND2_X1 U437 ( .A1(n388), .A2(n385), .ZN(n692) );
  NAND2_X1 U438 ( .A1(n356), .A2(n365), .ZN(n373) );
  NAND2_X1 U439 ( .A1(n367), .A2(n366), .ZN(n365) );
  NOR2_X1 U440 ( .A1(n602), .A2(n354), .ZN(n452) );
  INV_X1 U441 ( .A(KEYINPUT78), .ZN(n374) );
  XOR2_X1 U442 ( .A(KEYINPUT22), .B(KEYINPUT73), .Z(n600) );
  NOR2_X1 U443 ( .A1(n609), .A2(n608), .ZN(n611) );
  INV_X1 U444 ( .A(KEYINPUT1), .ZN(n567) );
  AND2_X2 U445 ( .A1(n405), .A2(n625), .ZN(n729) );
  XNOR2_X1 U446 ( .A(n448), .B(KEYINPUT64), .ZN(n405) );
  NAND2_X1 U447 ( .A1(n449), .A2(n624), .ZN(n448) );
  INV_X1 U448 ( .A(KEYINPUT85), .ZN(n430) );
  AND2_X1 U449 ( .A1(n416), .A2(n407), .ZN(n413) );
  INV_X1 U450 ( .A(KEYINPUT34), .ZN(n594) );
  INV_X1 U451 ( .A(G134), .ZN(n481) );
  NAND2_X1 U452 ( .A1(G237), .A2(G234), .ZN(n496) );
  AND2_X1 U453 ( .A1(n694), .A2(KEYINPUT41), .ZN(n387) );
  NAND2_X1 U454 ( .A1(n697), .A2(n391), .ZN(n390) );
  XNOR2_X1 U455 ( .A(n419), .B(n418), .ZN(n563) );
  INV_X1 U456 ( .A(KEYINPUT68), .ZN(n418) );
  NAND2_X1 U457 ( .A1(n351), .A2(n420), .ZN(n419) );
  OR2_X1 U458 ( .A1(G237), .A2(G902), .ZN(n493) );
  XNOR2_X1 U459 ( .A(n514), .B(n383), .ZN(n746) );
  XNOR2_X1 U460 ( .A(G128), .B(KEYINPUT94), .ZN(n516) );
  INV_X1 U461 ( .A(KEYINPUT23), .ZN(n518) );
  XNOR2_X1 U462 ( .A(G110), .B(G119), .ZN(n519) );
  XNOR2_X1 U463 ( .A(KEYINPUT7), .B(KEYINPUT9), .ZN(n535) );
  XNOR2_X1 U464 ( .A(n447), .B(n446), .ZN(n537) );
  INV_X1 U465 ( .A(KEYINPUT8), .ZN(n446) );
  NAND2_X1 U466 ( .A1(n754), .A2(G234), .ZN(n447) );
  AND2_X1 U467 ( .A1(n384), .A2(n360), .ZN(n400) );
  XNOR2_X1 U468 ( .A(n509), .B(n358), .ZN(n433) );
  XNOR2_X1 U469 ( .A(n395), .B(n479), .ZN(n717) );
  AND2_X1 U470 ( .A1(n752), .A2(n353), .ZN(n670) );
  NAND2_X1 U471 ( .A1(n609), .A2(n440), .ZN(n439) );
  AND2_X1 U472 ( .A1(n438), .A2(n437), .ZN(n436) );
  XNOR2_X1 U473 ( .A(KEYINPUT101), .B(G472), .ZN(n492) );
  INV_X1 U474 ( .A(KEYINPUT0), .ZN(n450) );
  BUF_X1 U475 ( .A(n562), .Z(n681) );
  XNOR2_X1 U476 ( .A(n377), .B(n453), .ZN(n363) );
  XNOR2_X1 U477 ( .A(n392), .B(KEYINPUT91), .ZN(n403) );
  XNOR2_X1 U478 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U479 ( .A(G122), .B(G104), .ZN(n463) );
  INV_X1 U480 ( .A(KEYINPUT42), .ZN(n443) );
  INV_X1 U481 ( .A(KEYINPUT35), .ZN(n370) );
  INV_X1 U482 ( .A(KEYINPUT32), .ZN(n451) );
  NAND2_X1 U483 ( .A1(n398), .A2(n397), .ZN(n411) );
  AND2_X1 U484 ( .A1(n452), .A2(n351), .ZN(n397) );
  XNOR2_X1 U485 ( .A(n611), .B(n610), .ZN(n612) );
  INV_X1 U486 ( .A(KEYINPUT86), .ZN(n610) );
  AND2_X1 U487 ( .A1(n641), .A2(n640), .ZN(n642) );
  XNOR2_X1 U488 ( .A(n407), .B(G140), .ZN(G42) );
  AND2_X1 U489 ( .A1(n364), .A2(KEYINPUT2), .ZN(n353) );
  XOR2_X1 U490 ( .A(n609), .B(n374), .Z(n354) );
  AND2_X1 U491 ( .A1(n621), .A2(n454), .ZN(n355) );
  AND2_X1 U492 ( .A1(n369), .A2(n368), .ZN(n356) );
  NAND2_X1 U493 ( .A1(G210), .A2(n493), .ZN(n357) );
  XOR2_X1 U494 ( .A(n504), .B(n515), .Z(n358) );
  OR2_X1 U495 ( .A1(n620), .A2(n619), .ZN(n359) );
  AND2_X1 U496 ( .A1(n432), .A2(n622), .ZN(n360) );
  XOR2_X1 U497 ( .A(KEYINPUT109), .B(n545), .Z(n361) );
  INV_X1 U498 ( .A(KEYINPUT41), .ZN(n391) );
  XNOR2_X1 U499 ( .A(KEYINPUT90), .B(n628), .ZN(n735) );
  XNOR2_X2 U500 ( .A(n362), .B(n361), .ZN(n375) );
  NAND2_X1 U501 ( .A1(n544), .A2(n659), .ZN(n362) );
  NAND2_X1 U502 ( .A1(n597), .A2(n386), .ZN(n385) );
  NAND2_X1 U503 ( .A1(n445), .A2(n574), .ZN(n444) );
  XNOR2_X1 U504 ( .A(n363), .B(n503), .ZN(n631) );
  NAND2_X1 U505 ( .A1(n400), .A2(n364), .ZN(n449) );
  NOR2_X1 U506 ( .A1(n364), .A2(n668), .ZN(n667) );
  NAND2_X1 U507 ( .A1(n364), .A2(n754), .ZN(n739) );
  XNOR2_X2 U508 ( .A(n402), .B(KEYINPUT45), .ZN(n364) );
  INV_X1 U509 ( .A(n613), .ZN(n366) );
  NAND2_X1 U510 ( .A1(n613), .A2(n594), .ZN(n369) );
  XNOR2_X2 U511 ( .A(n371), .B(n370), .ZN(n759) );
  NAND2_X1 U512 ( .A1(n373), .A2(n372), .ZN(n371) );
  INV_X1 U513 ( .A(n595), .ZN(n372) );
  NOR2_X2 U514 ( .A1(n375), .A2(n761), .ZN(n556) );
  XNOR2_X1 U515 ( .A(n375), .B(G131), .ZN(n760) );
  NAND2_X1 U516 ( .A1(n376), .A2(n695), .ZN(n530) );
  NAND2_X1 U517 ( .A1(n376), .A2(n408), .ZN(n559) );
  NOR2_X2 U518 ( .A1(n529), .A2(n528), .ZN(n376) );
  XNOR2_X1 U519 ( .A(n377), .B(n740), .ZN(n395) );
  NAND2_X1 U520 ( .A1(n657), .A2(n576), .ZN(n379) );
  NAND2_X1 U521 ( .A1(n578), .A2(n657), .ZN(n380) );
  XNOR2_X2 U522 ( .A(n575), .B(KEYINPUT79), .ZN(n657) );
  NOR2_X1 U523 ( .A1(n731), .A2(G902), .ZN(n527) );
  XNOR2_X1 U524 ( .A(n746), .B(n381), .ZN(n731) );
  XNOR2_X1 U525 ( .A(n382), .B(n522), .ZN(n381) );
  XNOR2_X1 U526 ( .A(n521), .B(n520), .ZN(n382) );
  INV_X1 U527 ( .A(n515), .ZN(n383) );
  AND2_X1 U528 ( .A1(n384), .A2(n432), .ZN(n752) );
  NAND2_X1 U529 ( .A1(n695), .A2(n694), .ZN(n698) );
  XNOR2_X2 U530 ( .A(n565), .B(KEYINPUT38), .ZN(n695) );
  NAND2_X1 U531 ( .A1(n698), .A2(n391), .ZN(n389) );
  AND2_X1 U532 ( .A1(n695), .A2(n387), .ZN(n386) );
  XNOR2_X2 U533 ( .A(G113), .B(KEYINPUT71), .ZN(n392) );
  NAND2_X1 U534 ( .A1(n393), .A2(n609), .ZN(n581) );
  NOR2_X1 U535 ( .A1(n394), .A2(n564), .ZN(n393) );
  NAND2_X1 U536 ( .A1(n563), .A2(n694), .ZN(n394) );
  NOR2_X1 U537 ( .A1(n608), .A2(n677), .ZN(n399) );
  AND2_X1 U538 ( .A1(n399), .A2(n410), .ZN(n653) );
  XNOR2_X2 U539 ( .A(n530), .B(KEYINPUT39), .ZN(n544) );
  NAND2_X1 U540 ( .A1(n571), .A2(n570), .ZN(n580) );
  XNOR2_X1 U541 ( .A(n626), .B(n627), .ZN(n629) );
  XNOR2_X1 U542 ( .A(n718), .B(n719), .ZN(n720) );
  NAND2_X1 U543 ( .A1(n759), .A2(n596), .ZN(n435) );
  NOR2_X2 U544 ( .A1(n762), .A2(n653), .ZN(n606) );
  OR2_X1 U545 ( .A1(n682), .A2(n351), .ZN(n406) );
  INV_X1 U546 ( .A(n408), .ZN(n565) );
  NAND2_X1 U547 ( .A1(n408), .A2(n694), .ZN(n573) );
  XNOR2_X2 U548 ( .A(n480), .B(n357), .ZN(n408) );
  OR2_X1 U549 ( .A1(n584), .A2(n408), .ZN(n407) );
  XNOR2_X1 U550 ( .A(n409), .B(n741), .ZN(n742) );
  NOR2_X1 U551 ( .A1(n682), .A2(n603), .ZN(n410) );
  NAND2_X1 U552 ( .A1(n579), .A2(KEYINPUT48), .ZN(n416) );
  NAND2_X1 U553 ( .A1(n414), .A2(n415), .ZN(n412) );
  NOR2_X1 U554 ( .A1(n579), .A2(KEYINPUT48), .ZN(n414) );
  INV_X1 U555 ( .A(n580), .ZN(n415) );
  NAND2_X1 U556 ( .A1(n580), .A2(KEYINPUT48), .ZN(n417) );
  XNOR2_X1 U557 ( .A(n547), .B(KEYINPUT69), .ZN(n420) );
  XNOR2_X2 U558 ( .A(n422), .B(n450), .ZN(n599) );
  XNOR2_X1 U559 ( .A(n606), .B(n427), .ZN(n426) );
  INV_X1 U560 ( .A(KEYINPUT87), .ZN(n427) );
  INV_X1 U561 ( .A(n656), .ZN(n428) );
  NAND2_X1 U562 ( .A1(n431), .A2(n569), .ZN(n665) );
  XNOR2_X1 U563 ( .A(n566), .B(KEYINPUT36), .ZN(n431) );
  XNOR2_X1 U564 ( .A(n433), .B(n503), .ZN(n723) );
  NAND2_X1 U565 ( .A1(n617), .A2(n442), .ZN(n437) );
  AND2_X1 U566 ( .A1(n682), .A2(n441), .ZN(n440) );
  INV_X1 U567 ( .A(n593), .ZN(n442) );
  INV_X1 U568 ( .A(n692), .ZN(n445) );
  XNOR2_X1 U569 ( .A(n554), .B(KEYINPUT108), .ZN(n574) );
  INV_X1 U570 ( .A(n599), .ZN(n613) );
  INV_X1 U571 ( .A(n670), .ZN(n625) );
  XOR2_X1 U572 ( .A(n491), .B(n490), .Z(n453) );
  AND2_X1 U573 ( .A1(n643), .A2(n359), .ZN(n454) );
  INV_X1 U574 ( .A(KEYINPUT107), .ZN(n548) );
  XNOR2_X1 U575 ( .A(n549), .B(n548), .ZN(n550) );
  XNOR2_X1 U576 ( .A(n519), .B(n518), .ZN(n520) );
  AND2_X1 U577 ( .A1(n597), .A2(n678), .ZN(n598) );
  XNOR2_X1 U578 ( .A(n466), .B(n465), .ZN(n531) );
  XNOR2_X1 U579 ( .A(n631), .B(n632), .ZN(n633) );
  XNOR2_X1 U580 ( .A(n733), .B(n732), .ZN(n734) );
  NAND2_X1 U581 ( .A1(n489), .A2(G214), .ZN(n455) );
  XNOR2_X1 U582 ( .A(n455), .B(n514), .ZN(n456) );
  XOR2_X1 U583 ( .A(KEYINPUT67), .B(G131), .Z(n486) );
  XOR2_X1 U584 ( .A(n456), .B(n486), .Z(n466) );
  XOR2_X1 U585 ( .A(KEYINPUT97), .B(G140), .Z(n458) );
  XNOR2_X1 U586 ( .A(n458), .B(n457), .ZN(n462) );
  XOR2_X1 U587 ( .A(KEYINPUT12), .B(KEYINPUT98), .Z(n460) );
  XNOR2_X1 U588 ( .A(KEYINPUT11), .B(KEYINPUT99), .ZN(n459) );
  XNOR2_X1 U589 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U590 ( .A(n462), .B(n461), .ZN(n464) );
  NAND2_X1 U591 ( .A1(KEYINPUT3), .A2(n467), .ZN(n470) );
  NAND2_X1 U592 ( .A1(n468), .A2(G119), .ZN(n469) );
  NAND2_X1 U593 ( .A1(n470), .A2(n469), .ZN(n471) );
  NAND2_X1 U594 ( .A1(G224), .A2(n754), .ZN(n472) );
  XNOR2_X1 U595 ( .A(n473), .B(n472), .ZN(n474) );
  XOR2_X1 U596 ( .A(n474), .B(KEYINPUT17), .Z(n478) );
  INV_X1 U597 ( .A(n475), .ZN(n476) );
  XNOR2_X1 U598 ( .A(n482), .B(n476), .ZN(n477) );
  XNOR2_X1 U599 ( .A(n478), .B(n477), .ZN(n479) );
  NAND2_X1 U600 ( .A1(n482), .A2(n481), .ZN(n485) );
  XNOR2_X1 U601 ( .A(G143), .B(G128), .ZN(n483) );
  NAND2_X1 U602 ( .A1(G134), .A2(n483), .ZN(n484) );
  NAND2_X1 U603 ( .A1(n485), .A2(n484), .ZN(n534) );
  XNOR2_X1 U604 ( .A(n488), .B(n487), .ZN(n491) );
  NAND2_X1 U605 ( .A1(n489), .A2(G210), .ZN(n490) );
  NOR2_X2 U606 ( .A1(G902), .A2(n631), .ZN(n561) );
  NAND2_X1 U607 ( .A1(G214), .A2(n493), .ZN(n694) );
  NAND2_X1 U608 ( .A1(n603), .A2(n694), .ZN(n495) );
  XOR2_X1 U609 ( .A(KEYINPUT30), .B(KEYINPUT104), .Z(n494) );
  XNOR2_X1 U610 ( .A(n495), .B(n494), .ZN(n502) );
  XNOR2_X1 U611 ( .A(n496), .B(KEYINPUT92), .ZN(n497) );
  XNOR2_X1 U612 ( .A(KEYINPUT14), .B(n497), .ZN(n499) );
  NAND2_X1 U613 ( .A1(G952), .A2(n499), .ZN(n709) );
  NOR2_X1 U614 ( .A1(G953), .A2(n709), .ZN(n498) );
  XNOR2_X1 U615 ( .A(KEYINPUT93), .B(n498), .ZN(n588) );
  NAND2_X1 U616 ( .A1(G902), .A2(n499), .ZN(n586) );
  NOR2_X1 U617 ( .A1(G900), .A2(n586), .ZN(n500) );
  NAND2_X1 U618 ( .A1(G953), .A2(n500), .ZN(n501) );
  NAND2_X1 U619 ( .A1(n588), .A2(n501), .ZN(n546) );
  NAND2_X1 U620 ( .A1(n502), .A2(n546), .ZN(n529) );
  NAND2_X1 U621 ( .A1(G227), .A2(n754), .ZN(n506) );
  XNOR2_X1 U622 ( .A(n508), .B(n507), .ZN(n509) );
  NOR2_X1 U623 ( .A1(G902), .A2(n723), .ZN(n511) );
  XNOR2_X1 U624 ( .A(KEYINPUT70), .B(G469), .ZN(n510) );
  NAND2_X1 U625 ( .A1(G234), .A2(n623), .ZN(n512) );
  XNOR2_X1 U626 ( .A(KEYINPUT20), .B(n512), .ZN(n523) );
  NAND2_X1 U627 ( .A1(G221), .A2(n523), .ZN(n513) );
  XOR2_X1 U628 ( .A(KEYINPUT21), .B(n513), .Z(n678) );
  NAND2_X1 U629 ( .A1(n537), .A2(G221), .ZN(n522) );
  XOR2_X1 U630 ( .A(KEYINPUT24), .B(KEYINPUT76), .Z(n517) );
  XNOR2_X1 U631 ( .A(n517), .B(n516), .ZN(n521) );
  XOR2_X1 U632 ( .A(KEYINPUT25), .B(KEYINPUT95), .Z(n525) );
  NAND2_X1 U633 ( .A1(n523), .A2(G217), .ZN(n524) );
  XNOR2_X1 U634 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U635 ( .A(n527), .B(n526), .ZN(n601) );
  NAND2_X1 U636 ( .A1(n678), .A2(n601), .ZN(n592) );
  NOR2_X1 U637 ( .A1(n568), .A2(n592), .ZN(n614) );
  XNOR2_X1 U638 ( .A(n614), .B(KEYINPUT103), .ZN(n528) );
  XNOR2_X1 U639 ( .A(KEYINPUT13), .B(G475), .ZN(n533) );
  NOR2_X1 U640 ( .A1(G902), .A2(n531), .ZN(n532) );
  XNOR2_X1 U641 ( .A(n533), .B(n532), .ZN(n555) );
  XNOR2_X1 U642 ( .A(n535), .B(KEYINPUT100), .ZN(n536) );
  XOR2_X1 U643 ( .A(n534), .B(n536), .Z(n539) );
  NAND2_X1 U644 ( .A1(G217), .A2(n537), .ZN(n538) );
  XNOR2_X1 U645 ( .A(n539), .B(n538), .ZN(n540) );
  XOR2_X1 U646 ( .A(n541), .B(n540), .Z(n637) );
  NOR2_X1 U647 ( .A1(n637), .A2(G902), .ZN(n542) );
  XNOR2_X1 U648 ( .A(G478), .B(n542), .ZN(n558) );
  NOR2_X1 U649 ( .A1(n555), .A2(n558), .ZN(n661) );
  NAND2_X1 U650 ( .A1(n544), .A2(n661), .ZN(n543) );
  XNOR2_X1 U651 ( .A(n543), .B(KEYINPUT111), .ZN(n758) );
  INV_X1 U652 ( .A(KEYINPUT84), .ZN(n585) );
  NAND2_X1 U653 ( .A1(n555), .A2(n558), .ZN(n564) );
  INV_X1 U654 ( .A(n564), .ZN(n659) );
  XOR2_X1 U655 ( .A(KEYINPUT110), .B(KEYINPUT40), .Z(n545) );
  NAND2_X1 U656 ( .A1(n546), .A2(n678), .ZN(n547) );
  INV_X1 U657 ( .A(KEYINPUT28), .ZN(n549) );
  XNOR2_X1 U658 ( .A(n551), .B(n550), .ZN(n553) );
  XNOR2_X1 U659 ( .A(n568), .B(KEYINPUT106), .ZN(n552) );
  NOR2_X1 U660 ( .A1(n553), .A2(n552), .ZN(n554) );
  INV_X1 U661 ( .A(n555), .ZN(n557) );
  NAND2_X1 U662 ( .A1(n558), .A2(n557), .ZN(n697) );
  XNOR2_X1 U663 ( .A(n556), .B(KEYINPUT46), .ZN(n571) );
  OR2_X1 U664 ( .A1(n558), .A2(n557), .ZN(n595) );
  XOR2_X1 U665 ( .A(KEYINPUT105), .B(n559), .Z(n560) );
  NOR2_X1 U666 ( .A1(n595), .A2(n560), .ZN(n656) );
  NOR2_X1 U667 ( .A1(n565), .A2(n581), .ZN(n566) );
  XNOR2_X2 U668 ( .A(n568), .B(n567), .ZN(n682) );
  INV_X1 U669 ( .A(n682), .ZN(n604) );
  XOR2_X1 U670 ( .A(KEYINPUT89), .B(n604), .Z(n602) );
  INV_X1 U671 ( .A(n602), .ZN(n569) );
  INV_X1 U672 ( .A(n699), .ZN(n576) );
  XOR2_X1 U673 ( .A(KEYINPUT19), .B(KEYINPUT65), .Z(n572) );
  NAND2_X1 U674 ( .A1(n574), .A2(n591), .ZN(n575) );
  XNOR2_X1 U675 ( .A(n699), .B(KEYINPUT82), .ZN(n620) );
  NOR2_X1 U676 ( .A1(KEYINPUT47), .A2(n620), .ZN(n577) );
  XNOR2_X1 U677 ( .A(KEYINPUT74), .B(n577), .ZN(n578) );
  XNOR2_X1 U678 ( .A(KEYINPUT102), .B(n581), .ZN(n582) );
  NOR2_X1 U679 ( .A1(n682), .A2(n582), .ZN(n583) );
  XNOR2_X1 U680 ( .A(n583), .B(KEYINPUT43), .ZN(n584) );
  NOR2_X1 U681 ( .A1(G898), .A2(n754), .ZN(n743) );
  INV_X1 U682 ( .A(n586), .ZN(n587) );
  NAND2_X1 U683 ( .A1(n743), .A2(n587), .ZN(n589) );
  NAND2_X1 U684 ( .A1(n589), .A2(n588), .ZN(n590) );
  INV_X1 U685 ( .A(n592), .ZN(n683) );
  XNOR2_X1 U686 ( .A(KEYINPUT33), .B(KEYINPUT72), .ZN(n593) );
  INV_X1 U687 ( .A(KEYINPUT44), .ZN(n596) );
  INV_X1 U688 ( .A(n697), .ZN(n597) );
  INV_X1 U689 ( .A(n351), .ZN(n677) );
  NAND2_X1 U690 ( .A1(n606), .A2(n759), .ZN(n607) );
  NAND2_X1 U691 ( .A1(n607), .A2(KEYINPUT44), .ZN(n621) );
  INV_X1 U692 ( .A(n681), .ZN(n616) );
  NAND2_X1 U693 ( .A1(n614), .A2(n366), .ZN(n615) );
  NOR2_X1 U694 ( .A1(n616), .A2(n615), .ZN(n648) );
  NOR2_X1 U695 ( .A1(n681), .A2(n617), .ZN(n688) );
  NAND2_X1 U696 ( .A1(n599), .A2(n688), .ZN(n618) );
  XNOR2_X1 U697 ( .A(n618), .B(KEYINPUT31), .ZN(n662) );
  NOR2_X1 U698 ( .A1(n648), .A2(n662), .ZN(n619) );
  INV_X1 U699 ( .A(KEYINPUT2), .ZN(n666) );
  OR2_X1 U700 ( .A1(n623), .A2(n666), .ZN(n624) );
  NAND2_X1 U701 ( .A1(n729), .A2(G475), .ZN(n626) );
  NOR2_X1 U702 ( .A1(G952), .A2(n754), .ZN(n628) );
  NOR2_X2 U703 ( .A1(n629), .A2(n735), .ZN(n630) );
  XNOR2_X1 U704 ( .A(n630), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U705 ( .A1(n729), .A2(G472), .ZN(n634) );
  XOR2_X1 U706 ( .A(KEYINPUT62), .B(KEYINPUT88), .Z(n632) );
  XNOR2_X1 U707 ( .A(n634), .B(n633), .ZN(n635) );
  NAND2_X1 U708 ( .A1(n635), .A2(n640), .ZN(n636) );
  XNOR2_X1 U709 ( .A(n636), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U710 ( .A1(G478), .A2(n729), .ZN(n639) );
  INV_X1 U711 ( .A(n637), .ZN(n638) );
  XNOR2_X1 U712 ( .A(n639), .B(n638), .ZN(n641) );
  INV_X1 U713 ( .A(n735), .ZN(n640) );
  XNOR2_X1 U714 ( .A(n642), .B(KEYINPUT124), .ZN(G63) );
  XNOR2_X1 U715 ( .A(G101), .B(KEYINPUT112), .ZN(n644) );
  XNOR2_X1 U716 ( .A(n644), .B(n643), .ZN(G3) );
  NAND2_X1 U717 ( .A1(n648), .A2(n659), .ZN(n645) );
  XNOR2_X1 U718 ( .A(n645), .B(G104), .ZN(G6) );
  XOR2_X1 U719 ( .A(KEYINPUT115), .B(KEYINPUT27), .Z(n647) );
  XNOR2_X1 U720 ( .A(KEYINPUT113), .B(KEYINPUT114), .ZN(n646) );
  XNOR2_X1 U721 ( .A(n647), .B(n646), .ZN(n652) );
  XNOR2_X1 U722 ( .A(G107), .B(KEYINPUT26), .ZN(n650) );
  NAND2_X1 U723 ( .A1(n661), .A2(n648), .ZN(n649) );
  XNOR2_X1 U724 ( .A(n650), .B(n649), .ZN(n651) );
  XNOR2_X1 U725 ( .A(n652), .B(n651), .ZN(G9) );
  XOR2_X1 U726 ( .A(G110), .B(n653), .Z(G12) );
  XOR2_X1 U727 ( .A(G128), .B(KEYINPUT29), .Z(n655) );
  NAND2_X1 U728 ( .A1(n657), .A2(n661), .ZN(n654) );
  XNOR2_X1 U729 ( .A(n655), .B(n654), .ZN(G30) );
  XOR2_X1 U730 ( .A(G143), .B(n656), .Z(G45) );
  NAND2_X1 U731 ( .A1(n659), .A2(n657), .ZN(n658) );
  XNOR2_X1 U732 ( .A(G146), .B(n658), .ZN(G48) );
  NAND2_X1 U733 ( .A1(n662), .A2(n659), .ZN(n660) );
  XNOR2_X1 U734 ( .A(n660), .B(G113), .ZN(G15) );
  NAND2_X1 U735 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U736 ( .A(n663), .B(G116), .ZN(G18) );
  XOR2_X1 U737 ( .A(G125), .B(KEYINPUT37), .Z(n664) );
  XNOR2_X1 U738 ( .A(n665), .B(n664), .ZN(G27) );
  XNOR2_X1 U739 ( .A(KEYINPUT81), .B(n666), .ZN(n668) );
  XNOR2_X1 U740 ( .A(n667), .B(KEYINPUT83), .ZN(n672) );
  NOR2_X1 U741 ( .A1(n752), .A2(n668), .ZN(n669) );
  NOR2_X1 U742 ( .A1(n670), .A2(n669), .ZN(n671) );
  NAND2_X1 U743 ( .A1(n672), .A2(n671), .ZN(n676) );
  NOR2_X1 U744 ( .A1(n704), .A2(n692), .ZN(n673) );
  XNOR2_X1 U745 ( .A(KEYINPUT120), .B(n673), .ZN(n674) );
  NOR2_X1 U746 ( .A1(G953), .A2(n674), .ZN(n675) );
  NAND2_X1 U747 ( .A1(n676), .A2(n675), .ZN(n712) );
  NOR2_X1 U748 ( .A1(n678), .A2(n677), .ZN(n679) );
  XNOR2_X1 U749 ( .A(n679), .B(KEYINPUT49), .ZN(n680) );
  NAND2_X1 U750 ( .A1(n681), .A2(n680), .ZN(n686) );
  NOR2_X1 U751 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X1 U752 ( .A(n684), .B(KEYINPUT50), .ZN(n685) );
  NOR2_X1 U753 ( .A1(n686), .A2(n685), .ZN(n687) );
  NOR2_X1 U754 ( .A1(n688), .A2(n687), .ZN(n689) );
  XOR2_X1 U755 ( .A(KEYINPUT51), .B(n689), .Z(n690) );
  XNOR2_X1 U756 ( .A(n690), .B(KEYINPUT116), .ZN(n691) );
  NOR2_X1 U757 ( .A1(n692), .A2(n691), .ZN(n693) );
  XOR2_X1 U758 ( .A(KEYINPUT117), .B(n693), .Z(n706) );
  NOR2_X1 U759 ( .A1(n695), .A2(n694), .ZN(n696) );
  NOR2_X1 U760 ( .A1(n697), .A2(n696), .ZN(n702) );
  NOR2_X1 U761 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U762 ( .A(n700), .B(KEYINPUT118), .ZN(n701) );
  NOR2_X1 U763 ( .A1(n702), .A2(n701), .ZN(n703) );
  NOR2_X1 U764 ( .A1(n704), .A2(n703), .ZN(n705) );
  NOR2_X1 U765 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U766 ( .A(n707), .B(KEYINPUT52), .ZN(n708) );
  NOR2_X1 U767 ( .A1(n709), .A2(n708), .ZN(n710) );
  XOR2_X1 U768 ( .A(KEYINPUT119), .B(n710), .Z(n711) );
  NOR2_X1 U769 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U770 ( .A(KEYINPUT53), .B(n713), .ZN(G75) );
  XOR2_X1 U771 ( .A(KEYINPUT80), .B(KEYINPUT55), .Z(n715) );
  XNOR2_X1 U772 ( .A(KEYINPUT121), .B(KEYINPUT54), .ZN(n714) );
  XNOR2_X1 U773 ( .A(n715), .B(n714), .ZN(n716) );
  XOR2_X1 U774 ( .A(n717), .B(n716), .Z(n719) );
  NAND2_X1 U775 ( .A1(n729), .A2(G210), .ZN(n718) );
  NOR2_X2 U776 ( .A1(n720), .A2(n735), .ZN(n722) );
  XNOR2_X1 U777 ( .A(KEYINPUT122), .B(KEYINPUT56), .ZN(n721) );
  XNOR2_X1 U778 ( .A(n722), .B(n721), .ZN(G51) );
  XOR2_X1 U779 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n725) );
  XNOR2_X1 U780 ( .A(n723), .B(KEYINPUT123), .ZN(n724) );
  XNOR2_X1 U781 ( .A(n725), .B(n724), .ZN(n727) );
  NAND2_X1 U782 ( .A1(n729), .A2(G469), .ZN(n726) );
  XOR2_X1 U783 ( .A(n727), .B(n726), .Z(n728) );
  NOR2_X1 U784 ( .A1(n735), .A2(n728), .ZN(G54) );
  NAND2_X1 U785 ( .A1(n729), .A2(G217), .ZN(n733) );
  INV_X1 U786 ( .A(KEYINPUT125), .ZN(n730) );
  XNOR2_X1 U787 ( .A(n731), .B(n730), .ZN(n732) );
  NOR2_X1 U788 ( .A1(n735), .A2(n734), .ZN(G66) );
  NAND2_X1 U789 ( .A1(G953), .A2(G224), .ZN(n736) );
  XNOR2_X1 U790 ( .A(KEYINPUT61), .B(n736), .ZN(n737) );
  NAND2_X1 U791 ( .A1(n737), .A2(G898), .ZN(n738) );
  NAND2_X1 U792 ( .A1(n739), .A2(n738), .ZN(n745) );
  XNOR2_X1 U793 ( .A(n740), .B(G101), .ZN(n741) );
  NOR2_X1 U794 ( .A1(n743), .A2(n742), .ZN(n744) );
  XNOR2_X1 U795 ( .A(n745), .B(n744), .ZN(G69) );
  XOR2_X1 U796 ( .A(KEYINPUT4), .B(n746), .Z(n747) );
  XOR2_X1 U797 ( .A(n748), .B(n747), .Z(n753) );
  XOR2_X1 U798 ( .A(n753), .B(KEYINPUT126), .Z(n749) );
  XNOR2_X1 U799 ( .A(G227), .B(n749), .ZN(n750) );
  NAND2_X1 U800 ( .A1(G900), .A2(n750), .ZN(n751) );
  NAND2_X1 U801 ( .A1(n751), .A2(G953), .ZN(n757) );
  XNOR2_X1 U802 ( .A(n753), .B(n752), .ZN(n755) );
  NAND2_X1 U803 ( .A1(n755), .A2(n754), .ZN(n756) );
  NAND2_X1 U804 ( .A1(n757), .A2(n756), .ZN(G72) );
  XOR2_X1 U805 ( .A(G134), .B(n758), .Z(G36) );
  XNOR2_X1 U806 ( .A(G122), .B(n759), .ZN(G24) );
  XNOR2_X1 U807 ( .A(n760), .B(KEYINPUT127), .ZN(G33) );
  XOR2_X1 U808 ( .A(n352), .B(G137), .Z(G39) );
  XOR2_X1 U809 ( .A(n762), .B(G119), .Z(G21) );
endmodule

